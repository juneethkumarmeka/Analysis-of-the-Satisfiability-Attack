module basic_500_3000_500_60_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_291,In_288);
nor U1 (N_1,In_417,In_92);
nor U2 (N_2,In_257,In_167);
nor U3 (N_3,In_168,In_388);
and U4 (N_4,In_426,In_409);
or U5 (N_5,In_278,In_85);
xnor U6 (N_6,In_470,In_196);
nor U7 (N_7,In_370,In_10);
nor U8 (N_8,In_82,In_272);
and U9 (N_9,In_390,In_343);
and U10 (N_10,In_428,In_50);
nand U11 (N_11,In_273,In_57);
nand U12 (N_12,In_58,In_33);
nor U13 (N_13,In_171,In_311);
xnor U14 (N_14,In_448,In_460);
xor U15 (N_15,In_125,In_115);
nand U16 (N_16,In_255,In_131);
and U17 (N_17,In_69,In_297);
and U18 (N_18,In_239,In_3);
or U19 (N_19,In_78,In_52);
or U20 (N_20,In_165,In_120);
or U21 (N_21,In_155,In_379);
and U22 (N_22,In_292,In_193);
or U23 (N_23,In_400,In_24);
nand U24 (N_24,In_175,In_478);
and U25 (N_25,In_84,In_282);
and U26 (N_26,In_399,In_389);
or U27 (N_27,In_124,In_268);
nor U28 (N_28,In_462,In_469);
nor U29 (N_29,In_453,In_35);
nor U30 (N_30,In_54,In_161);
nor U31 (N_31,In_75,In_364);
and U32 (N_32,In_422,In_396);
and U33 (N_33,In_67,In_227);
or U34 (N_34,In_357,In_318);
xor U35 (N_35,In_481,In_435);
nand U36 (N_36,In_283,In_112);
nor U37 (N_37,In_184,In_334);
and U38 (N_38,In_139,In_466);
or U39 (N_39,In_19,In_488);
nor U40 (N_40,In_181,In_247);
and U41 (N_41,In_178,In_95);
nand U42 (N_42,In_1,In_274);
and U43 (N_43,In_441,In_148);
or U44 (N_44,In_46,In_219);
nand U45 (N_45,In_495,In_89);
nor U46 (N_46,In_374,In_285);
nor U47 (N_47,In_208,In_450);
and U48 (N_48,In_499,In_60);
nand U49 (N_49,In_130,In_62);
or U50 (N_50,In_264,In_382);
nor U51 (N_51,In_313,N_35);
and U52 (N_52,In_280,N_28);
xnor U53 (N_53,In_375,In_156);
or U54 (N_54,N_46,In_98);
or U55 (N_55,In_380,In_126);
nor U56 (N_56,N_21,N_34);
or U57 (N_57,In_185,In_80);
and U58 (N_58,In_199,In_250);
or U59 (N_59,In_397,N_3);
nand U60 (N_60,In_29,In_197);
or U61 (N_61,N_29,N_31);
or U62 (N_62,In_147,In_214);
nor U63 (N_63,In_294,In_73);
nor U64 (N_64,N_49,In_203);
nand U65 (N_65,In_207,In_319);
or U66 (N_66,In_355,In_103);
and U67 (N_67,In_480,In_277);
or U68 (N_68,In_220,In_157);
and U69 (N_69,In_437,In_293);
or U70 (N_70,In_325,In_232);
xor U71 (N_71,In_238,In_320);
or U72 (N_72,N_33,In_408);
and U73 (N_73,In_217,In_300);
and U74 (N_74,In_269,In_496);
nor U75 (N_75,In_132,In_306);
or U76 (N_76,In_83,In_482);
nor U77 (N_77,In_43,In_471);
or U78 (N_78,In_420,In_473);
or U79 (N_79,In_424,In_252);
nand U80 (N_80,In_498,In_258);
nand U81 (N_81,In_403,In_367);
xnor U82 (N_82,In_218,In_129);
or U83 (N_83,In_114,In_472);
nor U84 (N_84,N_25,In_381);
and U85 (N_85,In_287,In_34);
nor U86 (N_86,In_198,In_106);
and U87 (N_87,In_241,In_51);
and U88 (N_88,N_45,In_386);
nand U89 (N_89,In_121,In_432);
nor U90 (N_90,In_180,In_192);
nor U91 (N_91,In_242,N_11);
nand U92 (N_92,In_378,In_463);
or U93 (N_93,In_225,In_135);
nor U94 (N_94,In_249,In_159);
and U95 (N_95,In_342,In_123);
nand U96 (N_96,In_117,In_359);
or U97 (N_97,In_183,In_410);
nand U98 (N_98,In_205,N_42);
nand U99 (N_99,In_2,In_200);
xor U100 (N_100,In_204,N_70);
and U101 (N_101,In_336,In_497);
nand U102 (N_102,In_284,In_385);
and U103 (N_103,In_328,In_394);
and U104 (N_104,In_493,In_245);
nand U105 (N_105,In_353,In_163);
nand U106 (N_106,In_93,In_454);
nand U107 (N_107,In_270,In_419);
nand U108 (N_108,In_455,In_337);
or U109 (N_109,In_63,In_8);
nand U110 (N_110,In_186,In_66);
nand U111 (N_111,In_362,N_60);
and U112 (N_112,In_392,In_363);
nand U113 (N_113,N_88,In_176);
nand U114 (N_114,In_369,In_254);
nor U115 (N_115,In_486,N_19);
nand U116 (N_116,N_89,N_95);
and U117 (N_117,In_201,In_423);
and U118 (N_118,In_299,N_10);
and U119 (N_119,N_27,In_36);
or U120 (N_120,N_90,In_136);
nor U121 (N_121,In_223,In_271);
nand U122 (N_122,In_345,N_0);
nand U123 (N_123,In_401,N_99);
nand U124 (N_124,N_20,In_23);
or U125 (N_125,N_69,In_308);
nor U126 (N_126,In_251,In_240);
nor U127 (N_127,In_301,In_231);
nor U128 (N_128,N_36,N_96);
nor U129 (N_129,In_206,In_361);
or U130 (N_130,In_338,In_351);
and U131 (N_131,In_0,In_279);
or U132 (N_132,In_86,In_489);
or U133 (N_133,In_237,In_28);
nor U134 (N_134,In_127,In_354);
and U135 (N_135,In_260,In_166);
and U136 (N_136,N_32,In_158);
and U137 (N_137,N_52,In_210);
and U138 (N_138,In_314,In_194);
nand U139 (N_139,In_25,In_31);
nand U140 (N_140,In_76,In_465);
or U141 (N_141,In_137,In_138);
nor U142 (N_142,N_63,N_26);
or U143 (N_143,In_53,In_246);
and U144 (N_144,In_302,In_459);
nand U145 (N_145,In_267,In_187);
nand U146 (N_146,In_87,N_71);
or U147 (N_147,N_57,N_81);
or U148 (N_148,In_234,N_6);
nand U149 (N_149,In_290,In_236);
or U150 (N_150,In_329,N_4);
or U151 (N_151,N_68,In_324);
nand U152 (N_152,In_235,In_474);
or U153 (N_153,N_147,N_98);
nor U154 (N_154,In_48,In_339);
or U155 (N_155,N_59,In_407);
nand U156 (N_156,In_310,In_341);
or U157 (N_157,In_105,N_116);
and U158 (N_158,In_377,In_326);
nand U159 (N_159,In_449,In_6);
nor U160 (N_160,N_104,In_169);
nand U161 (N_161,In_406,N_48);
nor U162 (N_162,In_384,N_91);
or U163 (N_163,In_261,In_77);
and U164 (N_164,N_73,In_321);
or U165 (N_165,N_114,N_144);
nor U166 (N_166,In_146,In_430);
nor U167 (N_167,N_117,In_366);
nor U168 (N_168,In_438,In_295);
nand U169 (N_169,In_412,N_133);
nor U170 (N_170,In_4,In_27);
nor U171 (N_171,In_42,N_37);
or U172 (N_172,In_492,In_13);
nor U173 (N_173,In_11,In_215);
nand U174 (N_174,In_372,In_228);
nand U175 (N_175,In_416,N_51);
nor U176 (N_176,In_134,N_94);
xnor U177 (N_177,In_40,In_177);
or U178 (N_178,N_138,In_212);
nor U179 (N_179,In_172,In_111);
nor U180 (N_180,In_26,In_104);
or U181 (N_181,In_477,In_182);
nand U182 (N_182,N_41,In_464);
nand U183 (N_183,In_128,In_70);
nor U184 (N_184,N_83,N_137);
and U185 (N_185,In_312,N_64);
nor U186 (N_186,In_356,In_61);
nor U187 (N_187,N_78,N_107);
or U188 (N_188,In_393,In_253);
or U189 (N_189,N_7,In_179);
xor U190 (N_190,In_335,In_444);
nor U191 (N_191,In_233,N_122);
and U192 (N_192,In_440,In_32);
or U193 (N_193,In_439,N_124);
and U194 (N_194,N_86,N_56);
and U195 (N_195,In_226,In_487);
nand U196 (N_196,N_47,In_445);
nor U197 (N_197,N_67,In_209);
or U198 (N_198,In_160,In_371);
nand U199 (N_199,N_128,In_222);
xnor U200 (N_200,In_350,In_485);
or U201 (N_201,N_40,N_76);
nor U202 (N_202,N_184,In_211);
and U203 (N_203,In_418,In_373);
or U204 (N_204,In_387,In_262);
nand U205 (N_205,In_88,In_309);
nor U206 (N_206,In_140,In_44);
and U207 (N_207,N_139,N_166);
or U208 (N_208,N_157,In_174);
or U209 (N_209,In_102,N_74);
nand U210 (N_210,In_59,In_479);
and U211 (N_211,In_447,N_97);
nand U212 (N_212,N_75,In_173);
nor U213 (N_213,N_53,In_298);
nor U214 (N_214,N_2,In_118);
nor U215 (N_215,N_87,In_243);
and U216 (N_216,N_119,N_143);
or U217 (N_217,In_344,In_376);
and U218 (N_218,In_276,N_177);
and U219 (N_219,N_171,N_188);
nor U220 (N_220,In_141,N_54);
nand U221 (N_221,N_131,In_368);
or U222 (N_222,In_39,In_195);
and U223 (N_223,In_151,In_49);
nor U224 (N_224,N_84,N_55);
nand U225 (N_225,In_286,In_16);
nand U226 (N_226,In_133,In_452);
and U227 (N_227,N_142,In_15);
and U228 (N_228,In_467,N_187);
nor U229 (N_229,N_165,In_433);
nor U230 (N_230,N_161,In_490);
xnor U231 (N_231,In_391,In_259);
nand U232 (N_232,In_427,N_180);
nor U233 (N_233,In_162,N_1);
nand U234 (N_234,In_109,In_152);
nand U235 (N_235,In_170,In_64);
nand U236 (N_236,N_162,N_113);
nor U237 (N_237,In_116,In_425);
nand U238 (N_238,In_107,In_451);
or U239 (N_239,N_155,N_38);
or U240 (N_240,N_39,In_21);
nand U241 (N_241,In_405,N_109);
nand U242 (N_242,N_18,In_414);
or U243 (N_243,N_135,In_14);
or U244 (N_244,N_154,In_189);
nand U245 (N_245,In_191,N_80);
or U246 (N_246,N_24,N_121);
xnor U247 (N_247,N_102,N_58);
or U248 (N_248,N_199,N_100);
nand U249 (N_249,N_141,In_110);
nand U250 (N_250,N_112,N_243);
or U251 (N_251,In_332,N_149);
or U252 (N_252,In_99,N_140);
nor U253 (N_253,N_111,In_244);
nand U254 (N_254,In_30,N_181);
nor U255 (N_255,N_220,In_296);
or U256 (N_256,In_383,N_125);
and U257 (N_257,N_193,In_164);
nor U258 (N_258,N_126,N_9);
and U259 (N_259,In_150,N_231);
and U260 (N_260,N_175,N_120);
and U261 (N_261,N_164,N_153);
nor U262 (N_262,N_85,In_365);
nor U263 (N_263,N_204,N_44);
and U264 (N_264,In_248,N_150);
nor U265 (N_265,In_402,In_434);
nor U266 (N_266,N_238,In_45);
or U267 (N_267,In_47,In_20);
or U268 (N_268,In_97,In_266);
or U269 (N_269,N_237,N_167);
nand U270 (N_270,N_207,N_196);
or U271 (N_271,N_213,N_210);
or U272 (N_272,In_316,N_13);
nor U273 (N_273,In_101,N_115);
nand U274 (N_274,In_456,N_14);
or U275 (N_275,In_340,N_156);
nor U276 (N_276,In_411,In_323);
nand U277 (N_277,In_330,N_173);
or U278 (N_278,N_118,In_349);
xor U279 (N_279,In_65,In_143);
nor U280 (N_280,N_195,In_216);
xor U281 (N_281,In_119,N_92);
and U282 (N_282,N_182,In_9);
or U283 (N_283,In_72,N_105);
or U284 (N_284,In_144,N_186);
and U285 (N_285,In_461,In_108);
nand U286 (N_286,N_8,N_219);
and U287 (N_287,In_188,N_163);
nor U288 (N_288,N_215,In_331);
nor U289 (N_289,In_395,In_446);
nand U290 (N_290,In_352,In_149);
and U291 (N_291,N_205,In_153);
nand U292 (N_292,In_436,In_281);
and U293 (N_293,N_72,N_235);
xnor U294 (N_294,N_15,In_347);
and U295 (N_295,N_108,N_216);
nor U296 (N_296,N_65,In_263);
nor U297 (N_297,N_211,N_249);
and U298 (N_298,N_229,N_234);
nor U299 (N_299,In_96,N_192);
or U300 (N_300,In_122,N_134);
and U301 (N_301,N_170,N_266);
and U302 (N_302,In_12,In_229);
nand U303 (N_303,N_260,N_256);
nand U304 (N_304,N_30,N_12);
or U305 (N_305,In_317,N_267);
xnor U306 (N_306,N_240,N_281);
or U307 (N_307,N_151,In_100);
nand U308 (N_308,In_303,N_244);
and U309 (N_309,N_241,N_282);
nand U310 (N_310,In_333,In_224);
and U311 (N_311,N_185,In_289);
nand U312 (N_312,N_178,In_443);
and U313 (N_313,In_145,N_103);
nand U314 (N_314,In_484,N_298);
nand U315 (N_315,N_130,N_190);
or U316 (N_316,In_327,N_291);
nor U317 (N_317,In_94,In_142);
and U318 (N_318,N_250,N_255);
xor U319 (N_319,N_245,In_398);
nand U320 (N_320,N_265,N_160);
nor U321 (N_321,N_236,In_475);
or U322 (N_322,N_168,N_101);
or U323 (N_323,N_189,N_208);
or U324 (N_324,N_127,N_194);
and U325 (N_325,N_242,N_286);
and U326 (N_326,In_307,N_200);
or U327 (N_327,In_358,N_252);
and U328 (N_328,N_289,N_293);
and U329 (N_329,In_41,N_50);
nor U330 (N_330,N_263,N_232);
and U331 (N_331,N_217,N_268);
nor U332 (N_332,N_259,In_190);
nand U333 (N_333,In_429,N_43);
or U334 (N_334,N_246,N_262);
xor U335 (N_335,N_148,N_272);
nand U336 (N_336,In_56,N_158);
or U337 (N_337,N_228,In_476);
nand U338 (N_338,N_225,N_273);
or U339 (N_339,N_145,N_62);
nand U340 (N_340,N_203,N_209);
nand U341 (N_341,N_261,In_305);
nor U342 (N_342,N_17,In_90);
nor U343 (N_343,N_110,N_23);
nor U344 (N_344,In_113,N_222);
nor U345 (N_345,N_79,N_223);
nor U346 (N_346,N_258,N_226);
nand U347 (N_347,N_218,N_82);
nand U348 (N_348,N_129,N_212);
and U349 (N_349,In_404,In_491);
xor U350 (N_350,N_333,N_201);
nand U351 (N_351,N_278,In_202);
or U352 (N_352,N_302,N_296);
nand U353 (N_353,N_279,N_290);
nor U354 (N_354,N_253,N_251);
nor U355 (N_355,In_346,N_331);
and U356 (N_356,N_319,In_275);
or U357 (N_357,In_17,In_442);
or U358 (N_358,N_254,N_338);
and U359 (N_359,N_335,N_330);
or U360 (N_360,N_197,N_304);
or U361 (N_361,N_224,N_317);
nor U362 (N_362,In_431,N_283);
nor U363 (N_363,N_349,N_306);
nor U364 (N_364,N_297,In_7);
and U365 (N_365,N_132,In_265);
or U366 (N_366,In_68,N_299);
nand U367 (N_367,In_494,N_311);
nor U368 (N_368,N_309,In_413);
nand U369 (N_369,N_276,N_301);
or U370 (N_370,In_37,N_314);
xor U371 (N_371,In_304,N_146);
and U372 (N_372,N_294,In_213);
nor U373 (N_373,N_123,N_275);
or U374 (N_374,N_308,N_280);
and U375 (N_375,N_176,N_315);
or U376 (N_376,In_38,In_230);
and U377 (N_377,N_345,N_221);
and U378 (N_378,In_81,N_93);
nor U379 (N_379,N_347,N_332);
or U380 (N_380,N_321,N_337);
nand U381 (N_381,N_22,N_277);
and U382 (N_382,In_22,In_91);
nor U383 (N_383,N_341,In_457);
nand U384 (N_384,N_16,N_324);
and U385 (N_385,N_152,N_172);
and U386 (N_386,N_318,N_305);
or U387 (N_387,N_292,N_227);
nand U388 (N_388,N_342,N_323);
and U389 (N_389,N_214,In_348);
or U390 (N_390,N_340,N_326);
nand U391 (N_391,N_274,N_329);
and U392 (N_392,N_346,N_284);
nor U393 (N_393,N_310,N_334);
nand U394 (N_394,N_327,N_61);
and U395 (N_395,In_71,N_77);
nand U396 (N_396,N_307,N_287);
and U397 (N_397,In_458,In_18);
nand U398 (N_398,N_248,N_285);
nor U399 (N_399,N_344,N_106);
nand U400 (N_400,N_336,N_394);
nand U401 (N_401,N_359,In_483);
nor U402 (N_402,N_316,N_198);
or U403 (N_403,N_398,N_300);
nor U404 (N_404,N_270,N_373);
nor U405 (N_405,N_384,N_202);
or U406 (N_406,N_370,N_395);
nand U407 (N_407,N_365,N_387);
and U408 (N_408,N_375,In_468);
and U409 (N_409,N_378,N_269);
and U410 (N_410,N_136,N_379);
and U411 (N_411,N_5,N_179);
or U412 (N_412,N_369,N_382);
and U413 (N_413,N_320,In_421);
or U414 (N_414,N_264,In_360);
nor U415 (N_415,N_390,N_230);
or U416 (N_416,N_396,In_79);
nor U417 (N_417,N_377,N_386);
and U418 (N_418,N_361,N_339);
nand U419 (N_419,N_368,N_391);
xnor U420 (N_420,N_364,N_354);
nor U421 (N_421,In_315,In_415);
nor U422 (N_422,N_191,In_5);
xnor U423 (N_423,N_322,N_353);
nand U424 (N_424,N_350,N_371);
and U425 (N_425,N_313,N_66);
nand U426 (N_426,N_399,N_352);
nor U427 (N_427,N_392,N_366);
nor U428 (N_428,In_322,N_183);
nor U429 (N_429,In_74,N_247);
nor U430 (N_430,N_288,N_343);
nand U431 (N_431,N_356,N_355);
nand U432 (N_432,In_221,N_380);
nand U433 (N_433,N_389,In_256);
or U434 (N_434,In_55,N_348);
nand U435 (N_435,N_174,N_159);
nand U436 (N_436,N_312,N_325);
or U437 (N_437,N_233,N_393);
or U438 (N_438,N_358,N_295);
nor U439 (N_439,N_383,N_363);
nand U440 (N_440,N_367,N_376);
and U441 (N_441,N_257,N_385);
and U442 (N_442,N_381,N_351);
nor U443 (N_443,N_169,N_303);
or U444 (N_444,N_372,N_239);
and U445 (N_445,N_360,N_328);
or U446 (N_446,N_397,In_154);
nand U447 (N_447,N_271,N_357);
nor U448 (N_448,N_362,N_388);
nand U449 (N_449,N_206,N_374);
or U450 (N_450,N_419,N_445);
nand U451 (N_451,N_443,N_415);
nand U452 (N_452,N_441,N_444);
and U453 (N_453,N_430,N_448);
nor U454 (N_454,N_418,N_423);
or U455 (N_455,N_429,N_400);
and U456 (N_456,N_413,N_440);
or U457 (N_457,N_407,N_426);
or U458 (N_458,N_446,N_412);
nor U459 (N_459,N_447,N_449);
xor U460 (N_460,N_421,N_439);
or U461 (N_461,N_431,N_410);
and U462 (N_462,N_402,N_409);
xnor U463 (N_463,N_405,N_416);
nor U464 (N_464,N_408,N_411);
nor U465 (N_465,N_424,N_403);
nor U466 (N_466,N_401,N_434);
and U467 (N_467,N_427,N_414);
and U468 (N_468,N_436,N_422);
and U469 (N_469,N_433,N_425);
and U470 (N_470,N_432,N_420);
and U471 (N_471,N_404,N_406);
nor U472 (N_472,N_428,N_442);
and U473 (N_473,N_438,N_417);
and U474 (N_474,N_437,N_435);
or U475 (N_475,N_425,N_400);
nand U476 (N_476,N_417,N_415);
and U477 (N_477,N_429,N_428);
xnor U478 (N_478,N_419,N_400);
nor U479 (N_479,N_426,N_449);
and U480 (N_480,N_441,N_410);
nand U481 (N_481,N_431,N_429);
nand U482 (N_482,N_422,N_400);
nand U483 (N_483,N_448,N_410);
nor U484 (N_484,N_419,N_405);
or U485 (N_485,N_424,N_431);
or U486 (N_486,N_414,N_445);
nand U487 (N_487,N_429,N_441);
nor U488 (N_488,N_404,N_434);
nor U489 (N_489,N_430,N_432);
nor U490 (N_490,N_414,N_441);
nor U491 (N_491,N_413,N_443);
nor U492 (N_492,N_420,N_415);
nor U493 (N_493,N_427,N_421);
and U494 (N_494,N_422,N_409);
or U495 (N_495,N_428,N_447);
nand U496 (N_496,N_432,N_439);
and U497 (N_497,N_430,N_428);
or U498 (N_498,N_423,N_436);
nand U499 (N_499,N_417,N_416);
xnor U500 (N_500,N_486,N_499);
nand U501 (N_501,N_498,N_491);
or U502 (N_502,N_463,N_466);
nand U503 (N_503,N_469,N_489);
or U504 (N_504,N_470,N_485);
or U505 (N_505,N_496,N_484);
and U506 (N_506,N_471,N_464);
and U507 (N_507,N_492,N_477);
nand U508 (N_508,N_451,N_452);
or U509 (N_509,N_460,N_495);
nor U510 (N_510,N_493,N_488);
nand U511 (N_511,N_459,N_468);
nand U512 (N_512,N_465,N_473);
and U513 (N_513,N_453,N_462);
or U514 (N_514,N_478,N_483);
nor U515 (N_515,N_490,N_454);
or U516 (N_516,N_457,N_482);
nand U517 (N_517,N_455,N_479);
or U518 (N_518,N_476,N_467);
xor U519 (N_519,N_475,N_480);
or U520 (N_520,N_458,N_497);
or U521 (N_521,N_472,N_456);
nand U522 (N_522,N_450,N_461);
nand U523 (N_523,N_494,N_474);
nand U524 (N_524,N_487,N_481);
and U525 (N_525,N_481,N_470);
xnor U526 (N_526,N_499,N_476);
nand U527 (N_527,N_493,N_483);
and U528 (N_528,N_453,N_479);
nand U529 (N_529,N_477,N_468);
nand U530 (N_530,N_466,N_472);
nor U531 (N_531,N_459,N_498);
or U532 (N_532,N_462,N_478);
or U533 (N_533,N_471,N_487);
and U534 (N_534,N_471,N_457);
and U535 (N_535,N_493,N_497);
and U536 (N_536,N_486,N_457);
nor U537 (N_537,N_469,N_452);
nand U538 (N_538,N_466,N_483);
and U539 (N_539,N_453,N_461);
and U540 (N_540,N_461,N_475);
and U541 (N_541,N_479,N_489);
nor U542 (N_542,N_465,N_454);
nand U543 (N_543,N_465,N_464);
nor U544 (N_544,N_475,N_479);
or U545 (N_545,N_497,N_495);
nor U546 (N_546,N_457,N_476);
nor U547 (N_547,N_452,N_458);
nand U548 (N_548,N_490,N_478);
nor U549 (N_549,N_461,N_494);
and U550 (N_550,N_511,N_549);
and U551 (N_551,N_515,N_527);
nor U552 (N_552,N_513,N_537);
nor U553 (N_553,N_503,N_533);
nor U554 (N_554,N_542,N_506);
or U555 (N_555,N_508,N_524);
nand U556 (N_556,N_514,N_532);
or U557 (N_557,N_539,N_520);
or U558 (N_558,N_546,N_517);
nand U559 (N_559,N_504,N_518);
nor U560 (N_560,N_522,N_509);
and U561 (N_561,N_530,N_536);
nor U562 (N_562,N_545,N_541);
nor U563 (N_563,N_523,N_505);
nor U564 (N_564,N_519,N_512);
nor U565 (N_565,N_507,N_534);
and U566 (N_566,N_501,N_528);
nor U567 (N_567,N_526,N_529);
nor U568 (N_568,N_516,N_543);
nor U569 (N_569,N_548,N_538);
or U570 (N_570,N_547,N_521);
xor U571 (N_571,N_531,N_525);
and U572 (N_572,N_500,N_544);
nand U573 (N_573,N_510,N_535);
nand U574 (N_574,N_540,N_502);
or U575 (N_575,N_548,N_537);
or U576 (N_576,N_517,N_519);
nor U577 (N_577,N_513,N_516);
or U578 (N_578,N_518,N_502);
nor U579 (N_579,N_534,N_506);
and U580 (N_580,N_543,N_513);
nor U581 (N_581,N_524,N_504);
nand U582 (N_582,N_500,N_537);
or U583 (N_583,N_521,N_544);
or U584 (N_584,N_504,N_509);
nor U585 (N_585,N_532,N_518);
nand U586 (N_586,N_509,N_501);
nand U587 (N_587,N_548,N_530);
or U588 (N_588,N_534,N_513);
and U589 (N_589,N_509,N_546);
and U590 (N_590,N_500,N_532);
or U591 (N_591,N_536,N_549);
nand U592 (N_592,N_526,N_536);
and U593 (N_593,N_539,N_549);
and U594 (N_594,N_522,N_528);
nor U595 (N_595,N_529,N_530);
nor U596 (N_596,N_542,N_539);
and U597 (N_597,N_504,N_533);
nand U598 (N_598,N_517,N_540);
nor U599 (N_599,N_525,N_517);
and U600 (N_600,N_580,N_572);
nor U601 (N_601,N_555,N_554);
or U602 (N_602,N_553,N_590);
and U603 (N_603,N_563,N_565);
nor U604 (N_604,N_557,N_561);
nand U605 (N_605,N_564,N_597);
nand U606 (N_606,N_551,N_592);
or U607 (N_607,N_591,N_550);
nor U608 (N_608,N_584,N_552);
nand U609 (N_609,N_569,N_560);
nand U610 (N_610,N_596,N_575);
nand U611 (N_611,N_574,N_587);
or U612 (N_612,N_581,N_578);
and U613 (N_613,N_582,N_599);
nor U614 (N_614,N_577,N_567);
or U615 (N_615,N_586,N_576);
nand U616 (N_616,N_589,N_568);
and U617 (N_617,N_556,N_585);
and U618 (N_618,N_558,N_559);
and U619 (N_619,N_579,N_583);
and U620 (N_620,N_594,N_588);
nand U621 (N_621,N_593,N_595);
nand U622 (N_622,N_598,N_570);
xnor U623 (N_623,N_566,N_571);
nor U624 (N_624,N_562,N_573);
xor U625 (N_625,N_553,N_593);
nand U626 (N_626,N_583,N_556);
and U627 (N_627,N_564,N_562);
nor U628 (N_628,N_557,N_574);
nor U629 (N_629,N_584,N_583);
nand U630 (N_630,N_566,N_579);
nand U631 (N_631,N_556,N_596);
or U632 (N_632,N_594,N_574);
xor U633 (N_633,N_595,N_587);
nor U634 (N_634,N_557,N_598);
nor U635 (N_635,N_571,N_558);
nand U636 (N_636,N_572,N_591);
or U637 (N_637,N_566,N_591);
or U638 (N_638,N_584,N_567);
nor U639 (N_639,N_565,N_557);
or U640 (N_640,N_569,N_584);
or U641 (N_641,N_559,N_557);
or U642 (N_642,N_567,N_592);
nor U643 (N_643,N_570,N_581);
or U644 (N_644,N_594,N_557);
nand U645 (N_645,N_586,N_593);
nor U646 (N_646,N_571,N_555);
or U647 (N_647,N_581,N_552);
or U648 (N_648,N_599,N_550);
and U649 (N_649,N_581,N_569);
nor U650 (N_650,N_648,N_633);
nand U651 (N_651,N_632,N_604);
or U652 (N_652,N_629,N_625);
nand U653 (N_653,N_605,N_620);
nand U654 (N_654,N_614,N_638);
nor U655 (N_655,N_631,N_626);
or U656 (N_656,N_621,N_617);
and U657 (N_657,N_635,N_619);
or U658 (N_658,N_644,N_630);
xnor U659 (N_659,N_606,N_642);
nor U660 (N_660,N_622,N_634);
nor U661 (N_661,N_647,N_645);
nand U662 (N_662,N_616,N_603);
xnor U663 (N_663,N_615,N_612);
nand U664 (N_664,N_649,N_611);
nand U665 (N_665,N_636,N_613);
nor U666 (N_666,N_600,N_618);
nand U667 (N_667,N_607,N_627);
or U668 (N_668,N_624,N_601);
nor U669 (N_669,N_609,N_623);
nand U670 (N_670,N_637,N_643);
nand U671 (N_671,N_602,N_641);
nor U672 (N_672,N_608,N_639);
or U673 (N_673,N_646,N_628);
xnor U674 (N_674,N_640,N_610);
and U675 (N_675,N_646,N_618);
nor U676 (N_676,N_631,N_646);
nand U677 (N_677,N_629,N_622);
nor U678 (N_678,N_642,N_643);
and U679 (N_679,N_641,N_611);
or U680 (N_680,N_647,N_627);
nand U681 (N_681,N_624,N_613);
nand U682 (N_682,N_641,N_628);
or U683 (N_683,N_639,N_634);
nor U684 (N_684,N_620,N_644);
or U685 (N_685,N_621,N_640);
or U686 (N_686,N_602,N_631);
and U687 (N_687,N_623,N_646);
nor U688 (N_688,N_610,N_606);
and U689 (N_689,N_632,N_645);
or U690 (N_690,N_612,N_604);
nand U691 (N_691,N_610,N_644);
and U692 (N_692,N_610,N_628);
nor U693 (N_693,N_606,N_612);
and U694 (N_694,N_615,N_639);
nor U695 (N_695,N_633,N_630);
or U696 (N_696,N_623,N_645);
or U697 (N_697,N_621,N_626);
nor U698 (N_698,N_601,N_621);
and U699 (N_699,N_639,N_618);
and U700 (N_700,N_661,N_651);
or U701 (N_701,N_698,N_669);
nand U702 (N_702,N_695,N_692);
or U703 (N_703,N_650,N_683);
nor U704 (N_704,N_665,N_671);
or U705 (N_705,N_660,N_693);
nor U706 (N_706,N_680,N_663);
and U707 (N_707,N_689,N_686);
nor U708 (N_708,N_687,N_675);
and U709 (N_709,N_668,N_699);
nand U710 (N_710,N_656,N_690);
nand U711 (N_711,N_666,N_691);
and U712 (N_712,N_684,N_670);
nand U713 (N_713,N_658,N_694);
nor U714 (N_714,N_678,N_664);
and U715 (N_715,N_652,N_654);
nor U716 (N_716,N_676,N_662);
or U717 (N_717,N_688,N_682);
nand U718 (N_718,N_657,N_681);
or U719 (N_719,N_659,N_667);
nand U720 (N_720,N_685,N_696);
and U721 (N_721,N_672,N_677);
and U722 (N_722,N_673,N_697);
nand U723 (N_723,N_679,N_655);
and U724 (N_724,N_674,N_653);
nand U725 (N_725,N_683,N_655);
and U726 (N_726,N_667,N_686);
and U727 (N_727,N_683,N_684);
or U728 (N_728,N_679,N_674);
and U729 (N_729,N_681,N_678);
or U730 (N_730,N_677,N_682);
and U731 (N_731,N_675,N_699);
nor U732 (N_732,N_651,N_669);
nand U733 (N_733,N_694,N_696);
and U734 (N_734,N_668,N_655);
xnor U735 (N_735,N_667,N_682);
nand U736 (N_736,N_652,N_698);
nand U737 (N_737,N_688,N_674);
or U738 (N_738,N_675,N_671);
or U739 (N_739,N_699,N_690);
nand U740 (N_740,N_651,N_677);
and U741 (N_741,N_662,N_670);
and U742 (N_742,N_659,N_656);
nor U743 (N_743,N_664,N_685);
or U744 (N_744,N_692,N_660);
or U745 (N_745,N_656,N_686);
and U746 (N_746,N_697,N_668);
or U747 (N_747,N_682,N_684);
nor U748 (N_748,N_663,N_686);
or U749 (N_749,N_678,N_672);
and U750 (N_750,N_727,N_718);
or U751 (N_751,N_744,N_707);
or U752 (N_752,N_711,N_733);
xnor U753 (N_753,N_701,N_748);
and U754 (N_754,N_724,N_725);
or U755 (N_755,N_742,N_743);
nor U756 (N_756,N_708,N_746);
nor U757 (N_757,N_716,N_709);
nand U758 (N_758,N_706,N_719);
nand U759 (N_759,N_738,N_732);
nor U760 (N_760,N_741,N_729);
nor U761 (N_761,N_717,N_704);
and U762 (N_762,N_713,N_710);
or U763 (N_763,N_739,N_740);
nand U764 (N_764,N_730,N_714);
and U765 (N_765,N_749,N_721);
nor U766 (N_766,N_726,N_734);
nor U767 (N_767,N_702,N_703);
and U768 (N_768,N_712,N_736);
and U769 (N_769,N_705,N_735);
and U770 (N_770,N_720,N_731);
nand U771 (N_771,N_737,N_747);
and U772 (N_772,N_728,N_700);
nand U773 (N_773,N_722,N_715);
or U774 (N_774,N_745,N_723);
xnor U775 (N_775,N_745,N_701);
and U776 (N_776,N_709,N_722);
nor U777 (N_777,N_727,N_733);
or U778 (N_778,N_715,N_717);
xor U779 (N_779,N_727,N_704);
nor U780 (N_780,N_711,N_720);
nor U781 (N_781,N_704,N_733);
nor U782 (N_782,N_728,N_749);
nand U783 (N_783,N_735,N_725);
nand U784 (N_784,N_722,N_703);
nand U785 (N_785,N_736,N_721);
nor U786 (N_786,N_721,N_747);
nand U787 (N_787,N_706,N_714);
or U788 (N_788,N_719,N_741);
or U789 (N_789,N_703,N_747);
or U790 (N_790,N_728,N_709);
nand U791 (N_791,N_721,N_718);
nor U792 (N_792,N_717,N_731);
or U793 (N_793,N_719,N_728);
and U794 (N_794,N_725,N_700);
and U795 (N_795,N_744,N_703);
or U796 (N_796,N_739,N_731);
nor U797 (N_797,N_734,N_719);
nor U798 (N_798,N_717,N_708);
nor U799 (N_799,N_725,N_737);
or U800 (N_800,N_790,N_753);
and U801 (N_801,N_797,N_765);
nand U802 (N_802,N_768,N_792);
and U803 (N_803,N_750,N_757);
xor U804 (N_804,N_760,N_794);
or U805 (N_805,N_762,N_755);
nor U806 (N_806,N_759,N_776);
and U807 (N_807,N_784,N_798);
nand U808 (N_808,N_781,N_773);
nor U809 (N_809,N_779,N_769);
nor U810 (N_810,N_752,N_763);
nor U811 (N_811,N_775,N_756);
and U812 (N_812,N_782,N_771);
or U813 (N_813,N_786,N_761);
and U814 (N_814,N_793,N_789);
nand U815 (N_815,N_772,N_795);
and U816 (N_816,N_770,N_799);
or U817 (N_817,N_796,N_764);
or U818 (N_818,N_780,N_767);
and U819 (N_819,N_787,N_758);
nand U820 (N_820,N_777,N_774);
or U821 (N_821,N_751,N_783);
nor U822 (N_822,N_766,N_785);
nor U823 (N_823,N_778,N_791);
nor U824 (N_824,N_754,N_788);
or U825 (N_825,N_775,N_751);
nor U826 (N_826,N_796,N_775);
nor U827 (N_827,N_789,N_775);
and U828 (N_828,N_763,N_782);
nand U829 (N_829,N_771,N_788);
or U830 (N_830,N_756,N_798);
or U831 (N_831,N_790,N_782);
nand U832 (N_832,N_768,N_795);
nor U833 (N_833,N_774,N_752);
and U834 (N_834,N_751,N_752);
xor U835 (N_835,N_778,N_752);
and U836 (N_836,N_773,N_782);
and U837 (N_837,N_761,N_755);
nand U838 (N_838,N_793,N_788);
and U839 (N_839,N_797,N_781);
or U840 (N_840,N_771,N_779);
and U841 (N_841,N_789,N_792);
or U842 (N_842,N_793,N_797);
and U843 (N_843,N_772,N_750);
nor U844 (N_844,N_785,N_756);
and U845 (N_845,N_769,N_785);
or U846 (N_846,N_779,N_786);
nor U847 (N_847,N_765,N_767);
and U848 (N_848,N_760,N_764);
nand U849 (N_849,N_768,N_770);
or U850 (N_850,N_819,N_827);
nor U851 (N_851,N_843,N_803);
or U852 (N_852,N_815,N_834);
or U853 (N_853,N_811,N_830);
nor U854 (N_854,N_802,N_809);
and U855 (N_855,N_822,N_845);
nor U856 (N_856,N_812,N_841);
nor U857 (N_857,N_806,N_835);
and U858 (N_858,N_821,N_824);
nand U859 (N_859,N_829,N_810);
nor U860 (N_860,N_828,N_818);
or U861 (N_861,N_816,N_833);
or U862 (N_862,N_813,N_826);
nand U863 (N_863,N_848,N_849);
or U864 (N_864,N_831,N_800);
nor U865 (N_865,N_814,N_823);
or U866 (N_866,N_801,N_820);
and U867 (N_867,N_825,N_805);
nor U868 (N_868,N_832,N_837);
and U869 (N_869,N_844,N_808);
or U870 (N_870,N_839,N_807);
or U871 (N_871,N_817,N_842);
and U872 (N_872,N_804,N_838);
nor U873 (N_873,N_840,N_846);
or U874 (N_874,N_847,N_836);
xnor U875 (N_875,N_807,N_801);
nand U876 (N_876,N_809,N_833);
nand U877 (N_877,N_817,N_821);
and U878 (N_878,N_844,N_833);
nor U879 (N_879,N_841,N_808);
nor U880 (N_880,N_826,N_830);
and U881 (N_881,N_837,N_838);
and U882 (N_882,N_802,N_808);
nor U883 (N_883,N_825,N_810);
nor U884 (N_884,N_807,N_820);
nand U885 (N_885,N_820,N_816);
xnor U886 (N_886,N_801,N_804);
and U887 (N_887,N_835,N_818);
or U888 (N_888,N_839,N_840);
and U889 (N_889,N_819,N_837);
or U890 (N_890,N_848,N_823);
or U891 (N_891,N_841,N_846);
or U892 (N_892,N_846,N_842);
and U893 (N_893,N_807,N_815);
nand U894 (N_894,N_805,N_818);
and U895 (N_895,N_828,N_849);
and U896 (N_896,N_802,N_845);
and U897 (N_897,N_813,N_810);
xnor U898 (N_898,N_808,N_830);
nand U899 (N_899,N_821,N_808);
and U900 (N_900,N_868,N_887);
and U901 (N_901,N_864,N_854);
nand U902 (N_902,N_889,N_856);
and U903 (N_903,N_851,N_872);
and U904 (N_904,N_893,N_878);
or U905 (N_905,N_884,N_885);
nor U906 (N_906,N_880,N_871);
xor U907 (N_907,N_898,N_857);
or U908 (N_908,N_891,N_860);
and U909 (N_909,N_866,N_874);
nand U910 (N_910,N_892,N_855);
nand U911 (N_911,N_859,N_877);
nand U912 (N_912,N_890,N_879);
and U913 (N_913,N_895,N_882);
nand U914 (N_914,N_896,N_850);
and U915 (N_915,N_894,N_858);
nor U916 (N_916,N_862,N_873);
xor U917 (N_917,N_876,N_853);
nand U918 (N_918,N_875,N_883);
and U919 (N_919,N_899,N_881);
nand U920 (N_920,N_869,N_870);
and U921 (N_921,N_863,N_867);
nand U922 (N_922,N_888,N_861);
or U923 (N_923,N_897,N_852);
xor U924 (N_924,N_886,N_865);
and U925 (N_925,N_872,N_866);
or U926 (N_926,N_893,N_867);
nand U927 (N_927,N_882,N_896);
nand U928 (N_928,N_887,N_893);
and U929 (N_929,N_865,N_878);
and U930 (N_930,N_881,N_873);
nand U931 (N_931,N_857,N_879);
nand U932 (N_932,N_896,N_862);
nand U933 (N_933,N_880,N_867);
nand U934 (N_934,N_891,N_868);
or U935 (N_935,N_854,N_897);
and U936 (N_936,N_856,N_875);
nand U937 (N_937,N_861,N_894);
nor U938 (N_938,N_887,N_874);
or U939 (N_939,N_869,N_887);
and U940 (N_940,N_863,N_858);
nor U941 (N_941,N_865,N_864);
or U942 (N_942,N_887,N_882);
nand U943 (N_943,N_860,N_875);
nand U944 (N_944,N_898,N_886);
or U945 (N_945,N_874,N_871);
or U946 (N_946,N_859,N_899);
nor U947 (N_947,N_854,N_878);
or U948 (N_948,N_896,N_866);
nand U949 (N_949,N_866,N_868);
and U950 (N_950,N_931,N_912);
nand U951 (N_951,N_929,N_900);
or U952 (N_952,N_908,N_947);
nor U953 (N_953,N_918,N_927);
nand U954 (N_954,N_941,N_921);
nor U955 (N_955,N_903,N_924);
nand U956 (N_956,N_930,N_944);
nand U957 (N_957,N_932,N_934);
and U958 (N_958,N_919,N_902);
nand U959 (N_959,N_938,N_905);
nand U960 (N_960,N_901,N_928);
or U961 (N_961,N_916,N_933);
nand U962 (N_962,N_911,N_906);
and U963 (N_963,N_907,N_945);
or U964 (N_964,N_936,N_926);
and U965 (N_965,N_935,N_943);
nor U966 (N_966,N_937,N_920);
nand U967 (N_967,N_922,N_946);
or U968 (N_968,N_909,N_913);
and U969 (N_969,N_904,N_939);
or U970 (N_970,N_915,N_917);
or U971 (N_971,N_949,N_923);
nor U972 (N_972,N_942,N_940);
nand U973 (N_973,N_925,N_910);
and U974 (N_974,N_948,N_914);
nand U975 (N_975,N_924,N_912);
nor U976 (N_976,N_928,N_909);
nand U977 (N_977,N_949,N_945);
nor U978 (N_978,N_902,N_905);
nand U979 (N_979,N_920,N_927);
nand U980 (N_980,N_923,N_911);
nand U981 (N_981,N_913,N_912);
or U982 (N_982,N_928,N_910);
and U983 (N_983,N_916,N_912);
nor U984 (N_984,N_949,N_939);
or U985 (N_985,N_904,N_929);
and U986 (N_986,N_942,N_944);
or U987 (N_987,N_943,N_945);
and U988 (N_988,N_943,N_928);
or U989 (N_989,N_908,N_946);
nor U990 (N_990,N_928,N_941);
nor U991 (N_991,N_929,N_942);
and U992 (N_992,N_920,N_946);
and U993 (N_993,N_906,N_912);
nand U994 (N_994,N_940,N_918);
and U995 (N_995,N_921,N_933);
nand U996 (N_996,N_943,N_948);
and U997 (N_997,N_915,N_923);
nand U998 (N_998,N_912,N_933);
and U999 (N_999,N_947,N_923);
or U1000 (N_1000,N_998,N_980);
nor U1001 (N_1001,N_959,N_978);
xnor U1002 (N_1002,N_974,N_962);
or U1003 (N_1003,N_975,N_990);
nor U1004 (N_1004,N_951,N_986);
or U1005 (N_1005,N_972,N_961);
and U1006 (N_1006,N_967,N_993);
nor U1007 (N_1007,N_991,N_982);
nand U1008 (N_1008,N_968,N_979);
or U1009 (N_1009,N_994,N_999);
and U1010 (N_1010,N_977,N_969);
nor U1011 (N_1011,N_989,N_988);
and U1012 (N_1012,N_964,N_983);
xnor U1013 (N_1013,N_971,N_956);
or U1014 (N_1014,N_996,N_966);
and U1015 (N_1015,N_963,N_960);
nor U1016 (N_1016,N_954,N_955);
and U1017 (N_1017,N_950,N_952);
and U1018 (N_1018,N_984,N_992);
or U1019 (N_1019,N_976,N_958);
or U1020 (N_1020,N_970,N_981);
or U1021 (N_1021,N_985,N_953);
nand U1022 (N_1022,N_987,N_997);
or U1023 (N_1023,N_957,N_973);
or U1024 (N_1024,N_965,N_995);
nor U1025 (N_1025,N_986,N_950);
nor U1026 (N_1026,N_960,N_995);
and U1027 (N_1027,N_952,N_980);
nor U1028 (N_1028,N_985,N_950);
or U1029 (N_1029,N_970,N_985);
and U1030 (N_1030,N_952,N_985);
nand U1031 (N_1031,N_964,N_974);
nor U1032 (N_1032,N_977,N_967);
and U1033 (N_1033,N_952,N_961);
nor U1034 (N_1034,N_961,N_957);
nor U1035 (N_1035,N_958,N_950);
nor U1036 (N_1036,N_991,N_970);
or U1037 (N_1037,N_988,N_984);
nand U1038 (N_1038,N_966,N_955);
nand U1039 (N_1039,N_957,N_974);
nor U1040 (N_1040,N_988,N_990);
or U1041 (N_1041,N_967,N_958);
and U1042 (N_1042,N_966,N_980);
nor U1043 (N_1043,N_988,N_972);
nand U1044 (N_1044,N_997,N_953);
and U1045 (N_1045,N_953,N_958);
nor U1046 (N_1046,N_974,N_955);
nor U1047 (N_1047,N_988,N_971);
nor U1048 (N_1048,N_975,N_974);
nand U1049 (N_1049,N_972,N_950);
or U1050 (N_1050,N_1000,N_1027);
nor U1051 (N_1051,N_1033,N_1019);
and U1052 (N_1052,N_1013,N_1010);
nor U1053 (N_1053,N_1009,N_1040);
nand U1054 (N_1054,N_1020,N_1048);
nor U1055 (N_1055,N_1042,N_1049);
nand U1056 (N_1056,N_1028,N_1018);
and U1057 (N_1057,N_1001,N_1006);
and U1058 (N_1058,N_1002,N_1011);
nand U1059 (N_1059,N_1030,N_1017);
and U1060 (N_1060,N_1034,N_1047);
or U1061 (N_1061,N_1035,N_1044);
and U1062 (N_1062,N_1039,N_1037);
or U1063 (N_1063,N_1021,N_1007);
nor U1064 (N_1064,N_1031,N_1041);
nor U1065 (N_1065,N_1038,N_1022);
nand U1066 (N_1066,N_1023,N_1015);
or U1067 (N_1067,N_1014,N_1016);
nand U1068 (N_1068,N_1036,N_1003);
nand U1069 (N_1069,N_1005,N_1004);
nor U1070 (N_1070,N_1032,N_1012);
nor U1071 (N_1071,N_1008,N_1024);
nor U1072 (N_1072,N_1025,N_1045);
nand U1073 (N_1073,N_1029,N_1026);
and U1074 (N_1074,N_1043,N_1046);
nand U1075 (N_1075,N_1023,N_1024);
nand U1076 (N_1076,N_1000,N_1026);
or U1077 (N_1077,N_1000,N_1039);
or U1078 (N_1078,N_1016,N_1026);
nand U1079 (N_1079,N_1001,N_1029);
nor U1080 (N_1080,N_1035,N_1004);
or U1081 (N_1081,N_1007,N_1033);
nor U1082 (N_1082,N_1047,N_1023);
nand U1083 (N_1083,N_1028,N_1043);
nor U1084 (N_1084,N_1010,N_1004);
and U1085 (N_1085,N_1002,N_1013);
and U1086 (N_1086,N_1004,N_1025);
nor U1087 (N_1087,N_1015,N_1032);
nand U1088 (N_1088,N_1024,N_1013);
nor U1089 (N_1089,N_1038,N_1017);
nand U1090 (N_1090,N_1045,N_1006);
or U1091 (N_1091,N_1007,N_1011);
or U1092 (N_1092,N_1042,N_1036);
nor U1093 (N_1093,N_1044,N_1011);
and U1094 (N_1094,N_1029,N_1002);
nand U1095 (N_1095,N_1000,N_1012);
and U1096 (N_1096,N_1038,N_1047);
and U1097 (N_1097,N_1009,N_1048);
and U1098 (N_1098,N_1015,N_1039);
nand U1099 (N_1099,N_1022,N_1028);
and U1100 (N_1100,N_1050,N_1099);
or U1101 (N_1101,N_1081,N_1078);
and U1102 (N_1102,N_1090,N_1059);
nor U1103 (N_1103,N_1052,N_1051);
nand U1104 (N_1104,N_1086,N_1080);
or U1105 (N_1105,N_1069,N_1060);
nor U1106 (N_1106,N_1071,N_1085);
or U1107 (N_1107,N_1087,N_1074);
nor U1108 (N_1108,N_1066,N_1063);
xnor U1109 (N_1109,N_1094,N_1088);
and U1110 (N_1110,N_1083,N_1076);
and U1111 (N_1111,N_1075,N_1053);
or U1112 (N_1112,N_1098,N_1064);
nor U1113 (N_1113,N_1062,N_1057);
nor U1114 (N_1114,N_1092,N_1073);
xnor U1115 (N_1115,N_1065,N_1096);
or U1116 (N_1116,N_1070,N_1072);
and U1117 (N_1117,N_1077,N_1056);
or U1118 (N_1118,N_1082,N_1068);
or U1119 (N_1119,N_1089,N_1054);
nor U1120 (N_1120,N_1079,N_1055);
and U1121 (N_1121,N_1061,N_1091);
xor U1122 (N_1122,N_1058,N_1097);
nor U1123 (N_1123,N_1093,N_1067);
and U1124 (N_1124,N_1084,N_1095);
or U1125 (N_1125,N_1055,N_1088);
and U1126 (N_1126,N_1051,N_1088);
nand U1127 (N_1127,N_1088,N_1072);
nor U1128 (N_1128,N_1066,N_1087);
nor U1129 (N_1129,N_1085,N_1055);
and U1130 (N_1130,N_1068,N_1084);
nor U1131 (N_1131,N_1063,N_1055);
or U1132 (N_1132,N_1094,N_1086);
and U1133 (N_1133,N_1069,N_1096);
nor U1134 (N_1134,N_1092,N_1070);
nand U1135 (N_1135,N_1081,N_1061);
nand U1136 (N_1136,N_1060,N_1057);
nand U1137 (N_1137,N_1083,N_1069);
nand U1138 (N_1138,N_1073,N_1077);
or U1139 (N_1139,N_1051,N_1068);
or U1140 (N_1140,N_1092,N_1088);
nor U1141 (N_1141,N_1054,N_1059);
and U1142 (N_1142,N_1054,N_1079);
or U1143 (N_1143,N_1095,N_1056);
nand U1144 (N_1144,N_1099,N_1056);
nor U1145 (N_1145,N_1097,N_1084);
nand U1146 (N_1146,N_1055,N_1054);
or U1147 (N_1147,N_1064,N_1078);
or U1148 (N_1148,N_1085,N_1099);
nor U1149 (N_1149,N_1052,N_1072);
nand U1150 (N_1150,N_1110,N_1147);
nor U1151 (N_1151,N_1114,N_1116);
nand U1152 (N_1152,N_1118,N_1149);
and U1153 (N_1153,N_1108,N_1129);
or U1154 (N_1154,N_1106,N_1135);
or U1155 (N_1155,N_1102,N_1137);
or U1156 (N_1156,N_1134,N_1117);
nor U1157 (N_1157,N_1131,N_1119);
nand U1158 (N_1158,N_1123,N_1140);
nand U1159 (N_1159,N_1144,N_1124);
nor U1160 (N_1160,N_1139,N_1132);
or U1161 (N_1161,N_1136,N_1145);
nand U1162 (N_1162,N_1112,N_1104);
nand U1163 (N_1163,N_1143,N_1111);
nor U1164 (N_1164,N_1113,N_1105);
nand U1165 (N_1165,N_1101,N_1103);
nand U1166 (N_1166,N_1141,N_1107);
nor U1167 (N_1167,N_1121,N_1120);
nand U1168 (N_1168,N_1130,N_1128);
nor U1169 (N_1169,N_1115,N_1127);
or U1170 (N_1170,N_1142,N_1109);
or U1171 (N_1171,N_1100,N_1146);
nand U1172 (N_1172,N_1148,N_1122);
and U1173 (N_1173,N_1126,N_1133);
nand U1174 (N_1174,N_1125,N_1138);
and U1175 (N_1175,N_1105,N_1117);
or U1176 (N_1176,N_1133,N_1124);
and U1177 (N_1177,N_1145,N_1108);
and U1178 (N_1178,N_1138,N_1122);
nand U1179 (N_1179,N_1109,N_1133);
nor U1180 (N_1180,N_1111,N_1146);
and U1181 (N_1181,N_1137,N_1139);
nand U1182 (N_1182,N_1117,N_1139);
nand U1183 (N_1183,N_1131,N_1107);
or U1184 (N_1184,N_1144,N_1135);
and U1185 (N_1185,N_1125,N_1117);
and U1186 (N_1186,N_1122,N_1139);
or U1187 (N_1187,N_1109,N_1111);
nand U1188 (N_1188,N_1118,N_1111);
and U1189 (N_1189,N_1142,N_1133);
nor U1190 (N_1190,N_1101,N_1144);
nand U1191 (N_1191,N_1134,N_1124);
nand U1192 (N_1192,N_1120,N_1138);
nand U1193 (N_1193,N_1118,N_1100);
and U1194 (N_1194,N_1142,N_1128);
nor U1195 (N_1195,N_1146,N_1107);
or U1196 (N_1196,N_1117,N_1102);
nor U1197 (N_1197,N_1107,N_1142);
nor U1198 (N_1198,N_1111,N_1144);
nor U1199 (N_1199,N_1123,N_1107);
nor U1200 (N_1200,N_1160,N_1172);
or U1201 (N_1201,N_1195,N_1156);
and U1202 (N_1202,N_1196,N_1180);
nand U1203 (N_1203,N_1165,N_1184);
nand U1204 (N_1204,N_1163,N_1150);
and U1205 (N_1205,N_1178,N_1192);
nand U1206 (N_1206,N_1170,N_1173);
nor U1207 (N_1207,N_1193,N_1169);
nand U1208 (N_1208,N_1158,N_1190);
or U1209 (N_1209,N_1188,N_1177);
nand U1210 (N_1210,N_1181,N_1168);
nor U1211 (N_1211,N_1189,N_1186);
and U1212 (N_1212,N_1187,N_1191);
nand U1213 (N_1213,N_1185,N_1154);
nand U1214 (N_1214,N_1159,N_1174);
or U1215 (N_1215,N_1198,N_1197);
or U1216 (N_1216,N_1194,N_1155);
and U1217 (N_1217,N_1151,N_1176);
and U1218 (N_1218,N_1153,N_1171);
nand U1219 (N_1219,N_1183,N_1167);
and U1220 (N_1220,N_1162,N_1164);
nand U1221 (N_1221,N_1199,N_1161);
nor U1222 (N_1222,N_1152,N_1166);
nor U1223 (N_1223,N_1175,N_1182);
and U1224 (N_1224,N_1179,N_1157);
nand U1225 (N_1225,N_1197,N_1169);
nor U1226 (N_1226,N_1172,N_1178);
or U1227 (N_1227,N_1184,N_1188);
nor U1228 (N_1228,N_1199,N_1166);
or U1229 (N_1229,N_1185,N_1192);
and U1230 (N_1230,N_1196,N_1155);
nor U1231 (N_1231,N_1169,N_1164);
or U1232 (N_1232,N_1198,N_1161);
nand U1233 (N_1233,N_1160,N_1178);
and U1234 (N_1234,N_1161,N_1173);
and U1235 (N_1235,N_1187,N_1176);
and U1236 (N_1236,N_1194,N_1161);
xnor U1237 (N_1237,N_1184,N_1183);
nand U1238 (N_1238,N_1182,N_1177);
or U1239 (N_1239,N_1158,N_1191);
nor U1240 (N_1240,N_1159,N_1184);
or U1241 (N_1241,N_1185,N_1199);
nor U1242 (N_1242,N_1171,N_1184);
nand U1243 (N_1243,N_1194,N_1169);
and U1244 (N_1244,N_1183,N_1187);
and U1245 (N_1245,N_1198,N_1175);
and U1246 (N_1246,N_1176,N_1168);
nor U1247 (N_1247,N_1156,N_1178);
nor U1248 (N_1248,N_1183,N_1197);
and U1249 (N_1249,N_1168,N_1193);
nor U1250 (N_1250,N_1215,N_1210);
nand U1251 (N_1251,N_1245,N_1242);
nand U1252 (N_1252,N_1247,N_1248);
nand U1253 (N_1253,N_1230,N_1223);
and U1254 (N_1254,N_1224,N_1235);
nand U1255 (N_1255,N_1219,N_1229);
nor U1256 (N_1256,N_1202,N_1200);
nor U1257 (N_1257,N_1208,N_1217);
nand U1258 (N_1258,N_1201,N_1211);
nand U1259 (N_1259,N_1213,N_1221);
or U1260 (N_1260,N_1238,N_1232);
nor U1261 (N_1261,N_1222,N_1214);
and U1262 (N_1262,N_1233,N_1234);
and U1263 (N_1263,N_1218,N_1244);
nand U1264 (N_1264,N_1207,N_1216);
nand U1265 (N_1265,N_1220,N_1227);
and U1266 (N_1266,N_1206,N_1225);
or U1267 (N_1267,N_1249,N_1212);
and U1268 (N_1268,N_1240,N_1241);
nor U1269 (N_1269,N_1209,N_1243);
nand U1270 (N_1270,N_1246,N_1203);
nor U1271 (N_1271,N_1239,N_1236);
and U1272 (N_1272,N_1226,N_1237);
and U1273 (N_1273,N_1204,N_1228);
nand U1274 (N_1274,N_1205,N_1231);
nand U1275 (N_1275,N_1206,N_1213);
or U1276 (N_1276,N_1227,N_1214);
and U1277 (N_1277,N_1239,N_1246);
nand U1278 (N_1278,N_1235,N_1232);
and U1279 (N_1279,N_1201,N_1227);
nand U1280 (N_1280,N_1214,N_1219);
nand U1281 (N_1281,N_1209,N_1223);
and U1282 (N_1282,N_1204,N_1236);
nor U1283 (N_1283,N_1228,N_1229);
xor U1284 (N_1284,N_1240,N_1233);
nor U1285 (N_1285,N_1246,N_1209);
or U1286 (N_1286,N_1224,N_1245);
and U1287 (N_1287,N_1209,N_1242);
and U1288 (N_1288,N_1242,N_1231);
or U1289 (N_1289,N_1221,N_1239);
nor U1290 (N_1290,N_1212,N_1204);
and U1291 (N_1291,N_1201,N_1213);
or U1292 (N_1292,N_1207,N_1221);
and U1293 (N_1293,N_1213,N_1224);
or U1294 (N_1294,N_1228,N_1217);
and U1295 (N_1295,N_1238,N_1208);
and U1296 (N_1296,N_1224,N_1205);
nor U1297 (N_1297,N_1244,N_1210);
and U1298 (N_1298,N_1231,N_1244);
nor U1299 (N_1299,N_1200,N_1209);
nor U1300 (N_1300,N_1268,N_1298);
and U1301 (N_1301,N_1250,N_1289);
or U1302 (N_1302,N_1272,N_1257);
nor U1303 (N_1303,N_1270,N_1290);
or U1304 (N_1304,N_1254,N_1251);
and U1305 (N_1305,N_1288,N_1275);
nor U1306 (N_1306,N_1252,N_1256);
and U1307 (N_1307,N_1253,N_1293);
nand U1308 (N_1308,N_1292,N_1280);
nor U1309 (N_1309,N_1263,N_1269);
and U1310 (N_1310,N_1283,N_1266);
and U1311 (N_1311,N_1264,N_1278);
nor U1312 (N_1312,N_1291,N_1282);
or U1313 (N_1313,N_1258,N_1297);
and U1314 (N_1314,N_1265,N_1296);
or U1315 (N_1315,N_1299,N_1267);
nand U1316 (N_1316,N_1277,N_1287);
nand U1317 (N_1317,N_1261,N_1262);
or U1318 (N_1318,N_1286,N_1281);
nand U1319 (N_1319,N_1255,N_1274);
nand U1320 (N_1320,N_1279,N_1276);
nor U1321 (N_1321,N_1259,N_1273);
nand U1322 (N_1322,N_1284,N_1294);
or U1323 (N_1323,N_1295,N_1285);
or U1324 (N_1324,N_1260,N_1271);
and U1325 (N_1325,N_1269,N_1264);
nand U1326 (N_1326,N_1293,N_1260);
or U1327 (N_1327,N_1261,N_1255);
nor U1328 (N_1328,N_1279,N_1281);
or U1329 (N_1329,N_1284,N_1290);
and U1330 (N_1330,N_1289,N_1298);
and U1331 (N_1331,N_1257,N_1295);
and U1332 (N_1332,N_1260,N_1257);
nand U1333 (N_1333,N_1296,N_1275);
nor U1334 (N_1334,N_1296,N_1288);
nand U1335 (N_1335,N_1293,N_1277);
nand U1336 (N_1336,N_1269,N_1295);
or U1337 (N_1337,N_1294,N_1297);
or U1338 (N_1338,N_1255,N_1292);
or U1339 (N_1339,N_1267,N_1250);
or U1340 (N_1340,N_1288,N_1287);
nor U1341 (N_1341,N_1287,N_1272);
nor U1342 (N_1342,N_1256,N_1299);
or U1343 (N_1343,N_1251,N_1281);
or U1344 (N_1344,N_1293,N_1254);
nand U1345 (N_1345,N_1261,N_1273);
or U1346 (N_1346,N_1293,N_1290);
xor U1347 (N_1347,N_1296,N_1282);
nor U1348 (N_1348,N_1254,N_1259);
nand U1349 (N_1349,N_1273,N_1264);
xor U1350 (N_1350,N_1301,N_1309);
nor U1351 (N_1351,N_1322,N_1304);
nor U1352 (N_1352,N_1346,N_1314);
nand U1353 (N_1353,N_1329,N_1313);
nand U1354 (N_1354,N_1342,N_1321);
and U1355 (N_1355,N_1311,N_1318);
or U1356 (N_1356,N_1325,N_1317);
or U1357 (N_1357,N_1327,N_1331);
nand U1358 (N_1358,N_1308,N_1312);
and U1359 (N_1359,N_1341,N_1328);
or U1360 (N_1360,N_1336,N_1340);
xor U1361 (N_1361,N_1338,N_1335);
nor U1362 (N_1362,N_1349,N_1343);
and U1363 (N_1363,N_1348,N_1316);
nor U1364 (N_1364,N_1310,N_1337);
or U1365 (N_1365,N_1344,N_1300);
and U1366 (N_1366,N_1302,N_1326);
and U1367 (N_1367,N_1345,N_1315);
nand U1368 (N_1368,N_1324,N_1320);
nand U1369 (N_1369,N_1307,N_1332);
nor U1370 (N_1370,N_1333,N_1339);
nor U1371 (N_1371,N_1319,N_1347);
nand U1372 (N_1372,N_1305,N_1323);
nor U1373 (N_1373,N_1334,N_1303);
and U1374 (N_1374,N_1330,N_1306);
or U1375 (N_1375,N_1327,N_1336);
nand U1376 (N_1376,N_1330,N_1339);
nand U1377 (N_1377,N_1337,N_1330);
or U1378 (N_1378,N_1304,N_1318);
and U1379 (N_1379,N_1316,N_1341);
nand U1380 (N_1380,N_1346,N_1329);
nor U1381 (N_1381,N_1342,N_1301);
or U1382 (N_1382,N_1339,N_1302);
nand U1383 (N_1383,N_1301,N_1331);
xor U1384 (N_1384,N_1326,N_1346);
nand U1385 (N_1385,N_1348,N_1338);
and U1386 (N_1386,N_1343,N_1329);
or U1387 (N_1387,N_1306,N_1344);
nor U1388 (N_1388,N_1300,N_1346);
nor U1389 (N_1389,N_1300,N_1327);
or U1390 (N_1390,N_1314,N_1310);
nand U1391 (N_1391,N_1308,N_1318);
xor U1392 (N_1392,N_1307,N_1303);
nor U1393 (N_1393,N_1305,N_1327);
nor U1394 (N_1394,N_1341,N_1301);
nor U1395 (N_1395,N_1338,N_1339);
or U1396 (N_1396,N_1324,N_1335);
and U1397 (N_1397,N_1325,N_1311);
nand U1398 (N_1398,N_1339,N_1325);
nand U1399 (N_1399,N_1307,N_1308);
and U1400 (N_1400,N_1398,N_1376);
or U1401 (N_1401,N_1350,N_1392);
or U1402 (N_1402,N_1368,N_1382);
or U1403 (N_1403,N_1386,N_1360);
nor U1404 (N_1404,N_1361,N_1357);
and U1405 (N_1405,N_1381,N_1351);
nor U1406 (N_1406,N_1390,N_1353);
nor U1407 (N_1407,N_1354,N_1363);
or U1408 (N_1408,N_1378,N_1377);
nor U1409 (N_1409,N_1389,N_1396);
nor U1410 (N_1410,N_1373,N_1399);
nand U1411 (N_1411,N_1370,N_1388);
nor U1412 (N_1412,N_1393,N_1395);
nor U1413 (N_1413,N_1372,N_1365);
nand U1414 (N_1414,N_1374,N_1369);
nand U1415 (N_1415,N_1384,N_1391);
or U1416 (N_1416,N_1358,N_1352);
or U1417 (N_1417,N_1364,N_1367);
nand U1418 (N_1418,N_1359,N_1394);
nor U1419 (N_1419,N_1385,N_1355);
nor U1420 (N_1420,N_1362,N_1379);
nand U1421 (N_1421,N_1366,N_1387);
nand U1422 (N_1422,N_1375,N_1397);
nand U1423 (N_1423,N_1356,N_1371);
or U1424 (N_1424,N_1383,N_1380);
nor U1425 (N_1425,N_1395,N_1359);
and U1426 (N_1426,N_1389,N_1390);
or U1427 (N_1427,N_1398,N_1382);
or U1428 (N_1428,N_1380,N_1367);
or U1429 (N_1429,N_1385,N_1381);
nor U1430 (N_1430,N_1364,N_1394);
or U1431 (N_1431,N_1359,N_1376);
nand U1432 (N_1432,N_1393,N_1388);
and U1433 (N_1433,N_1386,N_1384);
nor U1434 (N_1434,N_1385,N_1374);
and U1435 (N_1435,N_1373,N_1355);
nor U1436 (N_1436,N_1393,N_1365);
xor U1437 (N_1437,N_1388,N_1357);
nand U1438 (N_1438,N_1384,N_1372);
or U1439 (N_1439,N_1379,N_1386);
xor U1440 (N_1440,N_1366,N_1356);
and U1441 (N_1441,N_1394,N_1393);
nand U1442 (N_1442,N_1391,N_1387);
nor U1443 (N_1443,N_1364,N_1392);
and U1444 (N_1444,N_1380,N_1361);
nor U1445 (N_1445,N_1359,N_1355);
or U1446 (N_1446,N_1375,N_1385);
or U1447 (N_1447,N_1359,N_1356);
or U1448 (N_1448,N_1387,N_1369);
or U1449 (N_1449,N_1364,N_1352);
or U1450 (N_1450,N_1411,N_1403);
and U1451 (N_1451,N_1440,N_1421);
or U1452 (N_1452,N_1432,N_1444);
nand U1453 (N_1453,N_1424,N_1409);
and U1454 (N_1454,N_1420,N_1417);
nor U1455 (N_1455,N_1415,N_1405);
nand U1456 (N_1456,N_1449,N_1439);
and U1457 (N_1457,N_1418,N_1435);
nor U1458 (N_1458,N_1441,N_1404);
nand U1459 (N_1459,N_1428,N_1412);
nand U1460 (N_1460,N_1422,N_1429);
and U1461 (N_1461,N_1407,N_1443);
nand U1462 (N_1462,N_1426,N_1434);
nand U1463 (N_1463,N_1427,N_1425);
nand U1464 (N_1464,N_1447,N_1413);
and U1465 (N_1465,N_1446,N_1442);
and U1466 (N_1466,N_1438,N_1433);
nand U1467 (N_1467,N_1408,N_1416);
nand U1468 (N_1468,N_1431,N_1401);
and U1469 (N_1469,N_1423,N_1437);
and U1470 (N_1470,N_1436,N_1400);
and U1471 (N_1471,N_1430,N_1448);
or U1472 (N_1472,N_1402,N_1410);
nor U1473 (N_1473,N_1406,N_1414);
or U1474 (N_1474,N_1445,N_1419);
nor U1475 (N_1475,N_1404,N_1425);
and U1476 (N_1476,N_1406,N_1425);
and U1477 (N_1477,N_1400,N_1442);
or U1478 (N_1478,N_1419,N_1405);
and U1479 (N_1479,N_1423,N_1438);
and U1480 (N_1480,N_1421,N_1432);
nand U1481 (N_1481,N_1426,N_1420);
nor U1482 (N_1482,N_1443,N_1422);
nor U1483 (N_1483,N_1447,N_1422);
and U1484 (N_1484,N_1427,N_1406);
and U1485 (N_1485,N_1418,N_1410);
nor U1486 (N_1486,N_1413,N_1401);
and U1487 (N_1487,N_1420,N_1412);
xnor U1488 (N_1488,N_1434,N_1411);
and U1489 (N_1489,N_1427,N_1413);
and U1490 (N_1490,N_1433,N_1430);
or U1491 (N_1491,N_1409,N_1436);
xnor U1492 (N_1492,N_1436,N_1405);
or U1493 (N_1493,N_1424,N_1418);
and U1494 (N_1494,N_1436,N_1407);
or U1495 (N_1495,N_1427,N_1414);
or U1496 (N_1496,N_1400,N_1401);
and U1497 (N_1497,N_1404,N_1424);
nand U1498 (N_1498,N_1411,N_1409);
or U1499 (N_1499,N_1430,N_1447);
nand U1500 (N_1500,N_1486,N_1471);
and U1501 (N_1501,N_1465,N_1499);
and U1502 (N_1502,N_1487,N_1473);
or U1503 (N_1503,N_1458,N_1463);
and U1504 (N_1504,N_1460,N_1457);
nor U1505 (N_1505,N_1491,N_1459);
nand U1506 (N_1506,N_1488,N_1492);
nand U1507 (N_1507,N_1461,N_1477);
nor U1508 (N_1508,N_1476,N_1454);
nand U1509 (N_1509,N_1468,N_1470);
nand U1510 (N_1510,N_1484,N_1483);
nand U1511 (N_1511,N_1498,N_1494);
or U1512 (N_1512,N_1496,N_1467);
nand U1513 (N_1513,N_1456,N_1480);
and U1514 (N_1514,N_1472,N_1479);
nand U1515 (N_1515,N_1495,N_1475);
and U1516 (N_1516,N_1453,N_1490);
or U1517 (N_1517,N_1464,N_1485);
nor U1518 (N_1518,N_1489,N_1462);
nand U1519 (N_1519,N_1482,N_1493);
or U1520 (N_1520,N_1455,N_1469);
or U1521 (N_1521,N_1497,N_1466);
and U1522 (N_1522,N_1452,N_1474);
or U1523 (N_1523,N_1478,N_1451);
and U1524 (N_1524,N_1481,N_1450);
and U1525 (N_1525,N_1472,N_1457);
nand U1526 (N_1526,N_1454,N_1496);
nor U1527 (N_1527,N_1467,N_1469);
nand U1528 (N_1528,N_1471,N_1497);
nand U1529 (N_1529,N_1495,N_1454);
nand U1530 (N_1530,N_1451,N_1466);
nand U1531 (N_1531,N_1451,N_1493);
nand U1532 (N_1532,N_1451,N_1485);
or U1533 (N_1533,N_1477,N_1464);
and U1534 (N_1534,N_1465,N_1461);
and U1535 (N_1535,N_1499,N_1478);
nand U1536 (N_1536,N_1461,N_1467);
and U1537 (N_1537,N_1483,N_1499);
or U1538 (N_1538,N_1466,N_1498);
nor U1539 (N_1539,N_1485,N_1479);
nor U1540 (N_1540,N_1491,N_1465);
xor U1541 (N_1541,N_1473,N_1471);
xor U1542 (N_1542,N_1470,N_1476);
or U1543 (N_1543,N_1494,N_1461);
and U1544 (N_1544,N_1482,N_1470);
and U1545 (N_1545,N_1459,N_1463);
and U1546 (N_1546,N_1496,N_1473);
nand U1547 (N_1547,N_1453,N_1451);
nand U1548 (N_1548,N_1489,N_1491);
or U1549 (N_1549,N_1470,N_1457);
nand U1550 (N_1550,N_1516,N_1512);
and U1551 (N_1551,N_1515,N_1535);
or U1552 (N_1552,N_1503,N_1545);
nor U1553 (N_1553,N_1506,N_1538);
and U1554 (N_1554,N_1547,N_1532);
nand U1555 (N_1555,N_1530,N_1541);
nand U1556 (N_1556,N_1520,N_1527);
nand U1557 (N_1557,N_1513,N_1531);
or U1558 (N_1558,N_1518,N_1507);
nor U1559 (N_1559,N_1502,N_1508);
and U1560 (N_1560,N_1539,N_1548);
nor U1561 (N_1561,N_1542,N_1523);
and U1562 (N_1562,N_1525,N_1534);
or U1563 (N_1563,N_1511,N_1514);
or U1564 (N_1564,N_1529,N_1536);
and U1565 (N_1565,N_1549,N_1544);
or U1566 (N_1566,N_1522,N_1501);
or U1567 (N_1567,N_1546,N_1543);
or U1568 (N_1568,N_1528,N_1500);
and U1569 (N_1569,N_1517,N_1524);
and U1570 (N_1570,N_1504,N_1519);
or U1571 (N_1571,N_1505,N_1510);
or U1572 (N_1572,N_1509,N_1540);
or U1573 (N_1573,N_1521,N_1526);
nor U1574 (N_1574,N_1537,N_1533);
nor U1575 (N_1575,N_1511,N_1517);
and U1576 (N_1576,N_1532,N_1521);
nand U1577 (N_1577,N_1523,N_1511);
nand U1578 (N_1578,N_1536,N_1516);
or U1579 (N_1579,N_1519,N_1511);
or U1580 (N_1580,N_1525,N_1544);
nand U1581 (N_1581,N_1533,N_1511);
or U1582 (N_1582,N_1507,N_1515);
and U1583 (N_1583,N_1501,N_1547);
nand U1584 (N_1584,N_1502,N_1527);
nand U1585 (N_1585,N_1519,N_1506);
or U1586 (N_1586,N_1545,N_1531);
nor U1587 (N_1587,N_1509,N_1503);
nand U1588 (N_1588,N_1502,N_1500);
nor U1589 (N_1589,N_1512,N_1526);
or U1590 (N_1590,N_1502,N_1516);
and U1591 (N_1591,N_1512,N_1524);
and U1592 (N_1592,N_1531,N_1532);
and U1593 (N_1593,N_1503,N_1501);
or U1594 (N_1594,N_1544,N_1507);
and U1595 (N_1595,N_1516,N_1541);
nand U1596 (N_1596,N_1526,N_1523);
nor U1597 (N_1597,N_1528,N_1519);
nor U1598 (N_1598,N_1510,N_1517);
nand U1599 (N_1599,N_1527,N_1534);
nor U1600 (N_1600,N_1558,N_1582);
nor U1601 (N_1601,N_1590,N_1559);
nand U1602 (N_1602,N_1572,N_1551);
and U1603 (N_1603,N_1595,N_1567);
nor U1604 (N_1604,N_1597,N_1556);
and U1605 (N_1605,N_1565,N_1553);
nand U1606 (N_1606,N_1573,N_1552);
and U1607 (N_1607,N_1598,N_1574);
nand U1608 (N_1608,N_1563,N_1560);
and U1609 (N_1609,N_1566,N_1581);
nand U1610 (N_1610,N_1588,N_1592);
nand U1611 (N_1611,N_1569,N_1568);
or U1612 (N_1612,N_1555,N_1562);
and U1613 (N_1613,N_1586,N_1583);
nor U1614 (N_1614,N_1570,N_1580);
nand U1615 (N_1615,N_1587,N_1554);
or U1616 (N_1616,N_1575,N_1596);
nor U1617 (N_1617,N_1585,N_1591);
nand U1618 (N_1618,N_1576,N_1577);
and U1619 (N_1619,N_1561,N_1594);
and U1620 (N_1620,N_1589,N_1599);
and U1621 (N_1621,N_1578,N_1584);
nand U1622 (N_1622,N_1564,N_1571);
nand U1623 (N_1623,N_1593,N_1550);
nor U1624 (N_1624,N_1557,N_1579);
nand U1625 (N_1625,N_1585,N_1556);
nor U1626 (N_1626,N_1572,N_1596);
or U1627 (N_1627,N_1587,N_1550);
and U1628 (N_1628,N_1568,N_1577);
or U1629 (N_1629,N_1575,N_1598);
nor U1630 (N_1630,N_1598,N_1589);
nor U1631 (N_1631,N_1560,N_1599);
nor U1632 (N_1632,N_1566,N_1599);
nor U1633 (N_1633,N_1560,N_1580);
nor U1634 (N_1634,N_1588,N_1579);
and U1635 (N_1635,N_1580,N_1562);
or U1636 (N_1636,N_1564,N_1576);
nor U1637 (N_1637,N_1551,N_1594);
nand U1638 (N_1638,N_1556,N_1576);
xor U1639 (N_1639,N_1589,N_1569);
or U1640 (N_1640,N_1590,N_1552);
nor U1641 (N_1641,N_1590,N_1565);
nand U1642 (N_1642,N_1550,N_1581);
xnor U1643 (N_1643,N_1552,N_1597);
or U1644 (N_1644,N_1574,N_1576);
and U1645 (N_1645,N_1566,N_1571);
nor U1646 (N_1646,N_1599,N_1590);
nor U1647 (N_1647,N_1592,N_1596);
nand U1648 (N_1648,N_1592,N_1552);
and U1649 (N_1649,N_1580,N_1574);
and U1650 (N_1650,N_1606,N_1614);
nor U1651 (N_1651,N_1630,N_1603);
nor U1652 (N_1652,N_1628,N_1649);
nand U1653 (N_1653,N_1618,N_1605);
and U1654 (N_1654,N_1647,N_1642);
nand U1655 (N_1655,N_1632,N_1607);
nand U1656 (N_1656,N_1620,N_1616);
and U1657 (N_1657,N_1635,N_1631);
nor U1658 (N_1658,N_1636,N_1637);
and U1659 (N_1659,N_1608,N_1643);
or U1660 (N_1660,N_1609,N_1617);
and U1661 (N_1661,N_1646,N_1622);
nand U1662 (N_1662,N_1641,N_1623);
and U1663 (N_1663,N_1601,N_1634);
and U1664 (N_1664,N_1613,N_1611);
or U1665 (N_1665,N_1619,N_1612);
or U1666 (N_1666,N_1625,N_1633);
and U1667 (N_1667,N_1640,N_1602);
nand U1668 (N_1668,N_1629,N_1648);
or U1669 (N_1669,N_1644,N_1621);
or U1670 (N_1670,N_1624,N_1626);
or U1671 (N_1671,N_1604,N_1610);
nand U1672 (N_1672,N_1615,N_1638);
and U1673 (N_1673,N_1600,N_1627);
and U1674 (N_1674,N_1639,N_1645);
xor U1675 (N_1675,N_1612,N_1607);
and U1676 (N_1676,N_1632,N_1602);
nand U1677 (N_1677,N_1648,N_1604);
nor U1678 (N_1678,N_1619,N_1632);
and U1679 (N_1679,N_1619,N_1611);
nor U1680 (N_1680,N_1631,N_1612);
or U1681 (N_1681,N_1619,N_1605);
and U1682 (N_1682,N_1608,N_1602);
and U1683 (N_1683,N_1615,N_1635);
nand U1684 (N_1684,N_1601,N_1605);
nand U1685 (N_1685,N_1623,N_1606);
nor U1686 (N_1686,N_1641,N_1649);
nor U1687 (N_1687,N_1636,N_1633);
or U1688 (N_1688,N_1643,N_1614);
nand U1689 (N_1689,N_1626,N_1616);
or U1690 (N_1690,N_1603,N_1644);
and U1691 (N_1691,N_1615,N_1603);
nand U1692 (N_1692,N_1615,N_1618);
and U1693 (N_1693,N_1612,N_1630);
xor U1694 (N_1694,N_1638,N_1620);
nor U1695 (N_1695,N_1625,N_1619);
nand U1696 (N_1696,N_1602,N_1638);
and U1697 (N_1697,N_1643,N_1600);
and U1698 (N_1698,N_1630,N_1648);
nor U1699 (N_1699,N_1626,N_1628);
nand U1700 (N_1700,N_1673,N_1676);
nor U1701 (N_1701,N_1697,N_1678);
and U1702 (N_1702,N_1690,N_1670);
nor U1703 (N_1703,N_1671,N_1681);
and U1704 (N_1704,N_1665,N_1680);
xor U1705 (N_1705,N_1672,N_1684);
nor U1706 (N_1706,N_1699,N_1696);
and U1707 (N_1707,N_1653,N_1650);
nor U1708 (N_1708,N_1675,N_1666);
and U1709 (N_1709,N_1695,N_1683);
and U1710 (N_1710,N_1663,N_1688);
and U1711 (N_1711,N_1652,N_1668);
and U1712 (N_1712,N_1661,N_1654);
nor U1713 (N_1713,N_1656,N_1691);
or U1714 (N_1714,N_1698,N_1664);
nand U1715 (N_1715,N_1686,N_1687);
nor U1716 (N_1716,N_1689,N_1679);
nand U1717 (N_1717,N_1677,N_1694);
and U1718 (N_1718,N_1692,N_1662);
and U1719 (N_1719,N_1682,N_1657);
nor U1720 (N_1720,N_1674,N_1660);
or U1721 (N_1721,N_1693,N_1651);
nor U1722 (N_1722,N_1659,N_1655);
or U1723 (N_1723,N_1658,N_1667);
nand U1724 (N_1724,N_1669,N_1685);
or U1725 (N_1725,N_1689,N_1675);
or U1726 (N_1726,N_1656,N_1670);
nand U1727 (N_1727,N_1676,N_1693);
and U1728 (N_1728,N_1662,N_1660);
nand U1729 (N_1729,N_1668,N_1671);
nand U1730 (N_1730,N_1670,N_1688);
nor U1731 (N_1731,N_1669,N_1661);
and U1732 (N_1732,N_1683,N_1680);
or U1733 (N_1733,N_1683,N_1666);
nor U1734 (N_1734,N_1687,N_1671);
and U1735 (N_1735,N_1693,N_1673);
nor U1736 (N_1736,N_1667,N_1664);
and U1737 (N_1737,N_1687,N_1692);
nand U1738 (N_1738,N_1650,N_1664);
xor U1739 (N_1739,N_1699,N_1693);
or U1740 (N_1740,N_1669,N_1652);
nand U1741 (N_1741,N_1667,N_1697);
nor U1742 (N_1742,N_1662,N_1671);
or U1743 (N_1743,N_1651,N_1687);
nor U1744 (N_1744,N_1656,N_1662);
or U1745 (N_1745,N_1650,N_1668);
nand U1746 (N_1746,N_1658,N_1687);
and U1747 (N_1747,N_1651,N_1660);
or U1748 (N_1748,N_1655,N_1681);
or U1749 (N_1749,N_1684,N_1673);
nand U1750 (N_1750,N_1703,N_1706);
nand U1751 (N_1751,N_1708,N_1702);
nand U1752 (N_1752,N_1739,N_1721);
and U1753 (N_1753,N_1737,N_1713);
or U1754 (N_1754,N_1732,N_1719);
or U1755 (N_1755,N_1700,N_1727);
or U1756 (N_1756,N_1710,N_1718);
and U1757 (N_1757,N_1701,N_1742);
nor U1758 (N_1758,N_1745,N_1743);
nand U1759 (N_1759,N_1730,N_1728);
and U1760 (N_1760,N_1716,N_1705);
nand U1761 (N_1761,N_1740,N_1707);
xor U1762 (N_1762,N_1734,N_1744);
nand U1763 (N_1763,N_1715,N_1729);
nand U1764 (N_1764,N_1726,N_1738);
and U1765 (N_1765,N_1733,N_1720);
and U1766 (N_1766,N_1717,N_1747);
nor U1767 (N_1767,N_1711,N_1736);
nor U1768 (N_1768,N_1731,N_1725);
nor U1769 (N_1769,N_1714,N_1724);
and U1770 (N_1770,N_1749,N_1746);
nor U1771 (N_1771,N_1748,N_1709);
or U1772 (N_1772,N_1741,N_1712);
and U1773 (N_1773,N_1704,N_1722);
nor U1774 (N_1774,N_1735,N_1723);
and U1775 (N_1775,N_1724,N_1739);
nand U1776 (N_1776,N_1720,N_1725);
nand U1777 (N_1777,N_1734,N_1706);
and U1778 (N_1778,N_1712,N_1736);
nor U1779 (N_1779,N_1721,N_1705);
nor U1780 (N_1780,N_1746,N_1725);
xor U1781 (N_1781,N_1744,N_1736);
nand U1782 (N_1782,N_1717,N_1725);
or U1783 (N_1783,N_1737,N_1726);
nor U1784 (N_1784,N_1709,N_1749);
and U1785 (N_1785,N_1720,N_1748);
xor U1786 (N_1786,N_1725,N_1708);
nand U1787 (N_1787,N_1712,N_1743);
and U1788 (N_1788,N_1743,N_1724);
nor U1789 (N_1789,N_1723,N_1734);
and U1790 (N_1790,N_1721,N_1740);
xnor U1791 (N_1791,N_1705,N_1700);
and U1792 (N_1792,N_1725,N_1739);
nor U1793 (N_1793,N_1709,N_1716);
xor U1794 (N_1794,N_1742,N_1740);
nor U1795 (N_1795,N_1718,N_1702);
or U1796 (N_1796,N_1729,N_1726);
and U1797 (N_1797,N_1726,N_1710);
and U1798 (N_1798,N_1748,N_1706);
or U1799 (N_1799,N_1742,N_1712);
nor U1800 (N_1800,N_1756,N_1797);
or U1801 (N_1801,N_1798,N_1799);
and U1802 (N_1802,N_1778,N_1788);
nand U1803 (N_1803,N_1768,N_1760);
nand U1804 (N_1804,N_1791,N_1762);
and U1805 (N_1805,N_1771,N_1761);
nor U1806 (N_1806,N_1777,N_1764);
nand U1807 (N_1807,N_1759,N_1795);
nand U1808 (N_1808,N_1773,N_1769);
nand U1809 (N_1809,N_1775,N_1766);
nand U1810 (N_1810,N_1789,N_1770);
nand U1811 (N_1811,N_1767,N_1785);
nand U1812 (N_1812,N_1781,N_1763);
nor U1813 (N_1813,N_1755,N_1794);
and U1814 (N_1814,N_1772,N_1776);
or U1815 (N_1815,N_1779,N_1752);
or U1816 (N_1816,N_1783,N_1786);
nor U1817 (N_1817,N_1792,N_1750);
xor U1818 (N_1818,N_1757,N_1753);
nand U1819 (N_1819,N_1751,N_1774);
nand U1820 (N_1820,N_1754,N_1787);
nor U1821 (N_1821,N_1765,N_1784);
nor U1822 (N_1822,N_1790,N_1793);
nor U1823 (N_1823,N_1758,N_1796);
or U1824 (N_1824,N_1782,N_1780);
or U1825 (N_1825,N_1755,N_1788);
nand U1826 (N_1826,N_1768,N_1774);
and U1827 (N_1827,N_1781,N_1776);
and U1828 (N_1828,N_1798,N_1751);
or U1829 (N_1829,N_1772,N_1793);
xor U1830 (N_1830,N_1771,N_1770);
nand U1831 (N_1831,N_1772,N_1790);
or U1832 (N_1832,N_1764,N_1769);
and U1833 (N_1833,N_1768,N_1793);
nand U1834 (N_1834,N_1780,N_1787);
nand U1835 (N_1835,N_1773,N_1788);
nand U1836 (N_1836,N_1789,N_1782);
or U1837 (N_1837,N_1789,N_1779);
nor U1838 (N_1838,N_1794,N_1768);
or U1839 (N_1839,N_1761,N_1751);
or U1840 (N_1840,N_1757,N_1751);
nand U1841 (N_1841,N_1798,N_1771);
or U1842 (N_1842,N_1778,N_1757);
or U1843 (N_1843,N_1789,N_1771);
nand U1844 (N_1844,N_1762,N_1752);
nand U1845 (N_1845,N_1790,N_1754);
or U1846 (N_1846,N_1789,N_1786);
nand U1847 (N_1847,N_1786,N_1798);
or U1848 (N_1848,N_1771,N_1772);
xnor U1849 (N_1849,N_1761,N_1757);
or U1850 (N_1850,N_1821,N_1814);
or U1851 (N_1851,N_1820,N_1827);
xor U1852 (N_1852,N_1834,N_1816);
nand U1853 (N_1853,N_1839,N_1840);
nand U1854 (N_1854,N_1849,N_1801);
and U1855 (N_1855,N_1815,N_1832);
nand U1856 (N_1856,N_1843,N_1800);
nor U1857 (N_1857,N_1802,N_1841);
and U1858 (N_1858,N_1811,N_1804);
or U1859 (N_1859,N_1813,N_1846);
or U1860 (N_1860,N_1817,N_1845);
nand U1861 (N_1861,N_1829,N_1824);
nand U1862 (N_1862,N_1848,N_1809);
nor U1863 (N_1863,N_1803,N_1825);
nand U1864 (N_1864,N_1833,N_1818);
nor U1865 (N_1865,N_1805,N_1808);
nand U1866 (N_1866,N_1807,N_1826);
or U1867 (N_1867,N_1823,N_1844);
nor U1868 (N_1868,N_1830,N_1812);
or U1869 (N_1869,N_1806,N_1831);
nor U1870 (N_1870,N_1836,N_1810);
and U1871 (N_1871,N_1842,N_1847);
or U1872 (N_1872,N_1837,N_1819);
and U1873 (N_1873,N_1822,N_1835);
nand U1874 (N_1874,N_1828,N_1838);
nand U1875 (N_1875,N_1829,N_1807);
and U1876 (N_1876,N_1811,N_1813);
nor U1877 (N_1877,N_1831,N_1838);
and U1878 (N_1878,N_1819,N_1825);
nand U1879 (N_1879,N_1834,N_1848);
nand U1880 (N_1880,N_1838,N_1817);
and U1881 (N_1881,N_1819,N_1820);
and U1882 (N_1882,N_1817,N_1831);
or U1883 (N_1883,N_1849,N_1820);
and U1884 (N_1884,N_1815,N_1825);
or U1885 (N_1885,N_1847,N_1810);
nor U1886 (N_1886,N_1802,N_1830);
nand U1887 (N_1887,N_1830,N_1809);
or U1888 (N_1888,N_1811,N_1839);
nor U1889 (N_1889,N_1834,N_1823);
or U1890 (N_1890,N_1836,N_1822);
or U1891 (N_1891,N_1812,N_1822);
nor U1892 (N_1892,N_1842,N_1828);
nor U1893 (N_1893,N_1825,N_1831);
nor U1894 (N_1894,N_1844,N_1846);
nor U1895 (N_1895,N_1845,N_1828);
nand U1896 (N_1896,N_1844,N_1833);
nor U1897 (N_1897,N_1826,N_1821);
or U1898 (N_1898,N_1813,N_1815);
and U1899 (N_1899,N_1840,N_1831);
nor U1900 (N_1900,N_1882,N_1875);
nor U1901 (N_1901,N_1886,N_1860);
nor U1902 (N_1902,N_1868,N_1881);
nor U1903 (N_1903,N_1897,N_1877);
and U1904 (N_1904,N_1887,N_1858);
or U1905 (N_1905,N_1870,N_1891);
or U1906 (N_1906,N_1883,N_1871);
nor U1907 (N_1907,N_1865,N_1873);
nor U1908 (N_1908,N_1879,N_1859);
nor U1909 (N_1909,N_1880,N_1888);
nand U1910 (N_1910,N_1862,N_1895);
nand U1911 (N_1911,N_1854,N_1851);
or U1912 (N_1912,N_1899,N_1894);
and U1913 (N_1913,N_1869,N_1861);
nand U1914 (N_1914,N_1874,N_1866);
xor U1915 (N_1915,N_1876,N_1872);
or U1916 (N_1916,N_1857,N_1850);
or U1917 (N_1917,N_1852,N_1867);
and U1918 (N_1918,N_1893,N_1885);
nand U1919 (N_1919,N_1856,N_1855);
and U1920 (N_1920,N_1853,N_1896);
nor U1921 (N_1921,N_1884,N_1864);
and U1922 (N_1922,N_1898,N_1878);
or U1923 (N_1923,N_1889,N_1890);
and U1924 (N_1924,N_1892,N_1863);
and U1925 (N_1925,N_1861,N_1882);
nand U1926 (N_1926,N_1858,N_1873);
or U1927 (N_1927,N_1889,N_1857);
and U1928 (N_1928,N_1863,N_1877);
and U1929 (N_1929,N_1889,N_1853);
nand U1930 (N_1930,N_1889,N_1891);
nor U1931 (N_1931,N_1866,N_1893);
nor U1932 (N_1932,N_1863,N_1874);
and U1933 (N_1933,N_1872,N_1875);
nand U1934 (N_1934,N_1888,N_1876);
nor U1935 (N_1935,N_1874,N_1872);
and U1936 (N_1936,N_1850,N_1898);
nor U1937 (N_1937,N_1884,N_1858);
or U1938 (N_1938,N_1865,N_1856);
nor U1939 (N_1939,N_1859,N_1868);
nand U1940 (N_1940,N_1863,N_1859);
or U1941 (N_1941,N_1886,N_1854);
nor U1942 (N_1942,N_1898,N_1893);
nor U1943 (N_1943,N_1886,N_1884);
or U1944 (N_1944,N_1876,N_1881);
and U1945 (N_1945,N_1883,N_1893);
and U1946 (N_1946,N_1860,N_1852);
or U1947 (N_1947,N_1857,N_1870);
and U1948 (N_1948,N_1862,N_1850);
nand U1949 (N_1949,N_1898,N_1897);
nand U1950 (N_1950,N_1905,N_1929);
and U1951 (N_1951,N_1922,N_1933);
or U1952 (N_1952,N_1906,N_1917);
nand U1953 (N_1953,N_1935,N_1949);
nand U1954 (N_1954,N_1908,N_1938);
xnor U1955 (N_1955,N_1934,N_1911);
or U1956 (N_1956,N_1924,N_1930);
or U1957 (N_1957,N_1931,N_1919);
and U1958 (N_1958,N_1909,N_1928);
nor U1959 (N_1959,N_1920,N_1910);
or U1960 (N_1960,N_1903,N_1907);
nor U1961 (N_1961,N_1943,N_1925);
nand U1962 (N_1962,N_1904,N_1913);
or U1963 (N_1963,N_1916,N_1918);
nor U1964 (N_1964,N_1926,N_1932);
or U1965 (N_1965,N_1927,N_1941);
and U1966 (N_1966,N_1946,N_1901);
and U1967 (N_1967,N_1936,N_1921);
and U1968 (N_1968,N_1914,N_1937);
nor U1969 (N_1969,N_1923,N_1947);
nor U1970 (N_1970,N_1940,N_1939);
nor U1971 (N_1971,N_1900,N_1945);
nor U1972 (N_1972,N_1915,N_1912);
nand U1973 (N_1973,N_1942,N_1948);
nor U1974 (N_1974,N_1902,N_1944);
xor U1975 (N_1975,N_1935,N_1936);
nand U1976 (N_1976,N_1940,N_1943);
and U1977 (N_1977,N_1945,N_1917);
and U1978 (N_1978,N_1932,N_1901);
nand U1979 (N_1979,N_1931,N_1937);
nor U1980 (N_1980,N_1923,N_1949);
or U1981 (N_1981,N_1941,N_1902);
xnor U1982 (N_1982,N_1931,N_1910);
nor U1983 (N_1983,N_1925,N_1922);
nand U1984 (N_1984,N_1939,N_1922);
or U1985 (N_1985,N_1917,N_1932);
nor U1986 (N_1986,N_1907,N_1936);
nor U1987 (N_1987,N_1931,N_1944);
nand U1988 (N_1988,N_1913,N_1901);
nor U1989 (N_1989,N_1937,N_1947);
nand U1990 (N_1990,N_1913,N_1932);
nor U1991 (N_1991,N_1941,N_1923);
nand U1992 (N_1992,N_1906,N_1944);
or U1993 (N_1993,N_1924,N_1912);
nand U1994 (N_1994,N_1943,N_1935);
nand U1995 (N_1995,N_1902,N_1921);
and U1996 (N_1996,N_1930,N_1906);
and U1997 (N_1997,N_1928,N_1947);
or U1998 (N_1998,N_1900,N_1901);
nor U1999 (N_1999,N_1936,N_1903);
or U2000 (N_2000,N_1985,N_1988);
or U2001 (N_2001,N_1976,N_1957);
and U2002 (N_2002,N_1961,N_1954);
nand U2003 (N_2003,N_1953,N_1987);
or U2004 (N_2004,N_1964,N_1952);
or U2005 (N_2005,N_1950,N_1973);
nor U2006 (N_2006,N_1970,N_1968);
and U2007 (N_2007,N_1990,N_1992);
and U2008 (N_2008,N_1995,N_1963);
or U2009 (N_2009,N_1994,N_1997);
nor U2010 (N_2010,N_1977,N_1974);
or U2011 (N_2011,N_1978,N_1986);
nor U2012 (N_2012,N_1967,N_1980);
nor U2013 (N_2013,N_1989,N_1965);
or U2014 (N_2014,N_1993,N_1960);
or U2015 (N_2015,N_1996,N_1983);
xor U2016 (N_2016,N_1951,N_1982);
nand U2017 (N_2017,N_1981,N_1975);
and U2018 (N_2018,N_1984,N_1956);
nand U2019 (N_2019,N_1999,N_1998);
xnor U2020 (N_2020,N_1962,N_1958);
nor U2021 (N_2021,N_1991,N_1971);
or U2022 (N_2022,N_1959,N_1979);
and U2023 (N_2023,N_1972,N_1966);
xor U2024 (N_2024,N_1955,N_1969);
nand U2025 (N_2025,N_1976,N_1993);
nor U2026 (N_2026,N_1980,N_1982);
nor U2027 (N_2027,N_1976,N_1975);
nand U2028 (N_2028,N_1960,N_1989);
and U2029 (N_2029,N_1992,N_1977);
or U2030 (N_2030,N_1957,N_1955);
or U2031 (N_2031,N_1991,N_1985);
or U2032 (N_2032,N_1977,N_1998);
or U2033 (N_2033,N_1979,N_1960);
nor U2034 (N_2034,N_1988,N_1978);
xnor U2035 (N_2035,N_1983,N_1974);
nor U2036 (N_2036,N_1993,N_1977);
nand U2037 (N_2037,N_1989,N_1969);
nand U2038 (N_2038,N_1973,N_1963);
and U2039 (N_2039,N_1996,N_1969);
nor U2040 (N_2040,N_1991,N_1988);
nand U2041 (N_2041,N_1966,N_1964);
and U2042 (N_2042,N_1953,N_1952);
or U2043 (N_2043,N_1982,N_1955);
and U2044 (N_2044,N_1961,N_1995);
nor U2045 (N_2045,N_1955,N_1983);
or U2046 (N_2046,N_1972,N_1991);
and U2047 (N_2047,N_1958,N_1982);
or U2048 (N_2048,N_1964,N_1967);
nand U2049 (N_2049,N_1962,N_1967);
nor U2050 (N_2050,N_2024,N_2048);
nand U2051 (N_2051,N_2035,N_2031);
and U2052 (N_2052,N_2000,N_2002);
nand U2053 (N_2053,N_2023,N_2028);
nor U2054 (N_2054,N_2015,N_2004);
nand U2055 (N_2055,N_2038,N_2016);
and U2056 (N_2056,N_2025,N_2009);
nand U2057 (N_2057,N_2034,N_2026);
nand U2058 (N_2058,N_2032,N_2008);
nand U2059 (N_2059,N_2020,N_2041);
and U2060 (N_2060,N_2033,N_2012);
and U2061 (N_2061,N_2046,N_2039);
nor U2062 (N_2062,N_2027,N_2010);
or U2063 (N_2063,N_2017,N_2030);
or U2064 (N_2064,N_2018,N_2013);
or U2065 (N_2065,N_2003,N_2047);
nor U2066 (N_2066,N_2019,N_2045);
nand U2067 (N_2067,N_2001,N_2043);
and U2068 (N_2068,N_2044,N_2021);
or U2069 (N_2069,N_2022,N_2029);
or U2070 (N_2070,N_2036,N_2005);
or U2071 (N_2071,N_2037,N_2007);
nor U2072 (N_2072,N_2042,N_2011);
nand U2073 (N_2073,N_2014,N_2040);
nand U2074 (N_2074,N_2006,N_2049);
nand U2075 (N_2075,N_2024,N_2031);
or U2076 (N_2076,N_2005,N_2006);
nor U2077 (N_2077,N_2019,N_2010);
nand U2078 (N_2078,N_2014,N_2031);
nand U2079 (N_2079,N_2018,N_2024);
nand U2080 (N_2080,N_2016,N_2017);
nor U2081 (N_2081,N_2000,N_2017);
nor U2082 (N_2082,N_2022,N_2042);
nor U2083 (N_2083,N_2015,N_2035);
nand U2084 (N_2084,N_2025,N_2001);
or U2085 (N_2085,N_2009,N_2002);
nand U2086 (N_2086,N_2004,N_2017);
nor U2087 (N_2087,N_2015,N_2045);
nor U2088 (N_2088,N_2003,N_2027);
and U2089 (N_2089,N_2028,N_2042);
nor U2090 (N_2090,N_2038,N_2014);
nor U2091 (N_2091,N_2046,N_2023);
or U2092 (N_2092,N_2015,N_2017);
and U2093 (N_2093,N_2043,N_2007);
and U2094 (N_2094,N_2045,N_2034);
nor U2095 (N_2095,N_2047,N_2048);
and U2096 (N_2096,N_2024,N_2000);
nand U2097 (N_2097,N_2029,N_2032);
nor U2098 (N_2098,N_2008,N_2020);
or U2099 (N_2099,N_2031,N_2015);
nand U2100 (N_2100,N_2071,N_2092);
nand U2101 (N_2101,N_2077,N_2065);
and U2102 (N_2102,N_2083,N_2066);
nand U2103 (N_2103,N_2068,N_2094);
nor U2104 (N_2104,N_2084,N_2090);
or U2105 (N_2105,N_2054,N_2053);
or U2106 (N_2106,N_2073,N_2079);
xor U2107 (N_2107,N_2099,N_2088);
and U2108 (N_2108,N_2078,N_2060);
nand U2109 (N_2109,N_2058,N_2052);
nor U2110 (N_2110,N_2087,N_2081);
and U2111 (N_2111,N_2076,N_2056);
and U2112 (N_2112,N_2074,N_2064);
or U2113 (N_2113,N_2050,N_2085);
nor U2114 (N_2114,N_2069,N_2093);
or U2115 (N_2115,N_2059,N_2080);
nand U2116 (N_2116,N_2062,N_2096);
and U2117 (N_2117,N_2061,N_2051);
nor U2118 (N_2118,N_2072,N_2097);
nor U2119 (N_2119,N_2089,N_2055);
nand U2120 (N_2120,N_2095,N_2067);
or U2121 (N_2121,N_2057,N_2098);
or U2122 (N_2122,N_2063,N_2082);
nand U2123 (N_2123,N_2091,N_2075);
nand U2124 (N_2124,N_2086,N_2070);
nand U2125 (N_2125,N_2090,N_2083);
or U2126 (N_2126,N_2068,N_2052);
nor U2127 (N_2127,N_2051,N_2085);
and U2128 (N_2128,N_2099,N_2094);
nor U2129 (N_2129,N_2083,N_2055);
or U2130 (N_2130,N_2062,N_2059);
xnor U2131 (N_2131,N_2091,N_2087);
nand U2132 (N_2132,N_2071,N_2081);
and U2133 (N_2133,N_2053,N_2052);
or U2134 (N_2134,N_2054,N_2058);
nor U2135 (N_2135,N_2059,N_2095);
nor U2136 (N_2136,N_2050,N_2066);
nor U2137 (N_2137,N_2080,N_2085);
nand U2138 (N_2138,N_2062,N_2075);
or U2139 (N_2139,N_2077,N_2089);
or U2140 (N_2140,N_2062,N_2051);
nand U2141 (N_2141,N_2087,N_2084);
nand U2142 (N_2142,N_2062,N_2054);
or U2143 (N_2143,N_2086,N_2064);
and U2144 (N_2144,N_2052,N_2095);
nor U2145 (N_2145,N_2057,N_2090);
or U2146 (N_2146,N_2058,N_2082);
and U2147 (N_2147,N_2061,N_2057);
nand U2148 (N_2148,N_2055,N_2073);
nor U2149 (N_2149,N_2080,N_2057);
nand U2150 (N_2150,N_2144,N_2111);
nand U2151 (N_2151,N_2138,N_2146);
nor U2152 (N_2152,N_2126,N_2100);
nor U2153 (N_2153,N_2120,N_2109);
or U2154 (N_2154,N_2143,N_2134);
nand U2155 (N_2155,N_2114,N_2108);
or U2156 (N_2156,N_2147,N_2136);
or U2157 (N_2157,N_2149,N_2118);
and U2158 (N_2158,N_2110,N_2129);
nor U2159 (N_2159,N_2113,N_2132);
or U2160 (N_2160,N_2133,N_2123);
nand U2161 (N_2161,N_2140,N_2107);
and U2162 (N_2162,N_2105,N_2101);
and U2163 (N_2163,N_2128,N_2139);
or U2164 (N_2164,N_2119,N_2141);
or U2165 (N_2165,N_2125,N_2148);
and U2166 (N_2166,N_2104,N_2130);
nand U2167 (N_2167,N_2103,N_2112);
or U2168 (N_2168,N_2145,N_2131);
and U2169 (N_2169,N_2102,N_2124);
nand U2170 (N_2170,N_2135,N_2106);
nand U2171 (N_2171,N_2142,N_2121);
and U2172 (N_2172,N_2116,N_2122);
nor U2173 (N_2173,N_2115,N_2117);
or U2174 (N_2174,N_2127,N_2137);
nand U2175 (N_2175,N_2122,N_2133);
nand U2176 (N_2176,N_2106,N_2144);
nor U2177 (N_2177,N_2132,N_2129);
xor U2178 (N_2178,N_2135,N_2112);
nor U2179 (N_2179,N_2118,N_2112);
and U2180 (N_2180,N_2149,N_2104);
nor U2181 (N_2181,N_2126,N_2124);
or U2182 (N_2182,N_2131,N_2100);
nand U2183 (N_2183,N_2146,N_2128);
and U2184 (N_2184,N_2117,N_2106);
nand U2185 (N_2185,N_2145,N_2129);
nor U2186 (N_2186,N_2125,N_2133);
and U2187 (N_2187,N_2104,N_2121);
nor U2188 (N_2188,N_2128,N_2144);
nor U2189 (N_2189,N_2119,N_2148);
nand U2190 (N_2190,N_2108,N_2124);
nor U2191 (N_2191,N_2142,N_2100);
and U2192 (N_2192,N_2135,N_2142);
nor U2193 (N_2193,N_2101,N_2132);
or U2194 (N_2194,N_2132,N_2126);
and U2195 (N_2195,N_2129,N_2141);
or U2196 (N_2196,N_2144,N_2140);
xor U2197 (N_2197,N_2121,N_2129);
or U2198 (N_2198,N_2103,N_2115);
or U2199 (N_2199,N_2135,N_2126);
and U2200 (N_2200,N_2190,N_2191);
and U2201 (N_2201,N_2150,N_2174);
nand U2202 (N_2202,N_2193,N_2197);
nand U2203 (N_2203,N_2164,N_2153);
and U2204 (N_2204,N_2175,N_2188);
nand U2205 (N_2205,N_2184,N_2180);
and U2206 (N_2206,N_2194,N_2161);
nand U2207 (N_2207,N_2158,N_2166);
nand U2208 (N_2208,N_2170,N_2156);
nor U2209 (N_2209,N_2173,N_2176);
and U2210 (N_2210,N_2154,N_2179);
and U2211 (N_2211,N_2199,N_2198);
nand U2212 (N_2212,N_2155,N_2167);
and U2213 (N_2213,N_2171,N_2192);
nand U2214 (N_2214,N_2163,N_2152);
nor U2215 (N_2215,N_2187,N_2169);
and U2216 (N_2216,N_2182,N_2168);
nand U2217 (N_2217,N_2186,N_2189);
nor U2218 (N_2218,N_2162,N_2185);
nor U2219 (N_2219,N_2172,N_2195);
nand U2220 (N_2220,N_2151,N_2159);
and U2221 (N_2221,N_2183,N_2177);
and U2222 (N_2222,N_2157,N_2160);
and U2223 (N_2223,N_2181,N_2165);
and U2224 (N_2224,N_2178,N_2196);
nor U2225 (N_2225,N_2154,N_2182);
nand U2226 (N_2226,N_2156,N_2164);
or U2227 (N_2227,N_2172,N_2171);
and U2228 (N_2228,N_2190,N_2177);
or U2229 (N_2229,N_2199,N_2157);
and U2230 (N_2230,N_2150,N_2187);
nand U2231 (N_2231,N_2193,N_2171);
or U2232 (N_2232,N_2168,N_2155);
nor U2233 (N_2233,N_2198,N_2189);
nand U2234 (N_2234,N_2158,N_2151);
nand U2235 (N_2235,N_2160,N_2182);
nor U2236 (N_2236,N_2193,N_2175);
and U2237 (N_2237,N_2185,N_2179);
nand U2238 (N_2238,N_2165,N_2184);
nor U2239 (N_2239,N_2180,N_2175);
nor U2240 (N_2240,N_2159,N_2178);
nor U2241 (N_2241,N_2194,N_2199);
nor U2242 (N_2242,N_2198,N_2156);
nand U2243 (N_2243,N_2184,N_2150);
nor U2244 (N_2244,N_2150,N_2168);
xor U2245 (N_2245,N_2153,N_2197);
nor U2246 (N_2246,N_2164,N_2158);
or U2247 (N_2247,N_2157,N_2178);
nor U2248 (N_2248,N_2191,N_2169);
nand U2249 (N_2249,N_2183,N_2151);
nor U2250 (N_2250,N_2245,N_2243);
or U2251 (N_2251,N_2230,N_2229);
or U2252 (N_2252,N_2204,N_2249);
or U2253 (N_2253,N_2223,N_2236);
nor U2254 (N_2254,N_2218,N_2238);
and U2255 (N_2255,N_2233,N_2205);
or U2256 (N_2256,N_2206,N_2213);
or U2257 (N_2257,N_2207,N_2239);
or U2258 (N_2258,N_2219,N_2247);
nand U2259 (N_2259,N_2244,N_2240);
and U2260 (N_2260,N_2234,N_2212);
nor U2261 (N_2261,N_2201,N_2227);
and U2262 (N_2262,N_2235,N_2217);
or U2263 (N_2263,N_2232,N_2216);
and U2264 (N_2264,N_2214,N_2200);
or U2265 (N_2265,N_2215,N_2211);
or U2266 (N_2266,N_2208,N_2210);
and U2267 (N_2267,N_2202,N_2226);
and U2268 (N_2268,N_2224,N_2222);
or U2269 (N_2269,N_2203,N_2221);
or U2270 (N_2270,N_2248,N_2246);
nor U2271 (N_2271,N_2231,N_2220);
and U2272 (N_2272,N_2225,N_2228);
or U2273 (N_2273,N_2242,N_2237);
and U2274 (N_2274,N_2241,N_2209);
or U2275 (N_2275,N_2238,N_2230);
nand U2276 (N_2276,N_2236,N_2203);
or U2277 (N_2277,N_2214,N_2220);
and U2278 (N_2278,N_2230,N_2235);
or U2279 (N_2279,N_2249,N_2223);
or U2280 (N_2280,N_2203,N_2232);
and U2281 (N_2281,N_2220,N_2238);
or U2282 (N_2282,N_2236,N_2241);
or U2283 (N_2283,N_2225,N_2244);
or U2284 (N_2284,N_2229,N_2213);
and U2285 (N_2285,N_2247,N_2237);
or U2286 (N_2286,N_2230,N_2225);
xor U2287 (N_2287,N_2245,N_2246);
and U2288 (N_2288,N_2215,N_2235);
nand U2289 (N_2289,N_2220,N_2232);
and U2290 (N_2290,N_2228,N_2216);
or U2291 (N_2291,N_2244,N_2221);
nor U2292 (N_2292,N_2211,N_2209);
or U2293 (N_2293,N_2217,N_2211);
nand U2294 (N_2294,N_2217,N_2208);
or U2295 (N_2295,N_2209,N_2237);
nand U2296 (N_2296,N_2236,N_2232);
nand U2297 (N_2297,N_2200,N_2201);
nand U2298 (N_2298,N_2233,N_2240);
nor U2299 (N_2299,N_2226,N_2222);
nand U2300 (N_2300,N_2294,N_2276);
nand U2301 (N_2301,N_2258,N_2273);
nand U2302 (N_2302,N_2254,N_2280);
nand U2303 (N_2303,N_2293,N_2262);
or U2304 (N_2304,N_2297,N_2285);
and U2305 (N_2305,N_2261,N_2286);
and U2306 (N_2306,N_2270,N_2253);
nor U2307 (N_2307,N_2269,N_2274);
nand U2308 (N_2308,N_2296,N_2287);
nand U2309 (N_2309,N_2256,N_2277);
nor U2310 (N_2310,N_2257,N_2279);
or U2311 (N_2311,N_2299,N_2265);
or U2312 (N_2312,N_2292,N_2268);
nand U2313 (N_2313,N_2288,N_2260);
and U2314 (N_2314,N_2263,N_2264);
nor U2315 (N_2315,N_2251,N_2250);
nor U2316 (N_2316,N_2284,N_2272);
or U2317 (N_2317,N_2290,N_2295);
or U2318 (N_2318,N_2271,N_2255);
nand U2319 (N_2319,N_2289,N_2259);
or U2320 (N_2320,N_2282,N_2298);
or U2321 (N_2321,N_2275,N_2291);
or U2322 (N_2322,N_2281,N_2283);
or U2323 (N_2323,N_2278,N_2266);
and U2324 (N_2324,N_2252,N_2267);
or U2325 (N_2325,N_2276,N_2265);
or U2326 (N_2326,N_2294,N_2293);
and U2327 (N_2327,N_2274,N_2296);
or U2328 (N_2328,N_2293,N_2255);
nor U2329 (N_2329,N_2273,N_2278);
or U2330 (N_2330,N_2278,N_2289);
and U2331 (N_2331,N_2280,N_2262);
nand U2332 (N_2332,N_2287,N_2273);
and U2333 (N_2333,N_2277,N_2262);
nand U2334 (N_2334,N_2294,N_2288);
nand U2335 (N_2335,N_2287,N_2261);
nand U2336 (N_2336,N_2278,N_2275);
nor U2337 (N_2337,N_2271,N_2251);
and U2338 (N_2338,N_2252,N_2254);
and U2339 (N_2339,N_2298,N_2297);
nor U2340 (N_2340,N_2277,N_2276);
xnor U2341 (N_2341,N_2287,N_2298);
and U2342 (N_2342,N_2253,N_2293);
nand U2343 (N_2343,N_2263,N_2287);
and U2344 (N_2344,N_2290,N_2297);
nor U2345 (N_2345,N_2262,N_2257);
or U2346 (N_2346,N_2266,N_2262);
nand U2347 (N_2347,N_2266,N_2277);
nand U2348 (N_2348,N_2252,N_2265);
nand U2349 (N_2349,N_2267,N_2276);
nand U2350 (N_2350,N_2334,N_2310);
nor U2351 (N_2351,N_2309,N_2348);
nand U2352 (N_2352,N_2323,N_2301);
or U2353 (N_2353,N_2344,N_2345);
and U2354 (N_2354,N_2336,N_2335);
and U2355 (N_2355,N_2331,N_2326);
or U2356 (N_2356,N_2319,N_2318);
nand U2357 (N_2357,N_2349,N_2340);
nand U2358 (N_2358,N_2316,N_2300);
xnor U2359 (N_2359,N_2322,N_2337);
and U2360 (N_2360,N_2302,N_2315);
and U2361 (N_2361,N_2332,N_2343);
and U2362 (N_2362,N_2324,N_2306);
nand U2363 (N_2363,N_2307,N_2320);
nand U2364 (N_2364,N_2317,N_2304);
and U2365 (N_2365,N_2329,N_2325);
or U2366 (N_2366,N_2311,N_2339);
nand U2367 (N_2367,N_2346,N_2341);
or U2368 (N_2368,N_2321,N_2305);
nand U2369 (N_2369,N_2330,N_2327);
nand U2370 (N_2370,N_2342,N_2333);
nor U2371 (N_2371,N_2303,N_2312);
and U2372 (N_2372,N_2347,N_2338);
and U2373 (N_2373,N_2313,N_2328);
nand U2374 (N_2374,N_2308,N_2314);
nor U2375 (N_2375,N_2347,N_2340);
or U2376 (N_2376,N_2344,N_2321);
nor U2377 (N_2377,N_2313,N_2316);
nor U2378 (N_2378,N_2316,N_2306);
or U2379 (N_2379,N_2305,N_2340);
nor U2380 (N_2380,N_2317,N_2300);
or U2381 (N_2381,N_2317,N_2309);
nor U2382 (N_2382,N_2331,N_2323);
or U2383 (N_2383,N_2342,N_2331);
nor U2384 (N_2384,N_2347,N_2344);
xor U2385 (N_2385,N_2314,N_2348);
or U2386 (N_2386,N_2301,N_2347);
nand U2387 (N_2387,N_2319,N_2312);
nand U2388 (N_2388,N_2327,N_2328);
nor U2389 (N_2389,N_2315,N_2331);
or U2390 (N_2390,N_2302,N_2338);
or U2391 (N_2391,N_2342,N_2301);
or U2392 (N_2392,N_2335,N_2333);
nor U2393 (N_2393,N_2309,N_2305);
or U2394 (N_2394,N_2324,N_2328);
nor U2395 (N_2395,N_2346,N_2304);
nor U2396 (N_2396,N_2323,N_2337);
nand U2397 (N_2397,N_2331,N_2333);
nand U2398 (N_2398,N_2341,N_2300);
nor U2399 (N_2399,N_2340,N_2344);
nor U2400 (N_2400,N_2368,N_2363);
or U2401 (N_2401,N_2360,N_2390);
or U2402 (N_2402,N_2358,N_2379);
and U2403 (N_2403,N_2384,N_2375);
nand U2404 (N_2404,N_2364,N_2382);
or U2405 (N_2405,N_2391,N_2396);
and U2406 (N_2406,N_2393,N_2378);
nor U2407 (N_2407,N_2356,N_2370);
and U2408 (N_2408,N_2374,N_2380);
and U2409 (N_2409,N_2373,N_2365);
and U2410 (N_2410,N_2369,N_2376);
nand U2411 (N_2411,N_2377,N_2351);
nand U2412 (N_2412,N_2367,N_2372);
or U2413 (N_2413,N_2366,N_2350);
or U2414 (N_2414,N_2353,N_2386);
nor U2415 (N_2415,N_2389,N_2383);
or U2416 (N_2416,N_2392,N_2352);
or U2417 (N_2417,N_2397,N_2399);
or U2418 (N_2418,N_2395,N_2385);
and U2419 (N_2419,N_2398,N_2359);
and U2420 (N_2420,N_2357,N_2362);
nor U2421 (N_2421,N_2354,N_2387);
or U2422 (N_2422,N_2371,N_2394);
or U2423 (N_2423,N_2388,N_2381);
nor U2424 (N_2424,N_2355,N_2361);
or U2425 (N_2425,N_2383,N_2381);
and U2426 (N_2426,N_2362,N_2396);
and U2427 (N_2427,N_2350,N_2394);
and U2428 (N_2428,N_2363,N_2364);
nand U2429 (N_2429,N_2394,N_2399);
or U2430 (N_2430,N_2351,N_2376);
and U2431 (N_2431,N_2378,N_2350);
nor U2432 (N_2432,N_2382,N_2383);
nor U2433 (N_2433,N_2389,N_2392);
nor U2434 (N_2434,N_2385,N_2367);
and U2435 (N_2435,N_2361,N_2399);
or U2436 (N_2436,N_2398,N_2376);
nand U2437 (N_2437,N_2358,N_2360);
and U2438 (N_2438,N_2379,N_2394);
and U2439 (N_2439,N_2380,N_2381);
nor U2440 (N_2440,N_2387,N_2373);
nor U2441 (N_2441,N_2372,N_2394);
and U2442 (N_2442,N_2382,N_2353);
or U2443 (N_2443,N_2386,N_2364);
and U2444 (N_2444,N_2384,N_2361);
nor U2445 (N_2445,N_2365,N_2372);
and U2446 (N_2446,N_2387,N_2385);
nand U2447 (N_2447,N_2359,N_2377);
and U2448 (N_2448,N_2370,N_2354);
and U2449 (N_2449,N_2356,N_2386);
and U2450 (N_2450,N_2434,N_2422);
nand U2451 (N_2451,N_2418,N_2426);
and U2452 (N_2452,N_2414,N_2410);
and U2453 (N_2453,N_2448,N_2411);
and U2454 (N_2454,N_2436,N_2442);
or U2455 (N_2455,N_2446,N_2419);
nand U2456 (N_2456,N_2405,N_2424);
and U2457 (N_2457,N_2430,N_2416);
or U2458 (N_2458,N_2433,N_2441);
and U2459 (N_2459,N_2400,N_2404);
or U2460 (N_2460,N_2421,N_2402);
and U2461 (N_2461,N_2432,N_2415);
nand U2462 (N_2462,N_2413,N_2425);
nor U2463 (N_2463,N_2435,N_2444);
nand U2464 (N_2464,N_2412,N_2429);
and U2465 (N_2465,N_2449,N_2417);
and U2466 (N_2466,N_2437,N_2407);
and U2467 (N_2467,N_2447,N_2445);
nor U2468 (N_2468,N_2403,N_2428);
nor U2469 (N_2469,N_2420,N_2423);
nand U2470 (N_2470,N_2440,N_2401);
nand U2471 (N_2471,N_2406,N_2409);
or U2472 (N_2472,N_2439,N_2427);
or U2473 (N_2473,N_2438,N_2431);
nand U2474 (N_2474,N_2443,N_2408);
or U2475 (N_2475,N_2426,N_2416);
nand U2476 (N_2476,N_2405,N_2444);
and U2477 (N_2477,N_2428,N_2410);
nand U2478 (N_2478,N_2418,N_2412);
nor U2479 (N_2479,N_2403,N_2443);
nor U2480 (N_2480,N_2404,N_2413);
nor U2481 (N_2481,N_2404,N_2437);
nand U2482 (N_2482,N_2408,N_2430);
nor U2483 (N_2483,N_2424,N_2439);
nand U2484 (N_2484,N_2400,N_2420);
or U2485 (N_2485,N_2436,N_2422);
nor U2486 (N_2486,N_2423,N_2403);
and U2487 (N_2487,N_2439,N_2437);
or U2488 (N_2488,N_2435,N_2407);
or U2489 (N_2489,N_2444,N_2421);
nor U2490 (N_2490,N_2445,N_2422);
xnor U2491 (N_2491,N_2445,N_2434);
and U2492 (N_2492,N_2418,N_2416);
or U2493 (N_2493,N_2413,N_2408);
nor U2494 (N_2494,N_2412,N_2422);
and U2495 (N_2495,N_2425,N_2442);
and U2496 (N_2496,N_2446,N_2441);
and U2497 (N_2497,N_2400,N_2429);
and U2498 (N_2498,N_2418,N_2441);
nand U2499 (N_2499,N_2439,N_2429);
and U2500 (N_2500,N_2486,N_2491);
and U2501 (N_2501,N_2489,N_2472);
or U2502 (N_2502,N_2494,N_2452);
nor U2503 (N_2503,N_2496,N_2474);
and U2504 (N_2504,N_2460,N_2471);
nand U2505 (N_2505,N_2487,N_2475);
or U2506 (N_2506,N_2451,N_2457);
nor U2507 (N_2507,N_2459,N_2466);
nand U2508 (N_2508,N_2479,N_2495);
nor U2509 (N_2509,N_2464,N_2488);
and U2510 (N_2510,N_2454,N_2483);
nor U2511 (N_2511,N_2480,N_2465);
and U2512 (N_2512,N_2450,N_2462);
or U2513 (N_2513,N_2477,N_2481);
xor U2514 (N_2514,N_2453,N_2476);
nor U2515 (N_2515,N_2498,N_2490);
or U2516 (N_2516,N_2478,N_2468);
and U2517 (N_2517,N_2484,N_2499);
and U2518 (N_2518,N_2456,N_2482);
nand U2519 (N_2519,N_2470,N_2493);
nand U2520 (N_2520,N_2463,N_2461);
nor U2521 (N_2521,N_2485,N_2458);
nor U2522 (N_2522,N_2492,N_2467);
and U2523 (N_2523,N_2473,N_2497);
nand U2524 (N_2524,N_2455,N_2469);
and U2525 (N_2525,N_2459,N_2454);
nor U2526 (N_2526,N_2488,N_2494);
nand U2527 (N_2527,N_2460,N_2489);
and U2528 (N_2528,N_2470,N_2459);
or U2529 (N_2529,N_2468,N_2470);
and U2530 (N_2530,N_2454,N_2451);
or U2531 (N_2531,N_2499,N_2477);
nor U2532 (N_2532,N_2470,N_2453);
or U2533 (N_2533,N_2459,N_2494);
and U2534 (N_2534,N_2486,N_2481);
nand U2535 (N_2535,N_2481,N_2457);
and U2536 (N_2536,N_2471,N_2498);
or U2537 (N_2537,N_2465,N_2473);
or U2538 (N_2538,N_2495,N_2457);
and U2539 (N_2539,N_2451,N_2453);
nor U2540 (N_2540,N_2493,N_2450);
or U2541 (N_2541,N_2473,N_2499);
or U2542 (N_2542,N_2480,N_2477);
xnor U2543 (N_2543,N_2466,N_2489);
and U2544 (N_2544,N_2480,N_2476);
nor U2545 (N_2545,N_2462,N_2486);
nor U2546 (N_2546,N_2455,N_2459);
and U2547 (N_2547,N_2457,N_2489);
nand U2548 (N_2548,N_2496,N_2455);
nor U2549 (N_2549,N_2496,N_2460);
nor U2550 (N_2550,N_2536,N_2542);
and U2551 (N_2551,N_2526,N_2535);
nand U2552 (N_2552,N_2525,N_2522);
nor U2553 (N_2553,N_2543,N_2501);
nor U2554 (N_2554,N_2502,N_2537);
nor U2555 (N_2555,N_2534,N_2509);
and U2556 (N_2556,N_2539,N_2515);
or U2557 (N_2557,N_2506,N_2511);
and U2558 (N_2558,N_2529,N_2544);
nor U2559 (N_2559,N_2507,N_2500);
or U2560 (N_2560,N_2520,N_2533);
nand U2561 (N_2561,N_2514,N_2503);
nor U2562 (N_2562,N_2512,N_2523);
and U2563 (N_2563,N_2546,N_2505);
nand U2564 (N_2564,N_2538,N_2541);
nor U2565 (N_2565,N_2510,N_2519);
nand U2566 (N_2566,N_2528,N_2504);
or U2567 (N_2567,N_2516,N_2508);
nand U2568 (N_2568,N_2547,N_2517);
nor U2569 (N_2569,N_2531,N_2513);
nor U2570 (N_2570,N_2527,N_2545);
and U2571 (N_2571,N_2548,N_2540);
nand U2572 (N_2572,N_2521,N_2518);
nand U2573 (N_2573,N_2532,N_2530);
nor U2574 (N_2574,N_2549,N_2524);
or U2575 (N_2575,N_2530,N_2527);
and U2576 (N_2576,N_2531,N_2527);
and U2577 (N_2577,N_2543,N_2502);
or U2578 (N_2578,N_2533,N_2549);
nor U2579 (N_2579,N_2548,N_2524);
nor U2580 (N_2580,N_2538,N_2528);
and U2581 (N_2581,N_2517,N_2531);
or U2582 (N_2582,N_2512,N_2517);
nand U2583 (N_2583,N_2515,N_2509);
nand U2584 (N_2584,N_2528,N_2533);
nor U2585 (N_2585,N_2513,N_2535);
nor U2586 (N_2586,N_2522,N_2519);
nand U2587 (N_2587,N_2500,N_2543);
or U2588 (N_2588,N_2535,N_2549);
and U2589 (N_2589,N_2510,N_2538);
nor U2590 (N_2590,N_2529,N_2521);
and U2591 (N_2591,N_2525,N_2549);
or U2592 (N_2592,N_2512,N_2535);
nor U2593 (N_2593,N_2515,N_2527);
nor U2594 (N_2594,N_2535,N_2538);
and U2595 (N_2595,N_2513,N_2539);
nand U2596 (N_2596,N_2511,N_2501);
or U2597 (N_2597,N_2512,N_2505);
nor U2598 (N_2598,N_2510,N_2505);
nor U2599 (N_2599,N_2535,N_2515);
nor U2600 (N_2600,N_2586,N_2561);
and U2601 (N_2601,N_2576,N_2593);
nand U2602 (N_2602,N_2557,N_2569);
nand U2603 (N_2603,N_2556,N_2558);
or U2604 (N_2604,N_2599,N_2587);
nand U2605 (N_2605,N_2598,N_2595);
or U2606 (N_2606,N_2563,N_2578);
nor U2607 (N_2607,N_2566,N_2567);
and U2608 (N_2608,N_2584,N_2580);
and U2609 (N_2609,N_2551,N_2594);
nand U2610 (N_2610,N_2574,N_2553);
nand U2611 (N_2611,N_2582,N_2577);
nand U2612 (N_2612,N_2589,N_2562);
nor U2613 (N_2613,N_2554,N_2575);
nand U2614 (N_2614,N_2560,N_2570);
or U2615 (N_2615,N_2583,N_2581);
nand U2616 (N_2616,N_2596,N_2550);
nor U2617 (N_2617,N_2573,N_2579);
and U2618 (N_2618,N_2592,N_2588);
nor U2619 (N_2619,N_2564,N_2571);
and U2620 (N_2620,N_2591,N_2555);
nand U2621 (N_2621,N_2568,N_2552);
or U2622 (N_2622,N_2597,N_2572);
or U2623 (N_2623,N_2590,N_2559);
and U2624 (N_2624,N_2585,N_2565);
nor U2625 (N_2625,N_2597,N_2588);
nand U2626 (N_2626,N_2559,N_2597);
or U2627 (N_2627,N_2558,N_2581);
and U2628 (N_2628,N_2572,N_2599);
or U2629 (N_2629,N_2576,N_2556);
nor U2630 (N_2630,N_2560,N_2580);
and U2631 (N_2631,N_2580,N_2573);
or U2632 (N_2632,N_2586,N_2580);
and U2633 (N_2633,N_2574,N_2586);
nand U2634 (N_2634,N_2554,N_2588);
nor U2635 (N_2635,N_2589,N_2554);
nor U2636 (N_2636,N_2576,N_2597);
or U2637 (N_2637,N_2566,N_2585);
nor U2638 (N_2638,N_2574,N_2583);
nand U2639 (N_2639,N_2587,N_2558);
nor U2640 (N_2640,N_2577,N_2570);
nor U2641 (N_2641,N_2591,N_2592);
or U2642 (N_2642,N_2557,N_2597);
nand U2643 (N_2643,N_2553,N_2566);
or U2644 (N_2644,N_2587,N_2580);
or U2645 (N_2645,N_2562,N_2565);
nor U2646 (N_2646,N_2590,N_2595);
nor U2647 (N_2647,N_2598,N_2575);
nand U2648 (N_2648,N_2583,N_2585);
nor U2649 (N_2649,N_2592,N_2578);
or U2650 (N_2650,N_2610,N_2615);
or U2651 (N_2651,N_2634,N_2631);
or U2652 (N_2652,N_2648,N_2637);
or U2653 (N_2653,N_2638,N_2625);
xnor U2654 (N_2654,N_2624,N_2649);
nand U2655 (N_2655,N_2605,N_2600);
or U2656 (N_2656,N_2633,N_2627);
and U2657 (N_2657,N_2611,N_2612);
nor U2658 (N_2658,N_2601,N_2606);
or U2659 (N_2659,N_2602,N_2642);
and U2660 (N_2660,N_2622,N_2623);
nor U2661 (N_2661,N_2628,N_2620);
nand U2662 (N_2662,N_2603,N_2609);
nand U2663 (N_2663,N_2613,N_2604);
nor U2664 (N_2664,N_2632,N_2626);
nand U2665 (N_2665,N_2614,N_2619);
nand U2666 (N_2666,N_2617,N_2630);
nand U2667 (N_2667,N_2647,N_2616);
and U2668 (N_2668,N_2646,N_2645);
nor U2669 (N_2669,N_2608,N_2643);
and U2670 (N_2670,N_2607,N_2618);
or U2671 (N_2671,N_2635,N_2641);
or U2672 (N_2672,N_2629,N_2639);
and U2673 (N_2673,N_2644,N_2640);
or U2674 (N_2674,N_2621,N_2636);
or U2675 (N_2675,N_2602,N_2604);
nand U2676 (N_2676,N_2640,N_2630);
nor U2677 (N_2677,N_2631,N_2629);
or U2678 (N_2678,N_2602,N_2647);
nor U2679 (N_2679,N_2612,N_2621);
nand U2680 (N_2680,N_2645,N_2633);
nand U2681 (N_2681,N_2635,N_2602);
and U2682 (N_2682,N_2637,N_2624);
nand U2683 (N_2683,N_2629,N_2610);
nand U2684 (N_2684,N_2638,N_2627);
nor U2685 (N_2685,N_2632,N_2644);
or U2686 (N_2686,N_2609,N_2634);
nand U2687 (N_2687,N_2612,N_2600);
or U2688 (N_2688,N_2604,N_2619);
and U2689 (N_2689,N_2631,N_2624);
or U2690 (N_2690,N_2632,N_2640);
and U2691 (N_2691,N_2626,N_2622);
nor U2692 (N_2692,N_2626,N_2604);
nor U2693 (N_2693,N_2647,N_2610);
or U2694 (N_2694,N_2628,N_2601);
nand U2695 (N_2695,N_2612,N_2632);
or U2696 (N_2696,N_2633,N_2613);
nor U2697 (N_2697,N_2624,N_2648);
nor U2698 (N_2698,N_2606,N_2614);
nor U2699 (N_2699,N_2635,N_2626);
and U2700 (N_2700,N_2665,N_2697);
or U2701 (N_2701,N_2683,N_2684);
nand U2702 (N_2702,N_2693,N_2676);
and U2703 (N_2703,N_2671,N_2677);
nand U2704 (N_2704,N_2696,N_2692);
nand U2705 (N_2705,N_2655,N_2666);
or U2706 (N_2706,N_2673,N_2653);
or U2707 (N_2707,N_2654,N_2651);
nand U2708 (N_2708,N_2662,N_2667);
nand U2709 (N_2709,N_2687,N_2698);
and U2710 (N_2710,N_2663,N_2672);
or U2711 (N_2711,N_2674,N_2670);
and U2712 (N_2712,N_2695,N_2668);
nand U2713 (N_2713,N_2652,N_2690);
and U2714 (N_2714,N_2682,N_2661);
nor U2715 (N_2715,N_2650,N_2688);
nor U2716 (N_2716,N_2685,N_2664);
and U2717 (N_2717,N_2669,N_2659);
or U2718 (N_2718,N_2699,N_2660);
or U2719 (N_2719,N_2658,N_2679);
nor U2720 (N_2720,N_2691,N_2656);
nand U2721 (N_2721,N_2681,N_2657);
nor U2722 (N_2722,N_2675,N_2680);
or U2723 (N_2723,N_2689,N_2694);
nor U2724 (N_2724,N_2678,N_2686);
or U2725 (N_2725,N_2670,N_2698);
xor U2726 (N_2726,N_2682,N_2665);
nor U2727 (N_2727,N_2666,N_2695);
nand U2728 (N_2728,N_2697,N_2660);
and U2729 (N_2729,N_2668,N_2670);
nand U2730 (N_2730,N_2693,N_2653);
and U2731 (N_2731,N_2652,N_2650);
or U2732 (N_2732,N_2686,N_2665);
nand U2733 (N_2733,N_2680,N_2667);
or U2734 (N_2734,N_2663,N_2699);
nor U2735 (N_2735,N_2686,N_2680);
nand U2736 (N_2736,N_2652,N_2676);
nor U2737 (N_2737,N_2662,N_2669);
nand U2738 (N_2738,N_2678,N_2667);
nand U2739 (N_2739,N_2653,N_2666);
or U2740 (N_2740,N_2697,N_2676);
nand U2741 (N_2741,N_2668,N_2677);
and U2742 (N_2742,N_2676,N_2678);
or U2743 (N_2743,N_2655,N_2658);
nor U2744 (N_2744,N_2661,N_2694);
nor U2745 (N_2745,N_2690,N_2656);
nor U2746 (N_2746,N_2676,N_2692);
or U2747 (N_2747,N_2694,N_2662);
nor U2748 (N_2748,N_2661,N_2688);
nor U2749 (N_2749,N_2657,N_2683);
nand U2750 (N_2750,N_2744,N_2745);
and U2751 (N_2751,N_2743,N_2703);
or U2752 (N_2752,N_2721,N_2737);
nand U2753 (N_2753,N_2718,N_2729);
or U2754 (N_2754,N_2706,N_2701);
and U2755 (N_2755,N_2702,N_2728);
nor U2756 (N_2756,N_2735,N_2716);
or U2757 (N_2757,N_2730,N_2727);
nor U2758 (N_2758,N_2738,N_2715);
and U2759 (N_2759,N_2746,N_2719);
nand U2760 (N_2760,N_2710,N_2714);
nand U2761 (N_2761,N_2749,N_2740);
or U2762 (N_2762,N_2732,N_2720);
nor U2763 (N_2763,N_2700,N_2708);
nor U2764 (N_2764,N_2711,N_2705);
nor U2765 (N_2765,N_2739,N_2742);
or U2766 (N_2766,N_2722,N_2712);
and U2767 (N_2767,N_2733,N_2713);
and U2768 (N_2768,N_2747,N_2726);
or U2769 (N_2769,N_2704,N_2717);
nand U2770 (N_2770,N_2748,N_2707);
and U2771 (N_2771,N_2709,N_2741);
nand U2772 (N_2772,N_2724,N_2725);
or U2773 (N_2773,N_2736,N_2731);
xor U2774 (N_2774,N_2734,N_2723);
and U2775 (N_2775,N_2741,N_2720);
and U2776 (N_2776,N_2736,N_2733);
or U2777 (N_2777,N_2746,N_2748);
and U2778 (N_2778,N_2708,N_2720);
nand U2779 (N_2779,N_2739,N_2730);
or U2780 (N_2780,N_2748,N_2725);
or U2781 (N_2781,N_2725,N_2735);
nor U2782 (N_2782,N_2747,N_2742);
and U2783 (N_2783,N_2724,N_2740);
and U2784 (N_2784,N_2711,N_2700);
or U2785 (N_2785,N_2731,N_2729);
and U2786 (N_2786,N_2707,N_2725);
nor U2787 (N_2787,N_2734,N_2703);
and U2788 (N_2788,N_2711,N_2732);
and U2789 (N_2789,N_2731,N_2705);
and U2790 (N_2790,N_2745,N_2728);
nand U2791 (N_2791,N_2739,N_2714);
nand U2792 (N_2792,N_2718,N_2707);
nor U2793 (N_2793,N_2703,N_2712);
xor U2794 (N_2794,N_2707,N_2712);
and U2795 (N_2795,N_2749,N_2722);
and U2796 (N_2796,N_2702,N_2722);
and U2797 (N_2797,N_2749,N_2700);
and U2798 (N_2798,N_2711,N_2708);
nand U2799 (N_2799,N_2732,N_2746);
nand U2800 (N_2800,N_2763,N_2755);
or U2801 (N_2801,N_2779,N_2759);
and U2802 (N_2802,N_2798,N_2781);
or U2803 (N_2803,N_2782,N_2769);
nand U2804 (N_2804,N_2786,N_2762);
nor U2805 (N_2805,N_2751,N_2777);
nor U2806 (N_2806,N_2785,N_2752);
nand U2807 (N_2807,N_2760,N_2773);
or U2808 (N_2808,N_2758,N_2795);
and U2809 (N_2809,N_2776,N_2799);
or U2810 (N_2810,N_2793,N_2797);
nor U2811 (N_2811,N_2767,N_2753);
xnor U2812 (N_2812,N_2764,N_2750);
or U2813 (N_2813,N_2757,N_2771);
nand U2814 (N_2814,N_2784,N_2770);
nor U2815 (N_2815,N_2765,N_2761);
nor U2816 (N_2816,N_2794,N_2792);
nand U2817 (N_2817,N_2754,N_2788);
nand U2818 (N_2818,N_2775,N_2768);
xor U2819 (N_2819,N_2790,N_2756);
and U2820 (N_2820,N_2783,N_2789);
nor U2821 (N_2821,N_2780,N_2774);
or U2822 (N_2822,N_2787,N_2772);
nor U2823 (N_2823,N_2796,N_2791);
nor U2824 (N_2824,N_2778,N_2766);
or U2825 (N_2825,N_2781,N_2797);
nand U2826 (N_2826,N_2786,N_2781);
or U2827 (N_2827,N_2799,N_2780);
nor U2828 (N_2828,N_2752,N_2754);
nand U2829 (N_2829,N_2775,N_2778);
nor U2830 (N_2830,N_2797,N_2782);
and U2831 (N_2831,N_2797,N_2787);
and U2832 (N_2832,N_2780,N_2766);
nor U2833 (N_2833,N_2782,N_2793);
or U2834 (N_2834,N_2785,N_2774);
nor U2835 (N_2835,N_2797,N_2767);
xnor U2836 (N_2836,N_2788,N_2756);
or U2837 (N_2837,N_2765,N_2799);
nor U2838 (N_2838,N_2784,N_2769);
and U2839 (N_2839,N_2767,N_2769);
and U2840 (N_2840,N_2769,N_2788);
nand U2841 (N_2841,N_2797,N_2770);
nor U2842 (N_2842,N_2757,N_2786);
nand U2843 (N_2843,N_2784,N_2758);
and U2844 (N_2844,N_2785,N_2764);
nand U2845 (N_2845,N_2773,N_2767);
and U2846 (N_2846,N_2771,N_2773);
or U2847 (N_2847,N_2796,N_2754);
nor U2848 (N_2848,N_2782,N_2770);
and U2849 (N_2849,N_2790,N_2793);
nand U2850 (N_2850,N_2843,N_2822);
and U2851 (N_2851,N_2839,N_2806);
nand U2852 (N_2852,N_2802,N_2841);
nor U2853 (N_2853,N_2819,N_2845);
nand U2854 (N_2854,N_2834,N_2830);
nand U2855 (N_2855,N_2844,N_2848);
nor U2856 (N_2856,N_2832,N_2829);
or U2857 (N_2857,N_2814,N_2820);
nor U2858 (N_2858,N_2831,N_2800);
and U2859 (N_2859,N_2810,N_2833);
nor U2860 (N_2860,N_2824,N_2808);
nand U2861 (N_2861,N_2838,N_2821);
nand U2862 (N_2862,N_2840,N_2837);
or U2863 (N_2863,N_2828,N_2818);
nor U2864 (N_2864,N_2807,N_2836);
and U2865 (N_2865,N_2826,N_2809);
or U2866 (N_2866,N_2805,N_2811);
or U2867 (N_2867,N_2847,N_2801);
or U2868 (N_2868,N_2823,N_2816);
nand U2869 (N_2869,N_2812,N_2825);
or U2870 (N_2870,N_2835,N_2803);
nand U2871 (N_2871,N_2842,N_2846);
xnor U2872 (N_2872,N_2849,N_2804);
nor U2873 (N_2873,N_2817,N_2827);
nand U2874 (N_2874,N_2813,N_2815);
and U2875 (N_2875,N_2816,N_2827);
and U2876 (N_2876,N_2835,N_2840);
and U2877 (N_2877,N_2820,N_2804);
nand U2878 (N_2878,N_2833,N_2805);
nand U2879 (N_2879,N_2816,N_2802);
or U2880 (N_2880,N_2848,N_2847);
nand U2881 (N_2881,N_2841,N_2833);
or U2882 (N_2882,N_2806,N_2821);
or U2883 (N_2883,N_2814,N_2831);
and U2884 (N_2884,N_2804,N_2814);
and U2885 (N_2885,N_2848,N_2830);
and U2886 (N_2886,N_2831,N_2809);
or U2887 (N_2887,N_2801,N_2805);
and U2888 (N_2888,N_2830,N_2842);
nor U2889 (N_2889,N_2818,N_2837);
or U2890 (N_2890,N_2809,N_2806);
nor U2891 (N_2891,N_2831,N_2845);
nand U2892 (N_2892,N_2818,N_2826);
or U2893 (N_2893,N_2841,N_2827);
and U2894 (N_2894,N_2839,N_2808);
nor U2895 (N_2895,N_2839,N_2840);
and U2896 (N_2896,N_2812,N_2831);
or U2897 (N_2897,N_2837,N_2838);
and U2898 (N_2898,N_2838,N_2832);
and U2899 (N_2899,N_2814,N_2848);
nand U2900 (N_2900,N_2869,N_2855);
xnor U2901 (N_2901,N_2872,N_2866);
nor U2902 (N_2902,N_2876,N_2882);
and U2903 (N_2903,N_2892,N_2887);
nand U2904 (N_2904,N_2868,N_2894);
or U2905 (N_2905,N_2858,N_2874);
nand U2906 (N_2906,N_2877,N_2881);
nor U2907 (N_2907,N_2857,N_2896);
or U2908 (N_2908,N_2862,N_2898);
nor U2909 (N_2909,N_2861,N_2854);
and U2910 (N_2910,N_2867,N_2873);
nand U2911 (N_2911,N_2852,N_2895);
and U2912 (N_2912,N_2893,N_2883);
nor U2913 (N_2913,N_2879,N_2853);
or U2914 (N_2914,N_2897,N_2880);
and U2915 (N_2915,N_2870,N_2860);
and U2916 (N_2916,N_2871,N_2864);
and U2917 (N_2917,N_2885,N_2859);
nand U2918 (N_2918,N_2888,N_2890);
nand U2919 (N_2919,N_2863,N_2850);
or U2920 (N_2920,N_2889,N_2891);
or U2921 (N_2921,N_2875,N_2899);
and U2922 (N_2922,N_2878,N_2865);
or U2923 (N_2923,N_2851,N_2886);
nor U2924 (N_2924,N_2884,N_2856);
xor U2925 (N_2925,N_2870,N_2895);
nand U2926 (N_2926,N_2868,N_2879);
nor U2927 (N_2927,N_2868,N_2859);
and U2928 (N_2928,N_2858,N_2889);
and U2929 (N_2929,N_2874,N_2863);
or U2930 (N_2930,N_2875,N_2893);
nor U2931 (N_2931,N_2866,N_2852);
and U2932 (N_2932,N_2869,N_2856);
and U2933 (N_2933,N_2867,N_2878);
nor U2934 (N_2934,N_2851,N_2895);
nand U2935 (N_2935,N_2851,N_2883);
or U2936 (N_2936,N_2884,N_2887);
nor U2937 (N_2937,N_2851,N_2891);
or U2938 (N_2938,N_2888,N_2897);
nor U2939 (N_2939,N_2870,N_2852);
xor U2940 (N_2940,N_2894,N_2859);
or U2941 (N_2941,N_2862,N_2897);
or U2942 (N_2942,N_2889,N_2899);
nor U2943 (N_2943,N_2868,N_2871);
and U2944 (N_2944,N_2889,N_2879);
or U2945 (N_2945,N_2878,N_2896);
and U2946 (N_2946,N_2884,N_2897);
and U2947 (N_2947,N_2860,N_2865);
nor U2948 (N_2948,N_2861,N_2862);
and U2949 (N_2949,N_2898,N_2896);
or U2950 (N_2950,N_2911,N_2925);
nor U2951 (N_2951,N_2908,N_2935);
or U2952 (N_2952,N_2945,N_2914);
xnor U2953 (N_2953,N_2900,N_2946);
nor U2954 (N_2954,N_2903,N_2902);
nor U2955 (N_2955,N_2931,N_2912);
or U2956 (N_2956,N_2927,N_2943);
nor U2957 (N_2957,N_2909,N_2907);
and U2958 (N_2958,N_2923,N_2933);
or U2959 (N_2959,N_2916,N_2939);
nor U2960 (N_2960,N_2928,N_2940);
and U2961 (N_2961,N_2901,N_2913);
nor U2962 (N_2962,N_2922,N_2937);
nor U2963 (N_2963,N_2944,N_2906);
nand U2964 (N_2964,N_2942,N_2949);
nor U2965 (N_2965,N_2919,N_2947);
nor U2966 (N_2966,N_2926,N_2905);
nor U2967 (N_2967,N_2936,N_2910);
and U2968 (N_2968,N_2904,N_2921);
or U2969 (N_2969,N_2941,N_2924);
nand U2970 (N_2970,N_2934,N_2920);
nand U2971 (N_2971,N_2929,N_2938);
nor U2972 (N_2972,N_2917,N_2918);
and U2973 (N_2973,N_2948,N_2915);
nand U2974 (N_2974,N_2932,N_2930);
and U2975 (N_2975,N_2926,N_2925);
or U2976 (N_2976,N_2944,N_2938);
and U2977 (N_2977,N_2940,N_2905);
nor U2978 (N_2978,N_2930,N_2924);
nand U2979 (N_2979,N_2942,N_2946);
and U2980 (N_2980,N_2947,N_2949);
nand U2981 (N_2981,N_2931,N_2903);
and U2982 (N_2982,N_2942,N_2941);
and U2983 (N_2983,N_2906,N_2914);
nand U2984 (N_2984,N_2949,N_2928);
nor U2985 (N_2985,N_2900,N_2904);
nand U2986 (N_2986,N_2926,N_2936);
nor U2987 (N_2987,N_2933,N_2931);
nor U2988 (N_2988,N_2911,N_2939);
or U2989 (N_2989,N_2900,N_2949);
or U2990 (N_2990,N_2937,N_2939);
or U2991 (N_2991,N_2929,N_2926);
and U2992 (N_2992,N_2942,N_2938);
or U2993 (N_2993,N_2907,N_2912);
or U2994 (N_2994,N_2946,N_2914);
xor U2995 (N_2995,N_2909,N_2930);
and U2996 (N_2996,N_2921,N_2915);
nor U2997 (N_2997,N_2903,N_2910);
and U2998 (N_2998,N_2911,N_2913);
xnor U2999 (N_2999,N_2943,N_2909);
nand UO_0 (O_0,N_2994,N_2985);
nand UO_1 (O_1,N_2965,N_2968);
or UO_2 (O_2,N_2961,N_2960);
nand UO_3 (O_3,N_2975,N_2987);
nand UO_4 (O_4,N_2998,N_2980);
or UO_5 (O_5,N_2972,N_2969);
nand UO_6 (O_6,N_2981,N_2966);
or UO_7 (O_7,N_2958,N_2974);
and UO_8 (O_8,N_2992,N_2962);
xor UO_9 (O_9,N_2952,N_2983);
or UO_10 (O_10,N_2988,N_2954);
nor UO_11 (O_11,N_2991,N_2976);
nor UO_12 (O_12,N_2999,N_2964);
nor UO_13 (O_13,N_2996,N_2979);
nor UO_14 (O_14,N_2957,N_2973);
and UO_15 (O_15,N_2995,N_2953);
and UO_16 (O_16,N_2990,N_2951);
nand UO_17 (O_17,N_2950,N_2982);
nor UO_18 (O_18,N_2959,N_2993);
or UO_19 (O_19,N_2986,N_2978);
nand UO_20 (O_20,N_2967,N_2970);
and UO_21 (O_21,N_2955,N_2997);
nand UO_22 (O_22,N_2984,N_2977);
nand UO_23 (O_23,N_2956,N_2963);
nor UO_24 (O_24,N_2989,N_2971);
nor UO_25 (O_25,N_2966,N_2978);
nor UO_26 (O_26,N_2975,N_2979);
or UO_27 (O_27,N_2977,N_2995);
nand UO_28 (O_28,N_2990,N_2966);
nand UO_29 (O_29,N_2951,N_2950);
nand UO_30 (O_30,N_2951,N_2976);
nand UO_31 (O_31,N_2966,N_2974);
nor UO_32 (O_32,N_2950,N_2998);
xor UO_33 (O_33,N_2961,N_2954);
nand UO_34 (O_34,N_2973,N_2986);
or UO_35 (O_35,N_2995,N_2982);
or UO_36 (O_36,N_2975,N_2950);
xor UO_37 (O_37,N_2954,N_2991);
or UO_38 (O_38,N_2979,N_2953);
and UO_39 (O_39,N_2959,N_2953);
nor UO_40 (O_40,N_2988,N_2997);
nand UO_41 (O_41,N_2957,N_2958);
nor UO_42 (O_42,N_2994,N_2970);
nand UO_43 (O_43,N_2969,N_2981);
or UO_44 (O_44,N_2952,N_2980);
nor UO_45 (O_45,N_2963,N_2995);
and UO_46 (O_46,N_2951,N_2992);
nor UO_47 (O_47,N_2953,N_2974);
and UO_48 (O_48,N_2973,N_2991);
nand UO_49 (O_49,N_2970,N_2955);
nor UO_50 (O_50,N_2976,N_2974);
nand UO_51 (O_51,N_2956,N_2970);
or UO_52 (O_52,N_2995,N_2998);
or UO_53 (O_53,N_2993,N_2953);
nand UO_54 (O_54,N_2979,N_2997);
or UO_55 (O_55,N_2964,N_2972);
or UO_56 (O_56,N_2999,N_2956);
and UO_57 (O_57,N_2996,N_2998);
xnor UO_58 (O_58,N_2988,N_2960);
and UO_59 (O_59,N_2964,N_2995);
xor UO_60 (O_60,N_2994,N_2953);
nor UO_61 (O_61,N_2994,N_2964);
nand UO_62 (O_62,N_2951,N_2978);
and UO_63 (O_63,N_2992,N_2982);
or UO_64 (O_64,N_2952,N_2964);
nor UO_65 (O_65,N_2974,N_2982);
nor UO_66 (O_66,N_2975,N_2997);
and UO_67 (O_67,N_2989,N_2952);
nand UO_68 (O_68,N_2958,N_2963);
or UO_69 (O_69,N_2956,N_2985);
or UO_70 (O_70,N_2967,N_2950);
and UO_71 (O_71,N_2968,N_2985);
and UO_72 (O_72,N_2959,N_2996);
nand UO_73 (O_73,N_2954,N_2972);
nand UO_74 (O_74,N_2981,N_2975);
and UO_75 (O_75,N_2974,N_2973);
nor UO_76 (O_76,N_2956,N_2984);
or UO_77 (O_77,N_2957,N_2972);
and UO_78 (O_78,N_2952,N_2999);
nor UO_79 (O_79,N_2979,N_2984);
nor UO_80 (O_80,N_2977,N_2983);
or UO_81 (O_81,N_2959,N_2991);
nor UO_82 (O_82,N_2984,N_2997);
and UO_83 (O_83,N_2964,N_2950);
nand UO_84 (O_84,N_2990,N_2965);
and UO_85 (O_85,N_2963,N_2967);
nand UO_86 (O_86,N_2996,N_2989);
nand UO_87 (O_87,N_2963,N_2977);
nand UO_88 (O_88,N_2981,N_2996);
or UO_89 (O_89,N_2964,N_2993);
nor UO_90 (O_90,N_2956,N_2965);
nand UO_91 (O_91,N_2996,N_2994);
or UO_92 (O_92,N_2992,N_2998);
and UO_93 (O_93,N_2960,N_2982);
nand UO_94 (O_94,N_2974,N_2990);
and UO_95 (O_95,N_2955,N_2986);
nor UO_96 (O_96,N_2953,N_2975);
or UO_97 (O_97,N_2971,N_2972);
nand UO_98 (O_98,N_2967,N_2973);
and UO_99 (O_99,N_2983,N_2981);
and UO_100 (O_100,N_2991,N_2978);
or UO_101 (O_101,N_2976,N_2973);
and UO_102 (O_102,N_2953,N_2969);
and UO_103 (O_103,N_2951,N_2975);
nand UO_104 (O_104,N_2959,N_2967);
nand UO_105 (O_105,N_2990,N_2995);
and UO_106 (O_106,N_2976,N_2993);
or UO_107 (O_107,N_2982,N_2953);
nand UO_108 (O_108,N_2987,N_2963);
and UO_109 (O_109,N_2984,N_2988);
nand UO_110 (O_110,N_2997,N_2954);
nand UO_111 (O_111,N_2972,N_2965);
nor UO_112 (O_112,N_2982,N_2967);
or UO_113 (O_113,N_2990,N_2994);
or UO_114 (O_114,N_2978,N_2984);
nor UO_115 (O_115,N_2989,N_2997);
nor UO_116 (O_116,N_2961,N_2950);
and UO_117 (O_117,N_2972,N_2993);
nand UO_118 (O_118,N_2976,N_2961);
and UO_119 (O_119,N_2975,N_2969);
nor UO_120 (O_120,N_2969,N_2952);
nor UO_121 (O_121,N_2950,N_2989);
and UO_122 (O_122,N_2995,N_2997);
nor UO_123 (O_123,N_2964,N_2958);
nand UO_124 (O_124,N_2988,N_2950);
or UO_125 (O_125,N_2970,N_2990);
or UO_126 (O_126,N_2952,N_2961);
or UO_127 (O_127,N_2997,N_2961);
and UO_128 (O_128,N_2981,N_2980);
nor UO_129 (O_129,N_2971,N_2994);
nor UO_130 (O_130,N_2973,N_2965);
and UO_131 (O_131,N_2982,N_2969);
or UO_132 (O_132,N_2955,N_2980);
nor UO_133 (O_133,N_2983,N_2984);
nor UO_134 (O_134,N_2970,N_2972);
nor UO_135 (O_135,N_2991,N_2993);
nor UO_136 (O_136,N_2975,N_2966);
nand UO_137 (O_137,N_2953,N_2966);
nand UO_138 (O_138,N_2992,N_2960);
nor UO_139 (O_139,N_2976,N_2980);
nand UO_140 (O_140,N_2950,N_2993);
or UO_141 (O_141,N_2960,N_2968);
or UO_142 (O_142,N_2975,N_2961);
and UO_143 (O_143,N_2962,N_2994);
and UO_144 (O_144,N_2975,N_2954);
nand UO_145 (O_145,N_2957,N_2994);
xor UO_146 (O_146,N_2957,N_2996);
or UO_147 (O_147,N_2954,N_2971);
nand UO_148 (O_148,N_2971,N_2957);
nor UO_149 (O_149,N_2972,N_2963);
nand UO_150 (O_150,N_2996,N_2999);
or UO_151 (O_151,N_2972,N_2976);
nand UO_152 (O_152,N_2960,N_2999);
nor UO_153 (O_153,N_2972,N_2979);
and UO_154 (O_154,N_2971,N_2960);
or UO_155 (O_155,N_2981,N_2985);
nor UO_156 (O_156,N_2977,N_2979);
nor UO_157 (O_157,N_2954,N_2994);
and UO_158 (O_158,N_2965,N_2967);
nand UO_159 (O_159,N_2955,N_2983);
nand UO_160 (O_160,N_2965,N_2989);
or UO_161 (O_161,N_2968,N_2998);
nand UO_162 (O_162,N_2954,N_2987);
nand UO_163 (O_163,N_2988,N_2964);
and UO_164 (O_164,N_2996,N_2978);
nand UO_165 (O_165,N_2998,N_2956);
nor UO_166 (O_166,N_2965,N_2992);
nand UO_167 (O_167,N_2997,N_2962);
nor UO_168 (O_168,N_2979,N_2955);
nand UO_169 (O_169,N_2996,N_2952);
or UO_170 (O_170,N_2973,N_2953);
nand UO_171 (O_171,N_2951,N_2957);
and UO_172 (O_172,N_2969,N_2996);
and UO_173 (O_173,N_2957,N_2977);
nand UO_174 (O_174,N_2960,N_2956);
nor UO_175 (O_175,N_2982,N_2991);
nand UO_176 (O_176,N_2987,N_2996);
and UO_177 (O_177,N_2996,N_2997);
and UO_178 (O_178,N_2991,N_2994);
nand UO_179 (O_179,N_2964,N_2985);
nand UO_180 (O_180,N_2960,N_2972);
nor UO_181 (O_181,N_2988,N_2956);
or UO_182 (O_182,N_2989,N_2992);
nand UO_183 (O_183,N_2951,N_2961);
nand UO_184 (O_184,N_2954,N_2951);
and UO_185 (O_185,N_2967,N_2958);
or UO_186 (O_186,N_2990,N_2999);
and UO_187 (O_187,N_2954,N_2964);
and UO_188 (O_188,N_2984,N_2996);
and UO_189 (O_189,N_2958,N_2978);
and UO_190 (O_190,N_2964,N_2990);
nand UO_191 (O_191,N_2999,N_2984);
nor UO_192 (O_192,N_2963,N_2979);
nor UO_193 (O_193,N_2965,N_2950);
or UO_194 (O_194,N_2962,N_2990);
and UO_195 (O_195,N_2991,N_2984);
and UO_196 (O_196,N_2965,N_2979);
or UO_197 (O_197,N_2974,N_2960);
nor UO_198 (O_198,N_2984,N_2970);
or UO_199 (O_199,N_2987,N_2972);
nand UO_200 (O_200,N_2967,N_2955);
nor UO_201 (O_201,N_2973,N_2997);
nor UO_202 (O_202,N_2979,N_2957);
nand UO_203 (O_203,N_2955,N_2978);
or UO_204 (O_204,N_2986,N_2961);
and UO_205 (O_205,N_2966,N_2951);
or UO_206 (O_206,N_2960,N_2967);
and UO_207 (O_207,N_2995,N_2975);
nand UO_208 (O_208,N_2987,N_2997);
and UO_209 (O_209,N_2965,N_2951);
nand UO_210 (O_210,N_2985,N_2970);
nand UO_211 (O_211,N_2974,N_2970);
or UO_212 (O_212,N_2963,N_2973);
or UO_213 (O_213,N_2952,N_2978);
and UO_214 (O_214,N_2965,N_2971);
nor UO_215 (O_215,N_2985,N_2965);
and UO_216 (O_216,N_2972,N_2952);
and UO_217 (O_217,N_2976,N_2959);
or UO_218 (O_218,N_2962,N_2973);
nand UO_219 (O_219,N_2988,N_2971);
nand UO_220 (O_220,N_2992,N_2967);
and UO_221 (O_221,N_2951,N_2952);
nor UO_222 (O_222,N_2978,N_2957);
nor UO_223 (O_223,N_2973,N_2982);
and UO_224 (O_224,N_2974,N_2956);
and UO_225 (O_225,N_2969,N_2971);
or UO_226 (O_226,N_2991,N_2980);
and UO_227 (O_227,N_2952,N_2990);
nor UO_228 (O_228,N_2986,N_2962);
and UO_229 (O_229,N_2994,N_2986);
and UO_230 (O_230,N_2991,N_2967);
or UO_231 (O_231,N_2982,N_2976);
and UO_232 (O_232,N_2987,N_2958);
and UO_233 (O_233,N_2994,N_2975);
nor UO_234 (O_234,N_2977,N_2999);
nor UO_235 (O_235,N_2963,N_2968);
nand UO_236 (O_236,N_2979,N_2981);
nand UO_237 (O_237,N_2995,N_2978);
and UO_238 (O_238,N_2981,N_2964);
or UO_239 (O_239,N_2963,N_2991);
nand UO_240 (O_240,N_2992,N_2961);
nand UO_241 (O_241,N_2990,N_2992);
nor UO_242 (O_242,N_2983,N_2968);
or UO_243 (O_243,N_2993,N_2998);
and UO_244 (O_244,N_2986,N_2977);
and UO_245 (O_245,N_2960,N_2964);
nand UO_246 (O_246,N_2984,N_2992);
nand UO_247 (O_247,N_2967,N_2972);
and UO_248 (O_248,N_2971,N_2996);
nor UO_249 (O_249,N_2971,N_2981);
and UO_250 (O_250,N_2980,N_2983);
and UO_251 (O_251,N_2977,N_2994);
or UO_252 (O_252,N_2953,N_2985);
xnor UO_253 (O_253,N_2958,N_2993);
nor UO_254 (O_254,N_2997,N_2968);
or UO_255 (O_255,N_2965,N_2978);
and UO_256 (O_256,N_2953,N_2950);
and UO_257 (O_257,N_2955,N_2992);
or UO_258 (O_258,N_2992,N_2978);
or UO_259 (O_259,N_2977,N_2980);
nor UO_260 (O_260,N_2959,N_2987);
nand UO_261 (O_261,N_2960,N_2993);
nor UO_262 (O_262,N_2954,N_2973);
and UO_263 (O_263,N_2993,N_2992);
nor UO_264 (O_264,N_2959,N_2986);
or UO_265 (O_265,N_2974,N_2989);
nand UO_266 (O_266,N_2994,N_2967);
nand UO_267 (O_267,N_2990,N_2988);
nor UO_268 (O_268,N_2999,N_2991);
nand UO_269 (O_269,N_2973,N_2975);
nor UO_270 (O_270,N_2958,N_2997);
xor UO_271 (O_271,N_2987,N_2964);
or UO_272 (O_272,N_2977,N_2955);
nand UO_273 (O_273,N_2991,N_2952);
or UO_274 (O_274,N_2963,N_2969);
nor UO_275 (O_275,N_2962,N_2974);
nand UO_276 (O_276,N_2972,N_2983);
or UO_277 (O_277,N_2977,N_2960);
nor UO_278 (O_278,N_2975,N_2952);
and UO_279 (O_279,N_2952,N_2995);
and UO_280 (O_280,N_2999,N_2974);
or UO_281 (O_281,N_2958,N_2985);
nand UO_282 (O_282,N_2969,N_2978);
nand UO_283 (O_283,N_2984,N_2980);
nand UO_284 (O_284,N_2985,N_2973);
nor UO_285 (O_285,N_2978,N_2977);
or UO_286 (O_286,N_2980,N_2954);
and UO_287 (O_287,N_2995,N_2983);
and UO_288 (O_288,N_2964,N_2970);
or UO_289 (O_289,N_2999,N_2959);
or UO_290 (O_290,N_2999,N_2962);
xor UO_291 (O_291,N_2963,N_2959);
nand UO_292 (O_292,N_2993,N_2982);
nor UO_293 (O_293,N_2987,N_2955);
nand UO_294 (O_294,N_2983,N_2951);
nor UO_295 (O_295,N_2990,N_2971);
and UO_296 (O_296,N_2996,N_2973);
xor UO_297 (O_297,N_2956,N_2958);
nand UO_298 (O_298,N_2974,N_2993);
nor UO_299 (O_299,N_2977,N_2992);
or UO_300 (O_300,N_2989,N_2985);
nand UO_301 (O_301,N_2968,N_2950);
nor UO_302 (O_302,N_2986,N_2990);
or UO_303 (O_303,N_2985,N_2978);
xor UO_304 (O_304,N_2955,N_2990);
nand UO_305 (O_305,N_2997,N_2982);
or UO_306 (O_306,N_2951,N_2982);
or UO_307 (O_307,N_2965,N_2975);
xnor UO_308 (O_308,N_2996,N_2977);
and UO_309 (O_309,N_2971,N_2986);
nor UO_310 (O_310,N_2976,N_2975);
and UO_311 (O_311,N_2998,N_2982);
and UO_312 (O_312,N_2972,N_2998);
xor UO_313 (O_313,N_2955,N_2994);
and UO_314 (O_314,N_2995,N_2965);
nor UO_315 (O_315,N_2991,N_2964);
nand UO_316 (O_316,N_2965,N_2964);
or UO_317 (O_317,N_2951,N_2993);
nor UO_318 (O_318,N_2952,N_2976);
nor UO_319 (O_319,N_2968,N_2953);
or UO_320 (O_320,N_2950,N_2990);
or UO_321 (O_321,N_2994,N_2981);
and UO_322 (O_322,N_2957,N_2954);
and UO_323 (O_323,N_2984,N_2957);
nor UO_324 (O_324,N_2976,N_2971);
nand UO_325 (O_325,N_2966,N_2962);
or UO_326 (O_326,N_2962,N_2980);
and UO_327 (O_327,N_2960,N_2965);
or UO_328 (O_328,N_2988,N_2999);
and UO_329 (O_329,N_2972,N_2978);
and UO_330 (O_330,N_2982,N_2978);
nor UO_331 (O_331,N_2981,N_2965);
and UO_332 (O_332,N_2978,N_2956);
or UO_333 (O_333,N_2983,N_2954);
xor UO_334 (O_334,N_2976,N_2966);
and UO_335 (O_335,N_2979,N_2969);
or UO_336 (O_336,N_2981,N_2953);
nand UO_337 (O_337,N_2962,N_2951);
nor UO_338 (O_338,N_2993,N_2961);
nor UO_339 (O_339,N_2952,N_2981);
nand UO_340 (O_340,N_2987,N_2970);
and UO_341 (O_341,N_2987,N_2957);
nand UO_342 (O_342,N_2979,N_2987);
or UO_343 (O_343,N_2987,N_2974);
xnor UO_344 (O_344,N_2965,N_2966);
nand UO_345 (O_345,N_2980,N_2965);
nand UO_346 (O_346,N_2965,N_2983);
or UO_347 (O_347,N_2989,N_2988);
and UO_348 (O_348,N_2987,N_2961);
nand UO_349 (O_349,N_2973,N_2971);
nor UO_350 (O_350,N_2960,N_2984);
nor UO_351 (O_351,N_2962,N_2963);
nor UO_352 (O_352,N_2988,N_2998);
and UO_353 (O_353,N_2969,N_2985);
nor UO_354 (O_354,N_2983,N_2993);
or UO_355 (O_355,N_2973,N_2972);
nor UO_356 (O_356,N_2966,N_2959);
nor UO_357 (O_357,N_2981,N_2967);
or UO_358 (O_358,N_2991,N_2970);
and UO_359 (O_359,N_2979,N_2962);
nor UO_360 (O_360,N_2964,N_2961);
or UO_361 (O_361,N_2969,N_2965);
and UO_362 (O_362,N_2997,N_2969);
nor UO_363 (O_363,N_2954,N_2999);
or UO_364 (O_364,N_2975,N_2989);
and UO_365 (O_365,N_2954,N_2990);
or UO_366 (O_366,N_2975,N_2999);
nor UO_367 (O_367,N_2970,N_2951);
nor UO_368 (O_368,N_2961,N_2995);
nor UO_369 (O_369,N_2956,N_2954);
nor UO_370 (O_370,N_2994,N_2963);
or UO_371 (O_371,N_2966,N_2989);
nor UO_372 (O_372,N_2983,N_2967);
or UO_373 (O_373,N_2955,N_2950);
nand UO_374 (O_374,N_2965,N_2955);
or UO_375 (O_375,N_2992,N_2986);
or UO_376 (O_376,N_2984,N_2959);
nor UO_377 (O_377,N_2989,N_2999);
nand UO_378 (O_378,N_2970,N_2993);
nand UO_379 (O_379,N_2961,N_2962);
nor UO_380 (O_380,N_2963,N_2954);
nand UO_381 (O_381,N_2968,N_2971);
and UO_382 (O_382,N_2998,N_2965);
nand UO_383 (O_383,N_2990,N_2998);
nand UO_384 (O_384,N_2960,N_2957);
or UO_385 (O_385,N_2970,N_2959);
and UO_386 (O_386,N_2978,N_2983);
nor UO_387 (O_387,N_2962,N_2967);
nand UO_388 (O_388,N_2960,N_2979);
nor UO_389 (O_389,N_2999,N_2992);
nand UO_390 (O_390,N_2995,N_2959);
nor UO_391 (O_391,N_2989,N_2951);
nor UO_392 (O_392,N_2978,N_2974);
and UO_393 (O_393,N_2976,N_2979);
xnor UO_394 (O_394,N_2991,N_2972);
nor UO_395 (O_395,N_2960,N_2987);
and UO_396 (O_396,N_2955,N_2985);
and UO_397 (O_397,N_2990,N_2958);
or UO_398 (O_398,N_2963,N_2985);
and UO_399 (O_399,N_2968,N_2976);
nor UO_400 (O_400,N_2964,N_2976);
nor UO_401 (O_401,N_2971,N_2974);
and UO_402 (O_402,N_2984,N_2974);
or UO_403 (O_403,N_2981,N_2987);
nor UO_404 (O_404,N_2985,N_2951);
nand UO_405 (O_405,N_2962,N_2953);
nand UO_406 (O_406,N_2999,N_2957);
nand UO_407 (O_407,N_2955,N_2957);
nand UO_408 (O_408,N_2990,N_2993);
or UO_409 (O_409,N_2991,N_2979);
or UO_410 (O_410,N_2953,N_2965);
and UO_411 (O_411,N_2956,N_2996);
nand UO_412 (O_412,N_2993,N_2997);
and UO_413 (O_413,N_2993,N_2968);
nand UO_414 (O_414,N_2955,N_2956);
nor UO_415 (O_415,N_2998,N_2986);
nor UO_416 (O_416,N_2950,N_2976);
and UO_417 (O_417,N_2998,N_2994);
nand UO_418 (O_418,N_2955,N_2974);
nor UO_419 (O_419,N_2969,N_2994);
and UO_420 (O_420,N_2994,N_2965);
or UO_421 (O_421,N_2964,N_2953);
nor UO_422 (O_422,N_2984,N_2982);
nand UO_423 (O_423,N_2963,N_2955);
or UO_424 (O_424,N_2957,N_2993);
or UO_425 (O_425,N_2989,N_2979);
and UO_426 (O_426,N_2970,N_2997);
or UO_427 (O_427,N_2954,N_2986);
or UO_428 (O_428,N_2977,N_2970);
or UO_429 (O_429,N_2974,N_2950);
nand UO_430 (O_430,N_2955,N_2958);
or UO_431 (O_431,N_2996,N_2954);
nor UO_432 (O_432,N_2977,N_2958);
nor UO_433 (O_433,N_2955,N_2988);
or UO_434 (O_434,N_2975,N_2964);
or UO_435 (O_435,N_2973,N_2952);
or UO_436 (O_436,N_2993,N_2986);
and UO_437 (O_437,N_2979,N_2980);
or UO_438 (O_438,N_2971,N_2951);
nand UO_439 (O_439,N_2994,N_2966);
nor UO_440 (O_440,N_2994,N_2992);
xnor UO_441 (O_441,N_2987,N_2998);
nor UO_442 (O_442,N_2950,N_2954);
nand UO_443 (O_443,N_2969,N_2999);
nand UO_444 (O_444,N_2995,N_2974);
nor UO_445 (O_445,N_2958,N_2954);
and UO_446 (O_446,N_2969,N_2984);
and UO_447 (O_447,N_2997,N_2950);
and UO_448 (O_448,N_2986,N_2975);
and UO_449 (O_449,N_2973,N_2988);
or UO_450 (O_450,N_2960,N_2973);
nor UO_451 (O_451,N_2997,N_2992);
nand UO_452 (O_452,N_2971,N_2985);
or UO_453 (O_453,N_2958,N_2951);
and UO_454 (O_454,N_2962,N_2985);
nor UO_455 (O_455,N_2991,N_2992);
and UO_456 (O_456,N_2980,N_2975);
nor UO_457 (O_457,N_2998,N_2999);
or UO_458 (O_458,N_2955,N_2971);
nand UO_459 (O_459,N_2950,N_2994);
and UO_460 (O_460,N_2973,N_2987);
nor UO_461 (O_461,N_2960,N_2975);
nor UO_462 (O_462,N_2967,N_2985);
and UO_463 (O_463,N_2961,N_2963);
nor UO_464 (O_464,N_2985,N_2987);
or UO_465 (O_465,N_2961,N_2999);
nand UO_466 (O_466,N_2982,N_2964);
nor UO_467 (O_467,N_2996,N_2958);
or UO_468 (O_468,N_2983,N_2996);
nand UO_469 (O_469,N_2980,N_2950);
nand UO_470 (O_470,N_2984,N_2995);
nand UO_471 (O_471,N_2972,N_2966);
and UO_472 (O_472,N_2963,N_2988);
or UO_473 (O_473,N_2974,N_2964);
nor UO_474 (O_474,N_2959,N_2960);
or UO_475 (O_475,N_2995,N_2966);
nor UO_476 (O_476,N_2986,N_2995);
nand UO_477 (O_477,N_2992,N_2972);
and UO_478 (O_478,N_2978,N_2999);
nor UO_479 (O_479,N_2965,N_2963);
nor UO_480 (O_480,N_2956,N_2962);
and UO_481 (O_481,N_2988,N_2979);
nor UO_482 (O_482,N_2955,N_2968);
nand UO_483 (O_483,N_2995,N_2962);
or UO_484 (O_484,N_2957,N_2956);
or UO_485 (O_485,N_2973,N_2968);
nor UO_486 (O_486,N_2990,N_2961);
nor UO_487 (O_487,N_2997,N_2977);
or UO_488 (O_488,N_2973,N_2969);
nor UO_489 (O_489,N_2968,N_2992);
nor UO_490 (O_490,N_2960,N_2996);
nor UO_491 (O_491,N_2976,N_2992);
nand UO_492 (O_492,N_2968,N_2981);
and UO_493 (O_493,N_2961,N_2973);
and UO_494 (O_494,N_2966,N_2956);
and UO_495 (O_495,N_2980,N_2951);
or UO_496 (O_496,N_2990,N_2979);
nor UO_497 (O_497,N_2959,N_2962);
or UO_498 (O_498,N_2969,N_2998);
or UO_499 (O_499,N_2956,N_2971);
endmodule