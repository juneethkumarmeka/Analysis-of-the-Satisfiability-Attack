module basic_1500_15000_2000_3_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10002,N_10003,N_10004,N_10006,N_10007,N_10009,N_10010,N_10011,N_10012,N_10014,N_10015,N_10016,N_10018,N_10022,N_10023,N_10024,N_10027,N_10028,N_10030,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10042,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10053,N_10056,N_10057,N_10058,N_10059,N_10060,N_10062,N_10063,N_10064,N_10066,N_10068,N_10069,N_10070,N_10071,N_10072,N_10074,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10099,N_10100,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10116,N_10117,N_10118,N_10119,N_10120,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10139,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10161,N_10162,N_10163,N_10164,N_10166,N_10168,N_10169,N_10170,N_10171,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10186,N_10188,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10209,N_10210,N_10211,N_10212,N_10213,N_10218,N_10220,N_10221,N_10223,N_10224,N_10225,N_10227,N_10228,N_10230,N_10233,N_10235,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10248,N_10249,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10259,N_10260,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10273,N_10274,N_10275,N_10276,N_10277,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10329,N_10330,N_10333,N_10334,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10345,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10354,N_10355,N_10356,N_10358,N_10360,N_10363,N_10366,N_10367,N_10368,N_10369,N_10370,N_10372,N_10373,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10410,N_10412,N_10413,N_10414,N_10416,N_10418,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10428,N_10429,N_10430,N_10431,N_10432,N_10435,N_10437,N_10438,N_10439,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10451,N_10453,N_10455,N_10456,N_10458,N_10459,N_10461,N_10463,N_10465,N_10466,N_10468,N_10469,N_10470,N_10471,N_10472,N_10474,N_10475,N_10476,N_10478,N_10480,N_10481,N_10482,N_10483,N_10485,N_10486,N_10487,N_10489,N_10490,N_10492,N_10493,N_10494,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10506,N_10507,N_10509,N_10510,N_10512,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10525,N_10527,N_10528,N_10530,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10547,N_10548,N_10549,N_10550,N_10552,N_10554,N_10555,N_10556,N_10557,N_10558,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10587,N_10588,N_10589,N_10590,N_10591,N_10593,N_10594,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10607,N_10608,N_10609,N_10610,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10620,N_10621,N_10622,N_10623,N_10626,N_10627,N_10628,N_10629,N_10631,N_10633,N_10635,N_10636,N_10637,N_10639,N_10640,N_10641,N_10642,N_10644,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10670,N_10672,N_10673,N_10674,N_10677,N_10679,N_10680,N_10681,N_10685,N_10687,N_10688,N_10690,N_10691,N_10694,N_10695,N_10696,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10724,N_10726,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10737,N_10738,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10751,N_10752,N_10754,N_10755,N_10756,N_10758,N_10759,N_10760,N_10761,N_10762,N_10765,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10788,N_10790,N_10792,N_10793,N_10794,N_10795,N_10796,N_10798,N_10799,N_10800,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10814,N_10815,N_10816,N_10817,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10843,N_10844,N_10845,N_10846,N_10847,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10862,N_10863,N_10864,N_10865,N_10867,N_10869,N_10870,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10881,N_10882,N_10883,N_10884,N_10886,N_10887,N_10888,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10904,N_10905,N_10906,N_10907,N_10909,N_10910,N_10911,N_10913,N_10914,N_10915,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10932,N_10933,N_10935,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10959,N_10960,N_10961,N_10964,N_10965,N_10966,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10979,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10991,N_10992,N_10994,N_10995,N_10996,N_10997,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11006,N_11007,N_11009,N_11010,N_11011,N_11012,N_11013,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11031,N_11034,N_11035,N_11036,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11045,N_11046,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11056,N_11058,N_11059,N_11060,N_11062,N_11063,N_11065,N_11066,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11075,N_11076,N_11077,N_11078,N_11079,N_11081,N_11082,N_11083,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11095,N_11098,N_11099,N_11100,N_11101,N_11102,N_11104,N_11105,N_11107,N_11108,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11121,N_11122,N_11123,N_11124,N_11125,N_11127,N_11130,N_11131,N_11135,N_11136,N_11137,N_11139,N_11140,N_11141,N_11143,N_11145,N_11146,N_11147,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11158,N_11160,N_11161,N_11162,N_11164,N_11165,N_11166,N_11168,N_11169,N_11171,N_11172,N_11173,N_11174,N_11175,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11216,N_11217,N_11218,N_11219,N_11221,N_11222,N_11224,N_11226,N_11227,N_11228,N_11229,N_11231,N_11233,N_11235,N_11237,N_11239,N_11240,N_11241,N_11242,N_11243,N_11245,N_11246,N_11247,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11266,N_11267,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11284,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11313,N_11314,N_11315,N_11316,N_11317,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11330,N_11332,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11348,N_11350,N_11351,N_11352,N_11353,N_11356,N_11358,N_11359,N_11360,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11371,N_11372,N_11373,N_11374,N_11376,N_11377,N_11378,N_11379,N_11381,N_11382,N_11384,N_11385,N_11386,N_11387,N_11389,N_11390,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11402,N_11403,N_11404,N_11405,N_11408,N_11410,N_11411,N_11414,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11425,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11446,N_11448,N_11449,N_11450,N_11451,N_11453,N_11454,N_11455,N_11457,N_11459,N_11460,N_11464,N_11465,N_11467,N_11468,N_11469,N_11471,N_11472,N_11473,N_11475,N_11477,N_11478,N_11479,N_11480,N_11481,N_11483,N_11484,N_11485,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11497,N_11498,N_11499,N_11500,N_11501,N_11503,N_11504,N_11505,N_11507,N_11508,N_11509,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11525,N_11526,N_11527,N_11528,N_11530,N_11531,N_11532,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11542,N_11543,N_11544,N_11547,N_11548,N_11549,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11558,N_11560,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11583,N_11584,N_11585,N_11586,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11619,N_11620,N_11621,N_11624,N_11625,N_11626,N_11627,N_11628,N_11630,N_11631,N_11633,N_11634,N_11636,N_11637,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11651,N_11652,N_11653,N_11655,N_11657,N_11658,N_11659,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11671,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11680,N_11682,N_11683,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11694,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11707,N_11708,N_11710,N_11711,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11748,N_11749,N_11751,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11765,N_11766,N_11767,N_11768,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11822,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11831,N_11832,N_11833,N_11834,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11867,N_11868,N_11870,N_11871,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11893,N_11894,N_11895,N_11897,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11906,N_11908,N_11910,N_11911,N_11912,N_11913,N_11914,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11926,N_11927,N_11928,N_11929,N_11931,N_11932,N_11933,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11945,N_11946,N_11947,N_11949,N_11950,N_11951,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11967,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12058,N_12059,N_12060,N_12063,N_12065,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12080,N_12081,N_12082,N_12083,N_12084,N_12087,N_12088,N_12089,N_12090,N_12091,N_12094,N_12095,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12116,N_12118,N_12119,N_12121,N_12123,N_12124,N_12125,N_12126,N_12127,N_12129,N_12130,N_12131,N_12133,N_12134,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12163,N_12164,N_12165,N_12166,N_12167,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12177,N_12179,N_12181,N_12182,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12192,N_12194,N_12195,N_12196,N_12198,N_12199,N_12200,N_12201,N_12202,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12216,N_12217,N_12218,N_12219,N_12221,N_12222,N_12223,N_12224,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12264,N_12265,N_12266,N_12269,N_12270,N_12272,N_12273,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12318,N_12321,N_12323,N_12324,N_12325,N_12326,N_12328,N_12330,N_12331,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12374,N_12376,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12391,N_12394,N_12395,N_12396,N_12398,N_12399,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12408,N_12409,N_12410,N_12412,N_12413,N_12414,N_12415,N_12416,N_12419,N_12420,N_12421,N_12422,N_12423,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12433,N_12434,N_12436,N_12437,N_12438,N_12439,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12456,N_12457,N_12458,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12493,N_12494,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12503,N_12504,N_12505,N_12507,N_12510,N_12511,N_12513,N_12514,N_12515,N_12516,N_12517,N_12519,N_12520,N_12521,N_12523,N_12524,N_12526,N_12528,N_12529,N_12530,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12548,N_12549,N_12550,N_12551,N_12552,N_12556,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12593,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12607,N_12609,N_12612,N_12613,N_12614,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12625,N_12628,N_12629,N_12630,N_12631,N_12632,N_12635,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12654,N_12655,N_12656,N_12658,N_12659,N_12662,N_12663,N_12665,N_12666,N_12667,N_12670,N_12671,N_12672,N_12673,N_12674,N_12676,N_12677,N_12678,N_12679,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12693,N_12694,N_12697,N_12698,N_12699,N_12700,N_12702,N_12704,N_12705,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12732,N_12733,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12751,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12761,N_12762,N_12764,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12785,N_12787,N_12789,N_12790,N_12791,N_12793,N_12795,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12807,N_12808,N_12809,N_12810,N_12812,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12823,N_12826,N_12827,N_12828,N_12830,N_12831,N_12832,N_12834,N_12836,N_12837,N_12838,N_12839,N_12841,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12863,N_12864,N_12865,N_12867,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12877,N_12878,N_12880,N_12881,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12890,N_12892,N_12893,N_12895,N_12896,N_12899,N_12900,N_12901,N_12902,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12937,N_12938,N_12940,N_12942,N_12943,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12954,N_12955,N_12956,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12981,N_12982,N_12983,N_12984,N_12985,N_12987,N_12989,N_12990,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13004,N_13005,N_13006,N_13008,N_13009,N_13010,N_13011,N_13013,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13025,N_13027,N_13028,N_13029,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13039,N_13040,N_13041,N_13042,N_13044,N_13045,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13076,N_13077,N_13080,N_13081,N_13082,N_13083,N_13084,N_13086,N_13087,N_13089,N_13090,N_13091,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13111,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13123,N_13125,N_13126,N_13127,N_13128,N_13130,N_13131,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13151,N_13152,N_13153,N_13154,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13169,N_13170,N_13171,N_13172,N_13173,N_13175,N_13177,N_13178,N_13179,N_13183,N_13185,N_13186,N_13187,N_13188,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13198,N_13199,N_13201,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13210,N_13212,N_13213,N_13215,N_13216,N_13217,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13235,N_13236,N_13238,N_13239,N_13241,N_13242,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13266,N_13267,N_13268,N_13269,N_13271,N_13273,N_13274,N_13275,N_13276,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13293,N_13294,N_13295,N_13296,N_13299,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13313,N_13314,N_13315,N_13318,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13333,N_13334,N_13335,N_13336,N_13339,N_13340,N_13341,N_13342,N_13345,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13355,N_13356,N_13357,N_13358,N_13359,N_13361,N_13362,N_13363,N_13364,N_13365,N_13367,N_13368,N_13370,N_13371,N_13372,N_13374,N_13376,N_13377,N_13379,N_13380,N_13382,N_13383,N_13384,N_13385,N_13386,N_13388,N_13389,N_13391,N_13392,N_13393,N_13394,N_13395,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13426,N_13427,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13447,N_13448,N_13449,N_13450,N_13452,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13476,N_13477,N_13478,N_13480,N_13481,N_13482,N_13483,N_13485,N_13486,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13501,N_13502,N_13503,N_13504,N_13506,N_13507,N_13509,N_13510,N_13511,N_13512,N_13513,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13523,N_13525,N_13526,N_13527,N_13528,N_13529,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13568,N_13571,N_13572,N_13573,N_13574,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13585,N_13586,N_13588,N_13590,N_13591,N_13593,N_13594,N_13595,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13630,N_13632,N_13633,N_13634,N_13635,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13645,N_13646,N_13647,N_13649,N_13650,N_13651,N_13652,N_13655,N_13656,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13678,N_13679,N_13680,N_13681,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13693,N_13694,N_13695,N_13696,N_13698,N_13700,N_13701,N_13702,N_13703,N_13704,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13716,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13731,N_13733,N_13734,N_13736,N_13740,N_13741,N_13742,N_13743,N_13745,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13757,N_13758,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13779,N_13780,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13790,N_13791,N_13792,N_13795,N_13796,N_13797,N_13798,N_13799,N_13801,N_13802,N_13803,N_13806,N_13807,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13820,N_13821,N_13823,N_13825,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13837,N_13840,N_13841,N_13842,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13869,N_13870,N_13871,N_13872,N_13873,N_13878,N_13879,N_13880,N_13881,N_13882,N_13884,N_13885,N_13886,N_13887,N_13889,N_13890,N_13892,N_13894,N_13895,N_13896,N_13900,N_13901,N_13904,N_13906,N_13907,N_13908,N_13910,N_13911,N_13913,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13930,N_13931,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13942,N_13944,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13965,N_13967,N_13968,N_13969,N_13970,N_13972,N_13973,N_13974,N_13975,N_13976,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13995,N_13996,N_13997,N_13998,N_13999,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14009,N_14010,N_14011,N_14012,N_14013,N_14016,N_14017,N_14018,N_14019,N_14021,N_14022,N_14023,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14044,N_14045,N_14046,N_14047,N_14049,N_14050,N_14051,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14063,N_14064,N_14065,N_14066,N_14067,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14076,N_14077,N_14079,N_14082,N_14083,N_14084,N_14085,N_14086,N_14088,N_14089,N_14090,N_14091,N_14092,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14117,N_14118,N_14119,N_14120,N_14121,N_14123,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14143,N_14145,N_14146,N_14147,N_14148,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14201,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14213,N_14214,N_14215,N_14217,N_14218,N_14219,N_14221,N_14225,N_14226,N_14227,N_14231,N_14232,N_14233,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14242,N_14243,N_14247,N_14248,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14263,N_14264,N_14266,N_14267,N_14268,N_14269,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14281,N_14282,N_14283,N_14284,N_14286,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14298,N_14299,N_14300,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14323,N_14324,N_14325,N_14327,N_14328,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14353,N_14354,N_14355,N_14356,N_14357,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14368,N_14369,N_14370,N_14372,N_14373,N_14374,N_14375,N_14377,N_14378,N_14380,N_14382,N_14383,N_14384,N_14386,N_14387,N_14388,N_14389,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14409,N_14410,N_14411,N_14412,N_14414,N_14415,N_14417,N_14419,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14450,N_14452,N_14453,N_14455,N_14456,N_14457,N_14458,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14467,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14501,N_14502,N_14503,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14530,N_14531,N_14532,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14546,N_14548,N_14549,N_14550,N_14551,N_14553,N_14554,N_14555,N_14556,N_14558,N_14559,N_14560,N_14561,N_14563,N_14564,N_14566,N_14567,N_14568,N_14569,N_14570,N_14572,N_14573,N_14574,N_14575,N_14576,N_14578,N_14579,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14602,N_14603,N_14604,N_14605,N_14606,N_14608,N_14609,N_14610,N_14611,N_14612,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14640,N_14641,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14672,N_14673,N_14674,N_14675,N_14676,N_14678,N_14680,N_14681,N_14682,N_14683,N_14684,N_14686,N_14687,N_14689,N_14690,N_14691,N_14692,N_14693,N_14695,N_14696,N_14697,N_14698,N_14700,N_14701,N_14702,N_14704,N_14705,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14714,N_14715,N_14716,N_14718,N_14723,N_14724,N_14725,N_14728,N_14729,N_14730,N_14731,N_14732,N_14735,N_14736,N_14737,N_14738,N_14739,N_14742,N_14743,N_14745,N_14746,N_14748,N_14749,N_14750,N_14751,N_14753,N_14754,N_14755,N_14757,N_14758,N_14759,N_14760,N_14763,N_14764,N_14766,N_14767,N_14768,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14779,N_14780,N_14781,N_14782,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14866,N_14868,N_14870,N_14871,N_14873,N_14874,N_14875,N_14876,N_14878,N_14879,N_14880,N_14881,N_14883,N_14884,N_14886,N_14887,N_14888,N_14889,N_14890,N_14893,N_14894,N_14895,N_14896,N_14897,N_14899,N_14900,N_14901,N_14902,N_14904,N_14905,N_14906,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14916,N_14917,N_14918,N_14920,N_14921,N_14922,N_14925,N_14926,N_14927,N_14928,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14953,N_14954,N_14955,N_14957,N_14959,N_14960,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14969,N_14970,N_14972,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1415,In_1240);
nand U1 (N_1,In_553,In_1274);
nand U2 (N_2,In_911,In_1160);
xnor U3 (N_3,In_653,In_276);
nand U4 (N_4,In_177,In_257);
nor U5 (N_5,In_756,In_1393);
and U6 (N_6,In_362,In_285);
xnor U7 (N_7,In_44,In_1477);
nor U8 (N_8,In_1287,In_839);
xnor U9 (N_9,In_422,In_1437);
and U10 (N_10,In_678,In_880);
and U11 (N_11,In_1243,In_154);
nor U12 (N_12,In_1245,In_1443);
nor U13 (N_13,In_1368,In_353);
and U14 (N_14,In_1339,In_235);
xnor U15 (N_15,In_1398,In_225);
nor U16 (N_16,In_987,In_575);
xor U17 (N_17,In_93,In_110);
nor U18 (N_18,In_397,In_32);
xor U19 (N_19,In_1221,In_238);
xor U20 (N_20,In_446,In_356);
or U21 (N_21,In_1338,In_569);
and U22 (N_22,In_1340,In_414);
or U23 (N_23,In_461,In_564);
nand U24 (N_24,In_760,In_803);
nor U25 (N_25,In_557,In_635);
and U26 (N_26,In_814,In_490);
or U27 (N_27,In_492,In_1344);
nor U28 (N_28,In_361,In_368);
xor U29 (N_29,In_301,In_1422);
xnor U30 (N_30,In_853,In_174);
nand U31 (N_31,In_1222,In_271);
nand U32 (N_32,In_1011,In_1029);
or U33 (N_33,In_943,In_1182);
or U34 (N_34,In_1329,In_722);
xnor U35 (N_35,In_1311,In_775);
xnor U36 (N_36,In_873,In_1291);
nor U37 (N_37,In_1288,In_950);
or U38 (N_38,In_907,In_1041);
or U39 (N_39,In_945,In_738);
nor U40 (N_40,In_1408,In_662);
and U41 (N_41,In_1219,In_1172);
nand U42 (N_42,In_532,In_26);
nand U43 (N_43,In_516,In_523);
and U44 (N_44,In_654,In_473);
and U45 (N_45,In_169,In_545);
nor U46 (N_46,In_1301,In_1430);
nor U47 (N_47,In_981,In_230);
nand U48 (N_48,In_1060,In_164);
nand U49 (N_49,In_11,In_1120);
xor U50 (N_50,In_588,In_268);
xnor U51 (N_51,In_940,In_53);
xnor U52 (N_52,In_1295,In_968);
xnor U53 (N_53,In_404,In_1103);
xnor U54 (N_54,In_596,In_568);
nor U55 (N_55,In_369,In_994);
nand U56 (N_56,In_410,In_1105);
xnor U57 (N_57,In_1350,In_672);
nor U58 (N_58,In_1209,In_69);
and U59 (N_59,In_65,In_1457);
xnor U60 (N_60,In_340,In_871);
xnor U61 (N_61,In_71,In_455);
nand U62 (N_62,In_1231,In_425);
nor U63 (N_63,In_609,In_24);
or U64 (N_64,In_903,In_72);
or U65 (N_65,In_424,In_1224);
xnor U66 (N_66,In_1284,In_1450);
nor U67 (N_67,In_1062,In_622);
xor U68 (N_68,In_142,In_891);
xnor U69 (N_69,In_148,In_339);
or U70 (N_70,In_354,In_636);
nor U71 (N_71,In_121,In_1346);
nand U72 (N_72,In_1214,In_1180);
and U73 (N_73,In_474,In_377);
nand U74 (N_74,In_909,In_211);
and U75 (N_75,In_953,In_1199);
nor U76 (N_76,In_76,In_453);
xor U77 (N_77,In_694,In_702);
nand U78 (N_78,In_212,In_1249);
nand U79 (N_79,In_1235,In_1205);
nor U80 (N_80,In_1002,In_777);
xnor U81 (N_81,In_639,In_979);
and U82 (N_82,In_638,In_1316);
xnor U83 (N_83,In_548,In_280);
and U84 (N_84,In_542,In_315);
or U85 (N_85,In_753,In_1232);
xnor U86 (N_86,In_868,In_107);
and U87 (N_87,In_1386,In_1006);
nor U88 (N_88,In_1404,In_888);
and U89 (N_89,In_398,In_84);
xor U90 (N_90,In_1061,In_677);
and U91 (N_91,In_196,In_1091);
or U92 (N_92,In_795,In_996);
nor U93 (N_93,In_912,In_367);
xnor U94 (N_94,In_927,In_1435);
xor U95 (N_95,In_949,In_746);
and U96 (N_96,In_854,In_580);
or U97 (N_97,In_432,In_1347);
or U98 (N_98,In_1446,In_780);
and U99 (N_99,In_1442,In_224);
nand U100 (N_100,In_37,In_203);
or U101 (N_101,In_1043,In_1434);
and U102 (N_102,In_403,In_1161);
and U103 (N_103,In_436,In_1376);
and U104 (N_104,In_965,In_842);
xor U105 (N_105,In_882,In_723);
and U106 (N_106,In_117,In_320);
or U107 (N_107,In_748,In_102);
xor U108 (N_108,In_657,In_974);
xor U109 (N_109,In_1330,In_326);
nor U110 (N_110,In_1036,In_525);
xor U111 (N_111,In_438,In_1271);
or U112 (N_112,In_159,In_1119);
nand U113 (N_113,In_852,In_952);
nand U114 (N_114,In_1387,In_1471);
or U115 (N_115,In_876,In_192);
nand U116 (N_116,In_380,In_845);
or U117 (N_117,In_787,In_337);
nand U118 (N_118,In_561,In_1308);
or U119 (N_119,In_329,In_449);
and U120 (N_120,In_566,In_623);
nor U121 (N_121,In_1290,In_769);
nand U122 (N_122,In_563,In_496);
xnor U123 (N_123,In_1109,In_1144);
xnor U124 (N_124,In_524,In_45);
nor U125 (N_125,In_1298,In_584);
or U126 (N_126,In_520,In_123);
nand U127 (N_127,In_939,In_386);
nor U128 (N_128,In_1012,In_560);
xor U129 (N_129,In_298,In_1448);
nor U130 (N_130,In_1454,In_1055);
xor U131 (N_131,In_1260,In_1263);
or U132 (N_132,In_799,In_665);
nor U133 (N_133,In_143,In_334);
xor U134 (N_134,In_1239,In_9);
nand U135 (N_135,In_254,In_1265);
or U136 (N_136,In_593,In_1475);
or U137 (N_137,In_883,In_1299);
nor U138 (N_138,In_1374,In_460);
or U139 (N_139,In_201,In_1065);
or U140 (N_140,In_183,In_1273);
or U141 (N_141,In_1303,In_620);
xnor U142 (N_142,In_381,In_1162);
and U143 (N_143,In_1035,In_155);
nand U144 (N_144,In_830,In_886);
xnor U145 (N_145,In_1497,In_942);
and U146 (N_146,In_1039,In_416);
nand U147 (N_147,In_364,In_1115);
and U148 (N_148,In_1028,In_15);
nor U149 (N_149,In_714,In_1075);
xor U150 (N_150,In_162,In_1013);
xnor U151 (N_151,In_816,In_1394);
or U152 (N_152,In_679,In_1428);
xnor U153 (N_153,In_605,In_969);
nor U154 (N_154,In_286,In_1466);
nand U155 (N_155,In_558,In_972);
or U156 (N_156,In_926,In_675);
nand U157 (N_157,In_1348,In_721);
nand U158 (N_158,In_152,In_388);
nand U159 (N_159,In_629,In_101);
xnor U160 (N_160,In_1268,In_1355);
xnor U161 (N_161,In_779,In_772);
xnor U162 (N_162,In_1197,In_713);
nand U163 (N_163,In_1112,In_744);
and U164 (N_164,In_1072,In_433);
or U165 (N_165,In_385,In_437);
nor U166 (N_166,In_917,In_1001);
nand U167 (N_167,In_505,In_223);
nor U168 (N_168,In_897,In_934);
nor U169 (N_169,In_1229,In_796);
nor U170 (N_170,In_111,In_1085);
nor U171 (N_171,In_597,In_113);
nand U172 (N_172,In_218,In_322);
xor U173 (N_173,In_935,In_592);
xnor U174 (N_174,In_1238,In_961);
or U175 (N_175,In_293,In_1022);
or U176 (N_176,In_791,In_1280);
or U177 (N_177,In_1345,In_944);
and U178 (N_178,In_80,In_1191);
xnor U179 (N_179,In_992,In_234);
xor U180 (N_180,In_144,In_468);
nor U181 (N_181,In_606,In_401);
nand U182 (N_182,In_242,In_1048);
and U183 (N_183,In_1370,In_712);
nor U184 (N_184,In_331,In_175);
xnor U185 (N_185,In_745,In_332);
and U186 (N_186,In_1285,In_846);
nand U187 (N_187,In_669,In_265);
or U188 (N_188,In_1196,In_13);
and U189 (N_189,In_1272,In_439);
and U190 (N_190,In_1320,In_156);
or U191 (N_191,In_1147,In_682);
or U192 (N_192,In_1116,In_408);
and U193 (N_193,In_5,In_179);
and U194 (N_194,In_749,In_956);
or U195 (N_195,In_1401,In_739);
nand U196 (N_196,In_241,In_1490);
nor U197 (N_197,In_633,In_836);
nand U198 (N_198,In_920,In_627);
or U199 (N_199,In_1210,In_829);
nor U200 (N_200,In_1121,In_614);
nand U201 (N_201,In_826,In_719);
nand U202 (N_202,In_452,In_1233);
xnor U203 (N_203,In_23,In_879);
nor U204 (N_204,In_12,In_57);
nand U205 (N_205,In_374,In_498);
and U206 (N_206,In_812,In_861);
xnor U207 (N_207,In_1194,In_287);
and U208 (N_208,In_1066,In_428);
nor U209 (N_209,In_890,In_1409);
nand U210 (N_210,In_948,In_1079);
or U211 (N_211,In_172,In_790);
xnor U212 (N_212,In_783,In_83);
xnor U213 (N_213,In_108,In_1436);
nor U214 (N_214,In_124,In_134);
and U215 (N_215,In_1252,In_1292);
nor U216 (N_216,In_366,In_877);
and U217 (N_217,In_458,In_199);
nand U218 (N_218,In_325,In_1247);
xnor U219 (N_219,In_1123,In_1126);
nor U220 (N_220,In_1007,In_1171);
or U221 (N_221,In_1014,In_549);
nand U222 (N_222,In_720,In_918);
nor U223 (N_223,In_774,In_690);
or U224 (N_224,In_762,In_1094);
xnor U225 (N_225,In_1371,In_1474);
or U226 (N_226,In_973,In_1410);
nand U227 (N_227,In_1318,In_922);
nand U228 (N_228,In_409,In_48);
xnor U229 (N_229,In_770,In_878);
and U230 (N_230,In_151,In_1143);
nand U231 (N_231,In_63,In_991);
nor U232 (N_232,In_650,In_1419);
and U233 (N_233,In_256,In_1080);
and U234 (N_234,In_3,In_92);
nor U235 (N_235,In_841,In_349);
and U236 (N_236,In_264,In_711);
xor U237 (N_237,In_365,In_1153);
nor U238 (N_238,In_881,In_1372);
and U239 (N_239,In_278,In_1176);
nor U240 (N_240,In_689,In_914);
or U241 (N_241,In_1195,In_1369);
and U242 (N_242,In_615,In_699);
xor U243 (N_243,In_247,In_249);
and U244 (N_244,In_344,In_1468);
or U245 (N_245,In_1418,In_273);
nor U246 (N_246,In_1325,In_798);
nor U247 (N_247,In_1237,In_288);
or U248 (N_248,In_1354,In_1148);
and U249 (N_249,In_493,In_801);
nand U250 (N_250,In_1278,In_915);
nand U251 (N_251,In_98,In_208);
nor U252 (N_252,In_114,In_1244);
and U253 (N_253,In_1360,In_58);
nor U254 (N_254,In_28,In_500);
or U255 (N_255,In_571,In_697);
nand U256 (N_256,In_1008,In_724);
nand U257 (N_257,In_316,In_1017);
and U258 (N_258,In_1300,In_467);
nand U259 (N_259,In_901,In_1154);
nor U260 (N_260,In_962,In_259);
nor U261 (N_261,In_239,In_34);
nor U262 (N_262,In_1169,In_105);
or U263 (N_263,In_1015,In_685);
xnor U264 (N_264,In_91,In_87);
nor U265 (N_265,In_1441,In_1269);
nor U266 (N_266,In_363,In_640);
xnor U267 (N_267,In_370,In_1070);
and U268 (N_268,In_715,In_181);
or U269 (N_269,In_1484,In_243);
xor U270 (N_270,In_1362,In_462);
nand U271 (N_271,In_378,In_999);
and U272 (N_272,In_180,In_550);
and U273 (N_273,In_747,In_1351);
and U274 (N_274,In_1411,In_663);
xnor U275 (N_275,In_1444,In_501);
xnor U276 (N_276,In_1420,In_691);
nand U277 (N_277,In_450,In_1117);
nand U278 (N_278,In_487,In_552);
nand U279 (N_279,In_863,In_1439);
nor U280 (N_280,In_499,In_1433);
or U281 (N_281,In_1107,In_413);
nor U282 (N_282,In_522,In_843);
xor U283 (N_283,In_305,In_734);
xor U284 (N_284,In_1204,In_391);
or U285 (N_285,In_910,In_383);
nand U286 (N_286,In_921,In_1451);
nand U287 (N_287,In_1499,In_488);
or U288 (N_288,In_309,In_209);
and U289 (N_289,In_1257,In_819);
and U290 (N_290,In_335,In_61);
nor U291 (N_291,In_1098,In_1077);
or U292 (N_292,In_1495,In_1138);
and U293 (N_293,In_621,In_125);
xor U294 (N_294,In_806,In_825);
or U295 (N_295,In_430,In_191);
and U296 (N_296,In_497,In_900);
nand U297 (N_297,In_1425,In_476);
and U298 (N_298,In_975,In_1128);
xnor U299 (N_299,In_1220,In_1053);
nand U300 (N_300,In_1076,In_1395);
xnor U301 (N_301,In_22,In_618);
nor U302 (N_302,In_521,In_735);
nand U303 (N_303,In_572,In_6);
nor U304 (N_304,In_214,In_630);
and U305 (N_305,In_740,In_1203);
xnor U306 (N_306,In_707,In_7);
or U307 (N_307,In_634,In_1492);
nand U308 (N_308,In_185,In_384);
or U309 (N_309,In_481,In_1491);
nand U310 (N_310,In_463,In_1163);
and U311 (N_311,In_684,In_423);
xnor U312 (N_312,In_1302,In_303);
and U313 (N_313,In_717,In_1262);
nand U314 (N_314,In_360,In_984);
nand U315 (N_315,In_632,In_1294);
nand U316 (N_316,In_10,In_1152);
nand U317 (N_317,In_986,In_392);
or U318 (N_318,In_127,In_170);
nand U319 (N_319,In_867,In_415);
nand U320 (N_320,In_1242,In_1040);
or U321 (N_321,In_793,In_947);
xor U322 (N_322,In_872,In_1289);
xor U323 (N_323,In_1184,In_1432);
and U324 (N_324,In_1092,In_262);
nand U325 (N_325,In_1321,In_628);
or U326 (N_326,In_706,In_565);
nand U327 (N_327,In_1248,In_275);
or U328 (N_328,In_421,In_14);
nor U329 (N_329,In_1025,In_1423);
xor U330 (N_330,In_1429,In_692);
xor U331 (N_331,In_937,In_959);
or U332 (N_332,In_456,In_1267);
or U333 (N_333,In_120,In_300);
nor U334 (N_334,In_808,In_1057);
nand U335 (N_335,In_279,In_1113);
or U336 (N_336,In_1174,In_1133);
nor U337 (N_337,In_1337,In_556);
and U338 (N_338,In_989,In_1306);
or U339 (N_339,In_296,In_133);
nor U340 (N_340,In_40,In_246);
and U341 (N_341,In_479,In_850);
xnor U342 (N_342,In_171,In_1390);
nand U343 (N_343,In_1333,In_393);
nand U344 (N_344,In_631,In_35);
or U345 (N_345,In_1122,In_1037);
nor U346 (N_346,In_411,In_138);
or U347 (N_347,In_1421,In_312);
nor U348 (N_348,In_1190,In_1464);
nor U349 (N_349,In_182,In_670);
and U350 (N_350,In_824,In_905);
and U351 (N_351,In_1286,In_495);
or U352 (N_352,In_119,In_274);
nor U353 (N_353,In_1101,In_1427);
and U354 (N_354,In_166,In_4);
nor U355 (N_355,In_232,In_1391);
nand U356 (N_356,In_1185,In_815);
or U357 (N_357,In_158,In_587);
nor U358 (N_358,In_874,In_1255);
xor U359 (N_359,In_782,In_604);
and U360 (N_360,In_1198,In_931);
nand U361 (N_361,In_104,In_444);
nand U362 (N_362,In_176,In_810);
nand U363 (N_363,In_695,In_625);
xnor U364 (N_364,In_38,In_1124);
xor U365 (N_365,In_851,In_135);
or U366 (N_366,In_544,In_792);
and U367 (N_367,In_660,In_1259);
or U368 (N_368,In_645,In_115);
xor U369 (N_369,In_431,In_323);
or U370 (N_370,In_1137,In_902);
nand U371 (N_371,In_673,In_1149);
and U372 (N_372,In_817,In_537);
nor U373 (N_373,In_1131,In_1151);
nand U374 (N_374,In_758,In_160);
and U375 (N_375,In_283,In_1335);
xnor U376 (N_376,In_1032,In_567);
nor U377 (N_377,In_708,In_1050);
or U378 (N_378,In_1047,In_1296);
nor U379 (N_379,In_1207,In_390);
and U380 (N_380,In_1465,In_586);
or U381 (N_381,In_674,In_194);
nor U382 (N_382,In_686,In_341);
and U383 (N_383,In_530,In_8);
xnor U384 (N_384,In_804,In_1168);
xor U385 (N_385,In_743,In_616);
nand U386 (N_386,In_237,In_844);
xnor U387 (N_387,In_261,In_290);
nor U388 (N_388,In_348,In_1087);
xnor U389 (N_389,In_598,In_993);
and U390 (N_390,In_1187,In_1241);
xnor U391 (N_391,In_17,In_1389);
nand U392 (N_392,In_465,In_146);
or U393 (N_393,In_215,In_840);
nor U394 (N_394,In_1108,In_297);
or U395 (N_395,In_884,In_612);
xor U396 (N_396,In_129,In_70);
nand U397 (N_397,In_574,In_1414);
nor U398 (N_398,In_269,In_1254);
nor U399 (N_399,In_150,In_304);
or U400 (N_400,In_681,In_190);
nor U401 (N_401,In_1166,In_81);
and U402 (N_402,In_1253,In_767);
nand U403 (N_403,In_318,In_195);
nand U404 (N_404,In_1445,In_372);
nand U405 (N_405,In_1096,In_1358);
nor U406 (N_406,In_1323,In_750);
nor U407 (N_407,In_887,In_106);
or U408 (N_408,In_1402,In_602);
nor U409 (N_409,In_579,In_668);
and U410 (N_410,In_1230,In_821);
nor U411 (N_411,In_1353,In_357);
xnor U412 (N_412,In_1326,In_95);
xnor U413 (N_413,In_188,In_894);
nand U414 (N_414,In_96,In_785);
xnor U415 (N_415,In_1357,In_88);
nor U416 (N_416,In_531,In_1063);
nand U417 (N_417,In_732,In_977);
xor U418 (N_418,In_420,In_227);
nor U419 (N_419,In_206,In_729);
nor U420 (N_420,In_1216,In_228);
nor U421 (N_421,In_517,In_1426);
nand U422 (N_422,In_519,In_60);
or U423 (N_423,In_59,In_2);
nor U424 (N_424,In_219,In_1307);
or U425 (N_425,In_608,In_1413);
nor U426 (N_426,In_1250,In_50);
nor U427 (N_427,In_330,In_1095);
and U428 (N_428,In_1074,In_1139);
and U429 (N_429,In_916,In_737);
nor U430 (N_430,In_539,In_1334);
or U431 (N_431,In_149,In_47);
or U432 (N_432,In_302,In_41);
and U433 (N_433,In_1481,In_857);
or U434 (N_434,In_1375,In_1155);
and U435 (N_435,In_1042,In_99);
nand U436 (N_436,In_1383,In_957);
nor U437 (N_437,In_471,In_1488);
nor U438 (N_438,In_763,In_941);
nor U439 (N_439,In_314,In_585);
or U440 (N_440,In_213,In_1038);
nor U441 (N_441,In_1156,In_379);
xnor U442 (N_442,In_137,In_570);
and U443 (N_443,In_533,In_656);
nand U444 (N_444,In_595,In_387);
or U445 (N_445,In_295,In_328);
xnor U446 (N_446,In_33,In_742);
or U447 (N_447,In_1382,In_862);
or U448 (N_448,In_1217,In_103);
or U449 (N_449,In_260,In_781);
and U450 (N_450,In_1396,In_908);
nand U451 (N_451,In_866,In_680);
nor U452 (N_452,In_658,In_983);
nor U453 (N_453,In_794,In_1211);
and U454 (N_454,In_896,In_875);
and U455 (N_455,In_641,In_577);
nor U456 (N_456,In_1336,In_526);
nor U457 (N_457,In_895,In_42);
or U458 (N_458,In_1343,In_1331);
xnor U459 (N_459,In_1416,In_966);
xnor U460 (N_460,In_502,In_637);
and U461 (N_461,In_1246,In_30);
nand U462 (N_462,In_145,In_1165);
nor U463 (N_463,In_1084,In_18);
or U464 (N_464,In_599,In_997);
nand U465 (N_465,In_833,In_1082);
or U466 (N_466,In_1310,In_1406);
or U467 (N_467,In_74,In_333);
and U468 (N_468,In_998,In_725);
xor U469 (N_469,In_1052,In_484);
and U470 (N_470,In_178,In_193);
nand U471 (N_471,In_62,In_507);
or U472 (N_472,In_1498,In_186);
nor U473 (N_473,In_967,In_643);
xor U474 (N_474,In_971,In_1478);
xor U475 (N_475,In_1483,In_405);
xor U476 (N_476,In_64,In_263);
xor U477 (N_477,In_168,In_1349);
nand U478 (N_478,In_210,In_1073);
nor U479 (N_479,In_299,In_510);
nand U480 (N_480,In_1030,In_683);
and U481 (N_481,In_813,In_250);
nand U482 (N_482,In_1069,In_1218);
and U483 (N_483,In_688,In_778);
nor U484 (N_484,In_786,In_1472);
xnor U485 (N_485,In_906,In_78);
nand U486 (N_486,In_427,In_776);
nand U487 (N_487,In_759,In_1297);
and U488 (N_488,In_1407,In_583);
xor U489 (N_489,In_1258,In_768);
nand U490 (N_490,In_820,In_1090);
and U491 (N_491,In_848,In_1227);
nand U492 (N_492,In_429,In_1200);
and U493 (N_493,In_435,In_1261);
nor U494 (N_494,In_978,In_406);
xor U495 (N_495,In_29,In_582);
or U496 (N_496,In_282,In_761);
or U497 (N_497,In_1226,In_1064);
and U498 (N_498,In_659,In_251);
and U499 (N_499,In_970,In_1431);
or U500 (N_500,In_655,In_229);
nand U501 (N_501,In_49,In_202);
or U502 (N_502,In_1141,In_562);
nor U503 (N_503,In_336,In_417);
nor U504 (N_504,In_1045,In_1438);
nand U505 (N_505,In_395,In_818);
and U506 (N_506,In_198,In_434);
and U507 (N_507,In_147,In_1283);
nor U508 (N_508,In_1317,In_506);
nor U509 (N_509,In_245,In_607);
or U510 (N_510,In_1225,In_837);
or U511 (N_511,In_847,In_855);
and U512 (N_512,In_1489,In_766);
or U513 (N_513,In_1208,In_1118);
nor U514 (N_514,In_75,In_1363);
nor U515 (N_515,In_371,In_1134);
or U516 (N_516,In_1016,In_928);
nand U517 (N_517,In_716,In_730);
nand U518 (N_518,In_963,In_396);
nor U519 (N_519,In_1356,In_67);
nand U520 (N_520,In_534,In_741);
and U521 (N_521,In_25,In_489);
nor U522 (N_522,In_1480,In_703);
xnor U523 (N_523,In_600,In_1322);
and U524 (N_524,In_1275,In_252);
xor U525 (N_525,In_827,In_112);
nor U526 (N_526,In_1452,In_823);
xnor U527 (N_527,In_1145,In_893);
or U528 (N_528,In_1212,In_617);
and U529 (N_529,In_511,In_1388);
and U530 (N_530,In_649,In_613);
and U531 (N_531,In_131,In_1021);
xnor U532 (N_532,In_345,In_126);
xnor U533 (N_533,In_652,In_899);
xnor U534 (N_534,In_407,In_1164);
and U535 (N_535,In_1315,In_1167);
nor U536 (N_536,In_929,In_94);
xnor U537 (N_537,In_267,In_1367);
and U538 (N_538,In_1461,In_581);
nand U539 (N_539,In_1193,In_594);
nand U540 (N_540,In_1201,In_442);
nand U541 (N_541,In_1373,In_1058);
nand U542 (N_542,In_253,In_508);
nand U543 (N_543,In_624,In_394);
and U544 (N_544,In_1485,In_376);
xnor U545 (N_545,In_964,In_709);
or U546 (N_546,In_1493,In_687);
nor U547 (N_547,In_359,In_355);
nand U548 (N_548,In_1234,In_885);
nor U549 (N_549,In_1186,In_1110);
nor U550 (N_550,In_418,In_448);
xor U551 (N_551,In_109,In_400);
nand U552 (N_552,In_313,In_457);
and U553 (N_553,In_1304,In_136);
nor U554 (N_554,In_412,In_1276);
or U555 (N_555,In_68,In_189);
nand U556 (N_556,In_754,In_1056);
nor U557 (N_557,In_504,In_535);
nand U558 (N_558,In_860,In_373);
nor U559 (N_559,In_832,In_1359);
xor U560 (N_560,In_513,In_1470);
xor U561 (N_561,In_350,In_73);
and U562 (N_562,In_163,In_701);
nor U563 (N_563,In_705,In_1405);
xor U564 (N_564,In_289,In_419);
and U565 (N_565,In_512,In_122);
nor U566 (N_566,In_1044,In_573);
nor U567 (N_567,In_1277,In_789);
or U568 (N_568,In_27,In_140);
nand U569 (N_569,In_291,In_1236);
nand U570 (N_570,In_1130,In_1463);
and U571 (N_571,In_1397,In_52);
xor U572 (N_572,In_733,In_277);
and U573 (N_573,In_1093,In_726);
or U574 (N_574,In_644,In_591);
or U575 (N_575,In_204,In_248);
nor U576 (N_576,In_1486,In_1157);
xor U577 (N_577,In_1440,In_475);
and U578 (N_578,In_1412,In_1459);
xnor U579 (N_579,In_757,In_859);
and U580 (N_580,In_578,In_831);
xor U581 (N_581,In_1293,In_470);
and U582 (N_582,In_727,In_951);
nor U583 (N_583,In_822,In_515);
nor U584 (N_584,In_514,In_1086);
nor U585 (N_585,In_469,In_666);
and U586 (N_586,In_555,In_811);
and U587 (N_587,In_161,In_16);
nor U588 (N_588,In_1469,In_477);
xor U589 (N_589,In_946,In_1365);
or U590 (N_590,In_1479,In_834);
xnor U591 (N_591,In_1158,In_116);
or U592 (N_592,In_346,In_441);
nor U593 (N_593,In_1059,In_486);
xnor U594 (N_594,In_491,In_601);
nand U595 (N_595,In_1173,In_667);
nand U596 (N_596,In_1106,In_485);
nor U597 (N_597,In_576,In_389);
or U598 (N_598,In_559,In_1027);
nor U599 (N_599,In_459,In_1377);
and U600 (N_600,In_693,In_1380);
xor U601 (N_601,In_982,In_292);
nand U602 (N_602,In_590,In_1179);
or U603 (N_603,In_529,In_51);
nand U604 (N_604,In_445,In_626);
nor U605 (N_605,In_141,In_509);
xnor U606 (N_606,In_1379,In_1496);
nand U607 (N_607,In_1181,In_1136);
or U608 (N_608,In_1381,In_220);
or U609 (N_609,In_764,In_710);
nand U610 (N_610,In_236,In_1305);
nor U611 (N_611,In_985,In_1324);
xnor U612 (N_612,In_1281,In_56);
or U613 (N_613,In_165,In_89);
or U614 (N_614,In_718,In_835);
or U615 (N_615,In_311,In_216);
nand U616 (N_616,In_1256,In_938);
xor U617 (N_617,In_980,In_1051);
or U618 (N_618,In_642,In_1111);
xnor U619 (N_619,In_118,In_1399);
xor U620 (N_620,In_321,In_97);
nand U621 (N_621,In_1213,In_802);
xnor U622 (N_622,In_132,In_1019);
or U623 (N_623,In_955,In_1279);
nor U624 (N_624,In_1400,In_503);
xor U625 (N_625,In_936,In_85);
xnor U626 (N_626,In_454,In_1455);
xor U627 (N_627,In_1004,In_347);
xnor U628 (N_628,In_809,In_1392);
or U629 (N_629,In_805,In_19);
nand U630 (N_630,In_784,In_919);
nor U631 (N_631,In_661,In_466);
or U632 (N_632,In_46,In_1366);
nand U633 (N_633,In_157,In_547);
or U634 (N_634,In_1332,In_1482);
xor U635 (N_635,In_1342,In_1494);
nand U636 (N_636,In_0,In_924);
xnor U637 (N_637,In_308,In_651);
nand U638 (N_638,In_898,In_1178);
nor U639 (N_639,In_1309,In_139);
and U640 (N_640,In_1175,In_31);
nor U641 (N_641,In_226,In_1026);
nor U642 (N_642,In_327,In_736);
xor U643 (N_643,In_1088,In_1146);
and U644 (N_644,In_1097,In_800);
nor U645 (N_645,In_1083,In_1476);
nor U646 (N_646,In_205,In_82);
nor U647 (N_647,In_231,In_1081);
or U648 (N_648,In_1424,In_913);
and U649 (N_649,In_1099,In_1313);
xor U650 (N_650,In_671,In_352);
nor U651 (N_651,In_1403,In_1031);
and U652 (N_652,In_1319,In_36);
and U653 (N_653,In_1135,In_925);
xor U654 (N_654,In_244,In_258);
and U655 (N_655,In_307,In_1328);
or U656 (N_656,In_255,In_284);
nor U657 (N_657,In_528,In_1018);
or U658 (N_658,In_281,In_79);
nand U659 (N_659,In_527,In_1177);
xnor U660 (N_660,In_1005,In_995);
or U661 (N_661,In_306,In_1009);
xnor U662 (N_662,In_478,In_1312);
nor U663 (N_663,In_807,In_39);
nor U664 (N_664,In_294,In_1378);
and U665 (N_665,In_1024,In_541);
xnor U666 (N_666,In_731,In_43);
nand U667 (N_667,In_1462,In_187);
nand U668 (N_668,In_755,In_1460);
and U669 (N_669,In_1000,In_1127);
nand U670 (N_670,In_838,In_954);
nand U671 (N_671,In_610,In_100);
and U672 (N_672,In_319,In_338);
nor U673 (N_673,In_1327,In_1189);
or U674 (N_674,In_54,In_184);
nor U675 (N_675,In_128,In_464);
nand U676 (N_676,In_546,In_603);
and U677 (N_677,In_1054,In_1251);
xnor U678 (N_678,In_55,In_1264);
xor U679 (N_679,In_66,In_864);
nor U680 (N_680,In_426,In_233);
and U681 (N_681,In_90,In_696);
or U682 (N_682,In_480,In_1129);
and U683 (N_683,In_1100,In_647);
nor U684 (N_684,In_1266,In_173);
xor U685 (N_685,In_1114,In_771);
nand U686 (N_686,In_856,In_1449);
xnor U687 (N_687,In_240,In_1467);
and U688 (N_688,In_217,In_1150);
xnor U689 (N_689,In_538,In_1473);
nand U690 (N_690,In_1192,In_167);
and U691 (N_691,In_646,In_700);
nand U692 (N_692,In_865,In_933);
or U693 (N_693,In_494,In_988);
xor U694 (N_694,In_324,In_1023);
or U695 (N_695,In_1034,In_698);
nor U696 (N_696,In_447,In_375);
and U697 (N_697,In_1033,In_1453);
nor U698 (N_698,In_1314,In_664);
nor U699 (N_699,In_648,In_540);
and U700 (N_700,In_676,In_197);
nor U701 (N_701,In_1089,In_1067);
or U702 (N_702,In_1384,In_1364);
and U703 (N_703,In_1068,In_858);
nand U704 (N_704,In_1183,In_1458);
and U705 (N_705,In_342,In_317);
and U706 (N_706,In_1020,In_1102);
or U707 (N_707,In_1049,In_77);
and U708 (N_708,In_207,In_222);
nor U709 (N_709,In_889,In_200);
nand U710 (N_710,In_1270,In_589);
nand U711 (N_711,In_849,In_1140);
nand U712 (N_712,In_892,In_153);
xor U713 (N_713,In_869,In_1361);
nand U714 (N_714,In_1456,In_958);
nor U715 (N_715,In_765,In_751);
or U716 (N_716,In_1341,In_382);
nand U717 (N_717,In_20,In_932);
nand U718 (N_718,In_1003,In_483);
or U719 (N_719,In_1,In_611);
nor U720 (N_720,In_1046,In_440);
nor U721 (N_721,In_543,In_1170);
and U722 (N_722,In_976,In_266);
and U723 (N_723,In_443,In_960);
or U724 (N_724,In_536,In_343);
or U725 (N_725,In_270,In_1078);
nand U726 (N_726,In_870,In_1228);
nor U727 (N_727,In_310,In_752);
nand U728 (N_728,In_619,In_773);
nor U729 (N_729,In_402,In_518);
xor U730 (N_730,In_797,In_1385);
xnor U731 (N_731,In_1352,In_1188);
xor U732 (N_732,In_1487,In_551);
nor U733 (N_733,In_1125,In_1223);
xor U734 (N_734,In_482,In_451);
and U735 (N_735,In_930,In_1417);
nor U736 (N_736,In_221,In_788);
nand U737 (N_737,In_272,In_1132);
nand U738 (N_738,In_1215,In_828);
nor U739 (N_739,In_1071,In_1010);
or U740 (N_740,In_358,In_704);
or U741 (N_741,In_1202,In_904);
nand U742 (N_742,In_554,In_1159);
nor U743 (N_743,In_21,In_351);
and U744 (N_744,In_1282,In_1447);
or U745 (N_745,In_130,In_86);
nand U746 (N_746,In_472,In_1142);
nand U747 (N_747,In_399,In_1104);
nand U748 (N_748,In_923,In_990);
and U749 (N_749,In_728,In_1206);
and U750 (N_750,In_962,In_311);
or U751 (N_751,In_1108,In_1236);
nor U752 (N_752,In_787,In_561);
and U753 (N_753,In_263,In_420);
nand U754 (N_754,In_634,In_1161);
and U755 (N_755,In_1418,In_50);
nand U756 (N_756,In_993,In_812);
nor U757 (N_757,In_662,In_1133);
nand U758 (N_758,In_714,In_72);
nor U759 (N_759,In_72,In_849);
or U760 (N_760,In_295,In_346);
xor U761 (N_761,In_820,In_932);
xnor U762 (N_762,In_673,In_867);
xnor U763 (N_763,In_406,In_120);
or U764 (N_764,In_1073,In_1267);
or U765 (N_765,In_568,In_1405);
nor U766 (N_766,In_458,In_900);
xor U767 (N_767,In_259,In_114);
xor U768 (N_768,In_1293,In_254);
nand U769 (N_769,In_1329,In_6);
xor U770 (N_770,In_402,In_1306);
nor U771 (N_771,In_571,In_168);
nor U772 (N_772,In_606,In_1244);
nand U773 (N_773,In_889,In_506);
and U774 (N_774,In_359,In_1212);
xnor U775 (N_775,In_787,In_809);
or U776 (N_776,In_501,In_578);
or U777 (N_777,In_549,In_808);
nand U778 (N_778,In_530,In_285);
nand U779 (N_779,In_644,In_114);
nor U780 (N_780,In_588,In_99);
and U781 (N_781,In_104,In_530);
xor U782 (N_782,In_493,In_643);
and U783 (N_783,In_997,In_1319);
and U784 (N_784,In_1036,In_1056);
nor U785 (N_785,In_43,In_502);
and U786 (N_786,In_722,In_852);
and U787 (N_787,In_314,In_1277);
and U788 (N_788,In_562,In_207);
nor U789 (N_789,In_1067,In_233);
xor U790 (N_790,In_502,In_658);
xnor U791 (N_791,In_311,In_512);
or U792 (N_792,In_756,In_552);
and U793 (N_793,In_912,In_43);
and U794 (N_794,In_1205,In_699);
nand U795 (N_795,In_934,In_911);
xnor U796 (N_796,In_847,In_1155);
nor U797 (N_797,In_240,In_774);
xor U798 (N_798,In_746,In_545);
or U799 (N_799,In_850,In_1129);
or U800 (N_800,In_791,In_1396);
nor U801 (N_801,In_648,In_670);
and U802 (N_802,In_555,In_1246);
nor U803 (N_803,In_533,In_635);
and U804 (N_804,In_58,In_1402);
nor U805 (N_805,In_1404,In_964);
xor U806 (N_806,In_73,In_967);
or U807 (N_807,In_387,In_410);
and U808 (N_808,In_892,In_742);
nor U809 (N_809,In_449,In_384);
xor U810 (N_810,In_611,In_1434);
and U811 (N_811,In_822,In_1335);
nor U812 (N_812,In_1438,In_432);
nor U813 (N_813,In_21,In_729);
nand U814 (N_814,In_803,In_603);
and U815 (N_815,In_473,In_522);
xor U816 (N_816,In_772,In_1263);
or U817 (N_817,In_932,In_1223);
nand U818 (N_818,In_348,In_466);
and U819 (N_819,In_585,In_406);
nand U820 (N_820,In_1489,In_530);
or U821 (N_821,In_907,In_222);
xnor U822 (N_822,In_941,In_979);
xor U823 (N_823,In_1210,In_1488);
nor U824 (N_824,In_1132,In_1372);
nor U825 (N_825,In_612,In_1260);
and U826 (N_826,In_1406,In_812);
nor U827 (N_827,In_117,In_563);
nand U828 (N_828,In_791,In_918);
nor U829 (N_829,In_586,In_419);
nand U830 (N_830,In_1348,In_1490);
nand U831 (N_831,In_762,In_86);
nand U832 (N_832,In_1242,In_959);
xor U833 (N_833,In_6,In_343);
nand U834 (N_834,In_801,In_38);
and U835 (N_835,In_837,In_764);
nor U836 (N_836,In_1346,In_1292);
xnor U837 (N_837,In_853,In_1087);
or U838 (N_838,In_1293,In_1428);
nor U839 (N_839,In_1282,In_228);
and U840 (N_840,In_641,In_1046);
xor U841 (N_841,In_361,In_39);
nor U842 (N_842,In_1168,In_1026);
and U843 (N_843,In_1039,In_64);
and U844 (N_844,In_167,In_96);
or U845 (N_845,In_1083,In_695);
xnor U846 (N_846,In_450,In_756);
nor U847 (N_847,In_608,In_1081);
and U848 (N_848,In_816,In_228);
nor U849 (N_849,In_450,In_497);
or U850 (N_850,In_1488,In_1261);
or U851 (N_851,In_1367,In_1064);
nand U852 (N_852,In_624,In_881);
xor U853 (N_853,In_1292,In_551);
xor U854 (N_854,In_959,In_625);
xnor U855 (N_855,In_1165,In_1239);
or U856 (N_856,In_422,In_1166);
and U857 (N_857,In_305,In_1426);
nor U858 (N_858,In_788,In_1191);
xor U859 (N_859,In_677,In_332);
nor U860 (N_860,In_957,In_721);
and U861 (N_861,In_354,In_1033);
xor U862 (N_862,In_772,In_480);
nor U863 (N_863,In_94,In_126);
nor U864 (N_864,In_983,In_180);
and U865 (N_865,In_956,In_50);
or U866 (N_866,In_1161,In_215);
xor U867 (N_867,In_1442,In_1214);
xor U868 (N_868,In_1212,In_1399);
xnor U869 (N_869,In_1105,In_1369);
nor U870 (N_870,In_463,In_1466);
or U871 (N_871,In_254,In_225);
nand U872 (N_872,In_1419,In_715);
nand U873 (N_873,In_1116,In_314);
or U874 (N_874,In_1475,In_1103);
or U875 (N_875,In_751,In_37);
and U876 (N_876,In_688,In_1194);
and U877 (N_877,In_388,In_518);
and U878 (N_878,In_361,In_404);
and U879 (N_879,In_634,In_686);
nand U880 (N_880,In_655,In_1331);
xor U881 (N_881,In_131,In_518);
and U882 (N_882,In_1042,In_1113);
nor U883 (N_883,In_1341,In_161);
and U884 (N_884,In_540,In_324);
nand U885 (N_885,In_692,In_781);
or U886 (N_886,In_443,In_392);
nor U887 (N_887,In_1275,In_6);
or U888 (N_888,In_1460,In_192);
nand U889 (N_889,In_955,In_1188);
xor U890 (N_890,In_1468,In_432);
and U891 (N_891,In_1464,In_573);
nand U892 (N_892,In_1082,In_1381);
or U893 (N_893,In_1454,In_644);
and U894 (N_894,In_485,In_1269);
nor U895 (N_895,In_1165,In_485);
nor U896 (N_896,In_1212,In_1113);
or U897 (N_897,In_652,In_85);
nor U898 (N_898,In_1427,In_545);
or U899 (N_899,In_1354,In_1431);
xor U900 (N_900,In_355,In_1492);
and U901 (N_901,In_194,In_1320);
nand U902 (N_902,In_165,In_1187);
nand U903 (N_903,In_119,In_1368);
xnor U904 (N_904,In_741,In_557);
nand U905 (N_905,In_848,In_679);
and U906 (N_906,In_1103,In_1317);
nand U907 (N_907,In_1404,In_1037);
xor U908 (N_908,In_344,In_401);
nand U909 (N_909,In_1010,In_41);
xnor U910 (N_910,In_1086,In_357);
nand U911 (N_911,In_912,In_170);
and U912 (N_912,In_568,In_1356);
xnor U913 (N_913,In_86,In_1060);
nand U914 (N_914,In_753,In_350);
nand U915 (N_915,In_1003,In_1163);
xor U916 (N_916,In_1390,In_226);
and U917 (N_917,In_938,In_269);
xnor U918 (N_918,In_111,In_1069);
xnor U919 (N_919,In_367,In_842);
nor U920 (N_920,In_983,In_1444);
and U921 (N_921,In_855,In_883);
or U922 (N_922,In_949,In_938);
nor U923 (N_923,In_1002,In_136);
nor U924 (N_924,In_1001,In_368);
or U925 (N_925,In_521,In_57);
or U926 (N_926,In_120,In_88);
xnor U927 (N_927,In_165,In_679);
xnor U928 (N_928,In_454,In_1171);
and U929 (N_929,In_1407,In_1337);
nand U930 (N_930,In_127,In_1290);
nor U931 (N_931,In_1395,In_668);
and U932 (N_932,In_847,In_322);
nor U933 (N_933,In_969,In_994);
xnor U934 (N_934,In_269,In_1246);
xor U935 (N_935,In_306,In_800);
and U936 (N_936,In_287,In_221);
nor U937 (N_937,In_21,In_1301);
and U938 (N_938,In_1065,In_1478);
and U939 (N_939,In_951,In_247);
xor U940 (N_940,In_537,In_69);
xor U941 (N_941,In_1373,In_548);
or U942 (N_942,In_280,In_0);
nor U943 (N_943,In_978,In_34);
nand U944 (N_944,In_658,In_1319);
nand U945 (N_945,In_703,In_1258);
nor U946 (N_946,In_777,In_1056);
or U947 (N_947,In_408,In_1455);
or U948 (N_948,In_155,In_773);
nor U949 (N_949,In_486,In_336);
or U950 (N_950,In_651,In_110);
and U951 (N_951,In_530,In_1313);
nor U952 (N_952,In_125,In_199);
nor U953 (N_953,In_169,In_842);
or U954 (N_954,In_1045,In_1439);
nand U955 (N_955,In_1242,In_487);
nor U956 (N_956,In_101,In_720);
nand U957 (N_957,In_314,In_1120);
and U958 (N_958,In_1240,In_478);
nor U959 (N_959,In_1207,In_788);
and U960 (N_960,In_1430,In_1454);
nand U961 (N_961,In_1113,In_1164);
and U962 (N_962,In_101,In_184);
nand U963 (N_963,In_1379,In_501);
nor U964 (N_964,In_413,In_239);
nand U965 (N_965,In_1446,In_186);
nor U966 (N_966,In_643,In_437);
nor U967 (N_967,In_1043,In_711);
and U968 (N_968,In_344,In_484);
and U969 (N_969,In_949,In_919);
xnor U970 (N_970,In_778,In_281);
or U971 (N_971,In_1078,In_375);
or U972 (N_972,In_546,In_413);
nand U973 (N_973,In_1125,In_850);
xor U974 (N_974,In_184,In_1203);
nor U975 (N_975,In_1300,In_529);
or U976 (N_976,In_712,In_1389);
or U977 (N_977,In_1487,In_849);
xor U978 (N_978,In_1190,In_882);
and U979 (N_979,In_765,In_340);
and U980 (N_980,In_933,In_482);
and U981 (N_981,In_66,In_217);
xnor U982 (N_982,In_661,In_1296);
nor U983 (N_983,In_1447,In_1050);
nand U984 (N_984,In_430,In_799);
nor U985 (N_985,In_1285,In_74);
xnor U986 (N_986,In_499,In_1499);
and U987 (N_987,In_1125,In_495);
xnor U988 (N_988,In_470,In_781);
or U989 (N_989,In_269,In_1158);
nand U990 (N_990,In_329,In_317);
nor U991 (N_991,In_1321,In_1364);
nor U992 (N_992,In_1398,In_877);
and U993 (N_993,In_543,In_1176);
nand U994 (N_994,In_765,In_30);
and U995 (N_995,In_1450,In_1354);
nand U996 (N_996,In_1084,In_159);
nand U997 (N_997,In_378,In_383);
nand U998 (N_998,In_640,In_1319);
nor U999 (N_999,In_681,In_13);
nor U1000 (N_1000,In_1064,In_613);
nand U1001 (N_1001,In_214,In_450);
or U1002 (N_1002,In_81,In_885);
or U1003 (N_1003,In_72,In_1288);
nor U1004 (N_1004,In_500,In_1402);
or U1005 (N_1005,In_1470,In_1443);
nand U1006 (N_1006,In_1029,In_1003);
nor U1007 (N_1007,In_1383,In_147);
and U1008 (N_1008,In_1190,In_209);
and U1009 (N_1009,In_1026,In_858);
nand U1010 (N_1010,In_1206,In_787);
nor U1011 (N_1011,In_378,In_1237);
nand U1012 (N_1012,In_871,In_245);
nand U1013 (N_1013,In_602,In_272);
nor U1014 (N_1014,In_474,In_970);
or U1015 (N_1015,In_424,In_1395);
and U1016 (N_1016,In_807,In_111);
or U1017 (N_1017,In_1368,In_685);
xor U1018 (N_1018,In_161,In_170);
nand U1019 (N_1019,In_101,In_1393);
xnor U1020 (N_1020,In_455,In_1438);
xor U1021 (N_1021,In_1334,In_1435);
and U1022 (N_1022,In_102,In_1396);
and U1023 (N_1023,In_181,In_93);
nand U1024 (N_1024,In_1073,In_53);
nor U1025 (N_1025,In_1353,In_545);
and U1026 (N_1026,In_966,In_760);
or U1027 (N_1027,In_1279,In_837);
nand U1028 (N_1028,In_891,In_1473);
and U1029 (N_1029,In_731,In_213);
and U1030 (N_1030,In_317,In_515);
nand U1031 (N_1031,In_1431,In_170);
and U1032 (N_1032,In_176,In_715);
nand U1033 (N_1033,In_345,In_35);
or U1034 (N_1034,In_351,In_1376);
and U1035 (N_1035,In_1,In_889);
xnor U1036 (N_1036,In_797,In_751);
or U1037 (N_1037,In_1209,In_1160);
nor U1038 (N_1038,In_484,In_131);
nor U1039 (N_1039,In_84,In_823);
nor U1040 (N_1040,In_284,In_1337);
and U1041 (N_1041,In_79,In_981);
xnor U1042 (N_1042,In_293,In_893);
and U1043 (N_1043,In_868,In_1067);
and U1044 (N_1044,In_174,In_1337);
xnor U1045 (N_1045,In_1459,In_1317);
and U1046 (N_1046,In_854,In_1436);
and U1047 (N_1047,In_19,In_943);
or U1048 (N_1048,In_883,In_842);
or U1049 (N_1049,In_601,In_777);
nand U1050 (N_1050,In_782,In_91);
xor U1051 (N_1051,In_393,In_1159);
xnor U1052 (N_1052,In_988,In_286);
nor U1053 (N_1053,In_137,In_370);
xor U1054 (N_1054,In_137,In_267);
nor U1055 (N_1055,In_125,In_122);
or U1056 (N_1056,In_235,In_788);
and U1057 (N_1057,In_1404,In_108);
nand U1058 (N_1058,In_1494,In_850);
or U1059 (N_1059,In_812,In_196);
nand U1060 (N_1060,In_1417,In_1192);
nand U1061 (N_1061,In_843,In_1473);
nand U1062 (N_1062,In_327,In_1044);
xor U1063 (N_1063,In_872,In_64);
nor U1064 (N_1064,In_1405,In_967);
nor U1065 (N_1065,In_917,In_1305);
or U1066 (N_1066,In_375,In_625);
nor U1067 (N_1067,In_8,In_867);
nor U1068 (N_1068,In_602,In_920);
xor U1069 (N_1069,In_1174,In_934);
nand U1070 (N_1070,In_161,In_993);
and U1071 (N_1071,In_569,In_1048);
or U1072 (N_1072,In_850,In_928);
or U1073 (N_1073,In_1360,In_682);
or U1074 (N_1074,In_1057,In_379);
and U1075 (N_1075,In_1405,In_349);
or U1076 (N_1076,In_32,In_291);
nor U1077 (N_1077,In_15,In_398);
and U1078 (N_1078,In_781,In_938);
nor U1079 (N_1079,In_662,In_1151);
and U1080 (N_1080,In_527,In_1309);
or U1081 (N_1081,In_685,In_557);
xor U1082 (N_1082,In_765,In_301);
nand U1083 (N_1083,In_1359,In_1333);
or U1084 (N_1084,In_104,In_1007);
nor U1085 (N_1085,In_42,In_541);
or U1086 (N_1086,In_856,In_367);
nor U1087 (N_1087,In_300,In_793);
nand U1088 (N_1088,In_993,In_539);
or U1089 (N_1089,In_346,In_1498);
and U1090 (N_1090,In_593,In_1461);
xor U1091 (N_1091,In_319,In_1035);
xnor U1092 (N_1092,In_557,In_622);
nand U1093 (N_1093,In_951,In_763);
nor U1094 (N_1094,In_462,In_269);
and U1095 (N_1095,In_478,In_167);
xnor U1096 (N_1096,In_323,In_1476);
xor U1097 (N_1097,In_1148,In_308);
or U1098 (N_1098,In_595,In_1442);
or U1099 (N_1099,In_724,In_1413);
or U1100 (N_1100,In_1361,In_503);
and U1101 (N_1101,In_1329,In_720);
nor U1102 (N_1102,In_697,In_89);
nand U1103 (N_1103,In_136,In_215);
or U1104 (N_1104,In_1091,In_1295);
xnor U1105 (N_1105,In_927,In_1217);
and U1106 (N_1106,In_787,In_336);
or U1107 (N_1107,In_14,In_11);
nand U1108 (N_1108,In_389,In_276);
or U1109 (N_1109,In_26,In_1216);
nand U1110 (N_1110,In_643,In_1000);
xor U1111 (N_1111,In_589,In_1353);
xor U1112 (N_1112,In_1027,In_1349);
nand U1113 (N_1113,In_788,In_1438);
or U1114 (N_1114,In_473,In_486);
nor U1115 (N_1115,In_32,In_1441);
nand U1116 (N_1116,In_457,In_1440);
or U1117 (N_1117,In_1175,In_836);
nand U1118 (N_1118,In_324,In_664);
or U1119 (N_1119,In_601,In_1150);
or U1120 (N_1120,In_42,In_740);
xor U1121 (N_1121,In_903,In_843);
xnor U1122 (N_1122,In_682,In_826);
nor U1123 (N_1123,In_879,In_100);
xor U1124 (N_1124,In_503,In_1272);
nand U1125 (N_1125,In_63,In_1013);
and U1126 (N_1126,In_552,In_1097);
nand U1127 (N_1127,In_1457,In_1357);
xor U1128 (N_1128,In_1259,In_401);
nor U1129 (N_1129,In_232,In_571);
nor U1130 (N_1130,In_30,In_617);
or U1131 (N_1131,In_843,In_250);
and U1132 (N_1132,In_759,In_540);
nand U1133 (N_1133,In_1250,In_64);
nor U1134 (N_1134,In_716,In_913);
or U1135 (N_1135,In_104,In_1311);
xnor U1136 (N_1136,In_1277,In_1142);
nand U1137 (N_1137,In_849,In_1117);
nand U1138 (N_1138,In_178,In_378);
nand U1139 (N_1139,In_966,In_1378);
or U1140 (N_1140,In_583,In_902);
nand U1141 (N_1141,In_403,In_986);
nor U1142 (N_1142,In_237,In_1175);
and U1143 (N_1143,In_686,In_575);
or U1144 (N_1144,In_674,In_1064);
xnor U1145 (N_1145,In_239,In_332);
xnor U1146 (N_1146,In_1100,In_1237);
or U1147 (N_1147,In_1118,In_910);
and U1148 (N_1148,In_1060,In_147);
or U1149 (N_1149,In_1303,In_1050);
nor U1150 (N_1150,In_705,In_715);
and U1151 (N_1151,In_705,In_1253);
or U1152 (N_1152,In_54,In_461);
nor U1153 (N_1153,In_551,In_294);
nand U1154 (N_1154,In_1116,In_1192);
nor U1155 (N_1155,In_1148,In_1144);
or U1156 (N_1156,In_1,In_697);
or U1157 (N_1157,In_569,In_602);
nand U1158 (N_1158,In_304,In_522);
or U1159 (N_1159,In_656,In_1448);
nand U1160 (N_1160,In_708,In_799);
and U1161 (N_1161,In_1243,In_69);
nor U1162 (N_1162,In_30,In_41);
or U1163 (N_1163,In_301,In_1380);
nand U1164 (N_1164,In_1313,In_1135);
and U1165 (N_1165,In_711,In_1049);
nand U1166 (N_1166,In_95,In_685);
and U1167 (N_1167,In_1299,In_73);
and U1168 (N_1168,In_510,In_249);
nand U1169 (N_1169,In_1489,In_1040);
and U1170 (N_1170,In_983,In_847);
xnor U1171 (N_1171,In_1127,In_1092);
xnor U1172 (N_1172,In_182,In_723);
or U1173 (N_1173,In_438,In_1104);
xnor U1174 (N_1174,In_338,In_160);
and U1175 (N_1175,In_1306,In_1178);
nand U1176 (N_1176,In_1178,In_234);
xor U1177 (N_1177,In_697,In_437);
xnor U1178 (N_1178,In_734,In_751);
xnor U1179 (N_1179,In_743,In_309);
or U1180 (N_1180,In_539,In_349);
nor U1181 (N_1181,In_941,In_510);
xor U1182 (N_1182,In_75,In_1027);
or U1183 (N_1183,In_712,In_873);
nor U1184 (N_1184,In_1046,In_1382);
nor U1185 (N_1185,In_1247,In_7);
and U1186 (N_1186,In_51,In_920);
or U1187 (N_1187,In_615,In_102);
xor U1188 (N_1188,In_1059,In_183);
or U1189 (N_1189,In_1418,In_140);
nor U1190 (N_1190,In_1390,In_652);
nor U1191 (N_1191,In_1013,In_872);
xnor U1192 (N_1192,In_207,In_62);
and U1193 (N_1193,In_835,In_1474);
and U1194 (N_1194,In_736,In_1322);
nand U1195 (N_1195,In_133,In_641);
nand U1196 (N_1196,In_1158,In_1152);
and U1197 (N_1197,In_1332,In_1132);
nor U1198 (N_1198,In_141,In_1474);
or U1199 (N_1199,In_1490,In_294);
nand U1200 (N_1200,In_958,In_721);
nor U1201 (N_1201,In_1233,In_207);
or U1202 (N_1202,In_684,In_1281);
nor U1203 (N_1203,In_1141,In_341);
nand U1204 (N_1204,In_917,In_929);
and U1205 (N_1205,In_640,In_829);
nand U1206 (N_1206,In_1084,In_777);
and U1207 (N_1207,In_136,In_635);
or U1208 (N_1208,In_1426,In_678);
or U1209 (N_1209,In_1068,In_593);
or U1210 (N_1210,In_1045,In_762);
nor U1211 (N_1211,In_412,In_1347);
or U1212 (N_1212,In_635,In_929);
nor U1213 (N_1213,In_1276,In_1193);
nor U1214 (N_1214,In_981,In_1447);
nor U1215 (N_1215,In_427,In_449);
nand U1216 (N_1216,In_481,In_154);
nand U1217 (N_1217,In_703,In_1290);
xnor U1218 (N_1218,In_739,In_939);
nor U1219 (N_1219,In_404,In_1224);
nor U1220 (N_1220,In_1212,In_1265);
and U1221 (N_1221,In_783,In_555);
or U1222 (N_1222,In_430,In_1462);
nor U1223 (N_1223,In_200,In_65);
nor U1224 (N_1224,In_949,In_804);
or U1225 (N_1225,In_1089,In_877);
xnor U1226 (N_1226,In_1421,In_135);
and U1227 (N_1227,In_1150,In_210);
nand U1228 (N_1228,In_740,In_747);
nor U1229 (N_1229,In_1416,In_619);
nand U1230 (N_1230,In_715,In_1182);
xnor U1231 (N_1231,In_512,In_644);
nand U1232 (N_1232,In_1232,In_1251);
or U1233 (N_1233,In_1276,In_1489);
or U1234 (N_1234,In_72,In_899);
nor U1235 (N_1235,In_1464,In_1114);
or U1236 (N_1236,In_1216,In_808);
or U1237 (N_1237,In_1030,In_1087);
and U1238 (N_1238,In_237,In_236);
nor U1239 (N_1239,In_920,In_1396);
nand U1240 (N_1240,In_262,In_53);
and U1241 (N_1241,In_1143,In_1236);
or U1242 (N_1242,In_880,In_22);
and U1243 (N_1243,In_990,In_1003);
nand U1244 (N_1244,In_665,In_578);
nand U1245 (N_1245,In_1029,In_215);
and U1246 (N_1246,In_867,In_55);
nand U1247 (N_1247,In_850,In_483);
and U1248 (N_1248,In_945,In_1416);
xnor U1249 (N_1249,In_1273,In_692);
nand U1250 (N_1250,In_739,In_517);
or U1251 (N_1251,In_1014,In_1345);
nor U1252 (N_1252,In_1279,In_747);
nor U1253 (N_1253,In_1026,In_1474);
nand U1254 (N_1254,In_930,In_387);
and U1255 (N_1255,In_672,In_1056);
and U1256 (N_1256,In_541,In_1328);
or U1257 (N_1257,In_625,In_716);
nand U1258 (N_1258,In_55,In_553);
nand U1259 (N_1259,In_231,In_605);
nor U1260 (N_1260,In_1260,In_970);
nor U1261 (N_1261,In_824,In_842);
and U1262 (N_1262,In_53,In_152);
xor U1263 (N_1263,In_905,In_592);
and U1264 (N_1264,In_104,In_404);
xor U1265 (N_1265,In_685,In_137);
or U1266 (N_1266,In_701,In_391);
and U1267 (N_1267,In_918,In_790);
and U1268 (N_1268,In_460,In_423);
nor U1269 (N_1269,In_1426,In_1163);
nor U1270 (N_1270,In_221,In_46);
and U1271 (N_1271,In_1227,In_1043);
nor U1272 (N_1272,In_434,In_1473);
nand U1273 (N_1273,In_313,In_1002);
and U1274 (N_1274,In_1152,In_163);
or U1275 (N_1275,In_1443,In_385);
nor U1276 (N_1276,In_38,In_762);
or U1277 (N_1277,In_651,In_1063);
xnor U1278 (N_1278,In_1142,In_1149);
and U1279 (N_1279,In_1067,In_766);
or U1280 (N_1280,In_1125,In_1376);
nor U1281 (N_1281,In_1350,In_1493);
and U1282 (N_1282,In_239,In_713);
or U1283 (N_1283,In_845,In_127);
nor U1284 (N_1284,In_1362,In_430);
and U1285 (N_1285,In_121,In_663);
xnor U1286 (N_1286,In_1061,In_490);
or U1287 (N_1287,In_575,In_1121);
and U1288 (N_1288,In_1142,In_148);
or U1289 (N_1289,In_1069,In_931);
nor U1290 (N_1290,In_438,In_874);
nand U1291 (N_1291,In_207,In_841);
xnor U1292 (N_1292,In_268,In_1397);
and U1293 (N_1293,In_922,In_608);
nand U1294 (N_1294,In_345,In_1193);
or U1295 (N_1295,In_788,In_256);
nor U1296 (N_1296,In_675,In_640);
and U1297 (N_1297,In_163,In_72);
nand U1298 (N_1298,In_736,In_1386);
xnor U1299 (N_1299,In_679,In_554);
xor U1300 (N_1300,In_925,In_939);
nand U1301 (N_1301,In_1010,In_832);
or U1302 (N_1302,In_1077,In_1296);
nand U1303 (N_1303,In_829,In_1142);
nand U1304 (N_1304,In_95,In_954);
and U1305 (N_1305,In_40,In_200);
and U1306 (N_1306,In_243,In_197);
or U1307 (N_1307,In_550,In_1335);
or U1308 (N_1308,In_505,In_1444);
or U1309 (N_1309,In_1086,In_438);
nor U1310 (N_1310,In_33,In_681);
nor U1311 (N_1311,In_532,In_881);
or U1312 (N_1312,In_1058,In_1431);
or U1313 (N_1313,In_101,In_674);
nand U1314 (N_1314,In_1069,In_590);
xor U1315 (N_1315,In_820,In_1387);
nand U1316 (N_1316,In_1337,In_136);
nor U1317 (N_1317,In_343,In_702);
and U1318 (N_1318,In_1431,In_139);
nor U1319 (N_1319,In_708,In_346);
xnor U1320 (N_1320,In_765,In_814);
nor U1321 (N_1321,In_1360,In_31);
nor U1322 (N_1322,In_139,In_285);
xor U1323 (N_1323,In_1138,In_291);
xnor U1324 (N_1324,In_331,In_554);
and U1325 (N_1325,In_1190,In_526);
or U1326 (N_1326,In_434,In_436);
or U1327 (N_1327,In_553,In_1081);
xor U1328 (N_1328,In_425,In_447);
xor U1329 (N_1329,In_1096,In_161);
nor U1330 (N_1330,In_723,In_679);
and U1331 (N_1331,In_676,In_64);
nand U1332 (N_1332,In_788,In_587);
xor U1333 (N_1333,In_539,In_930);
or U1334 (N_1334,In_388,In_443);
nand U1335 (N_1335,In_1149,In_1460);
nor U1336 (N_1336,In_269,In_1365);
nand U1337 (N_1337,In_1252,In_1438);
nor U1338 (N_1338,In_663,In_720);
and U1339 (N_1339,In_158,In_250);
xor U1340 (N_1340,In_1355,In_1446);
nand U1341 (N_1341,In_908,In_784);
nor U1342 (N_1342,In_189,In_620);
nand U1343 (N_1343,In_1155,In_700);
or U1344 (N_1344,In_56,In_348);
or U1345 (N_1345,In_1406,In_426);
and U1346 (N_1346,In_601,In_1498);
xnor U1347 (N_1347,In_1305,In_691);
or U1348 (N_1348,In_1146,In_1487);
and U1349 (N_1349,In_106,In_559);
nor U1350 (N_1350,In_1416,In_931);
xnor U1351 (N_1351,In_560,In_663);
and U1352 (N_1352,In_1147,In_1195);
nor U1353 (N_1353,In_784,In_1050);
and U1354 (N_1354,In_445,In_1080);
xor U1355 (N_1355,In_415,In_1424);
nand U1356 (N_1356,In_778,In_982);
nand U1357 (N_1357,In_481,In_1436);
nor U1358 (N_1358,In_865,In_432);
nand U1359 (N_1359,In_1374,In_1095);
nor U1360 (N_1360,In_90,In_989);
xnor U1361 (N_1361,In_559,In_950);
and U1362 (N_1362,In_17,In_100);
or U1363 (N_1363,In_1318,In_1432);
xor U1364 (N_1364,In_4,In_684);
and U1365 (N_1365,In_628,In_1143);
nor U1366 (N_1366,In_553,In_1103);
and U1367 (N_1367,In_530,In_522);
nor U1368 (N_1368,In_1300,In_832);
nand U1369 (N_1369,In_163,In_834);
nor U1370 (N_1370,In_892,In_958);
nand U1371 (N_1371,In_1257,In_682);
xnor U1372 (N_1372,In_33,In_1237);
xor U1373 (N_1373,In_970,In_273);
or U1374 (N_1374,In_26,In_106);
and U1375 (N_1375,In_252,In_431);
or U1376 (N_1376,In_1336,In_22);
nand U1377 (N_1377,In_1350,In_142);
xnor U1378 (N_1378,In_1132,In_882);
nand U1379 (N_1379,In_314,In_546);
xor U1380 (N_1380,In_4,In_1112);
or U1381 (N_1381,In_181,In_41);
xor U1382 (N_1382,In_597,In_36);
nor U1383 (N_1383,In_1372,In_1428);
or U1384 (N_1384,In_1480,In_481);
and U1385 (N_1385,In_1049,In_1117);
nand U1386 (N_1386,In_380,In_432);
and U1387 (N_1387,In_963,In_489);
or U1388 (N_1388,In_368,In_225);
or U1389 (N_1389,In_953,In_854);
nand U1390 (N_1390,In_1367,In_272);
and U1391 (N_1391,In_895,In_1125);
nand U1392 (N_1392,In_511,In_458);
nor U1393 (N_1393,In_218,In_1176);
xor U1394 (N_1394,In_668,In_1104);
and U1395 (N_1395,In_1477,In_575);
nor U1396 (N_1396,In_1205,In_644);
xnor U1397 (N_1397,In_646,In_909);
nor U1398 (N_1398,In_1372,In_288);
nor U1399 (N_1399,In_129,In_528);
nor U1400 (N_1400,In_882,In_475);
nor U1401 (N_1401,In_1070,In_1274);
nor U1402 (N_1402,In_1120,In_957);
xnor U1403 (N_1403,In_1273,In_1262);
nand U1404 (N_1404,In_386,In_1284);
nor U1405 (N_1405,In_1070,In_576);
and U1406 (N_1406,In_134,In_1476);
or U1407 (N_1407,In_1469,In_1363);
nor U1408 (N_1408,In_1201,In_288);
nor U1409 (N_1409,In_1154,In_1349);
nor U1410 (N_1410,In_172,In_840);
and U1411 (N_1411,In_1498,In_86);
xnor U1412 (N_1412,In_1234,In_74);
and U1413 (N_1413,In_327,In_739);
xor U1414 (N_1414,In_468,In_1083);
nor U1415 (N_1415,In_1091,In_1082);
or U1416 (N_1416,In_17,In_732);
or U1417 (N_1417,In_610,In_1150);
nand U1418 (N_1418,In_643,In_1306);
nor U1419 (N_1419,In_1291,In_1455);
xnor U1420 (N_1420,In_504,In_664);
nor U1421 (N_1421,In_1055,In_130);
and U1422 (N_1422,In_956,In_703);
and U1423 (N_1423,In_765,In_496);
xnor U1424 (N_1424,In_228,In_310);
nor U1425 (N_1425,In_1461,In_665);
nor U1426 (N_1426,In_319,In_622);
and U1427 (N_1427,In_145,In_1132);
nand U1428 (N_1428,In_1482,In_57);
or U1429 (N_1429,In_340,In_698);
nor U1430 (N_1430,In_875,In_993);
nor U1431 (N_1431,In_361,In_1239);
and U1432 (N_1432,In_946,In_445);
and U1433 (N_1433,In_475,In_637);
or U1434 (N_1434,In_688,In_1412);
xnor U1435 (N_1435,In_500,In_760);
and U1436 (N_1436,In_563,In_1275);
nor U1437 (N_1437,In_1456,In_730);
or U1438 (N_1438,In_1417,In_382);
and U1439 (N_1439,In_1054,In_75);
nor U1440 (N_1440,In_1072,In_983);
nor U1441 (N_1441,In_779,In_1044);
xor U1442 (N_1442,In_441,In_736);
or U1443 (N_1443,In_1451,In_1084);
nand U1444 (N_1444,In_568,In_1026);
xnor U1445 (N_1445,In_577,In_451);
or U1446 (N_1446,In_509,In_427);
xor U1447 (N_1447,In_1445,In_1226);
xnor U1448 (N_1448,In_1050,In_854);
and U1449 (N_1449,In_1086,In_1457);
xnor U1450 (N_1450,In_128,In_716);
and U1451 (N_1451,In_73,In_974);
and U1452 (N_1452,In_258,In_828);
nor U1453 (N_1453,In_513,In_1179);
nor U1454 (N_1454,In_1336,In_382);
and U1455 (N_1455,In_137,In_1321);
nor U1456 (N_1456,In_208,In_145);
and U1457 (N_1457,In_812,In_143);
nor U1458 (N_1458,In_820,In_65);
nand U1459 (N_1459,In_526,In_558);
and U1460 (N_1460,In_636,In_50);
nor U1461 (N_1461,In_392,In_833);
nand U1462 (N_1462,In_98,In_248);
nor U1463 (N_1463,In_1132,In_1131);
or U1464 (N_1464,In_145,In_735);
nand U1465 (N_1465,In_667,In_560);
nand U1466 (N_1466,In_1285,In_714);
or U1467 (N_1467,In_1128,In_341);
or U1468 (N_1468,In_888,In_901);
and U1469 (N_1469,In_652,In_191);
nor U1470 (N_1470,In_1481,In_904);
xor U1471 (N_1471,In_1059,In_426);
nand U1472 (N_1472,In_1097,In_144);
nand U1473 (N_1473,In_244,In_548);
xor U1474 (N_1474,In_936,In_1496);
xor U1475 (N_1475,In_1067,In_186);
xnor U1476 (N_1476,In_1435,In_695);
or U1477 (N_1477,In_1407,In_988);
xnor U1478 (N_1478,In_1250,In_15);
nand U1479 (N_1479,In_245,In_792);
or U1480 (N_1480,In_975,In_1461);
or U1481 (N_1481,In_300,In_650);
xnor U1482 (N_1482,In_450,In_1168);
nand U1483 (N_1483,In_278,In_386);
nor U1484 (N_1484,In_282,In_693);
xor U1485 (N_1485,In_1139,In_1481);
nor U1486 (N_1486,In_1367,In_1390);
or U1487 (N_1487,In_460,In_303);
nor U1488 (N_1488,In_200,In_538);
nand U1489 (N_1489,In_186,In_669);
or U1490 (N_1490,In_1233,In_1081);
xnor U1491 (N_1491,In_1095,In_1480);
nand U1492 (N_1492,In_935,In_614);
or U1493 (N_1493,In_583,In_711);
nand U1494 (N_1494,In_734,In_1304);
and U1495 (N_1495,In_1340,In_1040);
nand U1496 (N_1496,In_387,In_601);
xor U1497 (N_1497,In_277,In_784);
and U1498 (N_1498,In_580,In_965);
or U1499 (N_1499,In_159,In_1100);
or U1500 (N_1500,In_909,In_732);
nor U1501 (N_1501,In_761,In_626);
xnor U1502 (N_1502,In_712,In_219);
xnor U1503 (N_1503,In_832,In_499);
xnor U1504 (N_1504,In_327,In_1057);
and U1505 (N_1505,In_630,In_157);
nand U1506 (N_1506,In_916,In_428);
nand U1507 (N_1507,In_766,In_851);
or U1508 (N_1508,In_854,In_1153);
and U1509 (N_1509,In_978,In_768);
nand U1510 (N_1510,In_1461,In_323);
xor U1511 (N_1511,In_1237,In_1358);
or U1512 (N_1512,In_284,In_1212);
or U1513 (N_1513,In_1475,In_604);
and U1514 (N_1514,In_957,In_1034);
xnor U1515 (N_1515,In_1062,In_979);
xnor U1516 (N_1516,In_404,In_819);
nand U1517 (N_1517,In_1225,In_778);
and U1518 (N_1518,In_1007,In_625);
nor U1519 (N_1519,In_245,In_415);
nor U1520 (N_1520,In_1449,In_1388);
nor U1521 (N_1521,In_721,In_221);
nand U1522 (N_1522,In_1195,In_14);
or U1523 (N_1523,In_406,In_39);
nand U1524 (N_1524,In_447,In_74);
or U1525 (N_1525,In_1287,In_921);
nor U1526 (N_1526,In_517,In_1367);
nand U1527 (N_1527,In_574,In_1286);
nor U1528 (N_1528,In_1337,In_441);
nand U1529 (N_1529,In_1012,In_1434);
nand U1530 (N_1530,In_484,In_1209);
nor U1531 (N_1531,In_976,In_1400);
nor U1532 (N_1532,In_1450,In_891);
nand U1533 (N_1533,In_991,In_1403);
or U1534 (N_1534,In_640,In_1120);
nand U1535 (N_1535,In_1165,In_1244);
or U1536 (N_1536,In_308,In_377);
and U1537 (N_1537,In_4,In_198);
nor U1538 (N_1538,In_179,In_1496);
nand U1539 (N_1539,In_1457,In_1042);
and U1540 (N_1540,In_1427,In_76);
nor U1541 (N_1541,In_996,In_341);
or U1542 (N_1542,In_1413,In_417);
xor U1543 (N_1543,In_660,In_697);
xor U1544 (N_1544,In_1413,In_115);
and U1545 (N_1545,In_1212,In_1228);
nand U1546 (N_1546,In_719,In_900);
and U1547 (N_1547,In_1335,In_1488);
or U1548 (N_1548,In_900,In_309);
nand U1549 (N_1549,In_1435,In_565);
nand U1550 (N_1550,In_792,In_280);
nand U1551 (N_1551,In_1095,In_157);
or U1552 (N_1552,In_682,In_1266);
and U1553 (N_1553,In_259,In_1249);
xnor U1554 (N_1554,In_1350,In_507);
nor U1555 (N_1555,In_529,In_118);
and U1556 (N_1556,In_1478,In_1356);
and U1557 (N_1557,In_850,In_252);
and U1558 (N_1558,In_615,In_623);
and U1559 (N_1559,In_1475,In_94);
or U1560 (N_1560,In_1037,In_732);
xor U1561 (N_1561,In_1107,In_118);
xnor U1562 (N_1562,In_1179,In_1474);
nor U1563 (N_1563,In_1039,In_750);
and U1564 (N_1564,In_642,In_1228);
and U1565 (N_1565,In_1475,In_1307);
nor U1566 (N_1566,In_156,In_367);
or U1567 (N_1567,In_724,In_970);
xor U1568 (N_1568,In_84,In_1307);
nor U1569 (N_1569,In_807,In_1268);
xnor U1570 (N_1570,In_276,In_1457);
nand U1571 (N_1571,In_277,In_1345);
or U1572 (N_1572,In_483,In_32);
xnor U1573 (N_1573,In_1107,In_1205);
or U1574 (N_1574,In_74,In_1273);
nand U1575 (N_1575,In_1442,In_1124);
xor U1576 (N_1576,In_922,In_1103);
and U1577 (N_1577,In_761,In_630);
and U1578 (N_1578,In_1355,In_424);
nor U1579 (N_1579,In_262,In_66);
nand U1580 (N_1580,In_743,In_851);
or U1581 (N_1581,In_275,In_1422);
nor U1582 (N_1582,In_157,In_475);
or U1583 (N_1583,In_1277,In_59);
and U1584 (N_1584,In_363,In_87);
nor U1585 (N_1585,In_1389,In_61);
or U1586 (N_1586,In_1381,In_868);
xor U1587 (N_1587,In_1047,In_1474);
nand U1588 (N_1588,In_608,In_460);
nand U1589 (N_1589,In_978,In_333);
and U1590 (N_1590,In_1010,In_457);
or U1591 (N_1591,In_529,In_141);
nor U1592 (N_1592,In_1430,In_242);
nand U1593 (N_1593,In_1014,In_49);
xor U1594 (N_1594,In_1023,In_1048);
xnor U1595 (N_1595,In_1059,In_1382);
nor U1596 (N_1596,In_1300,In_1169);
nor U1597 (N_1597,In_800,In_1142);
and U1598 (N_1598,In_925,In_760);
nand U1599 (N_1599,In_1374,In_1002);
and U1600 (N_1600,In_1246,In_1172);
or U1601 (N_1601,In_580,In_1467);
nor U1602 (N_1602,In_375,In_468);
or U1603 (N_1603,In_1283,In_800);
nand U1604 (N_1604,In_1035,In_1121);
and U1605 (N_1605,In_547,In_611);
or U1606 (N_1606,In_1350,In_1393);
nand U1607 (N_1607,In_1205,In_1473);
nand U1608 (N_1608,In_331,In_679);
and U1609 (N_1609,In_1081,In_424);
xor U1610 (N_1610,In_807,In_1264);
and U1611 (N_1611,In_1110,In_883);
nor U1612 (N_1612,In_519,In_1456);
and U1613 (N_1613,In_1146,In_1207);
xnor U1614 (N_1614,In_1403,In_899);
nand U1615 (N_1615,In_1301,In_480);
nor U1616 (N_1616,In_578,In_900);
or U1617 (N_1617,In_825,In_1244);
and U1618 (N_1618,In_1098,In_379);
nand U1619 (N_1619,In_967,In_137);
and U1620 (N_1620,In_1183,In_1065);
or U1621 (N_1621,In_904,In_38);
nand U1622 (N_1622,In_956,In_814);
nor U1623 (N_1623,In_496,In_1417);
nand U1624 (N_1624,In_1361,In_1357);
xor U1625 (N_1625,In_1380,In_513);
nor U1626 (N_1626,In_14,In_944);
nand U1627 (N_1627,In_562,In_581);
and U1628 (N_1628,In_1092,In_1097);
nor U1629 (N_1629,In_915,In_348);
nor U1630 (N_1630,In_1355,In_81);
and U1631 (N_1631,In_823,In_1197);
and U1632 (N_1632,In_511,In_112);
and U1633 (N_1633,In_708,In_219);
xnor U1634 (N_1634,In_110,In_494);
or U1635 (N_1635,In_132,In_877);
nor U1636 (N_1636,In_795,In_1269);
nor U1637 (N_1637,In_1308,In_637);
xnor U1638 (N_1638,In_102,In_200);
nand U1639 (N_1639,In_1097,In_499);
xor U1640 (N_1640,In_692,In_540);
xor U1641 (N_1641,In_1157,In_57);
xor U1642 (N_1642,In_345,In_93);
xnor U1643 (N_1643,In_1327,In_299);
nor U1644 (N_1644,In_787,In_611);
and U1645 (N_1645,In_1294,In_1385);
xor U1646 (N_1646,In_1206,In_1119);
xor U1647 (N_1647,In_667,In_435);
and U1648 (N_1648,In_1462,In_727);
or U1649 (N_1649,In_647,In_630);
and U1650 (N_1650,In_109,In_1036);
and U1651 (N_1651,In_684,In_1125);
xor U1652 (N_1652,In_1422,In_362);
xor U1653 (N_1653,In_1493,In_503);
xor U1654 (N_1654,In_1206,In_353);
and U1655 (N_1655,In_1478,In_1072);
or U1656 (N_1656,In_397,In_351);
nor U1657 (N_1657,In_1074,In_774);
nand U1658 (N_1658,In_266,In_259);
or U1659 (N_1659,In_389,In_1349);
nand U1660 (N_1660,In_1452,In_489);
or U1661 (N_1661,In_342,In_1006);
nand U1662 (N_1662,In_1046,In_249);
xor U1663 (N_1663,In_621,In_554);
nand U1664 (N_1664,In_643,In_1244);
xor U1665 (N_1665,In_1102,In_1479);
nand U1666 (N_1666,In_1124,In_165);
nor U1667 (N_1667,In_1339,In_427);
or U1668 (N_1668,In_910,In_817);
nand U1669 (N_1669,In_1116,In_1265);
xnor U1670 (N_1670,In_651,In_520);
xnor U1671 (N_1671,In_837,In_300);
or U1672 (N_1672,In_939,In_355);
xnor U1673 (N_1673,In_1314,In_985);
and U1674 (N_1674,In_101,In_1273);
xnor U1675 (N_1675,In_1229,In_1407);
nor U1676 (N_1676,In_174,In_375);
xor U1677 (N_1677,In_1181,In_586);
or U1678 (N_1678,In_785,In_844);
nand U1679 (N_1679,In_357,In_262);
and U1680 (N_1680,In_83,In_1049);
nor U1681 (N_1681,In_965,In_1219);
xor U1682 (N_1682,In_28,In_1234);
nand U1683 (N_1683,In_594,In_116);
xnor U1684 (N_1684,In_273,In_735);
nor U1685 (N_1685,In_398,In_395);
nand U1686 (N_1686,In_1283,In_431);
or U1687 (N_1687,In_348,In_1072);
nand U1688 (N_1688,In_868,In_1051);
and U1689 (N_1689,In_183,In_1067);
nand U1690 (N_1690,In_264,In_1474);
and U1691 (N_1691,In_1063,In_1340);
or U1692 (N_1692,In_946,In_974);
and U1693 (N_1693,In_1355,In_207);
xor U1694 (N_1694,In_1393,In_614);
and U1695 (N_1695,In_925,In_223);
or U1696 (N_1696,In_1390,In_715);
or U1697 (N_1697,In_412,In_1305);
nor U1698 (N_1698,In_1427,In_219);
nor U1699 (N_1699,In_186,In_782);
or U1700 (N_1700,In_438,In_43);
nand U1701 (N_1701,In_1028,In_960);
nor U1702 (N_1702,In_711,In_802);
nand U1703 (N_1703,In_132,In_66);
and U1704 (N_1704,In_1031,In_781);
and U1705 (N_1705,In_696,In_104);
nor U1706 (N_1706,In_464,In_1385);
nor U1707 (N_1707,In_116,In_1085);
and U1708 (N_1708,In_738,In_287);
nand U1709 (N_1709,In_1289,In_1383);
nand U1710 (N_1710,In_553,In_1285);
nor U1711 (N_1711,In_918,In_694);
and U1712 (N_1712,In_198,In_702);
and U1713 (N_1713,In_1306,In_1451);
or U1714 (N_1714,In_214,In_768);
nor U1715 (N_1715,In_665,In_655);
and U1716 (N_1716,In_1351,In_503);
nand U1717 (N_1717,In_726,In_1343);
nor U1718 (N_1718,In_1328,In_1271);
xnor U1719 (N_1719,In_207,In_776);
and U1720 (N_1720,In_590,In_815);
nor U1721 (N_1721,In_1199,In_184);
nand U1722 (N_1722,In_152,In_156);
xor U1723 (N_1723,In_1316,In_1456);
or U1724 (N_1724,In_451,In_513);
or U1725 (N_1725,In_60,In_173);
xor U1726 (N_1726,In_1085,In_75);
or U1727 (N_1727,In_129,In_596);
nor U1728 (N_1728,In_318,In_564);
nand U1729 (N_1729,In_178,In_363);
or U1730 (N_1730,In_29,In_1279);
or U1731 (N_1731,In_1338,In_516);
nand U1732 (N_1732,In_60,In_84);
nand U1733 (N_1733,In_1179,In_960);
xor U1734 (N_1734,In_825,In_1308);
or U1735 (N_1735,In_816,In_120);
nor U1736 (N_1736,In_1221,In_810);
and U1737 (N_1737,In_718,In_1323);
nor U1738 (N_1738,In_927,In_397);
nand U1739 (N_1739,In_755,In_392);
nand U1740 (N_1740,In_653,In_1225);
xnor U1741 (N_1741,In_971,In_1340);
nor U1742 (N_1742,In_325,In_813);
nand U1743 (N_1743,In_915,In_1111);
xnor U1744 (N_1744,In_1110,In_1098);
xor U1745 (N_1745,In_990,In_818);
xor U1746 (N_1746,In_1389,In_640);
and U1747 (N_1747,In_964,In_199);
nand U1748 (N_1748,In_951,In_529);
or U1749 (N_1749,In_990,In_1496);
xnor U1750 (N_1750,In_1048,In_187);
or U1751 (N_1751,In_256,In_610);
or U1752 (N_1752,In_693,In_1182);
and U1753 (N_1753,In_234,In_139);
nor U1754 (N_1754,In_108,In_662);
xor U1755 (N_1755,In_1350,In_554);
nand U1756 (N_1756,In_1212,In_268);
nand U1757 (N_1757,In_644,In_1332);
and U1758 (N_1758,In_1237,In_307);
nor U1759 (N_1759,In_956,In_1493);
and U1760 (N_1760,In_578,In_997);
nor U1761 (N_1761,In_802,In_418);
or U1762 (N_1762,In_712,In_1134);
or U1763 (N_1763,In_307,In_1088);
nand U1764 (N_1764,In_1199,In_346);
xnor U1765 (N_1765,In_154,In_1271);
nor U1766 (N_1766,In_566,In_681);
nand U1767 (N_1767,In_673,In_1077);
and U1768 (N_1768,In_182,In_1137);
nor U1769 (N_1769,In_1064,In_280);
and U1770 (N_1770,In_1167,In_320);
and U1771 (N_1771,In_252,In_1353);
or U1772 (N_1772,In_602,In_1071);
xor U1773 (N_1773,In_345,In_1074);
and U1774 (N_1774,In_690,In_409);
nand U1775 (N_1775,In_3,In_648);
xor U1776 (N_1776,In_36,In_1206);
or U1777 (N_1777,In_229,In_1380);
or U1778 (N_1778,In_656,In_676);
or U1779 (N_1779,In_1430,In_65);
nand U1780 (N_1780,In_0,In_1147);
or U1781 (N_1781,In_610,In_1004);
xnor U1782 (N_1782,In_31,In_37);
xor U1783 (N_1783,In_1151,In_139);
nand U1784 (N_1784,In_1365,In_363);
nor U1785 (N_1785,In_1080,In_1336);
xor U1786 (N_1786,In_912,In_903);
nor U1787 (N_1787,In_481,In_516);
xnor U1788 (N_1788,In_924,In_431);
and U1789 (N_1789,In_60,In_93);
or U1790 (N_1790,In_636,In_456);
nand U1791 (N_1791,In_671,In_128);
nor U1792 (N_1792,In_52,In_866);
nor U1793 (N_1793,In_57,In_538);
xnor U1794 (N_1794,In_429,In_318);
or U1795 (N_1795,In_409,In_3);
xnor U1796 (N_1796,In_1333,In_931);
nor U1797 (N_1797,In_161,In_1437);
or U1798 (N_1798,In_1454,In_1168);
nor U1799 (N_1799,In_41,In_183);
or U1800 (N_1800,In_258,In_430);
xor U1801 (N_1801,In_274,In_1090);
nor U1802 (N_1802,In_881,In_959);
nand U1803 (N_1803,In_698,In_235);
nor U1804 (N_1804,In_474,In_614);
nand U1805 (N_1805,In_628,In_1255);
and U1806 (N_1806,In_469,In_931);
or U1807 (N_1807,In_374,In_434);
nor U1808 (N_1808,In_515,In_46);
xnor U1809 (N_1809,In_1199,In_607);
or U1810 (N_1810,In_1153,In_1150);
nand U1811 (N_1811,In_533,In_1000);
nor U1812 (N_1812,In_612,In_182);
nor U1813 (N_1813,In_702,In_1447);
and U1814 (N_1814,In_1451,In_955);
or U1815 (N_1815,In_1316,In_1369);
nand U1816 (N_1816,In_486,In_158);
nand U1817 (N_1817,In_87,In_1298);
nand U1818 (N_1818,In_1046,In_1210);
nand U1819 (N_1819,In_1230,In_327);
nor U1820 (N_1820,In_1340,In_431);
xnor U1821 (N_1821,In_990,In_214);
nand U1822 (N_1822,In_203,In_1102);
or U1823 (N_1823,In_1020,In_1159);
nor U1824 (N_1824,In_1106,In_643);
nor U1825 (N_1825,In_1328,In_49);
xnor U1826 (N_1826,In_543,In_632);
xor U1827 (N_1827,In_1214,In_758);
nor U1828 (N_1828,In_429,In_1108);
nand U1829 (N_1829,In_1201,In_200);
and U1830 (N_1830,In_725,In_1436);
nand U1831 (N_1831,In_670,In_406);
xor U1832 (N_1832,In_1286,In_624);
xnor U1833 (N_1833,In_1169,In_684);
and U1834 (N_1834,In_494,In_833);
nand U1835 (N_1835,In_1296,In_405);
xnor U1836 (N_1836,In_717,In_1415);
or U1837 (N_1837,In_138,In_214);
or U1838 (N_1838,In_1300,In_635);
and U1839 (N_1839,In_1200,In_637);
nor U1840 (N_1840,In_706,In_1073);
xor U1841 (N_1841,In_1206,In_339);
nor U1842 (N_1842,In_652,In_506);
xnor U1843 (N_1843,In_947,In_145);
or U1844 (N_1844,In_862,In_191);
and U1845 (N_1845,In_631,In_320);
or U1846 (N_1846,In_274,In_37);
or U1847 (N_1847,In_429,In_939);
xor U1848 (N_1848,In_1373,In_203);
xor U1849 (N_1849,In_934,In_619);
and U1850 (N_1850,In_1258,In_925);
nand U1851 (N_1851,In_352,In_1395);
and U1852 (N_1852,In_1442,In_811);
nor U1853 (N_1853,In_1063,In_217);
nor U1854 (N_1854,In_521,In_462);
xor U1855 (N_1855,In_423,In_784);
xnor U1856 (N_1856,In_520,In_629);
xnor U1857 (N_1857,In_1372,In_95);
nor U1858 (N_1858,In_516,In_1476);
and U1859 (N_1859,In_1011,In_237);
and U1860 (N_1860,In_428,In_961);
or U1861 (N_1861,In_1051,In_1173);
xnor U1862 (N_1862,In_717,In_1461);
nor U1863 (N_1863,In_459,In_1343);
nor U1864 (N_1864,In_1123,In_1060);
or U1865 (N_1865,In_946,In_105);
or U1866 (N_1866,In_657,In_34);
or U1867 (N_1867,In_397,In_894);
nor U1868 (N_1868,In_1449,In_1267);
xnor U1869 (N_1869,In_848,In_112);
xnor U1870 (N_1870,In_1335,In_466);
xnor U1871 (N_1871,In_1262,In_1409);
nand U1872 (N_1872,In_429,In_1495);
or U1873 (N_1873,In_1225,In_1444);
nor U1874 (N_1874,In_82,In_1035);
and U1875 (N_1875,In_1449,In_138);
nor U1876 (N_1876,In_625,In_1357);
and U1877 (N_1877,In_530,In_604);
nor U1878 (N_1878,In_241,In_442);
and U1879 (N_1879,In_1325,In_1307);
xnor U1880 (N_1880,In_470,In_874);
xor U1881 (N_1881,In_1285,In_123);
xor U1882 (N_1882,In_430,In_603);
nor U1883 (N_1883,In_74,In_758);
nor U1884 (N_1884,In_472,In_1028);
nor U1885 (N_1885,In_1225,In_236);
or U1886 (N_1886,In_247,In_1314);
nor U1887 (N_1887,In_142,In_279);
xor U1888 (N_1888,In_919,In_785);
xnor U1889 (N_1889,In_847,In_1201);
and U1890 (N_1890,In_737,In_997);
nor U1891 (N_1891,In_1416,In_879);
xor U1892 (N_1892,In_393,In_929);
and U1893 (N_1893,In_742,In_1230);
nand U1894 (N_1894,In_1115,In_1499);
and U1895 (N_1895,In_1212,In_1118);
nand U1896 (N_1896,In_599,In_223);
xor U1897 (N_1897,In_549,In_1431);
xnor U1898 (N_1898,In_1464,In_1158);
nand U1899 (N_1899,In_596,In_797);
nand U1900 (N_1900,In_1334,In_646);
xor U1901 (N_1901,In_1018,In_597);
nor U1902 (N_1902,In_553,In_937);
xnor U1903 (N_1903,In_864,In_426);
nand U1904 (N_1904,In_927,In_13);
nand U1905 (N_1905,In_1042,In_7);
nor U1906 (N_1906,In_905,In_251);
or U1907 (N_1907,In_679,In_1200);
and U1908 (N_1908,In_443,In_195);
or U1909 (N_1909,In_1289,In_444);
and U1910 (N_1910,In_453,In_863);
nor U1911 (N_1911,In_1276,In_685);
nand U1912 (N_1912,In_1279,In_529);
or U1913 (N_1913,In_268,In_1420);
or U1914 (N_1914,In_1481,In_372);
nand U1915 (N_1915,In_912,In_920);
and U1916 (N_1916,In_1411,In_1014);
nand U1917 (N_1917,In_1447,In_379);
and U1918 (N_1918,In_582,In_836);
nor U1919 (N_1919,In_1352,In_1230);
nor U1920 (N_1920,In_1407,In_238);
xnor U1921 (N_1921,In_414,In_1081);
and U1922 (N_1922,In_288,In_1269);
and U1923 (N_1923,In_877,In_966);
nand U1924 (N_1924,In_1446,In_1208);
nand U1925 (N_1925,In_1356,In_564);
nand U1926 (N_1926,In_432,In_1428);
and U1927 (N_1927,In_986,In_849);
nand U1928 (N_1928,In_1349,In_1392);
nor U1929 (N_1929,In_1268,In_218);
or U1930 (N_1930,In_1305,In_690);
xnor U1931 (N_1931,In_1105,In_77);
and U1932 (N_1932,In_353,In_1033);
and U1933 (N_1933,In_1258,In_1071);
nand U1934 (N_1934,In_1218,In_1127);
nand U1935 (N_1935,In_858,In_1019);
nor U1936 (N_1936,In_218,In_1124);
or U1937 (N_1937,In_1000,In_518);
and U1938 (N_1938,In_1421,In_956);
and U1939 (N_1939,In_1399,In_503);
xnor U1940 (N_1940,In_905,In_490);
nand U1941 (N_1941,In_997,In_1493);
or U1942 (N_1942,In_1173,In_1472);
or U1943 (N_1943,In_735,In_194);
and U1944 (N_1944,In_739,In_85);
nor U1945 (N_1945,In_1315,In_337);
nand U1946 (N_1946,In_1458,In_1035);
and U1947 (N_1947,In_229,In_1001);
nor U1948 (N_1948,In_404,In_1321);
nand U1949 (N_1949,In_1390,In_1337);
or U1950 (N_1950,In_963,In_1153);
xnor U1951 (N_1951,In_675,In_210);
nor U1952 (N_1952,In_25,In_886);
xnor U1953 (N_1953,In_186,In_93);
xnor U1954 (N_1954,In_595,In_986);
nor U1955 (N_1955,In_361,In_635);
or U1956 (N_1956,In_957,In_1077);
nand U1957 (N_1957,In_115,In_267);
and U1958 (N_1958,In_1145,In_738);
xor U1959 (N_1959,In_1298,In_634);
nand U1960 (N_1960,In_849,In_613);
and U1961 (N_1961,In_109,In_505);
nor U1962 (N_1962,In_598,In_1154);
nor U1963 (N_1963,In_659,In_632);
or U1964 (N_1964,In_699,In_237);
nor U1965 (N_1965,In_1164,In_758);
or U1966 (N_1966,In_838,In_1308);
nor U1967 (N_1967,In_95,In_313);
nand U1968 (N_1968,In_235,In_318);
or U1969 (N_1969,In_1432,In_1477);
xor U1970 (N_1970,In_681,In_837);
nor U1971 (N_1971,In_1084,In_431);
nand U1972 (N_1972,In_1358,In_326);
nand U1973 (N_1973,In_79,In_51);
or U1974 (N_1974,In_109,In_51);
xor U1975 (N_1975,In_1205,In_188);
xnor U1976 (N_1976,In_538,In_521);
xnor U1977 (N_1977,In_1123,In_688);
nand U1978 (N_1978,In_276,In_1238);
nor U1979 (N_1979,In_1125,In_1050);
nor U1980 (N_1980,In_1093,In_417);
or U1981 (N_1981,In_243,In_823);
or U1982 (N_1982,In_833,In_252);
and U1983 (N_1983,In_134,In_210);
nand U1984 (N_1984,In_813,In_114);
or U1985 (N_1985,In_107,In_831);
nand U1986 (N_1986,In_1250,In_52);
nand U1987 (N_1987,In_1362,In_0);
xor U1988 (N_1988,In_28,In_1315);
nor U1989 (N_1989,In_1202,In_399);
nor U1990 (N_1990,In_1292,In_231);
and U1991 (N_1991,In_1061,In_745);
or U1992 (N_1992,In_856,In_1203);
nand U1993 (N_1993,In_1247,In_1001);
nor U1994 (N_1994,In_1146,In_344);
nor U1995 (N_1995,In_687,In_880);
or U1996 (N_1996,In_353,In_266);
nor U1997 (N_1997,In_991,In_243);
nand U1998 (N_1998,In_1,In_329);
nor U1999 (N_1999,In_1289,In_1156);
and U2000 (N_2000,In_1375,In_426);
or U2001 (N_2001,In_1007,In_133);
nand U2002 (N_2002,In_320,In_1307);
xor U2003 (N_2003,In_213,In_1427);
or U2004 (N_2004,In_120,In_1349);
nand U2005 (N_2005,In_136,In_1178);
nand U2006 (N_2006,In_1012,In_164);
nand U2007 (N_2007,In_1098,In_654);
nand U2008 (N_2008,In_541,In_1359);
nand U2009 (N_2009,In_1145,In_242);
xor U2010 (N_2010,In_500,In_521);
xor U2011 (N_2011,In_1479,In_1105);
nor U2012 (N_2012,In_379,In_439);
or U2013 (N_2013,In_605,In_243);
nand U2014 (N_2014,In_957,In_601);
xor U2015 (N_2015,In_804,In_351);
or U2016 (N_2016,In_473,In_1368);
and U2017 (N_2017,In_768,In_839);
and U2018 (N_2018,In_8,In_930);
nand U2019 (N_2019,In_1108,In_909);
and U2020 (N_2020,In_95,In_1044);
xnor U2021 (N_2021,In_350,In_1084);
and U2022 (N_2022,In_918,In_20);
nand U2023 (N_2023,In_837,In_558);
nor U2024 (N_2024,In_1256,In_941);
or U2025 (N_2025,In_905,In_434);
and U2026 (N_2026,In_896,In_1406);
nor U2027 (N_2027,In_1339,In_761);
nor U2028 (N_2028,In_1482,In_72);
or U2029 (N_2029,In_1495,In_1234);
or U2030 (N_2030,In_915,In_1130);
nor U2031 (N_2031,In_189,In_800);
nand U2032 (N_2032,In_760,In_209);
nor U2033 (N_2033,In_571,In_990);
xor U2034 (N_2034,In_294,In_1377);
xor U2035 (N_2035,In_162,In_1486);
nand U2036 (N_2036,In_797,In_597);
and U2037 (N_2037,In_1096,In_180);
and U2038 (N_2038,In_440,In_170);
nand U2039 (N_2039,In_1176,In_1072);
nor U2040 (N_2040,In_261,In_740);
and U2041 (N_2041,In_968,In_1339);
nand U2042 (N_2042,In_1002,In_609);
nor U2043 (N_2043,In_1418,In_1145);
nor U2044 (N_2044,In_304,In_831);
nand U2045 (N_2045,In_1341,In_1116);
and U2046 (N_2046,In_604,In_1350);
nor U2047 (N_2047,In_536,In_892);
nand U2048 (N_2048,In_745,In_608);
and U2049 (N_2049,In_652,In_554);
or U2050 (N_2050,In_842,In_341);
xnor U2051 (N_2051,In_1385,In_1291);
and U2052 (N_2052,In_1355,In_1229);
nand U2053 (N_2053,In_528,In_140);
xor U2054 (N_2054,In_1314,In_823);
nor U2055 (N_2055,In_53,In_403);
or U2056 (N_2056,In_904,In_1306);
xor U2057 (N_2057,In_1374,In_1161);
nand U2058 (N_2058,In_1466,In_460);
nand U2059 (N_2059,In_1081,In_898);
or U2060 (N_2060,In_1431,In_981);
nand U2061 (N_2061,In_595,In_413);
or U2062 (N_2062,In_1258,In_138);
nor U2063 (N_2063,In_1385,In_660);
nor U2064 (N_2064,In_1243,In_1232);
and U2065 (N_2065,In_312,In_649);
xnor U2066 (N_2066,In_98,In_407);
or U2067 (N_2067,In_445,In_590);
xnor U2068 (N_2068,In_540,In_210);
xor U2069 (N_2069,In_1138,In_895);
or U2070 (N_2070,In_534,In_1084);
and U2071 (N_2071,In_473,In_506);
or U2072 (N_2072,In_1169,In_1199);
or U2073 (N_2073,In_752,In_870);
xor U2074 (N_2074,In_1115,In_669);
and U2075 (N_2075,In_1101,In_857);
and U2076 (N_2076,In_491,In_637);
and U2077 (N_2077,In_560,In_1170);
and U2078 (N_2078,In_1375,In_1328);
and U2079 (N_2079,In_78,In_936);
or U2080 (N_2080,In_701,In_583);
and U2081 (N_2081,In_1446,In_518);
nor U2082 (N_2082,In_950,In_1014);
nand U2083 (N_2083,In_1081,In_7);
or U2084 (N_2084,In_320,In_855);
and U2085 (N_2085,In_1476,In_495);
nor U2086 (N_2086,In_1445,In_110);
nor U2087 (N_2087,In_1175,In_871);
or U2088 (N_2088,In_76,In_944);
nor U2089 (N_2089,In_756,In_483);
or U2090 (N_2090,In_868,In_1474);
xor U2091 (N_2091,In_410,In_550);
and U2092 (N_2092,In_240,In_441);
and U2093 (N_2093,In_1061,In_638);
and U2094 (N_2094,In_774,In_45);
and U2095 (N_2095,In_417,In_1325);
and U2096 (N_2096,In_245,In_195);
and U2097 (N_2097,In_539,In_568);
xnor U2098 (N_2098,In_358,In_169);
nor U2099 (N_2099,In_622,In_106);
nor U2100 (N_2100,In_1190,In_40);
nand U2101 (N_2101,In_1492,In_590);
xor U2102 (N_2102,In_1434,In_1090);
xnor U2103 (N_2103,In_64,In_410);
and U2104 (N_2104,In_1258,In_256);
nand U2105 (N_2105,In_1333,In_1106);
and U2106 (N_2106,In_377,In_1307);
nor U2107 (N_2107,In_351,In_770);
and U2108 (N_2108,In_667,In_1295);
and U2109 (N_2109,In_1150,In_1210);
nand U2110 (N_2110,In_668,In_1129);
and U2111 (N_2111,In_1479,In_118);
nor U2112 (N_2112,In_1054,In_411);
nand U2113 (N_2113,In_1306,In_1039);
and U2114 (N_2114,In_546,In_709);
and U2115 (N_2115,In_70,In_81);
nor U2116 (N_2116,In_956,In_305);
nor U2117 (N_2117,In_664,In_349);
nor U2118 (N_2118,In_671,In_376);
nor U2119 (N_2119,In_1293,In_327);
nand U2120 (N_2120,In_1222,In_1233);
nand U2121 (N_2121,In_553,In_407);
and U2122 (N_2122,In_1392,In_83);
nor U2123 (N_2123,In_520,In_1062);
nor U2124 (N_2124,In_731,In_895);
and U2125 (N_2125,In_465,In_903);
xnor U2126 (N_2126,In_12,In_704);
nor U2127 (N_2127,In_428,In_804);
or U2128 (N_2128,In_210,In_549);
nor U2129 (N_2129,In_16,In_545);
nand U2130 (N_2130,In_491,In_1046);
and U2131 (N_2131,In_1476,In_1478);
or U2132 (N_2132,In_118,In_368);
xnor U2133 (N_2133,In_308,In_932);
nor U2134 (N_2134,In_401,In_839);
nand U2135 (N_2135,In_730,In_412);
xor U2136 (N_2136,In_1320,In_921);
nand U2137 (N_2137,In_1460,In_895);
nand U2138 (N_2138,In_1080,In_112);
nand U2139 (N_2139,In_608,In_515);
nor U2140 (N_2140,In_493,In_1173);
xnor U2141 (N_2141,In_1032,In_1084);
nor U2142 (N_2142,In_1218,In_535);
nor U2143 (N_2143,In_922,In_1442);
nand U2144 (N_2144,In_1403,In_1140);
nor U2145 (N_2145,In_1372,In_1329);
or U2146 (N_2146,In_1457,In_1452);
or U2147 (N_2147,In_1465,In_1150);
nand U2148 (N_2148,In_822,In_642);
nor U2149 (N_2149,In_1372,In_470);
or U2150 (N_2150,In_391,In_857);
xor U2151 (N_2151,In_649,In_335);
and U2152 (N_2152,In_70,In_502);
nor U2153 (N_2153,In_914,In_20);
xnor U2154 (N_2154,In_11,In_918);
nor U2155 (N_2155,In_804,In_537);
nand U2156 (N_2156,In_1108,In_350);
nand U2157 (N_2157,In_318,In_113);
nand U2158 (N_2158,In_194,In_496);
nand U2159 (N_2159,In_742,In_465);
and U2160 (N_2160,In_412,In_1174);
nand U2161 (N_2161,In_1376,In_544);
nand U2162 (N_2162,In_1041,In_437);
or U2163 (N_2163,In_1200,In_1474);
nor U2164 (N_2164,In_929,In_51);
or U2165 (N_2165,In_120,In_749);
nor U2166 (N_2166,In_970,In_125);
nand U2167 (N_2167,In_838,In_1092);
or U2168 (N_2168,In_1474,In_610);
nor U2169 (N_2169,In_252,In_318);
nand U2170 (N_2170,In_1252,In_776);
and U2171 (N_2171,In_297,In_737);
and U2172 (N_2172,In_856,In_498);
nand U2173 (N_2173,In_980,In_787);
nor U2174 (N_2174,In_948,In_1187);
and U2175 (N_2175,In_619,In_462);
or U2176 (N_2176,In_743,In_549);
nor U2177 (N_2177,In_1207,In_49);
or U2178 (N_2178,In_459,In_291);
xor U2179 (N_2179,In_472,In_701);
xnor U2180 (N_2180,In_398,In_625);
nor U2181 (N_2181,In_911,In_732);
or U2182 (N_2182,In_1276,In_59);
nor U2183 (N_2183,In_654,In_651);
and U2184 (N_2184,In_963,In_1073);
or U2185 (N_2185,In_692,In_1271);
and U2186 (N_2186,In_717,In_89);
nor U2187 (N_2187,In_61,In_1466);
or U2188 (N_2188,In_1065,In_391);
or U2189 (N_2189,In_1420,In_762);
xor U2190 (N_2190,In_896,In_775);
nand U2191 (N_2191,In_1366,In_242);
nand U2192 (N_2192,In_550,In_252);
and U2193 (N_2193,In_369,In_609);
nor U2194 (N_2194,In_1453,In_429);
or U2195 (N_2195,In_884,In_1331);
or U2196 (N_2196,In_168,In_1456);
or U2197 (N_2197,In_1205,In_1402);
nor U2198 (N_2198,In_935,In_408);
xor U2199 (N_2199,In_1272,In_55);
or U2200 (N_2200,In_767,In_1361);
or U2201 (N_2201,In_1148,In_867);
nand U2202 (N_2202,In_1339,In_1297);
nor U2203 (N_2203,In_1258,In_111);
nand U2204 (N_2204,In_849,In_1169);
nand U2205 (N_2205,In_631,In_1366);
nand U2206 (N_2206,In_1492,In_60);
and U2207 (N_2207,In_165,In_578);
or U2208 (N_2208,In_273,In_1147);
xor U2209 (N_2209,In_638,In_520);
nand U2210 (N_2210,In_1352,In_651);
and U2211 (N_2211,In_770,In_299);
xor U2212 (N_2212,In_845,In_964);
nand U2213 (N_2213,In_795,In_343);
nor U2214 (N_2214,In_345,In_447);
nand U2215 (N_2215,In_449,In_6);
nand U2216 (N_2216,In_1367,In_825);
nand U2217 (N_2217,In_243,In_308);
and U2218 (N_2218,In_1024,In_1093);
or U2219 (N_2219,In_1381,In_1449);
and U2220 (N_2220,In_356,In_1065);
and U2221 (N_2221,In_1266,In_50);
or U2222 (N_2222,In_226,In_1438);
and U2223 (N_2223,In_76,In_1148);
xor U2224 (N_2224,In_415,In_135);
xnor U2225 (N_2225,In_1025,In_1031);
nand U2226 (N_2226,In_1173,In_1078);
nor U2227 (N_2227,In_1240,In_721);
nor U2228 (N_2228,In_1108,In_231);
xor U2229 (N_2229,In_1362,In_1481);
nor U2230 (N_2230,In_1332,In_817);
and U2231 (N_2231,In_596,In_721);
nand U2232 (N_2232,In_27,In_587);
xnor U2233 (N_2233,In_1486,In_715);
and U2234 (N_2234,In_356,In_962);
and U2235 (N_2235,In_966,In_565);
nor U2236 (N_2236,In_617,In_834);
and U2237 (N_2237,In_805,In_1010);
and U2238 (N_2238,In_1253,In_104);
nand U2239 (N_2239,In_1439,In_34);
and U2240 (N_2240,In_772,In_1217);
nor U2241 (N_2241,In_594,In_516);
xnor U2242 (N_2242,In_1435,In_1331);
and U2243 (N_2243,In_202,In_1484);
nor U2244 (N_2244,In_1303,In_1369);
and U2245 (N_2245,In_1257,In_640);
nand U2246 (N_2246,In_318,In_1488);
or U2247 (N_2247,In_356,In_87);
and U2248 (N_2248,In_918,In_987);
and U2249 (N_2249,In_352,In_642);
xor U2250 (N_2250,In_915,In_239);
and U2251 (N_2251,In_577,In_816);
or U2252 (N_2252,In_770,In_1356);
xor U2253 (N_2253,In_1175,In_431);
or U2254 (N_2254,In_1106,In_168);
nor U2255 (N_2255,In_1153,In_1355);
and U2256 (N_2256,In_278,In_813);
or U2257 (N_2257,In_618,In_12);
xor U2258 (N_2258,In_1212,In_239);
or U2259 (N_2259,In_77,In_860);
and U2260 (N_2260,In_412,In_689);
or U2261 (N_2261,In_88,In_1445);
nor U2262 (N_2262,In_684,In_939);
nand U2263 (N_2263,In_1013,In_595);
or U2264 (N_2264,In_519,In_601);
xnor U2265 (N_2265,In_931,In_751);
and U2266 (N_2266,In_740,In_1125);
nor U2267 (N_2267,In_1014,In_1368);
and U2268 (N_2268,In_158,In_427);
nor U2269 (N_2269,In_259,In_540);
xor U2270 (N_2270,In_601,In_1005);
nor U2271 (N_2271,In_809,In_495);
nand U2272 (N_2272,In_1078,In_731);
nand U2273 (N_2273,In_665,In_1366);
and U2274 (N_2274,In_1142,In_572);
and U2275 (N_2275,In_1462,In_1374);
and U2276 (N_2276,In_97,In_317);
and U2277 (N_2277,In_321,In_801);
nand U2278 (N_2278,In_1345,In_1389);
or U2279 (N_2279,In_1062,In_739);
nor U2280 (N_2280,In_19,In_711);
xnor U2281 (N_2281,In_1009,In_1152);
or U2282 (N_2282,In_1423,In_746);
and U2283 (N_2283,In_48,In_1055);
or U2284 (N_2284,In_1208,In_680);
and U2285 (N_2285,In_380,In_958);
nor U2286 (N_2286,In_687,In_994);
nand U2287 (N_2287,In_523,In_444);
nor U2288 (N_2288,In_1398,In_961);
nor U2289 (N_2289,In_540,In_1018);
or U2290 (N_2290,In_896,In_142);
nand U2291 (N_2291,In_513,In_98);
nand U2292 (N_2292,In_13,In_1287);
or U2293 (N_2293,In_387,In_1466);
nor U2294 (N_2294,In_255,In_1227);
or U2295 (N_2295,In_12,In_241);
or U2296 (N_2296,In_869,In_1437);
and U2297 (N_2297,In_964,In_998);
xor U2298 (N_2298,In_201,In_1128);
nand U2299 (N_2299,In_220,In_177);
xnor U2300 (N_2300,In_408,In_1433);
nor U2301 (N_2301,In_1389,In_419);
or U2302 (N_2302,In_1233,In_1440);
or U2303 (N_2303,In_932,In_781);
xnor U2304 (N_2304,In_335,In_298);
and U2305 (N_2305,In_510,In_70);
xor U2306 (N_2306,In_399,In_300);
nor U2307 (N_2307,In_1227,In_1142);
xnor U2308 (N_2308,In_1387,In_68);
nand U2309 (N_2309,In_550,In_165);
nand U2310 (N_2310,In_1142,In_623);
xnor U2311 (N_2311,In_416,In_1495);
and U2312 (N_2312,In_556,In_566);
xor U2313 (N_2313,In_998,In_1205);
or U2314 (N_2314,In_1482,In_213);
nand U2315 (N_2315,In_330,In_980);
xor U2316 (N_2316,In_1218,In_1203);
or U2317 (N_2317,In_559,In_395);
nand U2318 (N_2318,In_758,In_33);
and U2319 (N_2319,In_1090,In_968);
nand U2320 (N_2320,In_569,In_1389);
nor U2321 (N_2321,In_1340,In_313);
xnor U2322 (N_2322,In_376,In_583);
nor U2323 (N_2323,In_1268,In_801);
nor U2324 (N_2324,In_839,In_583);
or U2325 (N_2325,In_670,In_1332);
and U2326 (N_2326,In_1040,In_914);
nor U2327 (N_2327,In_799,In_1158);
xor U2328 (N_2328,In_40,In_916);
and U2329 (N_2329,In_1336,In_537);
or U2330 (N_2330,In_188,In_286);
and U2331 (N_2331,In_615,In_339);
nor U2332 (N_2332,In_1120,In_1042);
nor U2333 (N_2333,In_528,In_658);
nand U2334 (N_2334,In_1276,In_1005);
xor U2335 (N_2335,In_711,In_1119);
nand U2336 (N_2336,In_903,In_1282);
or U2337 (N_2337,In_553,In_1127);
nand U2338 (N_2338,In_1436,In_257);
nor U2339 (N_2339,In_258,In_969);
xor U2340 (N_2340,In_266,In_1349);
or U2341 (N_2341,In_469,In_1229);
nor U2342 (N_2342,In_849,In_321);
xor U2343 (N_2343,In_1370,In_143);
or U2344 (N_2344,In_577,In_1383);
nand U2345 (N_2345,In_660,In_728);
xnor U2346 (N_2346,In_929,In_1310);
and U2347 (N_2347,In_964,In_643);
nand U2348 (N_2348,In_933,In_1112);
or U2349 (N_2349,In_800,In_152);
xor U2350 (N_2350,In_40,In_508);
nand U2351 (N_2351,In_1466,In_37);
and U2352 (N_2352,In_348,In_798);
or U2353 (N_2353,In_261,In_1401);
nor U2354 (N_2354,In_178,In_847);
nor U2355 (N_2355,In_1448,In_401);
nor U2356 (N_2356,In_897,In_1270);
nand U2357 (N_2357,In_1089,In_370);
and U2358 (N_2358,In_349,In_937);
or U2359 (N_2359,In_1250,In_381);
nor U2360 (N_2360,In_1418,In_708);
nor U2361 (N_2361,In_203,In_253);
nand U2362 (N_2362,In_1236,In_614);
or U2363 (N_2363,In_52,In_253);
xnor U2364 (N_2364,In_938,In_770);
xor U2365 (N_2365,In_1067,In_117);
or U2366 (N_2366,In_1001,In_573);
nand U2367 (N_2367,In_192,In_5);
nand U2368 (N_2368,In_1310,In_849);
and U2369 (N_2369,In_840,In_460);
nor U2370 (N_2370,In_1040,In_199);
nor U2371 (N_2371,In_719,In_734);
xor U2372 (N_2372,In_880,In_100);
xnor U2373 (N_2373,In_476,In_454);
and U2374 (N_2374,In_215,In_152);
and U2375 (N_2375,In_206,In_990);
nand U2376 (N_2376,In_418,In_822);
or U2377 (N_2377,In_896,In_1055);
nor U2378 (N_2378,In_1436,In_1115);
nand U2379 (N_2379,In_175,In_988);
xor U2380 (N_2380,In_610,In_27);
nor U2381 (N_2381,In_142,In_1454);
and U2382 (N_2382,In_723,In_1027);
and U2383 (N_2383,In_345,In_907);
nand U2384 (N_2384,In_1034,In_803);
or U2385 (N_2385,In_28,In_1400);
nor U2386 (N_2386,In_860,In_887);
nand U2387 (N_2387,In_1406,In_856);
or U2388 (N_2388,In_482,In_95);
nand U2389 (N_2389,In_462,In_1109);
or U2390 (N_2390,In_191,In_120);
xor U2391 (N_2391,In_705,In_963);
nor U2392 (N_2392,In_1243,In_12);
nor U2393 (N_2393,In_676,In_166);
and U2394 (N_2394,In_115,In_841);
xor U2395 (N_2395,In_1190,In_1498);
nand U2396 (N_2396,In_1056,In_907);
or U2397 (N_2397,In_717,In_66);
and U2398 (N_2398,In_1447,In_294);
nor U2399 (N_2399,In_938,In_899);
xnor U2400 (N_2400,In_314,In_534);
or U2401 (N_2401,In_702,In_1422);
xnor U2402 (N_2402,In_819,In_143);
xnor U2403 (N_2403,In_689,In_1125);
and U2404 (N_2404,In_1495,In_109);
xnor U2405 (N_2405,In_362,In_249);
and U2406 (N_2406,In_468,In_1140);
nor U2407 (N_2407,In_1118,In_854);
nand U2408 (N_2408,In_594,In_775);
or U2409 (N_2409,In_873,In_1047);
or U2410 (N_2410,In_673,In_93);
nand U2411 (N_2411,In_921,In_1450);
nor U2412 (N_2412,In_413,In_278);
xor U2413 (N_2413,In_298,In_645);
and U2414 (N_2414,In_1499,In_24);
xnor U2415 (N_2415,In_48,In_382);
or U2416 (N_2416,In_975,In_961);
nor U2417 (N_2417,In_1171,In_663);
xnor U2418 (N_2418,In_473,In_765);
or U2419 (N_2419,In_104,In_965);
and U2420 (N_2420,In_344,In_640);
or U2421 (N_2421,In_679,In_411);
nor U2422 (N_2422,In_1156,In_1162);
and U2423 (N_2423,In_998,In_1392);
nand U2424 (N_2424,In_1002,In_1023);
nand U2425 (N_2425,In_768,In_1284);
nand U2426 (N_2426,In_597,In_359);
nor U2427 (N_2427,In_1033,In_80);
nor U2428 (N_2428,In_451,In_90);
nor U2429 (N_2429,In_805,In_452);
and U2430 (N_2430,In_202,In_902);
and U2431 (N_2431,In_1045,In_1426);
xnor U2432 (N_2432,In_163,In_1003);
nand U2433 (N_2433,In_748,In_1478);
or U2434 (N_2434,In_486,In_647);
nand U2435 (N_2435,In_437,In_98);
nand U2436 (N_2436,In_1207,In_1156);
or U2437 (N_2437,In_574,In_30);
xnor U2438 (N_2438,In_396,In_563);
or U2439 (N_2439,In_886,In_1472);
nor U2440 (N_2440,In_1498,In_509);
xnor U2441 (N_2441,In_551,In_1085);
and U2442 (N_2442,In_128,In_304);
xor U2443 (N_2443,In_556,In_616);
and U2444 (N_2444,In_776,In_637);
and U2445 (N_2445,In_1020,In_1285);
nor U2446 (N_2446,In_993,In_738);
xnor U2447 (N_2447,In_36,In_130);
and U2448 (N_2448,In_1280,In_276);
nor U2449 (N_2449,In_102,In_1277);
nor U2450 (N_2450,In_338,In_1067);
and U2451 (N_2451,In_337,In_1158);
and U2452 (N_2452,In_1346,In_868);
nor U2453 (N_2453,In_1274,In_215);
nand U2454 (N_2454,In_351,In_298);
xor U2455 (N_2455,In_1169,In_336);
nor U2456 (N_2456,In_274,In_1201);
or U2457 (N_2457,In_864,In_1217);
nand U2458 (N_2458,In_354,In_138);
nor U2459 (N_2459,In_38,In_1287);
nor U2460 (N_2460,In_773,In_1396);
nand U2461 (N_2461,In_331,In_826);
nor U2462 (N_2462,In_392,In_1492);
or U2463 (N_2463,In_792,In_476);
and U2464 (N_2464,In_333,In_205);
and U2465 (N_2465,In_1235,In_115);
and U2466 (N_2466,In_0,In_1076);
or U2467 (N_2467,In_512,In_357);
nand U2468 (N_2468,In_281,In_1184);
and U2469 (N_2469,In_99,In_64);
or U2470 (N_2470,In_215,In_1096);
and U2471 (N_2471,In_840,In_1356);
and U2472 (N_2472,In_484,In_318);
and U2473 (N_2473,In_237,In_70);
and U2474 (N_2474,In_1285,In_169);
xor U2475 (N_2475,In_722,In_644);
and U2476 (N_2476,In_260,In_470);
xnor U2477 (N_2477,In_380,In_578);
or U2478 (N_2478,In_858,In_446);
or U2479 (N_2479,In_666,In_58);
and U2480 (N_2480,In_820,In_1398);
or U2481 (N_2481,In_46,In_81);
nor U2482 (N_2482,In_1098,In_613);
xor U2483 (N_2483,In_389,In_1069);
or U2484 (N_2484,In_438,In_200);
nor U2485 (N_2485,In_326,In_735);
and U2486 (N_2486,In_96,In_642);
nor U2487 (N_2487,In_801,In_954);
nor U2488 (N_2488,In_1101,In_608);
xor U2489 (N_2489,In_492,In_84);
nor U2490 (N_2490,In_1037,In_1431);
xor U2491 (N_2491,In_891,In_1158);
nand U2492 (N_2492,In_606,In_904);
nand U2493 (N_2493,In_309,In_694);
xnor U2494 (N_2494,In_1334,In_1459);
xnor U2495 (N_2495,In_1100,In_994);
nor U2496 (N_2496,In_1161,In_1012);
or U2497 (N_2497,In_86,In_902);
or U2498 (N_2498,In_853,In_732);
nor U2499 (N_2499,In_889,In_329);
xnor U2500 (N_2500,In_1381,In_685);
nor U2501 (N_2501,In_410,In_876);
nand U2502 (N_2502,In_980,In_500);
and U2503 (N_2503,In_1066,In_922);
and U2504 (N_2504,In_933,In_493);
nor U2505 (N_2505,In_1480,In_1151);
nor U2506 (N_2506,In_970,In_33);
and U2507 (N_2507,In_632,In_562);
or U2508 (N_2508,In_715,In_523);
nand U2509 (N_2509,In_901,In_513);
and U2510 (N_2510,In_468,In_1438);
and U2511 (N_2511,In_1460,In_247);
nand U2512 (N_2512,In_489,In_715);
or U2513 (N_2513,In_1340,In_927);
and U2514 (N_2514,In_827,In_620);
nor U2515 (N_2515,In_792,In_352);
and U2516 (N_2516,In_495,In_1321);
xor U2517 (N_2517,In_38,In_687);
nand U2518 (N_2518,In_884,In_695);
and U2519 (N_2519,In_493,In_686);
and U2520 (N_2520,In_203,In_239);
nand U2521 (N_2521,In_660,In_1031);
and U2522 (N_2522,In_932,In_291);
or U2523 (N_2523,In_1369,In_1158);
and U2524 (N_2524,In_223,In_413);
nand U2525 (N_2525,In_205,In_757);
nand U2526 (N_2526,In_275,In_882);
nor U2527 (N_2527,In_601,In_762);
or U2528 (N_2528,In_1464,In_48);
nand U2529 (N_2529,In_943,In_1447);
and U2530 (N_2530,In_189,In_648);
nor U2531 (N_2531,In_1250,In_163);
xnor U2532 (N_2532,In_1445,In_1066);
and U2533 (N_2533,In_330,In_1004);
nand U2534 (N_2534,In_232,In_823);
xnor U2535 (N_2535,In_399,In_1284);
nor U2536 (N_2536,In_1354,In_838);
and U2537 (N_2537,In_482,In_858);
and U2538 (N_2538,In_827,In_1092);
xor U2539 (N_2539,In_252,In_777);
or U2540 (N_2540,In_63,In_1093);
nand U2541 (N_2541,In_390,In_315);
nand U2542 (N_2542,In_448,In_620);
nand U2543 (N_2543,In_1421,In_1223);
xnor U2544 (N_2544,In_1460,In_8);
nand U2545 (N_2545,In_1267,In_483);
xor U2546 (N_2546,In_778,In_276);
or U2547 (N_2547,In_464,In_974);
and U2548 (N_2548,In_1437,In_834);
and U2549 (N_2549,In_1136,In_47);
nand U2550 (N_2550,In_32,In_926);
and U2551 (N_2551,In_27,In_536);
xor U2552 (N_2552,In_1396,In_83);
nor U2553 (N_2553,In_844,In_640);
xnor U2554 (N_2554,In_314,In_1132);
and U2555 (N_2555,In_91,In_1094);
nand U2556 (N_2556,In_1475,In_534);
or U2557 (N_2557,In_1025,In_424);
xor U2558 (N_2558,In_667,In_96);
xnor U2559 (N_2559,In_1214,In_1124);
and U2560 (N_2560,In_829,In_175);
or U2561 (N_2561,In_1085,In_150);
nand U2562 (N_2562,In_776,In_538);
nor U2563 (N_2563,In_1069,In_1145);
and U2564 (N_2564,In_119,In_410);
nand U2565 (N_2565,In_1393,In_191);
and U2566 (N_2566,In_1117,In_1178);
xor U2567 (N_2567,In_55,In_743);
nand U2568 (N_2568,In_257,In_704);
xor U2569 (N_2569,In_759,In_308);
xor U2570 (N_2570,In_129,In_784);
or U2571 (N_2571,In_153,In_745);
xor U2572 (N_2572,In_160,In_447);
xor U2573 (N_2573,In_746,In_756);
nand U2574 (N_2574,In_651,In_1124);
xor U2575 (N_2575,In_347,In_162);
nand U2576 (N_2576,In_1153,In_54);
or U2577 (N_2577,In_1032,In_667);
nand U2578 (N_2578,In_393,In_1192);
or U2579 (N_2579,In_1001,In_447);
and U2580 (N_2580,In_1439,In_549);
and U2581 (N_2581,In_1191,In_583);
and U2582 (N_2582,In_1328,In_237);
nand U2583 (N_2583,In_294,In_955);
nand U2584 (N_2584,In_561,In_882);
or U2585 (N_2585,In_367,In_344);
nor U2586 (N_2586,In_642,In_610);
nand U2587 (N_2587,In_120,In_853);
nand U2588 (N_2588,In_1498,In_31);
and U2589 (N_2589,In_1157,In_97);
or U2590 (N_2590,In_1365,In_914);
or U2591 (N_2591,In_366,In_1272);
nor U2592 (N_2592,In_628,In_786);
nor U2593 (N_2593,In_1347,In_296);
xor U2594 (N_2594,In_1358,In_1249);
xor U2595 (N_2595,In_204,In_1468);
xnor U2596 (N_2596,In_139,In_1415);
or U2597 (N_2597,In_277,In_1167);
nor U2598 (N_2598,In_1344,In_655);
nor U2599 (N_2599,In_1490,In_535);
nor U2600 (N_2600,In_992,In_730);
xnor U2601 (N_2601,In_835,In_660);
and U2602 (N_2602,In_640,In_1294);
nand U2603 (N_2603,In_350,In_1018);
xor U2604 (N_2604,In_335,In_46);
and U2605 (N_2605,In_246,In_666);
or U2606 (N_2606,In_252,In_1407);
nand U2607 (N_2607,In_218,In_221);
nand U2608 (N_2608,In_88,In_1122);
nand U2609 (N_2609,In_302,In_546);
xor U2610 (N_2610,In_1341,In_1230);
nand U2611 (N_2611,In_885,In_1339);
nand U2612 (N_2612,In_17,In_941);
nor U2613 (N_2613,In_56,In_177);
nor U2614 (N_2614,In_6,In_48);
or U2615 (N_2615,In_1470,In_851);
nor U2616 (N_2616,In_799,In_768);
or U2617 (N_2617,In_518,In_1201);
nor U2618 (N_2618,In_1301,In_942);
or U2619 (N_2619,In_1080,In_1074);
xnor U2620 (N_2620,In_440,In_331);
or U2621 (N_2621,In_662,In_1119);
or U2622 (N_2622,In_529,In_48);
nor U2623 (N_2623,In_1136,In_310);
nand U2624 (N_2624,In_1273,In_589);
nand U2625 (N_2625,In_214,In_1210);
and U2626 (N_2626,In_737,In_821);
nor U2627 (N_2627,In_1415,In_1231);
nor U2628 (N_2628,In_767,In_288);
xor U2629 (N_2629,In_894,In_322);
or U2630 (N_2630,In_638,In_1449);
xor U2631 (N_2631,In_589,In_1366);
nor U2632 (N_2632,In_857,In_1456);
nand U2633 (N_2633,In_540,In_1053);
nand U2634 (N_2634,In_1238,In_801);
nor U2635 (N_2635,In_1235,In_387);
or U2636 (N_2636,In_805,In_848);
xor U2637 (N_2637,In_336,In_1455);
nor U2638 (N_2638,In_964,In_193);
nand U2639 (N_2639,In_915,In_702);
nand U2640 (N_2640,In_106,In_1225);
or U2641 (N_2641,In_553,In_716);
nor U2642 (N_2642,In_1132,In_775);
xnor U2643 (N_2643,In_404,In_352);
and U2644 (N_2644,In_948,In_291);
nand U2645 (N_2645,In_614,In_32);
or U2646 (N_2646,In_1220,In_235);
nand U2647 (N_2647,In_1251,In_1350);
nor U2648 (N_2648,In_1247,In_344);
nand U2649 (N_2649,In_1241,In_117);
nor U2650 (N_2650,In_661,In_704);
nor U2651 (N_2651,In_723,In_271);
and U2652 (N_2652,In_489,In_750);
nor U2653 (N_2653,In_1170,In_630);
xnor U2654 (N_2654,In_738,In_722);
nand U2655 (N_2655,In_1072,In_1457);
xnor U2656 (N_2656,In_345,In_12);
xor U2657 (N_2657,In_1229,In_1460);
xor U2658 (N_2658,In_882,In_236);
and U2659 (N_2659,In_1348,In_137);
nand U2660 (N_2660,In_940,In_831);
nor U2661 (N_2661,In_662,In_1178);
nor U2662 (N_2662,In_1153,In_789);
xnor U2663 (N_2663,In_627,In_630);
xor U2664 (N_2664,In_789,In_723);
or U2665 (N_2665,In_673,In_279);
nand U2666 (N_2666,In_894,In_181);
nand U2667 (N_2667,In_101,In_773);
xor U2668 (N_2668,In_973,In_1008);
or U2669 (N_2669,In_1286,In_306);
or U2670 (N_2670,In_161,In_704);
and U2671 (N_2671,In_326,In_30);
nand U2672 (N_2672,In_1382,In_1296);
and U2673 (N_2673,In_10,In_1416);
xnor U2674 (N_2674,In_858,In_1102);
nor U2675 (N_2675,In_1004,In_646);
nor U2676 (N_2676,In_310,In_1010);
nand U2677 (N_2677,In_1436,In_393);
and U2678 (N_2678,In_330,In_1312);
and U2679 (N_2679,In_1442,In_1180);
xnor U2680 (N_2680,In_748,In_838);
and U2681 (N_2681,In_718,In_256);
nand U2682 (N_2682,In_833,In_942);
nand U2683 (N_2683,In_1130,In_130);
or U2684 (N_2684,In_42,In_963);
and U2685 (N_2685,In_1235,In_1412);
or U2686 (N_2686,In_960,In_431);
xor U2687 (N_2687,In_216,In_48);
xor U2688 (N_2688,In_1387,In_1078);
nor U2689 (N_2689,In_749,In_299);
and U2690 (N_2690,In_732,In_1120);
nand U2691 (N_2691,In_1167,In_494);
nand U2692 (N_2692,In_1319,In_1280);
nor U2693 (N_2693,In_277,In_534);
and U2694 (N_2694,In_541,In_537);
nand U2695 (N_2695,In_345,In_142);
nor U2696 (N_2696,In_749,In_1162);
nand U2697 (N_2697,In_1478,In_379);
and U2698 (N_2698,In_938,In_334);
nor U2699 (N_2699,In_741,In_1421);
and U2700 (N_2700,In_1079,In_476);
nor U2701 (N_2701,In_300,In_1406);
nor U2702 (N_2702,In_87,In_57);
and U2703 (N_2703,In_846,In_1130);
nand U2704 (N_2704,In_1023,In_1178);
and U2705 (N_2705,In_1345,In_1369);
nand U2706 (N_2706,In_935,In_496);
or U2707 (N_2707,In_1133,In_423);
or U2708 (N_2708,In_426,In_1439);
xor U2709 (N_2709,In_363,In_1409);
nor U2710 (N_2710,In_647,In_1015);
or U2711 (N_2711,In_598,In_331);
nand U2712 (N_2712,In_401,In_319);
nor U2713 (N_2713,In_400,In_558);
nor U2714 (N_2714,In_775,In_573);
and U2715 (N_2715,In_328,In_384);
and U2716 (N_2716,In_1453,In_1117);
nor U2717 (N_2717,In_928,In_1224);
nor U2718 (N_2718,In_720,In_758);
nand U2719 (N_2719,In_183,In_1480);
and U2720 (N_2720,In_559,In_646);
nor U2721 (N_2721,In_275,In_528);
and U2722 (N_2722,In_1316,In_1051);
and U2723 (N_2723,In_1463,In_1358);
nor U2724 (N_2724,In_413,In_185);
xor U2725 (N_2725,In_308,In_1448);
and U2726 (N_2726,In_1182,In_79);
or U2727 (N_2727,In_749,In_1049);
nor U2728 (N_2728,In_1044,In_35);
nor U2729 (N_2729,In_916,In_1132);
nor U2730 (N_2730,In_602,In_587);
nand U2731 (N_2731,In_1398,In_79);
nand U2732 (N_2732,In_1157,In_782);
nand U2733 (N_2733,In_1492,In_1255);
or U2734 (N_2734,In_1262,In_1259);
xnor U2735 (N_2735,In_1357,In_1021);
nand U2736 (N_2736,In_452,In_912);
nor U2737 (N_2737,In_1449,In_1435);
nor U2738 (N_2738,In_1379,In_720);
nand U2739 (N_2739,In_571,In_1082);
nand U2740 (N_2740,In_1077,In_1394);
or U2741 (N_2741,In_96,In_1488);
nor U2742 (N_2742,In_724,In_197);
or U2743 (N_2743,In_646,In_1080);
xor U2744 (N_2744,In_174,In_958);
nand U2745 (N_2745,In_1196,In_667);
nand U2746 (N_2746,In_1437,In_1149);
or U2747 (N_2747,In_763,In_726);
or U2748 (N_2748,In_769,In_683);
nand U2749 (N_2749,In_1438,In_1083);
nor U2750 (N_2750,In_264,In_896);
and U2751 (N_2751,In_1240,In_336);
or U2752 (N_2752,In_341,In_895);
or U2753 (N_2753,In_351,In_1305);
nand U2754 (N_2754,In_1086,In_374);
nor U2755 (N_2755,In_293,In_390);
nand U2756 (N_2756,In_895,In_327);
and U2757 (N_2757,In_1353,In_106);
and U2758 (N_2758,In_296,In_1407);
nor U2759 (N_2759,In_201,In_207);
or U2760 (N_2760,In_1162,In_1060);
xor U2761 (N_2761,In_998,In_582);
nor U2762 (N_2762,In_618,In_56);
nand U2763 (N_2763,In_205,In_929);
xnor U2764 (N_2764,In_1348,In_504);
nand U2765 (N_2765,In_455,In_570);
xor U2766 (N_2766,In_841,In_1499);
or U2767 (N_2767,In_669,In_1048);
nor U2768 (N_2768,In_913,In_768);
nor U2769 (N_2769,In_662,In_1127);
nor U2770 (N_2770,In_329,In_355);
nand U2771 (N_2771,In_1426,In_1137);
nor U2772 (N_2772,In_640,In_419);
and U2773 (N_2773,In_1007,In_367);
xnor U2774 (N_2774,In_1111,In_945);
nand U2775 (N_2775,In_758,In_929);
nand U2776 (N_2776,In_523,In_861);
xor U2777 (N_2777,In_396,In_828);
or U2778 (N_2778,In_1224,In_219);
nor U2779 (N_2779,In_1215,In_454);
xor U2780 (N_2780,In_1046,In_753);
xor U2781 (N_2781,In_1251,In_1258);
xnor U2782 (N_2782,In_1458,In_1343);
nor U2783 (N_2783,In_931,In_645);
nand U2784 (N_2784,In_514,In_1145);
nor U2785 (N_2785,In_1483,In_330);
xnor U2786 (N_2786,In_29,In_1096);
and U2787 (N_2787,In_520,In_1165);
or U2788 (N_2788,In_30,In_434);
nand U2789 (N_2789,In_182,In_1265);
and U2790 (N_2790,In_330,In_1266);
and U2791 (N_2791,In_1022,In_128);
nor U2792 (N_2792,In_919,In_1051);
xnor U2793 (N_2793,In_1025,In_176);
nand U2794 (N_2794,In_808,In_1064);
nor U2795 (N_2795,In_930,In_1230);
nor U2796 (N_2796,In_410,In_1497);
xnor U2797 (N_2797,In_821,In_77);
and U2798 (N_2798,In_445,In_425);
nand U2799 (N_2799,In_966,In_905);
nand U2800 (N_2800,In_506,In_567);
xnor U2801 (N_2801,In_397,In_298);
or U2802 (N_2802,In_669,In_377);
nand U2803 (N_2803,In_72,In_673);
and U2804 (N_2804,In_196,In_936);
nand U2805 (N_2805,In_1467,In_685);
xor U2806 (N_2806,In_514,In_692);
nor U2807 (N_2807,In_979,In_1087);
and U2808 (N_2808,In_445,In_487);
nand U2809 (N_2809,In_622,In_304);
nand U2810 (N_2810,In_625,In_10);
xor U2811 (N_2811,In_638,In_196);
xnor U2812 (N_2812,In_687,In_1287);
xor U2813 (N_2813,In_958,In_229);
and U2814 (N_2814,In_1110,In_830);
xor U2815 (N_2815,In_259,In_225);
or U2816 (N_2816,In_39,In_706);
or U2817 (N_2817,In_1211,In_1220);
nor U2818 (N_2818,In_282,In_274);
and U2819 (N_2819,In_1318,In_345);
or U2820 (N_2820,In_240,In_171);
nand U2821 (N_2821,In_1345,In_932);
xnor U2822 (N_2822,In_701,In_929);
nor U2823 (N_2823,In_1103,In_1338);
xnor U2824 (N_2824,In_899,In_33);
nor U2825 (N_2825,In_1458,In_980);
and U2826 (N_2826,In_1478,In_372);
nand U2827 (N_2827,In_794,In_397);
nor U2828 (N_2828,In_429,In_420);
nor U2829 (N_2829,In_298,In_659);
nand U2830 (N_2830,In_663,In_917);
or U2831 (N_2831,In_822,In_1341);
nor U2832 (N_2832,In_602,In_75);
xnor U2833 (N_2833,In_1496,In_93);
or U2834 (N_2834,In_1413,In_1455);
xor U2835 (N_2835,In_654,In_1094);
nand U2836 (N_2836,In_675,In_672);
or U2837 (N_2837,In_1288,In_586);
nor U2838 (N_2838,In_695,In_301);
xor U2839 (N_2839,In_590,In_312);
nand U2840 (N_2840,In_1224,In_340);
or U2841 (N_2841,In_436,In_1251);
nand U2842 (N_2842,In_1157,In_796);
and U2843 (N_2843,In_1212,In_1347);
nor U2844 (N_2844,In_1090,In_560);
nor U2845 (N_2845,In_1263,In_656);
xnor U2846 (N_2846,In_1362,In_939);
nor U2847 (N_2847,In_605,In_1175);
xnor U2848 (N_2848,In_517,In_495);
xor U2849 (N_2849,In_197,In_787);
nor U2850 (N_2850,In_816,In_1014);
or U2851 (N_2851,In_146,In_1000);
xnor U2852 (N_2852,In_599,In_1033);
and U2853 (N_2853,In_481,In_564);
or U2854 (N_2854,In_147,In_32);
or U2855 (N_2855,In_589,In_1153);
and U2856 (N_2856,In_258,In_733);
nor U2857 (N_2857,In_579,In_95);
nor U2858 (N_2858,In_1356,In_1105);
and U2859 (N_2859,In_489,In_329);
nor U2860 (N_2860,In_954,In_646);
nor U2861 (N_2861,In_10,In_77);
nor U2862 (N_2862,In_1211,In_178);
nor U2863 (N_2863,In_808,In_1185);
xnor U2864 (N_2864,In_829,In_603);
and U2865 (N_2865,In_1316,In_131);
nand U2866 (N_2866,In_1205,In_740);
and U2867 (N_2867,In_296,In_1404);
or U2868 (N_2868,In_1307,In_1041);
or U2869 (N_2869,In_638,In_757);
nor U2870 (N_2870,In_527,In_1268);
xnor U2871 (N_2871,In_8,In_253);
xor U2872 (N_2872,In_758,In_827);
or U2873 (N_2873,In_599,In_694);
nor U2874 (N_2874,In_433,In_492);
xor U2875 (N_2875,In_1400,In_1310);
or U2876 (N_2876,In_901,In_1474);
or U2877 (N_2877,In_870,In_813);
and U2878 (N_2878,In_588,In_967);
nor U2879 (N_2879,In_257,In_660);
and U2880 (N_2880,In_1025,In_1164);
xor U2881 (N_2881,In_1205,In_1328);
nor U2882 (N_2882,In_36,In_1338);
and U2883 (N_2883,In_812,In_310);
nor U2884 (N_2884,In_12,In_702);
nand U2885 (N_2885,In_1341,In_757);
xor U2886 (N_2886,In_243,In_403);
and U2887 (N_2887,In_1161,In_14);
xor U2888 (N_2888,In_88,In_761);
nor U2889 (N_2889,In_721,In_232);
and U2890 (N_2890,In_1366,In_656);
xnor U2891 (N_2891,In_830,In_81);
or U2892 (N_2892,In_1403,In_308);
nand U2893 (N_2893,In_39,In_859);
xor U2894 (N_2894,In_126,In_1326);
nor U2895 (N_2895,In_27,In_833);
and U2896 (N_2896,In_733,In_62);
or U2897 (N_2897,In_1211,In_289);
nand U2898 (N_2898,In_801,In_804);
and U2899 (N_2899,In_137,In_901);
and U2900 (N_2900,In_58,In_128);
nor U2901 (N_2901,In_348,In_472);
nor U2902 (N_2902,In_277,In_182);
nor U2903 (N_2903,In_238,In_99);
nand U2904 (N_2904,In_519,In_466);
and U2905 (N_2905,In_1489,In_838);
nand U2906 (N_2906,In_749,In_32);
xnor U2907 (N_2907,In_49,In_432);
or U2908 (N_2908,In_769,In_437);
and U2909 (N_2909,In_543,In_1231);
xnor U2910 (N_2910,In_177,In_405);
nor U2911 (N_2911,In_912,In_208);
nand U2912 (N_2912,In_378,In_1105);
nor U2913 (N_2913,In_1290,In_619);
nand U2914 (N_2914,In_1099,In_206);
xnor U2915 (N_2915,In_175,In_484);
nor U2916 (N_2916,In_371,In_1369);
and U2917 (N_2917,In_855,In_1059);
xnor U2918 (N_2918,In_1204,In_947);
or U2919 (N_2919,In_179,In_932);
nand U2920 (N_2920,In_931,In_1405);
and U2921 (N_2921,In_684,In_128);
and U2922 (N_2922,In_1285,In_782);
and U2923 (N_2923,In_284,In_1403);
nor U2924 (N_2924,In_1231,In_1158);
xor U2925 (N_2925,In_26,In_711);
nand U2926 (N_2926,In_485,In_730);
nand U2927 (N_2927,In_1091,In_523);
and U2928 (N_2928,In_69,In_684);
nor U2929 (N_2929,In_1321,In_1338);
nor U2930 (N_2930,In_1121,In_747);
and U2931 (N_2931,In_1033,In_359);
nor U2932 (N_2932,In_1122,In_1051);
xor U2933 (N_2933,In_1327,In_1101);
and U2934 (N_2934,In_987,In_1367);
or U2935 (N_2935,In_1103,In_113);
xnor U2936 (N_2936,In_1076,In_397);
and U2937 (N_2937,In_214,In_431);
or U2938 (N_2938,In_54,In_523);
or U2939 (N_2939,In_66,In_469);
nor U2940 (N_2940,In_223,In_302);
nand U2941 (N_2941,In_937,In_436);
nor U2942 (N_2942,In_164,In_130);
nand U2943 (N_2943,In_368,In_222);
nand U2944 (N_2944,In_1303,In_872);
and U2945 (N_2945,In_384,In_950);
and U2946 (N_2946,In_308,In_275);
nand U2947 (N_2947,In_993,In_1378);
and U2948 (N_2948,In_605,In_1407);
nand U2949 (N_2949,In_1109,In_547);
nand U2950 (N_2950,In_1002,In_68);
nor U2951 (N_2951,In_610,In_888);
or U2952 (N_2952,In_1207,In_590);
nand U2953 (N_2953,In_824,In_1045);
and U2954 (N_2954,In_366,In_136);
nand U2955 (N_2955,In_226,In_381);
and U2956 (N_2956,In_1460,In_741);
nor U2957 (N_2957,In_632,In_1142);
and U2958 (N_2958,In_1013,In_21);
or U2959 (N_2959,In_135,In_1309);
nand U2960 (N_2960,In_430,In_755);
xor U2961 (N_2961,In_831,In_1114);
nand U2962 (N_2962,In_939,In_595);
nand U2963 (N_2963,In_770,In_1069);
or U2964 (N_2964,In_1169,In_112);
or U2965 (N_2965,In_574,In_285);
nand U2966 (N_2966,In_1155,In_609);
xnor U2967 (N_2967,In_1358,In_1356);
or U2968 (N_2968,In_632,In_1295);
xnor U2969 (N_2969,In_1277,In_456);
nor U2970 (N_2970,In_239,In_26);
or U2971 (N_2971,In_717,In_589);
nand U2972 (N_2972,In_598,In_1310);
nor U2973 (N_2973,In_11,In_835);
and U2974 (N_2974,In_977,In_1084);
and U2975 (N_2975,In_1167,In_1264);
nor U2976 (N_2976,In_707,In_610);
nor U2977 (N_2977,In_1061,In_741);
or U2978 (N_2978,In_342,In_1155);
nor U2979 (N_2979,In_245,In_149);
xnor U2980 (N_2980,In_189,In_1026);
or U2981 (N_2981,In_1441,In_357);
or U2982 (N_2982,In_1467,In_650);
nand U2983 (N_2983,In_1096,In_492);
nand U2984 (N_2984,In_1310,In_696);
nand U2985 (N_2985,In_812,In_1446);
nor U2986 (N_2986,In_1154,In_1055);
nand U2987 (N_2987,In_356,In_1170);
nor U2988 (N_2988,In_1105,In_1154);
nor U2989 (N_2989,In_825,In_269);
nand U2990 (N_2990,In_1392,In_1303);
xnor U2991 (N_2991,In_1320,In_961);
nor U2992 (N_2992,In_40,In_1063);
nor U2993 (N_2993,In_322,In_65);
xor U2994 (N_2994,In_57,In_1328);
or U2995 (N_2995,In_695,In_196);
or U2996 (N_2996,In_1082,In_714);
or U2997 (N_2997,In_1471,In_1394);
or U2998 (N_2998,In_646,In_131);
or U2999 (N_2999,In_688,In_1145);
or U3000 (N_3000,In_237,In_795);
or U3001 (N_3001,In_744,In_527);
or U3002 (N_3002,In_430,In_866);
or U3003 (N_3003,In_537,In_1019);
or U3004 (N_3004,In_844,In_527);
or U3005 (N_3005,In_301,In_274);
xnor U3006 (N_3006,In_774,In_545);
nand U3007 (N_3007,In_1486,In_1221);
xnor U3008 (N_3008,In_167,In_541);
xor U3009 (N_3009,In_829,In_1327);
and U3010 (N_3010,In_138,In_149);
nand U3011 (N_3011,In_850,In_1309);
or U3012 (N_3012,In_958,In_479);
nor U3013 (N_3013,In_359,In_783);
nor U3014 (N_3014,In_1224,In_41);
and U3015 (N_3015,In_1326,In_887);
nand U3016 (N_3016,In_724,In_1102);
nand U3017 (N_3017,In_620,In_1431);
nand U3018 (N_3018,In_189,In_175);
and U3019 (N_3019,In_144,In_268);
nor U3020 (N_3020,In_1197,In_336);
and U3021 (N_3021,In_798,In_325);
and U3022 (N_3022,In_34,In_339);
xor U3023 (N_3023,In_717,In_617);
or U3024 (N_3024,In_556,In_680);
or U3025 (N_3025,In_460,In_305);
and U3026 (N_3026,In_133,In_254);
nor U3027 (N_3027,In_913,In_995);
nor U3028 (N_3028,In_966,In_1236);
xor U3029 (N_3029,In_418,In_894);
and U3030 (N_3030,In_430,In_405);
xnor U3031 (N_3031,In_1260,In_64);
xnor U3032 (N_3032,In_145,In_990);
or U3033 (N_3033,In_570,In_101);
and U3034 (N_3034,In_329,In_770);
xnor U3035 (N_3035,In_1218,In_1409);
nand U3036 (N_3036,In_882,In_28);
nand U3037 (N_3037,In_796,In_52);
xnor U3038 (N_3038,In_205,In_1394);
nor U3039 (N_3039,In_1045,In_233);
and U3040 (N_3040,In_131,In_244);
and U3041 (N_3041,In_314,In_1098);
xnor U3042 (N_3042,In_378,In_468);
and U3043 (N_3043,In_1211,In_1048);
nand U3044 (N_3044,In_869,In_913);
nor U3045 (N_3045,In_158,In_815);
xor U3046 (N_3046,In_363,In_828);
and U3047 (N_3047,In_295,In_256);
nand U3048 (N_3048,In_1479,In_1250);
or U3049 (N_3049,In_1052,In_203);
and U3050 (N_3050,In_953,In_960);
xor U3051 (N_3051,In_166,In_1019);
nor U3052 (N_3052,In_322,In_10);
or U3053 (N_3053,In_1484,In_718);
or U3054 (N_3054,In_1006,In_1088);
and U3055 (N_3055,In_388,In_762);
xor U3056 (N_3056,In_392,In_1479);
or U3057 (N_3057,In_1117,In_250);
nor U3058 (N_3058,In_1052,In_178);
xnor U3059 (N_3059,In_46,In_1392);
or U3060 (N_3060,In_292,In_1374);
or U3061 (N_3061,In_502,In_1151);
and U3062 (N_3062,In_308,In_17);
nand U3063 (N_3063,In_762,In_842);
xnor U3064 (N_3064,In_316,In_651);
nand U3065 (N_3065,In_277,In_753);
xor U3066 (N_3066,In_399,In_1024);
or U3067 (N_3067,In_873,In_1243);
or U3068 (N_3068,In_833,In_1019);
and U3069 (N_3069,In_129,In_1029);
and U3070 (N_3070,In_1458,In_855);
or U3071 (N_3071,In_165,In_600);
nor U3072 (N_3072,In_608,In_929);
and U3073 (N_3073,In_686,In_66);
or U3074 (N_3074,In_504,In_567);
nor U3075 (N_3075,In_1401,In_616);
nand U3076 (N_3076,In_1382,In_611);
or U3077 (N_3077,In_916,In_1262);
xor U3078 (N_3078,In_520,In_963);
xnor U3079 (N_3079,In_1225,In_140);
or U3080 (N_3080,In_653,In_536);
and U3081 (N_3081,In_142,In_1346);
nor U3082 (N_3082,In_718,In_348);
nand U3083 (N_3083,In_197,In_733);
and U3084 (N_3084,In_274,In_1432);
nor U3085 (N_3085,In_1285,In_848);
nor U3086 (N_3086,In_1494,In_328);
nor U3087 (N_3087,In_1478,In_1450);
and U3088 (N_3088,In_360,In_1292);
nor U3089 (N_3089,In_810,In_449);
nor U3090 (N_3090,In_1179,In_224);
xor U3091 (N_3091,In_542,In_886);
or U3092 (N_3092,In_1455,In_1162);
xor U3093 (N_3093,In_770,In_1317);
and U3094 (N_3094,In_94,In_1175);
and U3095 (N_3095,In_457,In_40);
or U3096 (N_3096,In_714,In_201);
nor U3097 (N_3097,In_1398,In_52);
xnor U3098 (N_3098,In_491,In_68);
xor U3099 (N_3099,In_1103,In_420);
and U3100 (N_3100,In_297,In_10);
nand U3101 (N_3101,In_204,In_1463);
and U3102 (N_3102,In_14,In_1426);
nand U3103 (N_3103,In_927,In_1452);
nor U3104 (N_3104,In_682,In_456);
nor U3105 (N_3105,In_862,In_474);
or U3106 (N_3106,In_1137,In_796);
xnor U3107 (N_3107,In_193,In_1233);
or U3108 (N_3108,In_103,In_538);
nor U3109 (N_3109,In_345,In_691);
and U3110 (N_3110,In_1079,In_1477);
xor U3111 (N_3111,In_795,In_1330);
or U3112 (N_3112,In_555,In_992);
nand U3113 (N_3113,In_975,In_1110);
and U3114 (N_3114,In_1342,In_344);
xnor U3115 (N_3115,In_936,In_1154);
nor U3116 (N_3116,In_963,In_91);
nor U3117 (N_3117,In_1431,In_1064);
nor U3118 (N_3118,In_609,In_1268);
and U3119 (N_3119,In_1284,In_1464);
xor U3120 (N_3120,In_464,In_1211);
nor U3121 (N_3121,In_514,In_995);
and U3122 (N_3122,In_670,In_1020);
nand U3123 (N_3123,In_1132,In_269);
nor U3124 (N_3124,In_1499,In_849);
nand U3125 (N_3125,In_426,In_637);
or U3126 (N_3126,In_825,In_603);
or U3127 (N_3127,In_543,In_1483);
nor U3128 (N_3128,In_604,In_1020);
and U3129 (N_3129,In_476,In_741);
or U3130 (N_3130,In_306,In_1409);
nor U3131 (N_3131,In_489,In_1040);
nor U3132 (N_3132,In_319,In_1417);
nand U3133 (N_3133,In_1351,In_401);
xor U3134 (N_3134,In_833,In_248);
nand U3135 (N_3135,In_867,In_682);
and U3136 (N_3136,In_73,In_563);
and U3137 (N_3137,In_178,In_1041);
nor U3138 (N_3138,In_1383,In_1073);
nor U3139 (N_3139,In_1493,In_1260);
or U3140 (N_3140,In_1073,In_611);
nand U3141 (N_3141,In_632,In_1205);
nor U3142 (N_3142,In_972,In_429);
or U3143 (N_3143,In_1161,In_25);
nor U3144 (N_3144,In_555,In_1094);
and U3145 (N_3145,In_1372,In_52);
and U3146 (N_3146,In_1353,In_893);
and U3147 (N_3147,In_817,In_1283);
xnor U3148 (N_3148,In_599,In_288);
nand U3149 (N_3149,In_809,In_815);
nor U3150 (N_3150,In_1282,In_1422);
and U3151 (N_3151,In_1016,In_248);
or U3152 (N_3152,In_16,In_105);
xor U3153 (N_3153,In_661,In_614);
and U3154 (N_3154,In_590,In_1080);
or U3155 (N_3155,In_57,In_419);
or U3156 (N_3156,In_732,In_677);
xnor U3157 (N_3157,In_649,In_307);
nand U3158 (N_3158,In_1279,In_942);
or U3159 (N_3159,In_128,In_1271);
xor U3160 (N_3160,In_48,In_829);
nand U3161 (N_3161,In_995,In_152);
nand U3162 (N_3162,In_369,In_1078);
or U3163 (N_3163,In_734,In_1450);
and U3164 (N_3164,In_259,In_347);
nand U3165 (N_3165,In_999,In_991);
and U3166 (N_3166,In_302,In_1262);
nor U3167 (N_3167,In_1233,In_1106);
or U3168 (N_3168,In_280,In_1122);
or U3169 (N_3169,In_437,In_1284);
or U3170 (N_3170,In_271,In_1497);
or U3171 (N_3171,In_1463,In_1350);
xor U3172 (N_3172,In_240,In_1325);
xor U3173 (N_3173,In_455,In_382);
or U3174 (N_3174,In_190,In_1076);
nand U3175 (N_3175,In_903,In_221);
nand U3176 (N_3176,In_1344,In_672);
xnor U3177 (N_3177,In_1155,In_1234);
and U3178 (N_3178,In_838,In_615);
xnor U3179 (N_3179,In_254,In_1218);
nand U3180 (N_3180,In_1446,In_1041);
nor U3181 (N_3181,In_1355,In_951);
nand U3182 (N_3182,In_1403,In_179);
or U3183 (N_3183,In_724,In_871);
and U3184 (N_3184,In_947,In_1015);
nor U3185 (N_3185,In_1221,In_357);
or U3186 (N_3186,In_987,In_445);
xor U3187 (N_3187,In_386,In_936);
and U3188 (N_3188,In_702,In_1461);
and U3189 (N_3189,In_1405,In_551);
xor U3190 (N_3190,In_1055,In_915);
nand U3191 (N_3191,In_922,In_1017);
nor U3192 (N_3192,In_403,In_699);
and U3193 (N_3193,In_1299,In_1301);
nand U3194 (N_3194,In_88,In_1029);
nor U3195 (N_3195,In_183,In_675);
nor U3196 (N_3196,In_222,In_342);
or U3197 (N_3197,In_1466,In_6);
and U3198 (N_3198,In_1106,In_1050);
nand U3199 (N_3199,In_410,In_132);
nand U3200 (N_3200,In_1169,In_1164);
nand U3201 (N_3201,In_540,In_1125);
and U3202 (N_3202,In_1382,In_575);
or U3203 (N_3203,In_1309,In_114);
or U3204 (N_3204,In_503,In_747);
or U3205 (N_3205,In_186,In_535);
or U3206 (N_3206,In_491,In_688);
or U3207 (N_3207,In_1171,In_42);
xnor U3208 (N_3208,In_1431,In_1127);
nand U3209 (N_3209,In_1446,In_10);
nor U3210 (N_3210,In_485,In_918);
and U3211 (N_3211,In_359,In_1159);
nand U3212 (N_3212,In_1494,In_630);
or U3213 (N_3213,In_963,In_350);
and U3214 (N_3214,In_192,In_994);
nor U3215 (N_3215,In_1224,In_1469);
xnor U3216 (N_3216,In_20,In_955);
xor U3217 (N_3217,In_25,In_342);
or U3218 (N_3218,In_1331,In_1324);
and U3219 (N_3219,In_1233,In_1046);
xor U3220 (N_3220,In_574,In_192);
and U3221 (N_3221,In_814,In_19);
nand U3222 (N_3222,In_1172,In_134);
nor U3223 (N_3223,In_341,In_1212);
nand U3224 (N_3224,In_696,In_1308);
nand U3225 (N_3225,In_487,In_490);
and U3226 (N_3226,In_1070,In_785);
or U3227 (N_3227,In_983,In_685);
or U3228 (N_3228,In_964,In_994);
nand U3229 (N_3229,In_1075,In_1087);
xor U3230 (N_3230,In_668,In_410);
or U3231 (N_3231,In_840,In_1440);
or U3232 (N_3232,In_567,In_1381);
xnor U3233 (N_3233,In_56,In_170);
and U3234 (N_3234,In_750,In_879);
nor U3235 (N_3235,In_1356,In_519);
xnor U3236 (N_3236,In_1364,In_387);
or U3237 (N_3237,In_1188,In_971);
and U3238 (N_3238,In_830,In_247);
and U3239 (N_3239,In_11,In_1307);
xor U3240 (N_3240,In_1171,In_28);
and U3241 (N_3241,In_1328,In_882);
nor U3242 (N_3242,In_1317,In_581);
nor U3243 (N_3243,In_1395,In_1009);
and U3244 (N_3244,In_1123,In_278);
nand U3245 (N_3245,In_1281,In_896);
and U3246 (N_3246,In_918,In_1423);
nor U3247 (N_3247,In_979,In_618);
nor U3248 (N_3248,In_347,In_1097);
nand U3249 (N_3249,In_1302,In_670);
xnor U3250 (N_3250,In_1075,In_164);
nor U3251 (N_3251,In_1283,In_187);
or U3252 (N_3252,In_661,In_1061);
nor U3253 (N_3253,In_4,In_619);
nand U3254 (N_3254,In_1471,In_478);
xnor U3255 (N_3255,In_1274,In_1088);
xnor U3256 (N_3256,In_322,In_75);
xnor U3257 (N_3257,In_1268,In_520);
or U3258 (N_3258,In_1212,In_1474);
nor U3259 (N_3259,In_429,In_320);
or U3260 (N_3260,In_1359,In_872);
nor U3261 (N_3261,In_430,In_36);
nand U3262 (N_3262,In_768,In_1428);
nand U3263 (N_3263,In_491,In_434);
and U3264 (N_3264,In_650,In_186);
or U3265 (N_3265,In_106,In_1276);
nand U3266 (N_3266,In_132,In_914);
xnor U3267 (N_3267,In_1447,In_3);
nor U3268 (N_3268,In_205,In_256);
and U3269 (N_3269,In_352,In_1010);
nor U3270 (N_3270,In_599,In_1335);
nand U3271 (N_3271,In_1035,In_527);
nand U3272 (N_3272,In_343,In_475);
or U3273 (N_3273,In_1234,In_1444);
nor U3274 (N_3274,In_162,In_210);
nand U3275 (N_3275,In_220,In_60);
nor U3276 (N_3276,In_1068,In_878);
nor U3277 (N_3277,In_442,In_607);
and U3278 (N_3278,In_295,In_588);
and U3279 (N_3279,In_634,In_526);
and U3280 (N_3280,In_1337,In_208);
or U3281 (N_3281,In_1267,In_116);
nor U3282 (N_3282,In_1150,In_263);
nand U3283 (N_3283,In_1413,In_541);
and U3284 (N_3284,In_1266,In_388);
xor U3285 (N_3285,In_484,In_1336);
or U3286 (N_3286,In_1330,In_359);
nand U3287 (N_3287,In_572,In_1391);
nor U3288 (N_3288,In_981,In_980);
nor U3289 (N_3289,In_690,In_1274);
and U3290 (N_3290,In_964,In_300);
nand U3291 (N_3291,In_1134,In_794);
nor U3292 (N_3292,In_558,In_1445);
or U3293 (N_3293,In_828,In_1078);
nor U3294 (N_3294,In_1292,In_926);
xnor U3295 (N_3295,In_262,In_750);
nand U3296 (N_3296,In_522,In_109);
or U3297 (N_3297,In_1333,In_1087);
or U3298 (N_3298,In_60,In_397);
and U3299 (N_3299,In_1403,In_79);
or U3300 (N_3300,In_689,In_870);
nor U3301 (N_3301,In_1440,In_584);
nand U3302 (N_3302,In_523,In_1232);
and U3303 (N_3303,In_14,In_378);
nor U3304 (N_3304,In_594,In_1097);
and U3305 (N_3305,In_498,In_1050);
nand U3306 (N_3306,In_1018,In_404);
xor U3307 (N_3307,In_305,In_1160);
or U3308 (N_3308,In_536,In_1019);
and U3309 (N_3309,In_1065,In_433);
or U3310 (N_3310,In_1254,In_865);
and U3311 (N_3311,In_220,In_518);
and U3312 (N_3312,In_343,In_787);
xor U3313 (N_3313,In_879,In_429);
xnor U3314 (N_3314,In_1370,In_1477);
or U3315 (N_3315,In_42,In_974);
or U3316 (N_3316,In_295,In_739);
or U3317 (N_3317,In_1348,In_500);
nand U3318 (N_3318,In_214,In_474);
or U3319 (N_3319,In_920,In_356);
xor U3320 (N_3320,In_190,In_861);
and U3321 (N_3321,In_1191,In_790);
or U3322 (N_3322,In_174,In_49);
xnor U3323 (N_3323,In_1155,In_407);
and U3324 (N_3324,In_746,In_628);
or U3325 (N_3325,In_1231,In_685);
and U3326 (N_3326,In_1098,In_592);
and U3327 (N_3327,In_628,In_1105);
xnor U3328 (N_3328,In_607,In_457);
xnor U3329 (N_3329,In_231,In_545);
or U3330 (N_3330,In_459,In_1016);
nand U3331 (N_3331,In_310,In_405);
or U3332 (N_3332,In_899,In_436);
and U3333 (N_3333,In_735,In_1121);
xor U3334 (N_3334,In_653,In_355);
xnor U3335 (N_3335,In_1389,In_960);
nand U3336 (N_3336,In_1267,In_796);
and U3337 (N_3337,In_3,In_310);
xnor U3338 (N_3338,In_1173,In_1057);
xnor U3339 (N_3339,In_560,In_1476);
xor U3340 (N_3340,In_734,In_254);
and U3341 (N_3341,In_53,In_577);
nand U3342 (N_3342,In_493,In_105);
nor U3343 (N_3343,In_547,In_566);
or U3344 (N_3344,In_59,In_1005);
and U3345 (N_3345,In_41,In_307);
nor U3346 (N_3346,In_1292,In_304);
and U3347 (N_3347,In_1335,In_1140);
xnor U3348 (N_3348,In_992,In_1104);
or U3349 (N_3349,In_305,In_64);
nand U3350 (N_3350,In_1414,In_771);
and U3351 (N_3351,In_1441,In_1172);
nor U3352 (N_3352,In_884,In_1168);
or U3353 (N_3353,In_1013,In_1201);
xor U3354 (N_3354,In_1103,In_1222);
nor U3355 (N_3355,In_1218,In_1198);
or U3356 (N_3356,In_307,In_1392);
nand U3357 (N_3357,In_916,In_992);
xor U3358 (N_3358,In_62,In_654);
or U3359 (N_3359,In_1013,In_109);
nand U3360 (N_3360,In_349,In_665);
or U3361 (N_3361,In_633,In_1040);
xor U3362 (N_3362,In_1043,In_548);
or U3363 (N_3363,In_1305,In_638);
xor U3364 (N_3364,In_1457,In_1167);
nor U3365 (N_3365,In_241,In_1296);
and U3366 (N_3366,In_645,In_555);
nand U3367 (N_3367,In_447,In_1155);
or U3368 (N_3368,In_19,In_645);
nor U3369 (N_3369,In_1348,In_714);
and U3370 (N_3370,In_1184,In_516);
and U3371 (N_3371,In_1469,In_719);
xnor U3372 (N_3372,In_652,In_921);
nand U3373 (N_3373,In_394,In_44);
nor U3374 (N_3374,In_1422,In_1164);
xor U3375 (N_3375,In_334,In_199);
nand U3376 (N_3376,In_1075,In_1448);
or U3377 (N_3377,In_240,In_591);
and U3378 (N_3378,In_91,In_829);
nand U3379 (N_3379,In_1089,In_548);
or U3380 (N_3380,In_600,In_583);
nand U3381 (N_3381,In_362,In_450);
xnor U3382 (N_3382,In_1207,In_105);
nand U3383 (N_3383,In_204,In_1403);
xor U3384 (N_3384,In_329,In_1079);
nor U3385 (N_3385,In_1251,In_255);
or U3386 (N_3386,In_373,In_257);
xor U3387 (N_3387,In_1465,In_724);
or U3388 (N_3388,In_141,In_525);
nor U3389 (N_3389,In_1244,In_1380);
and U3390 (N_3390,In_472,In_1168);
or U3391 (N_3391,In_483,In_1387);
xnor U3392 (N_3392,In_452,In_1154);
and U3393 (N_3393,In_1334,In_57);
and U3394 (N_3394,In_675,In_1091);
or U3395 (N_3395,In_1473,In_1193);
or U3396 (N_3396,In_18,In_38);
or U3397 (N_3397,In_1429,In_345);
and U3398 (N_3398,In_174,In_646);
xor U3399 (N_3399,In_547,In_589);
nand U3400 (N_3400,In_88,In_323);
or U3401 (N_3401,In_850,In_1313);
nor U3402 (N_3402,In_646,In_1131);
nand U3403 (N_3403,In_606,In_1470);
and U3404 (N_3404,In_664,In_1410);
nor U3405 (N_3405,In_27,In_994);
nand U3406 (N_3406,In_961,In_1355);
nand U3407 (N_3407,In_1063,In_1148);
nor U3408 (N_3408,In_520,In_1295);
xor U3409 (N_3409,In_127,In_484);
nand U3410 (N_3410,In_1457,In_52);
nor U3411 (N_3411,In_91,In_1293);
or U3412 (N_3412,In_1250,In_44);
xnor U3413 (N_3413,In_1435,In_771);
nand U3414 (N_3414,In_905,In_786);
and U3415 (N_3415,In_874,In_339);
nand U3416 (N_3416,In_518,In_642);
nand U3417 (N_3417,In_10,In_1230);
and U3418 (N_3418,In_776,In_1024);
nand U3419 (N_3419,In_619,In_57);
xnor U3420 (N_3420,In_970,In_735);
nand U3421 (N_3421,In_275,In_907);
nand U3422 (N_3422,In_456,In_1127);
and U3423 (N_3423,In_1270,In_1009);
nor U3424 (N_3424,In_35,In_1285);
xnor U3425 (N_3425,In_1403,In_81);
and U3426 (N_3426,In_749,In_601);
nand U3427 (N_3427,In_1432,In_1093);
nand U3428 (N_3428,In_626,In_1360);
nor U3429 (N_3429,In_478,In_1074);
xor U3430 (N_3430,In_298,In_754);
nand U3431 (N_3431,In_302,In_1288);
and U3432 (N_3432,In_760,In_1155);
nand U3433 (N_3433,In_163,In_1395);
and U3434 (N_3434,In_85,In_1412);
nand U3435 (N_3435,In_208,In_1062);
and U3436 (N_3436,In_86,In_575);
xor U3437 (N_3437,In_448,In_541);
and U3438 (N_3438,In_609,In_555);
nand U3439 (N_3439,In_1488,In_359);
nor U3440 (N_3440,In_497,In_39);
xor U3441 (N_3441,In_880,In_753);
or U3442 (N_3442,In_173,In_918);
and U3443 (N_3443,In_699,In_950);
or U3444 (N_3444,In_1246,In_1129);
nand U3445 (N_3445,In_569,In_989);
xnor U3446 (N_3446,In_318,In_1315);
and U3447 (N_3447,In_261,In_389);
nor U3448 (N_3448,In_935,In_538);
xnor U3449 (N_3449,In_452,In_193);
and U3450 (N_3450,In_891,In_1044);
and U3451 (N_3451,In_967,In_816);
nand U3452 (N_3452,In_768,In_1419);
and U3453 (N_3453,In_833,In_1233);
or U3454 (N_3454,In_169,In_471);
or U3455 (N_3455,In_710,In_1236);
or U3456 (N_3456,In_80,In_104);
xnor U3457 (N_3457,In_445,In_1311);
and U3458 (N_3458,In_1478,In_823);
xor U3459 (N_3459,In_1068,In_237);
xor U3460 (N_3460,In_293,In_576);
and U3461 (N_3461,In_147,In_1085);
nand U3462 (N_3462,In_1096,In_145);
or U3463 (N_3463,In_528,In_1152);
or U3464 (N_3464,In_84,In_1037);
nand U3465 (N_3465,In_1167,In_851);
or U3466 (N_3466,In_677,In_400);
nand U3467 (N_3467,In_35,In_401);
nand U3468 (N_3468,In_1221,In_24);
nand U3469 (N_3469,In_430,In_1235);
or U3470 (N_3470,In_646,In_684);
xnor U3471 (N_3471,In_1009,In_1038);
xor U3472 (N_3472,In_519,In_739);
and U3473 (N_3473,In_728,In_139);
nor U3474 (N_3474,In_817,In_230);
and U3475 (N_3475,In_1232,In_968);
and U3476 (N_3476,In_1435,In_213);
and U3477 (N_3477,In_478,In_813);
nand U3478 (N_3478,In_520,In_454);
or U3479 (N_3479,In_651,In_986);
and U3480 (N_3480,In_218,In_598);
and U3481 (N_3481,In_1379,In_1433);
nor U3482 (N_3482,In_780,In_1026);
or U3483 (N_3483,In_531,In_96);
nor U3484 (N_3484,In_674,In_488);
and U3485 (N_3485,In_557,In_73);
nor U3486 (N_3486,In_1317,In_535);
and U3487 (N_3487,In_285,In_1233);
nand U3488 (N_3488,In_790,In_32);
nor U3489 (N_3489,In_611,In_975);
nand U3490 (N_3490,In_334,In_846);
xnor U3491 (N_3491,In_1200,In_673);
or U3492 (N_3492,In_1359,In_127);
or U3493 (N_3493,In_126,In_1213);
or U3494 (N_3494,In_72,In_882);
nor U3495 (N_3495,In_350,In_941);
nand U3496 (N_3496,In_48,In_321);
or U3497 (N_3497,In_65,In_444);
and U3498 (N_3498,In_1067,In_553);
and U3499 (N_3499,In_1035,In_978);
and U3500 (N_3500,In_551,In_759);
xor U3501 (N_3501,In_1006,In_144);
nor U3502 (N_3502,In_597,In_39);
or U3503 (N_3503,In_454,In_894);
nor U3504 (N_3504,In_755,In_102);
xor U3505 (N_3505,In_678,In_1435);
nand U3506 (N_3506,In_61,In_1082);
nand U3507 (N_3507,In_1227,In_1252);
nor U3508 (N_3508,In_383,In_1);
xor U3509 (N_3509,In_1466,In_234);
xnor U3510 (N_3510,In_1041,In_123);
xor U3511 (N_3511,In_840,In_203);
or U3512 (N_3512,In_1176,In_807);
xnor U3513 (N_3513,In_1405,In_179);
and U3514 (N_3514,In_38,In_797);
nor U3515 (N_3515,In_125,In_183);
nor U3516 (N_3516,In_1298,In_930);
or U3517 (N_3517,In_1021,In_1123);
nand U3518 (N_3518,In_635,In_142);
nor U3519 (N_3519,In_1262,In_1380);
and U3520 (N_3520,In_625,In_1387);
nor U3521 (N_3521,In_985,In_191);
nor U3522 (N_3522,In_1399,In_728);
or U3523 (N_3523,In_1291,In_446);
and U3524 (N_3524,In_253,In_289);
nor U3525 (N_3525,In_1477,In_416);
xnor U3526 (N_3526,In_376,In_1344);
xor U3527 (N_3527,In_101,In_759);
or U3528 (N_3528,In_1009,In_597);
xnor U3529 (N_3529,In_1428,In_216);
and U3530 (N_3530,In_1272,In_788);
nor U3531 (N_3531,In_244,In_10);
nor U3532 (N_3532,In_931,In_740);
nor U3533 (N_3533,In_288,In_573);
xnor U3534 (N_3534,In_598,In_1420);
and U3535 (N_3535,In_441,In_1003);
nor U3536 (N_3536,In_607,In_96);
nor U3537 (N_3537,In_28,In_433);
nand U3538 (N_3538,In_514,In_110);
nor U3539 (N_3539,In_430,In_569);
or U3540 (N_3540,In_269,In_1183);
or U3541 (N_3541,In_554,In_720);
and U3542 (N_3542,In_1094,In_657);
or U3543 (N_3543,In_893,In_25);
xnor U3544 (N_3544,In_943,In_920);
and U3545 (N_3545,In_1396,In_922);
and U3546 (N_3546,In_1173,In_1053);
xor U3547 (N_3547,In_903,In_408);
and U3548 (N_3548,In_273,In_1057);
xor U3549 (N_3549,In_410,In_1358);
xnor U3550 (N_3550,In_709,In_1042);
and U3551 (N_3551,In_495,In_1053);
or U3552 (N_3552,In_758,In_227);
nand U3553 (N_3553,In_520,In_1003);
xnor U3554 (N_3554,In_1002,In_431);
and U3555 (N_3555,In_574,In_680);
xnor U3556 (N_3556,In_1022,In_1066);
or U3557 (N_3557,In_203,In_1019);
and U3558 (N_3558,In_173,In_803);
nand U3559 (N_3559,In_694,In_13);
nand U3560 (N_3560,In_1489,In_697);
or U3561 (N_3561,In_815,In_1061);
nor U3562 (N_3562,In_240,In_955);
or U3563 (N_3563,In_51,In_183);
nand U3564 (N_3564,In_988,In_721);
xnor U3565 (N_3565,In_776,In_232);
nand U3566 (N_3566,In_536,In_8);
and U3567 (N_3567,In_786,In_1297);
nand U3568 (N_3568,In_1221,In_899);
or U3569 (N_3569,In_999,In_554);
nand U3570 (N_3570,In_400,In_729);
nand U3571 (N_3571,In_543,In_1174);
and U3572 (N_3572,In_1401,In_1280);
and U3573 (N_3573,In_942,In_716);
nor U3574 (N_3574,In_977,In_412);
nand U3575 (N_3575,In_509,In_779);
nand U3576 (N_3576,In_1403,In_1449);
nor U3577 (N_3577,In_957,In_1078);
xor U3578 (N_3578,In_657,In_1007);
or U3579 (N_3579,In_538,In_186);
and U3580 (N_3580,In_233,In_928);
xor U3581 (N_3581,In_1351,In_1352);
or U3582 (N_3582,In_1108,In_783);
or U3583 (N_3583,In_906,In_431);
nor U3584 (N_3584,In_699,In_1324);
nand U3585 (N_3585,In_416,In_499);
nand U3586 (N_3586,In_723,In_860);
nand U3587 (N_3587,In_655,In_49);
nand U3588 (N_3588,In_408,In_1370);
nor U3589 (N_3589,In_625,In_793);
xnor U3590 (N_3590,In_1108,In_870);
and U3591 (N_3591,In_285,In_477);
nand U3592 (N_3592,In_121,In_123);
xnor U3593 (N_3593,In_1342,In_553);
nor U3594 (N_3594,In_244,In_40);
nor U3595 (N_3595,In_1403,In_531);
nor U3596 (N_3596,In_281,In_354);
nor U3597 (N_3597,In_402,In_1226);
and U3598 (N_3598,In_445,In_822);
xor U3599 (N_3599,In_1041,In_431);
and U3600 (N_3600,In_990,In_1123);
or U3601 (N_3601,In_836,In_230);
and U3602 (N_3602,In_1062,In_813);
or U3603 (N_3603,In_1111,In_1456);
nor U3604 (N_3604,In_302,In_826);
or U3605 (N_3605,In_684,In_954);
nand U3606 (N_3606,In_1115,In_1394);
nor U3607 (N_3607,In_229,In_567);
nor U3608 (N_3608,In_67,In_128);
nand U3609 (N_3609,In_189,In_1099);
and U3610 (N_3610,In_1394,In_214);
or U3611 (N_3611,In_1084,In_101);
nand U3612 (N_3612,In_501,In_441);
nand U3613 (N_3613,In_645,In_1205);
nand U3614 (N_3614,In_1479,In_824);
nor U3615 (N_3615,In_1021,In_794);
and U3616 (N_3616,In_837,In_350);
xnor U3617 (N_3617,In_1081,In_1084);
xor U3618 (N_3618,In_640,In_456);
and U3619 (N_3619,In_1438,In_1240);
nand U3620 (N_3620,In_667,In_1140);
xnor U3621 (N_3621,In_527,In_1173);
and U3622 (N_3622,In_40,In_468);
nor U3623 (N_3623,In_987,In_719);
nor U3624 (N_3624,In_178,In_1293);
or U3625 (N_3625,In_533,In_1451);
or U3626 (N_3626,In_632,In_1217);
and U3627 (N_3627,In_1136,In_432);
or U3628 (N_3628,In_1136,In_1295);
and U3629 (N_3629,In_703,In_1102);
nand U3630 (N_3630,In_713,In_781);
xnor U3631 (N_3631,In_875,In_940);
and U3632 (N_3632,In_1399,In_775);
nand U3633 (N_3633,In_329,In_1402);
nor U3634 (N_3634,In_287,In_935);
nor U3635 (N_3635,In_177,In_157);
and U3636 (N_3636,In_220,In_74);
or U3637 (N_3637,In_300,In_349);
or U3638 (N_3638,In_249,In_875);
or U3639 (N_3639,In_276,In_931);
nor U3640 (N_3640,In_247,In_549);
or U3641 (N_3641,In_342,In_708);
nor U3642 (N_3642,In_147,In_806);
nand U3643 (N_3643,In_841,In_1452);
nor U3644 (N_3644,In_707,In_1219);
xnor U3645 (N_3645,In_1134,In_1176);
and U3646 (N_3646,In_516,In_785);
or U3647 (N_3647,In_503,In_361);
nor U3648 (N_3648,In_963,In_1187);
nand U3649 (N_3649,In_257,In_489);
xnor U3650 (N_3650,In_394,In_1336);
or U3651 (N_3651,In_1459,In_1164);
nand U3652 (N_3652,In_408,In_1448);
nand U3653 (N_3653,In_786,In_402);
or U3654 (N_3654,In_701,In_614);
and U3655 (N_3655,In_292,In_1116);
or U3656 (N_3656,In_1132,In_734);
and U3657 (N_3657,In_508,In_64);
nand U3658 (N_3658,In_991,In_1064);
nor U3659 (N_3659,In_499,In_200);
nor U3660 (N_3660,In_1451,In_91);
nand U3661 (N_3661,In_792,In_1354);
or U3662 (N_3662,In_373,In_994);
nand U3663 (N_3663,In_237,In_464);
or U3664 (N_3664,In_1042,In_1349);
and U3665 (N_3665,In_70,In_1288);
or U3666 (N_3666,In_550,In_1312);
or U3667 (N_3667,In_1142,In_493);
nand U3668 (N_3668,In_707,In_16);
nand U3669 (N_3669,In_203,In_210);
and U3670 (N_3670,In_389,In_726);
nand U3671 (N_3671,In_775,In_981);
or U3672 (N_3672,In_217,In_1357);
xor U3673 (N_3673,In_971,In_858);
nand U3674 (N_3674,In_56,In_517);
and U3675 (N_3675,In_1474,In_882);
xor U3676 (N_3676,In_140,In_358);
and U3677 (N_3677,In_1216,In_251);
or U3678 (N_3678,In_904,In_658);
nand U3679 (N_3679,In_215,In_308);
xnor U3680 (N_3680,In_354,In_1103);
xnor U3681 (N_3681,In_654,In_1475);
and U3682 (N_3682,In_442,In_974);
or U3683 (N_3683,In_287,In_79);
and U3684 (N_3684,In_264,In_775);
nor U3685 (N_3685,In_810,In_694);
or U3686 (N_3686,In_830,In_227);
nand U3687 (N_3687,In_533,In_1217);
nand U3688 (N_3688,In_610,In_852);
nand U3689 (N_3689,In_425,In_517);
xnor U3690 (N_3690,In_312,In_157);
or U3691 (N_3691,In_684,In_471);
xnor U3692 (N_3692,In_351,In_749);
nand U3693 (N_3693,In_444,In_392);
and U3694 (N_3694,In_935,In_539);
nand U3695 (N_3695,In_963,In_88);
nor U3696 (N_3696,In_816,In_984);
nand U3697 (N_3697,In_294,In_976);
or U3698 (N_3698,In_841,In_902);
or U3699 (N_3699,In_199,In_1383);
nor U3700 (N_3700,In_385,In_645);
nor U3701 (N_3701,In_177,In_1433);
nand U3702 (N_3702,In_24,In_1212);
nor U3703 (N_3703,In_1457,In_887);
or U3704 (N_3704,In_917,In_871);
or U3705 (N_3705,In_1127,In_937);
nand U3706 (N_3706,In_391,In_1322);
xor U3707 (N_3707,In_807,In_768);
nor U3708 (N_3708,In_1291,In_617);
and U3709 (N_3709,In_1421,In_735);
or U3710 (N_3710,In_868,In_1394);
or U3711 (N_3711,In_1427,In_82);
nor U3712 (N_3712,In_411,In_1239);
nor U3713 (N_3713,In_1338,In_324);
nand U3714 (N_3714,In_904,In_54);
nand U3715 (N_3715,In_1150,In_177);
or U3716 (N_3716,In_291,In_841);
nor U3717 (N_3717,In_800,In_426);
nand U3718 (N_3718,In_1334,In_1460);
nand U3719 (N_3719,In_1216,In_1365);
nor U3720 (N_3720,In_429,In_1232);
and U3721 (N_3721,In_1279,In_1370);
or U3722 (N_3722,In_587,In_918);
nor U3723 (N_3723,In_1246,In_919);
nor U3724 (N_3724,In_1469,In_210);
nor U3725 (N_3725,In_28,In_1187);
and U3726 (N_3726,In_1039,In_831);
and U3727 (N_3727,In_178,In_797);
and U3728 (N_3728,In_1033,In_746);
or U3729 (N_3729,In_1439,In_894);
or U3730 (N_3730,In_949,In_389);
or U3731 (N_3731,In_552,In_899);
nand U3732 (N_3732,In_766,In_332);
and U3733 (N_3733,In_941,In_104);
or U3734 (N_3734,In_419,In_657);
nor U3735 (N_3735,In_913,In_1399);
xnor U3736 (N_3736,In_376,In_752);
or U3737 (N_3737,In_176,In_958);
and U3738 (N_3738,In_159,In_879);
nand U3739 (N_3739,In_946,In_962);
nor U3740 (N_3740,In_969,In_1458);
or U3741 (N_3741,In_1385,In_1476);
and U3742 (N_3742,In_813,In_367);
and U3743 (N_3743,In_1273,In_941);
nor U3744 (N_3744,In_187,In_1190);
or U3745 (N_3745,In_686,In_761);
xnor U3746 (N_3746,In_102,In_307);
or U3747 (N_3747,In_1343,In_769);
and U3748 (N_3748,In_1068,In_397);
and U3749 (N_3749,In_910,In_1465);
or U3750 (N_3750,In_810,In_100);
nand U3751 (N_3751,In_364,In_748);
and U3752 (N_3752,In_1135,In_375);
and U3753 (N_3753,In_1398,In_1472);
nand U3754 (N_3754,In_758,In_1003);
or U3755 (N_3755,In_1480,In_1249);
nor U3756 (N_3756,In_92,In_735);
nor U3757 (N_3757,In_918,In_1069);
nor U3758 (N_3758,In_1299,In_729);
or U3759 (N_3759,In_1372,In_412);
xnor U3760 (N_3760,In_178,In_975);
nand U3761 (N_3761,In_579,In_366);
xnor U3762 (N_3762,In_333,In_701);
nand U3763 (N_3763,In_649,In_1268);
nand U3764 (N_3764,In_793,In_1456);
and U3765 (N_3765,In_361,In_553);
or U3766 (N_3766,In_1288,In_689);
nand U3767 (N_3767,In_794,In_190);
and U3768 (N_3768,In_647,In_530);
and U3769 (N_3769,In_1390,In_766);
nand U3770 (N_3770,In_1470,In_880);
nand U3771 (N_3771,In_1114,In_980);
and U3772 (N_3772,In_795,In_1382);
xor U3773 (N_3773,In_443,In_808);
nand U3774 (N_3774,In_1328,In_573);
or U3775 (N_3775,In_1156,In_598);
and U3776 (N_3776,In_1307,In_66);
or U3777 (N_3777,In_279,In_880);
nand U3778 (N_3778,In_366,In_1268);
nand U3779 (N_3779,In_1337,In_1104);
or U3780 (N_3780,In_452,In_300);
and U3781 (N_3781,In_1057,In_870);
nand U3782 (N_3782,In_1361,In_1305);
or U3783 (N_3783,In_1230,In_13);
nand U3784 (N_3784,In_615,In_1466);
nand U3785 (N_3785,In_318,In_902);
xor U3786 (N_3786,In_1086,In_172);
or U3787 (N_3787,In_728,In_1215);
nand U3788 (N_3788,In_1168,In_867);
nand U3789 (N_3789,In_1142,In_484);
nand U3790 (N_3790,In_1328,In_1452);
nor U3791 (N_3791,In_440,In_451);
nand U3792 (N_3792,In_1169,In_524);
nand U3793 (N_3793,In_915,In_1304);
xnor U3794 (N_3794,In_249,In_1084);
or U3795 (N_3795,In_1470,In_339);
and U3796 (N_3796,In_1242,In_194);
or U3797 (N_3797,In_402,In_738);
xnor U3798 (N_3798,In_896,In_715);
xor U3799 (N_3799,In_917,In_326);
nor U3800 (N_3800,In_186,In_830);
xor U3801 (N_3801,In_1174,In_1102);
nor U3802 (N_3802,In_1018,In_595);
nand U3803 (N_3803,In_1252,In_425);
and U3804 (N_3804,In_315,In_572);
or U3805 (N_3805,In_1038,In_1140);
nor U3806 (N_3806,In_257,In_75);
and U3807 (N_3807,In_1101,In_788);
and U3808 (N_3808,In_1468,In_1134);
or U3809 (N_3809,In_1098,In_182);
nor U3810 (N_3810,In_780,In_89);
nand U3811 (N_3811,In_535,In_245);
xnor U3812 (N_3812,In_478,In_1498);
and U3813 (N_3813,In_1031,In_79);
nand U3814 (N_3814,In_639,In_762);
nor U3815 (N_3815,In_1473,In_1036);
and U3816 (N_3816,In_1231,In_801);
and U3817 (N_3817,In_1215,In_406);
or U3818 (N_3818,In_1132,In_237);
xnor U3819 (N_3819,In_820,In_784);
and U3820 (N_3820,In_1475,In_1403);
nand U3821 (N_3821,In_993,In_434);
xnor U3822 (N_3822,In_545,In_1319);
nand U3823 (N_3823,In_1220,In_715);
or U3824 (N_3824,In_49,In_114);
and U3825 (N_3825,In_1400,In_1099);
nor U3826 (N_3826,In_597,In_954);
xor U3827 (N_3827,In_1174,In_617);
nand U3828 (N_3828,In_246,In_396);
or U3829 (N_3829,In_13,In_1098);
xor U3830 (N_3830,In_1092,In_342);
or U3831 (N_3831,In_175,In_1308);
or U3832 (N_3832,In_659,In_990);
xnor U3833 (N_3833,In_613,In_1314);
nand U3834 (N_3834,In_102,In_1137);
and U3835 (N_3835,In_1018,In_857);
and U3836 (N_3836,In_122,In_1130);
nor U3837 (N_3837,In_735,In_529);
nand U3838 (N_3838,In_1030,In_1180);
and U3839 (N_3839,In_624,In_1076);
nand U3840 (N_3840,In_859,In_212);
xor U3841 (N_3841,In_809,In_1263);
nand U3842 (N_3842,In_832,In_235);
or U3843 (N_3843,In_254,In_1075);
xnor U3844 (N_3844,In_956,In_926);
or U3845 (N_3845,In_91,In_492);
and U3846 (N_3846,In_517,In_977);
nor U3847 (N_3847,In_944,In_35);
xor U3848 (N_3848,In_677,In_1225);
nor U3849 (N_3849,In_102,In_886);
nand U3850 (N_3850,In_778,In_42);
or U3851 (N_3851,In_259,In_946);
nand U3852 (N_3852,In_842,In_904);
nand U3853 (N_3853,In_503,In_1223);
nor U3854 (N_3854,In_169,In_29);
and U3855 (N_3855,In_1266,In_492);
or U3856 (N_3856,In_1381,In_307);
nand U3857 (N_3857,In_839,In_1339);
or U3858 (N_3858,In_442,In_1338);
or U3859 (N_3859,In_939,In_320);
and U3860 (N_3860,In_672,In_172);
nand U3861 (N_3861,In_220,In_107);
or U3862 (N_3862,In_767,In_18);
xor U3863 (N_3863,In_136,In_56);
and U3864 (N_3864,In_854,In_722);
or U3865 (N_3865,In_1483,In_242);
nor U3866 (N_3866,In_1031,In_772);
or U3867 (N_3867,In_187,In_1067);
and U3868 (N_3868,In_195,In_1221);
nor U3869 (N_3869,In_704,In_604);
xor U3870 (N_3870,In_1330,In_1063);
and U3871 (N_3871,In_298,In_1223);
and U3872 (N_3872,In_288,In_1225);
xor U3873 (N_3873,In_1257,In_274);
or U3874 (N_3874,In_14,In_315);
xnor U3875 (N_3875,In_1252,In_1161);
nand U3876 (N_3876,In_283,In_453);
nand U3877 (N_3877,In_1439,In_554);
xnor U3878 (N_3878,In_592,In_1431);
nor U3879 (N_3879,In_1320,In_1410);
and U3880 (N_3880,In_453,In_233);
nor U3881 (N_3881,In_755,In_484);
nand U3882 (N_3882,In_1016,In_615);
nand U3883 (N_3883,In_403,In_809);
xnor U3884 (N_3884,In_187,In_1138);
nand U3885 (N_3885,In_1053,In_546);
xnor U3886 (N_3886,In_415,In_171);
nor U3887 (N_3887,In_979,In_1022);
nand U3888 (N_3888,In_353,In_1342);
or U3889 (N_3889,In_1002,In_114);
xnor U3890 (N_3890,In_1050,In_749);
nor U3891 (N_3891,In_1002,In_345);
nand U3892 (N_3892,In_684,In_414);
nor U3893 (N_3893,In_12,In_469);
or U3894 (N_3894,In_1343,In_963);
nor U3895 (N_3895,In_158,In_481);
and U3896 (N_3896,In_345,In_1026);
nor U3897 (N_3897,In_1152,In_455);
or U3898 (N_3898,In_1240,In_603);
xor U3899 (N_3899,In_1153,In_1075);
nand U3900 (N_3900,In_1086,In_698);
xor U3901 (N_3901,In_494,In_465);
and U3902 (N_3902,In_1029,In_1221);
nand U3903 (N_3903,In_1093,In_95);
and U3904 (N_3904,In_1336,In_1450);
nand U3905 (N_3905,In_1380,In_869);
nand U3906 (N_3906,In_401,In_755);
nand U3907 (N_3907,In_391,In_837);
or U3908 (N_3908,In_502,In_566);
xor U3909 (N_3909,In_1427,In_1325);
nand U3910 (N_3910,In_201,In_372);
nor U3911 (N_3911,In_907,In_1111);
and U3912 (N_3912,In_379,In_371);
xor U3913 (N_3913,In_14,In_1398);
nand U3914 (N_3914,In_1155,In_705);
xor U3915 (N_3915,In_216,In_293);
nand U3916 (N_3916,In_303,In_1449);
nor U3917 (N_3917,In_1024,In_108);
nand U3918 (N_3918,In_612,In_1384);
nor U3919 (N_3919,In_169,In_298);
or U3920 (N_3920,In_60,In_838);
and U3921 (N_3921,In_951,In_369);
and U3922 (N_3922,In_856,In_776);
and U3923 (N_3923,In_409,In_71);
or U3924 (N_3924,In_1182,In_687);
xor U3925 (N_3925,In_720,In_1473);
nand U3926 (N_3926,In_1123,In_479);
or U3927 (N_3927,In_742,In_945);
xor U3928 (N_3928,In_79,In_447);
nand U3929 (N_3929,In_1291,In_212);
or U3930 (N_3930,In_1114,In_328);
nor U3931 (N_3931,In_200,In_1222);
nor U3932 (N_3932,In_1073,In_145);
or U3933 (N_3933,In_1275,In_1197);
or U3934 (N_3934,In_315,In_1493);
nand U3935 (N_3935,In_643,In_506);
and U3936 (N_3936,In_605,In_517);
xor U3937 (N_3937,In_1449,In_1038);
nor U3938 (N_3938,In_1273,In_478);
and U3939 (N_3939,In_180,In_227);
xor U3940 (N_3940,In_992,In_61);
nor U3941 (N_3941,In_1298,In_430);
xor U3942 (N_3942,In_174,In_1421);
nor U3943 (N_3943,In_533,In_1457);
xnor U3944 (N_3944,In_375,In_691);
and U3945 (N_3945,In_1318,In_1340);
xor U3946 (N_3946,In_1203,In_6);
or U3947 (N_3947,In_1448,In_334);
nor U3948 (N_3948,In_363,In_1344);
or U3949 (N_3949,In_630,In_401);
nor U3950 (N_3950,In_52,In_207);
nor U3951 (N_3951,In_7,In_519);
xor U3952 (N_3952,In_1249,In_1456);
and U3953 (N_3953,In_434,In_242);
nand U3954 (N_3954,In_824,In_1115);
and U3955 (N_3955,In_508,In_948);
or U3956 (N_3956,In_432,In_1225);
nor U3957 (N_3957,In_328,In_579);
and U3958 (N_3958,In_195,In_947);
nand U3959 (N_3959,In_15,In_19);
or U3960 (N_3960,In_1489,In_668);
nor U3961 (N_3961,In_120,In_1436);
nor U3962 (N_3962,In_280,In_1237);
xnor U3963 (N_3963,In_1208,In_802);
nand U3964 (N_3964,In_500,In_1411);
xnor U3965 (N_3965,In_22,In_286);
or U3966 (N_3966,In_263,In_1036);
or U3967 (N_3967,In_1113,In_907);
and U3968 (N_3968,In_1087,In_648);
nand U3969 (N_3969,In_601,In_255);
and U3970 (N_3970,In_1122,In_7);
or U3971 (N_3971,In_184,In_1308);
and U3972 (N_3972,In_262,In_391);
nor U3973 (N_3973,In_516,In_1270);
or U3974 (N_3974,In_1308,In_789);
xor U3975 (N_3975,In_928,In_194);
nor U3976 (N_3976,In_1100,In_579);
and U3977 (N_3977,In_243,In_601);
and U3978 (N_3978,In_17,In_117);
or U3979 (N_3979,In_121,In_614);
nand U3980 (N_3980,In_1107,In_1115);
nor U3981 (N_3981,In_913,In_180);
nor U3982 (N_3982,In_1358,In_1271);
xor U3983 (N_3983,In_480,In_947);
and U3984 (N_3984,In_979,In_1461);
xor U3985 (N_3985,In_1232,In_583);
nor U3986 (N_3986,In_1308,In_1253);
and U3987 (N_3987,In_1205,In_277);
or U3988 (N_3988,In_730,In_668);
and U3989 (N_3989,In_955,In_711);
xor U3990 (N_3990,In_953,In_1457);
xnor U3991 (N_3991,In_120,In_19);
and U3992 (N_3992,In_298,In_121);
or U3993 (N_3993,In_516,In_1426);
and U3994 (N_3994,In_1162,In_1493);
xor U3995 (N_3995,In_927,In_652);
nor U3996 (N_3996,In_1414,In_495);
and U3997 (N_3997,In_45,In_781);
or U3998 (N_3998,In_688,In_572);
and U3999 (N_3999,In_294,In_532);
xnor U4000 (N_4000,In_104,In_913);
xnor U4001 (N_4001,In_543,In_1451);
and U4002 (N_4002,In_521,In_1449);
and U4003 (N_4003,In_167,In_474);
or U4004 (N_4004,In_852,In_1409);
nand U4005 (N_4005,In_6,In_536);
and U4006 (N_4006,In_266,In_691);
or U4007 (N_4007,In_180,In_718);
xor U4008 (N_4008,In_1344,In_81);
and U4009 (N_4009,In_1127,In_228);
nand U4010 (N_4010,In_273,In_98);
nor U4011 (N_4011,In_942,In_717);
and U4012 (N_4012,In_428,In_101);
or U4013 (N_4013,In_1100,In_338);
nand U4014 (N_4014,In_8,In_128);
nand U4015 (N_4015,In_196,In_1168);
nand U4016 (N_4016,In_145,In_1373);
and U4017 (N_4017,In_80,In_1415);
xnor U4018 (N_4018,In_851,In_817);
xnor U4019 (N_4019,In_654,In_718);
and U4020 (N_4020,In_944,In_166);
xnor U4021 (N_4021,In_1417,In_1110);
and U4022 (N_4022,In_476,In_1067);
or U4023 (N_4023,In_709,In_1224);
and U4024 (N_4024,In_633,In_139);
nor U4025 (N_4025,In_304,In_1077);
nand U4026 (N_4026,In_292,In_391);
xnor U4027 (N_4027,In_474,In_881);
nand U4028 (N_4028,In_237,In_982);
or U4029 (N_4029,In_1257,In_1356);
xor U4030 (N_4030,In_248,In_109);
nor U4031 (N_4031,In_719,In_851);
nor U4032 (N_4032,In_431,In_254);
xor U4033 (N_4033,In_1182,In_382);
nor U4034 (N_4034,In_480,In_466);
xnor U4035 (N_4035,In_1153,In_1015);
xnor U4036 (N_4036,In_319,In_1486);
nand U4037 (N_4037,In_673,In_140);
xor U4038 (N_4038,In_752,In_100);
nand U4039 (N_4039,In_450,In_1032);
xor U4040 (N_4040,In_729,In_749);
xor U4041 (N_4041,In_1495,In_467);
xnor U4042 (N_4042,In_1239,In_1343);
nand U4043 (N_4043,In_781,In_108);
xor U4044 (N_4044,In_251,In_1292);
xor U4045 (N_4045,In_352,In_323);
nor U4046 (N_4046,In_1004,In_1279);
and U4047 (N_4047,In_166,In_434);
and U4048 (N_4048,In_611,In_319);
and U4049 (N_4049,In_561,In_1439);
nand U4050 (N_4050,In_878,In_418);
or U4051 (N_4051,In_1166,In_1404);
xor U4052 (N_4052,In_653,In_935);
nand U4053 (N_4053,In_738,In_1339);
and U4054 (N_4054,In_857,In_1001);
nor U4055 (N_4055,In_276,In_566);
xor U4056 (N_4056,In_1263,In_207);
xnor U4057 (N_4057,In_324,In_488);
and U4058 (N_4058,In_499,In_1094);
xnor U4059 (N_4059,In_1341,In_904);
and U4060 (N_4060,In_397,In_1112);
nor U4061 (N_4061,In_758,In_20);
or U4062 (N_4062,In_883,In_996);
nand U4063 (N_4063,In_425,In_316);
and U4064 (N_4064,In_361,In_970);
nor U4065 (N_4065,In_851,In_247);
nor U4066 (N_4066,In_1422,In_1047);
nand U4067 (N_4067,In_1383,In_875);
or U4068 (N_4068,In_1482,In_697);
or U4069 (N_4069,In_280,In_119);
and U4070 (N_4070,In_664,In_44);
and U4071 (N_4071,In_314,In_1381);
or U4072 (N_4072,In_96,In_1169);
nand U4073 (N_4073,In_370,In_1455);
and U4074 (N_4074,In_569,In_850);
nor U4075 (N_4075,In_1103,In_1055);
or U4076 (N_4076,In_773,In_700);
nand U4077 (N_4077,In_784,In_650);
nor U4078 (N_4078,In_1498,In_911);
nand U4079 (N_4079,In_257,In_220);
nor U4080 (N_4080,In_138,In_1176);
nor U4081 (N_4081,In_971,In_1001);
and U4082 (N_4082,In_479,In_784);
nor U4083 (N_4083,In_864,In_151);
xor U4084 (N_4084,In_1208,In_127);
xnor U4085 (N_4085,In_1448,In_370);
xnor U4086 (N_4086,In_994,In_818);
and U4087 (N_4087,In_432,In_2);
nand U4088 (N_4088,In_1188,In_415);
nand U4089 (N_4089,In_1459,In_1112);
or U4090 (N_4090,In_1073,In_166);
xnor U4091 (N_4091,In_142,In_892);
nor U4092 (N_4092,In_332,In_1377);
nor U4093 (N_4093,In_546,In_861);
or U4094 (N_4094,In_790,In_509);
or U4095 (N_4095,In_1281,In_41);
or U4096 (N_4096,In_18,In_299);
or U4097 (N_4097,In_871,In_1313);
and U4098 (N_4098,In_1190,In_825);
xnor U4099 (N_4099,In_170,In_1456);
or U4100 (N_4100,In_49,In_512);
or U4101 (N_4101,In_631,In_945);
and U4102 (N_4102,In_699,In_314);
nand U4103 (N_4103,In_678,In_687);
nor U4104 (N_4104,In_418,In_577);
xnor U4105 (N_4105,In_1096,In_989);
and U4106 (N_4106,In_165,In_511);
or U4107 (N_4107,In_1097,In_886);
nor U4108 (N_4108,In_392,In_1485);
nand U4109 (N_4109,In_1103,In_258);
nand U4110 (N_4110,In_1244,In_1444);
nand U4111 (N_4111,In_268,In_909);
xor U4112 (N_4112,In_954,In_608);
nand U4113 (N_4113,In_288,In_734);
or U4114 (N_4114,In_1381,In_661);
nand U4115 (N_4115,In_373,In_1138);
nor U4116 (N_4116,In_1307,In_807);
or U4117 (N_4117,In_940,In_523);
or U4118 (N_4118,In_284,In_761);
xnor U4119 (N_4119,In_1121,In_1319);
nor U4120 (N_4120,In_362,In_240);
nor U4121 (N_4121,In_935,In_676);
nand U4122 (N_4122,In_740,In_895);
nand U4123 (N_4123,In_517,In_689);
nand U4124 (N_4124,In_847,In_1372);
or U4125 (N_4125,In_628,In_629);
and U4126 (N_4126,In_5,In_1254);
nand U4127 (N_4127,In_1060,In_1478);
xnor U4128 (N_4128,In_930,In_913);
nor U4129 (N_4129,In_434,In_200);
nand U4130 (N_4130,In_13,In_1416);
or U4131 (N_4131,In_755,In_320);
and U4132 (N_4132,In_576,In_1468);
nor U4133 (N_4133,In_79,In_277);
xnor U4134 (N_4134,In_449,In_532);
nor U4135 (N_4135,In_888,In_119);
or U4136 (N_4136,In_80,In_1071);
xnor U4137 (N_4137,In_348,In_605);
nor U4138 (N_4138,In_140,In_694);
nor U4139 (N_4139,In_1425,In_363);
nand U4140 (N_4140,In_1340,In_1393);
nor U4141 (N_4141,In_462,In_1212);
xor U4142 (N_4142,In_89,In_1257);
nor U4143 (N_4143,In_1149,In_463);
and U4144 (N_4144,In_85,In_1437);
and U4145 (N_4145,In_539,In_316);
xnor U4146 (N_4146,In_1134,In_1127);
nand U4147 (N_4147,In_1189,In_1422);
nor U4148 (N_4148,In_362,In_691);
nand U4149 (N_4149,In_1429,In_1433);
xor U4150 (N_4150,In_173,In_1193);
and U4151 (N_4151,In_525,In_146);
or U4152 (N_4152,In_1139,In_916);
nand U4153 (N_4153,In_712,In_541);
nand U4154 (N_4154,In_562,In_1093);
and U4155 (N_4155,In_1238,In_409);
nand U4156 (N_4156,In_1282,In_969);
and U4157 (N_4157,In_1318,In_1103);
nor U4158 (N_4158,In_338,In_113);
nand U4159 (N_4159,In_849,In_902);
and U4160 (N_4160,In_67,In_555);
or U4161 (N_4161,In_968,In_470);
xnor U4162 (N_4162,In_137,In_10);
and U4163 (N_4163,In_1006,In_1264);
nand U4164 (N_4164,In_827,In_1435);
nor U4165 (N_4165,In_960,In_308);
nor U4166 (N_4166,In_962,In_247);
xor U4167 (N_4167,In_416,In_45);
xnor U4168 (N_4168,In_464,In_743);
and U4169 (N_4169,In_611,In_156);
xor U4170 (N_4170,In_546,In_2);
nand U4171 (N_4171,In_721,In_330);
nor U4172 (N_4172,In_1455,In_448);
nor U4173 (N_4173,In_1331,In_1081);
xor U4174 (N_4174,In_401,In_1369);
or U4175 (N_4175,In_1479,In_80);
nor U4176 (N_4176,In_660,In_470);
nand U4177 (N_4177,In_1333,In_998);
nor U4178 (N_4178,In_989,In_1195);
nand U4179 (N_4179,In_950,In_928);
and U4180 (N_4180,In_880,In_518);
nand U4181 (N_4181,In_1056,In_824);
nand U4182 (N_4182,In_514,In_454);
nor U4183 (N_4183,In_520,In_693);
nand U4184 (N_4184,In_210,In_937);
and U4185 (N_4185,In_1155,In_672);
or U4186 (N_4186,In_36,In_1183);
or U4187 (N_4187,In_896,In_760);
nand U4188 (N_4188,In_684,In_540);
or U4189 (N_4189,In_1271,In_243);
nor U4190 (N_4190,In_956,In_748);
nand U4191 (N_4191,In_676,In_63);
xor U4192 (N_4192,In_1114,In_1179);
xnor U4193 (N_4193,In_627,In_1109);
xor U4194 (N_4194,In_267,In_367);
or U4195 (N_4195,In_343,In_149);
nor U4196 (N_4196,In_1124,In_1163);
and U4197 (N_4197,In_1236,In_70);
nand U4198 (N_4198,In_1082,In_386);
and U4199 (N_4199,In_312,In_674);
nor U4200 (N_4200,In_977,In_664);
nor U4201 (N_4201,In_1434,In_1046);
or U4202 (N_4202,In_1247,In_140);
or U4203 (N_4203,In_671,In_884);
or U4204 (N_4204,In_1464,In_794);
xnor U4205 (N_4205,In_247,In_115);
nand U4206 (N_4206,In_1314,In_1315);
or U4207 (N_4207,In_36,In_122);
xnor U4208 (N_4208,In_971,In_282);
nor U4209 (N_4209,In_1261,In_122);
nand U4210 (N_4210,In_782,In_773);
nand U4211 (N_4211,In_117,In_380);
and U4212 (N_4212,In_1062,In_567);
and U4213 (N_4213,In_1369,In_1050);
nor U4214 (N_4214,In_86,In_543);
nor U4215 (N_4215,In_729,In_515);
xnor U4216 (N_4216,In_366,In_1399);
xnor U4217 (N_4217,In_203,In_1477);
nand U4218 (N_4218,In_554,In_1273);
nor U4219 (N_4219,In_1328,In_785);
or U4220 (N_4220,In_242,In_230);
nor U4221 (N_4221,In_870,In_52);
or U4222 (N_4222,In_231,In_964);
nor U4223 (N_4223,In_1438,In_1033);
or U4224 (N_4224,In_208,In_278);
and U4225 (N_4225,In_1149,In_702);
or U4226 (N_4226,In_28,In_167);
or U4227 (N_4227,In_213,In_165);
or U4228 (N_4228,In_721,In_205);
xor U4229 (N_4229,In_450,In_1162);
and U4230 (N_4230,In_179,In_962);
and U4231 (N_4231,In_267,In_138);
nor U4232 (N_4232,In_323,In_630);
xnor U4233 (N_4233,In_1497,In_1162);
xnor U4234 (N_4234,In_180,In_87);
and U4235 (N_4235,In_1154,In_528);
nor U4236 (N_4236,In_532,In_926);
nor U4237 (N_4237,In_306,In_184);
and U4238 (N_4238,In_498,In_1420);
and U4239 (N_4239,In_1390,In_744);
and U4240 (N_4240,In_927,In_684);
nor U4241 (N_4241,In_455,In_1184);
xnor U4242 (N_4242,In_187,In_84);
xnor U4243 (N_4243,In_1295,In_1498);
nand U4244 (N_4244,In_877,In_541);
or U4245 (N_4245,In_100,In_519);
or U4246 (N_4246,In_267,In_1102);
nand U4247 (N_4247,In_168,In_573);
xnor U4248 (N_4248,In_187,In_1477);
nor U4249 (N_4249,In_178,In_213);
or U4250 (N_4250,In_494,In_71);
nand U4251 (N_4251,In_221,In_589);
and U4252 (N_4252,In_57,In_1148);
or U4253 (N_4253,In_178,In_403);
nand U4254 (N_4254,In_228,In_327);
or U4255 (N_4255,In_1430,In_923);
or U4256 (N_4256,In_693,In_275);
nor U4257 (N_4257,In_1017,In_710);
or U4258 (N_4258,In_1271,In_1389);
nand U4259 (N_4259,In_1408,In_1428);
nand U4260 (N_4260,In_515,In_1022);
or U4261 (N_4261,In_855,In_1106);
or U4262 (N_4262,In_896,In_256);
xnor U4263 (N_4263,In_882,In_1003);
nand U4264 (N_4264,In_1400,In_126);
nor U4265 (N_4265,In_1398,In_482);
xnor U4266 (N_4266,In_966,In_48);
xnor U4267 (N_4267,In_1278,In_47);
nor U4268 (N_4268,In_139,In_1058);
nand U4269 (N_4269,In_1484,In_451);
nor U4270 (N_4270,In_1484,In_1066);
and U4271 (N_4271,In_1116,In_207);
xor U4272 (N_4272,In_1048,In_646);
nor U4273 (N_4273,In_728,In_106);
or U4274 (N_4274,In_311,In_1079);
nand U4275 (N_4275,In_1339,In_904);
nand U4276 (N_4276,In_389,In_823);
nor U4277 (N_4277,In_1412,In_239);
and U4278 (N_4278,In_406,In_710);
or U4279 (N_4279,In_638,In_707);
and U4280 (N_4280,In_1356,In_11);
or U4281 (N_4281,In_1287,In_825);
and U4282 (N_4282,In_1107,In_851);
or U4283 (N_4283,In_693,In_240);
xor U4284 (N_4284,In_116,In_390);
xor U4285 (N_4285,In_844,In_639);
and U4286 (N_4286,In_406,In_854);
or U4287 (N_4287,In_1457,In_829);
and U4288 (N_4288,In_944,In_1375);
nand U4289 (N_4289,In_1321,In_1339);
and U4290 (N_4290,In_364,In_758);
nor U4291 (N_4291,In_696,In_401);
or U4292 (N_4292,In_390,In_762);
nand U4293 (N_4293,In_562,In_143);
xnor U4294 (N_4294,In_790,In_58);
and U4295 (N_4295,In_936,In_876);
xor U4296 (N_4296,In_1304,In_1296);
nand U4297 (N_4297,In_105,In_804);
nand U4298 (N_4298,In_65,In_1121);
nand U4299 (N_4299,In_1265,In_829);
and U4300 (N_4300,In_989,In_108);
xor U4301 (N_4301,In_1109,In_1058);
nor U4302 (N_4302,In_476,In_1013);
and U4303 (N_4303,In_1014,In_325);
or U4304 (N_4304,In_866,In_1056);
or U4305 (N_4305,In_518,In_1029);
nor U4306 (N_4306,In_255,In_542);
nor U4307 (N_4307,In_206,In_897);
or U4308 (N_4308,In_109,In_270);
and U4309 (N_4309,In_230,In_153);
xor U4310 (N_4310,In_1434,In_646);
or U4311 (N_4311,In_879,In_1076);
nor U4312 (N_4312,In_308,In_774);
nand U4313 (N_4313,In_1062,In_947);
nand U4314 (N_4314,In_1268,In_667);
and U4315 (N_4315,In_257,In_18);
nand U4316 (N_4316,In_638,In_1489);
xor U4317 (N_4317,In_619,In_1163);
xnor U4318 (N_4318,In_389,In_440);
nand U4319 (N_4319,In_194,In_1275);
nor U4320 (N_4320,In_28,In_1018);
and U4321 (N_4321,In_98,In_1278);
or U4322 (N_4322,In_1008,In_516);
nand U4323 (N_4323,In_1478,In_976);
xnor U4324 (N_4324,In_1336,In_644);
or U4325 (N_4325,In_1419,In_751);
or U4326 (N_4326,In_1039,In_1423);
xor U4327 (N_4327,In_182,In_939);
nor U4328 (N_4328,In_454,In_1058);
nand U4329 (N_4329,In_355,In_949);
xnor U4330 (N_4330,In_1075,In_526);
nand U4331 (N_4331,In_913,In_463);
xnor U4332 (N_4332,In_717,In_159);
nor U4333 (N_4333,In_421,In_325);
nand U4334 (N_4334,In_575,In_120);
nand U4335 (N_4335,In_1044,In_1274);
and U4336 (N_4336,In_280,In_1106);
xnor U4337 (N_4337,In_613,In_766);
nor U4338 (N_4338,In_343,In_543);
nand U4339 (N_4339,In_1147,In_1434);
xnor U4340 (N_4340,In_1068,In_1243);
and U4341 (N_4341,In_1415,In_110);
xnor U4342 (N_4342,In_953,In_254);
or U4343 (N_4343,In_76,In_1059);
xor U4344 (N_4344,In_363,In_697);
nand U4345 (N_4345,In_743,In_175);
and U4346 (N_4346,In_1249,In_1156);
or U4347 (N_4347,In_1072,In_770);
nor U4348 (N_4348,In_24,In_136);
or U4349 (N_4349,In_1144,In_469);
nor U4350 (N_4350,In_795,In_165);
nand U4351 (N_4351,In_484,In_874);
nand U4352 (N_4352,In_199,In_48);
or U4353 (N_4353,In_1424,In_1389);
xor U4354 (N_4354,In_188,In_502);
xnor U4355 (N_4355,In_1163,In_395);
nor U4356 (N_4356,In_1124,In_290);
and U4357 (N_4357,In_158,In_507);
nor U4358 (N_4358,In_310,In_117);
or U4359 (N_4359,In_1161,In_374);
xnor U4360 (N_4360,In_107,In_1111);
nand U4361 (N_4361,In_513,In_48);
or U4362 (N_4362,In_1451,In_634);
nand U4363 (N_4363,In_1137,In_333);
nor U4364 (N_4364,In_955,In_1191);
xor U4365 (N_4365,In_1300,In_648);
nor U4366 (N_4366,In_1046,In_74);
and U4367 (N_4367,In_451,In_1130);
xor U4368 (N_4368,In_66,In_194);
or U4369 (N_4369,In_874,In_794);
nor U4370 (N_4370,In_1307,In_818);
xnor U4371 (N_4371,In_173,In_151);
or U4372 (N_4372,In_527,In_590);
or U4373 (N_4373,In_262,In_1283);
nor U4374 (N_4374,In_1353,In_124);
nor U4375 (N_4375,In_384,In_1461);
and U4376 (N_4376,In_1491,In_1162);
nor U4377 (N_4377,In_1236,In_678);
and U4378 (N_4378,In_957,In_624);
or U4379 (N_4379,In_1455,In_472);
xnor U4380 (N_4380,In_864,In_629);
xor U4381 (N_4381,In_494,In_105);
nor U4382 (N_4382,In_484,In_795);
or U4383 (N_4383,In_1216,In_1013);
or U4384 (N_4384,In_1265,In_751);
or U4385 (N_4385,In_1337,In_1456);
and U4386 (N_4386,In_682,In_236);
and U4387 (N_4387,In_474,In_122);
and U4388 (N_4388,In_830,In_147);
or U4389 (N_4389,In_1281,In_414);
and U4390 (N_4390,In_1147,In_561);
nor U4391 (N_4391,In_279,In_985);
nand U4392 (N_4392,In_258,In_247);
nor U4393 (N_4393,In_1495,In_1447);
and U4394 (N_4394,In_295,In_93);
nor U4395 (N_4395,In_1468,In_186);
and U4396 (N_4396,In_664,In_982);
and U4397 (N_4397,In_201,In_245);
or U4398 (N_4398,In_427,In_1333);
and U4399 (N_4399,In_1216,In_215);
nand U4400 (N_4400,In_20,In_1040);
and U4401 (N_4401,In_582,In_1388);
xnor U4402 (N_4402,In_17,In_722);
nor U4403 (N_4403,In_1199,In_741);
or U4404 (N_4404,In_560,In_469);
nor U4405 (N_4405,In_1468,In_843);
nor U4406 (N_4406,In_372,In_688);
nand U4407 (N_4407,In_598,In_352);
xor U4408 (N_4408,In_1260,In_321);
xor U4409 (N_4409,In_701,In_1203);
xor U4410 (N_4410,In_387,In_1413);
xnor U4411 (N_4411,In_340,In_1302);
xnor U4412 (N_4412,In_478,In_427);
or U4413 (N_4413,In_913,In_634);
nand U4414 (N_4414,In_1448,In_294);
nor U4415 (N_4415,In_1090,In_180);
xor U4416 (N_4416,In_1400,In_895);
nor U4417 (N_4417,In_1150,In_931);
nor U4418 (N_4418,In_1228,In_864);
and U4419 (N_4419,In_1397,In_136);
nand U4420 (N_4420,In_1005,In_1334);
or U4421 (N_4421,In_720,In_142);
nand U4422 (N_4422,In_1178,In_968);
or U4423 (N_4423,In_532,In_1088);
xnor U4424 (N_4424,In_1188,In_918);
or U4425 (N_4425,In_1425,In_471);
xnor U4426 (N_4426,In_1407,In_1065);
nand U4427 (N_4427,In_875,In_42);
or U4428 (N_4428,In_1158,In_586);
and U4429 (N_4429,In_1163,In_1149);
xnor U4430 (N_4430,In_952,In_543);
nand U4431 (N_4431,In_363,In_811);
and U4432 (N_4432,In_597,In_481);
nand U4433 (N_4433,In_853,In_1117);
or U4434 (N_4434,In_746,In_885);
nor U4435 (N_4435,In_1003,In_403);
nor U4436 (N_4436,In_845,In_1328);
xor U4437 (N_4437,In_600,In_468);
and U4438 (N_4438,In_384,In_921);
and U4439 (N_4439,In_543,In_12);
xor U4440 (N_4440,In_144,In_199);
and U4441 (N_4441,In_1047,In_981);
nor U4442 (N_4442,In_756,In_922);
or U4443 (N_4443,In_886,In_497);
xor U4444 (N_4444,In_785,In_610);
nand U4445 (N_4445,In_855,In_1020);
or U4446 (N_4446,In_1347,In_1259);
nand U4447 (N_4447,In_1192,In_770);
nor U4448 (N_4448,In_1235,In_895);
nor U4449 (N_4449,In_374,In_1013);
or U4450 (N_4450,In_114,In_948);
or U4451 (N_4451,In_728,In_1181);
nand U4452 (N_4452,In_522,In_1225);
xnor U4453 (N_4453,In_992,In_1230);
nand U4454 (N_4454,In_79,In_61);
xor U4455 (N_4455,In_343,In_814);
nor U4456 (N_4456,In_682,In_55);
xnor U4457 (N_4457,In_909,In_925);
or U4458 (N_4458,In_336,In_543);
nand U4459 (N_4459,In_667,In_162);
and U4460 (N_4460,In_1319,In_588);
or U4461 (N_4461,In_253,In_1228);
and U4462 (N_4462,In_215,In_1254);
or U4463 (N_4463,In_1227,In_1456);
or U4464 (N_4464,In_952,In_1186);
or U4465 (N_4465,In_731,In_198);
nand U4466 (N_4466,In_736,In_1030);
nor U4467 (N_4467,In_600,In_212);
nand U4468 (N_4468,In_1387,In_1022);
and U4469 (N_4469,In_512,In_912);
and U4470 (N_4470,In_1144,In_1408);
xor U4471 (N_4471,In_1084,In_1338);
nand U4472 (N_4472,In_1130,In_1281);
and U4473 (N_4473,In_1436,In_558);
nor U4474 (N_4474,In_203,In_370);
xor U4475 (N_4475,In_1442,In_1353);
or U4476 (N_4476,In_1313,In_25);
nand U4477 (N_4477,In_84,In_377);
and U4478 (N_4478,In_49,In_791);
xor U4479 (N_4479,In_792,In_591);
or U4480 (N_4480,In_108,In_1029);
and U4481 (N_4481,In_1008,In_378);
nor U4482 (N_4482,In_36,In_605);
nand U4483 (N_4483,In_1288,In_285);
nand U4484 (N_4484,In_462,In_638);
xor U4485 (N_4485,In_1492,In_965);
nand U4486 (N_4486,In_1163,In_558);
xnor U4487 (N_4487,In_185,In_1209);
xor U4488 (N_4488,In_645,In_1017);
and U4489 (N_4489,In_1403,In_766);
nand U4490 (N_4490,In_1278,In_502);
and U4491 (N_4491,In_387,In_1179);
or U4492 (N_4492,In_71,In_471);
xor U4493 (N_4493,In_384,In_325);
nor U4494 (N_4494,In_1268,In_1485);
and U4495 (N_4495,In_179,In_255);
xnor U4496 (N_4496,In_1049,In_508);
xnor U4497 (N_4497,In_974,In_294);
or U4498 (N_4498,In_1332,In_758);
and U4499 (N_4499,In_1411,In_472);
nor U4500 (N_4500,In_20,In_1139);
xor U4501 (N_4501,In_208,In_338);
nor U4502 (N_4502,In_1357,In_1189);
and U4503 (N_4503,In_411,In_1125);
nand U4504 (N_4504,In_118,In_202);
xnor U4505 (N_4505,In_256,In_560);
nor U4506 (N_4506,In_537,In_125);
nor U4507 (N_4507,In_1185,In_956);
xnor U4508 (N_4508,In_130,In_198);
xnor U4509 (N_4509,In_231,In_1017);
and U4510 (N_4510,In_412,In_565);
or U4511 (N_4511,In_136,In_1003);
nand U4512 (N_4512,In_1026,In_1283);
nand U4513 (N_4513,In_1463,In_858);
and U4514 (N_4514,In_330,In_1296);
or U4515 (N_4515,In_863,In_1139);
and U4516 (N_4516,In_1184,In_292);
or U4517 (N_4517,In_1322,In_1251);
or U4518 (N_4518,In_172,In_1099);
nor U4519 (N_4519,In_1187,In_788);
nor U4520 (N_4520,In_770,In_1285);
and U4521 (N_4521,In_568,In_1368);
xnor U4522 (N_4522,In_1374,In_1254);
and U4523 (N_4523,In_597,In_1486);
nor U4524 (N_4524,In_1478,In_1314);
xnor U4525 (N_4525,In_982,In_170);
and U4526 (N_4526,In_906,In_438);
nor U4527 (N_4527,In_512,In_1060);
and U4528 (N_4528,In_471,In_673);
nor U4529 (N_4529,In_1023,In_1346);
or U4530 (N_4530,In_706,In_1033);
and U4531 (N_4531,In_1330,In_897);
nand U4532 (N_4532,In_626,In_1111);
and U4533 (N_4533,In_792,In_349);
and U4534 (N_4534,In_1123,In_689);
nor U4535 (N_4535,In_38,In_590);
nor U4536 (N_4536,In_885,In_1435);
and U4537 (N_4537,In_1147,In_952);
nor U4538 (N_4538,In_1114,In_61);
nor U4539 (N_4539,In_1134,In_1291);
xnor U4540 (N_4540,In_1052,In_1125);
nor U4541 (N_4541,In_908,In_365);
and U4542 (N_4542,In_154,In_770);
xnor U4543 (N_4543,In_952,In_1077);
nand U4544 (N_4544,In_1092,In_1459);
or U4545 (N_4545,In_294,In_1176);
nor U4546 (N_4546,In_625,In_413);
xor U4547 (N_4547,In_648,In_1152);
and U4548 (N_4548,In_1427,In_184);
and U4549 (N_4549,In_1489,In_798);
or U4550 (N_4550,In_159,In_26);
nor U4551 (N_4551,In_665,In_789);
and U4552 (N_4552,In_1393,In_1228);
nor U4553 (N_4553,In_560,In_1338);
xor U4554 (N_4554,In_27,In_486);
and U4555 (N_4555,In_11,In_322);
nor U4556 (N_4556,In_396,In_561);
nor U4557 (N_4557,In_177,In_360);
nor U4558 (N_4558,In_433,In_410);
or U4559 (N_4559,In_582,In_322);
or U4560 (N_4560,In_1183,In_1417);
and U4561 (N_4561,In_131,In_922);
nor U4562 (N_4562,In_380,In_504);
nand U4563 (N_4563,In_203,In_85);
or U4564 (N_4564,In_681,In_521);
and U4565 (N_4565,In_133,In_370);
xnor U4566 (N_4566,In_986,In_720);
or U4567 (N_4567,In_336,In_432);
nand U4568 (N_4568,In_981,In_1495);
and U4569 (N_4569,In_1304,In_810);
nand U4570 (N_4570,In_954,In_1328);
and U4571 (N_4571,In_173,In_919);
or U4572 (N_4572,In_412,In_417);
and U4573 (N_4573,In_1074,In_1197);
and U4574 (N_4574,In_1424,In_93);
or U4575 (N_4575,In_1474,In_860);
and U4576 (N_4576,In_1197,In_1418);
or U4577 (N_4577,In_808,In_35);
or U4578 (N_4578,In_1126,In_107);
nand U4579 (N_4579,In_855,In_1064);
or U4580 (N_4580,In_73,In_249);
or U4581 (N_4581,In_105,In_1497);
and U4582 (N_4582,In_438,In_614);
nand U4583 (N_4583,In_1482,In_149);
xnor U4584 (N_4584,In_1261,In_817);
nand U4585 (N_4585,In_768,In_88);
and U4586 (N_4586,In_114,In_753);
or U4587 (N_4587,In_1469,In_237);
and U4588 (N_4588,In_878,In_476);
xnor U4589 (N_4589,In_632,In_410);
or U4590 (N_4590,In_1336,In_799);
nand U4591 (N_4591,In_478,In_1015);
or U4592 (N_4592,In_351,In_148);
nand U4593 (N_4593,In_1405,In_1143);
nand U4594 (N_4594,In_1284,In_197);
nand U4595 (N_4595,In_6,In_1485);
xnor U4596 (N_4596,In_82,In_189);
and U4597 (N_4597,In_1008,In_635);
or U4598 (N_4598,In_1161,In_1027);
or U4599 (N_4599,In_976,In_133);
nand U4600 (N_4600,In_1402,In_814);
nand U4601 (N_4601,In_1028,In_49);
or U4602 (N_4602,In_711,In_996);
nor U4603 (N_4603,In_1234,In_473);
and U4604 (N_4604,In_481,In_1052);
or U4605 (N_4605,In_188,In_1324);
xor U4606 (N_4606,In_1437,In_814);
xnor U4607 (N_4607,In_9,In_1109);
and U4608 (N_4608,In_46,In_1153);
nor U4609 (N_4609,In_83,In_969);
or U4610 (N_4610,In_722,In_579);
xor U4611 (N_4611,In_207,In_1292);
xnor U4612 (N_4612,In_861,In_1198);
nor U4613 (N_4613,In_1386,In_280);
nand U4614 (N_4614,In_1396,In_1228);
or U4615 (N_4615,In_998,In_231);
xnor U4616 (N_4616,In_1475,In_897);
nor U4617 (N_4617,In_187,In_838);
and U4618 (N_4618,In_823,In_1204);
and U4619 (N_4619,In_846,In_135);
xor U4620 (N_4620,In_633,In_78);
xor U4621 (N_4621,In_530,In_1351);
xnor U4622 (N_4622,In_897,In_1379);
or U4623 (N_4623,In_115,In_1441);
nor U4624 (N_4624,In_1394,In_1329);
xor U4625 (N_4625,In_793,In_39);
nand U4626 (N_4626,In_638,In_83);
or U4627 (N_4627,In_1233,In_507);
or U4628 (N_4628,In_1107,In_1347);
nor U4629 (N_4629,In_408,In_1494);
nand U4630 (N_4630,In_53,In_837);
nor U4631 (N_4631,In_707,In_417);
xor U4632 (N_4632,In_577,In_1317);
and U4633 (N_4633,In_1219,In_558);
nand U4634 (N_4634,In_345,In_973);
or U4635 (N_4635,In_1376,In_79);
nand U4636 (N_4636,In_825,In_158);
xor U4637 (N_4637,In_989,In_485);
and U4638 (N_4638,In_36,In_1452);
nand U4639 (N_4639,In_607,In_374);
xnor U4640 (N_4640,In_242,In_696);
nor U4641 (N_4641,In_1488,In_1112);
nand U4642 (N_4642,In_137,In_1342);
nor U4643 (N_4643,In_241,In_291);
and U4644 (N_4644,In_1092,In_54);
xor U4645 (N_4645,In_892,In_584);
nor U4646 (N_4646,In_264,In_635);
nor U4647 (N_4647,In_1244,In_1364);
nor U4648 (N_4648,In_1352,In_388);
nor U4649 (N_4649,In_404,In_396);
xor U4650 (N_4650,In_685,In_1262);
or U4651 (N_4651,In_1287,In_1187);
or U4652 (N_4652,In_1339,In_691);
and U4653 (N_4653,In_718,In_467);
xor U4654 (N_4654,In_1073,In_517);
xnor U4655 (N_4655,In_888,In_1475);
nor U4656 (N_4656,In_1472,In_840);
nor U4657 (N_4657,In_192,In_937);
nor U4658 (N_4658,In_592,In_1452);
and U4659 (N_4659,In_448,In_1469);
nand U4660 (N_4660,In_458,In_1396);
xnor U4661 (N_4661,In_1228,In_264);
nor U4662 (N_4662,In_795,In_1067);
nor U4663 (N_4663,In_1235,In_297);
or U4664 (N_4664,In_1140,In_164);
or U4665 (N_4665,In_1076,In_52);
xnor U4666 (N_4666,In_1132,In_122);
nand U4667 (N_4667,In_503,In_740);
and U4668 (N_4668,In_421,In_1390);
nand U4669 (N_4669,In_124,In_962);
xnor U4670 (N_4670,In_854,In_143);
nor U4671 (N_4671,In_941,In_570);
xor U4672 (N_4672,In_885,In_28);
or U4673 (N_4673,In_939,In_1482);
or U4674 (N_4674,In_171,In_1199);
xor U4675 (N_4675,In_470,In_936);
and U4676 (N_4676,In_1183,In_849);
xnor U4677 (N_4677,In_601,In_908);
nor U4678 (N_4678,In_1434,In_121);
xor U4679 (N_4679,In_1064,In_1056);
xor U4680 (N_4680,In_1045,In_1249);
nand U4681 (N_4681,In_369,In_597);
nand U4682 (N_4682,In_1413,In_461);
and U4683 (N_4683,In_1366,In_1321);
and U4684 (N_4684,In_1132,In_1116);
nand U4685 (N_4685,In_1244,In_1004);
nand U4686 (N_4686,In_922,In_1000);
nand U4687 (N_4687,In_368,In_11);
xor U4688 (N_4688,In_1475,In_1111);
and U4689 (N_4689,In_1269,In_1252);
or U4690 (N_4690,In_1034,In_850);
or U4691 (N_4691,In_431,In_1450);
nand U4692 (N_4692,In_1051,In_49);
nor U4693 (N_4693,In_1148,In_410);
nand U4694 (N_4694,In_1120,In_29);
or U4695 (N_4695,In_912,In_1096);
and U4696 (N_4696,In_1360,In_1098);
nor U4697 (N_4697,In_973,In_1407);
nand U4698 (N_4698,In_50,In_405);
or U4699 (N_4699,In_1456,In_1051);
nand U4700 (N_4700,In_983,In_763);
or U4701 (N_4701,In_212,In_200);
nor U4702 (N_4702,In_1135,In_1169);
or U4703 (N_4703,In_49,In_972);
nand U4704 (N_4704,In_1269,In_1389);
and U4705 (N_4705,In_663,In_1338);
or U4706 (N_4706,In_466,In_772);
xor U4707 (N_4707,In_714,In_1042);
nand U4708 (N_4708,In_1375,In_1444);
nand U4709 (N_4709,In_897,In_1137);
nand U4710 (N_4710,In_1349,In_1474);
xnor U4711 (N_4711,In_234,In_78);
and U4712 (N_4712,In_985,In_978);
or U4713 (N_4713,In_462,In_404);
or U4714 (N_4714,In_118,In_454);
xnor U4715 (N_4715,In_1203,In_1151);
xor U4716 (N_4716,In_1389,In_1428);
nor U4717 (N_4717,In_933,In_309);
and U4718 (N_4718,In_365,In_141);
nand U4719 (N_4719,In_1122,In_162);
nor U4720 (N_4720,In_1378,In_601);
nand U4721 (N_4721,In_174,In_1403);
or U4722 (N_4722,In_1096,In_729);
nor U4723 (N_4723,In_85,In_548);
and U4724 (N_4724,In_526,In_1289);
and U4725 (N_4725,In_909,In_707);
nor U4726 (N_4726,In_1088,In_246);
and U4727 (N_4727,In_411,In_1121);
xor U4728 (N_4728,In_1259,In_911);
and U4729 (N_4729,In_184,In_207);
xor U4730 (N_4730,In_688,In_824);
xnor U4731 (N_4731,In_649,In_208);
or U4732 (N_4732,In_965,In_437);
nor U4733 (N_4733,In_863,In_782);
nor U4734 (N_4734,In_1494,In_1186);
nor U4735 (N_4735,In_966,In_258);
xor U4736 (N_4736,In_586,In_104);
nand U4737 (N_4737,In_718,In_34);
xor U4738 (N_4738,In_1253,In_1083);
xor U4739 (N_4739,In_1010,In_1113);
or U4740 (N_4740,In_912,In_1130);
or U4741 (N_4741,In_824,In_790);
and U4742 (N_4742,In_376,In_1462);
and U4743 (N_4743,In_1427,In_625);
xnor U4744 (N_4744,In_675,In_1153);
nor U4745 (N_4745,In_679,In_1424);
nand U4746 (N_4746,In_1486,In_1183);
xor U4747 (N_4747,In_279,In_1415);
or U4748 (N_4748,In_563,In_1464);
and U4749 (N_4749,In_973,In_108);
xor U4750 (N_4750,In_894,In_982);
nand U4751 (N_4751,In_706,In_1481);
nor U4752 (N_4752,In_65,In_1471);
nor U4753 (N_4753,In_1327,In_1010);
or U4754 (N_4754,In_427,In_433);
nor U4755 (N_4755,In_1050,In_205);
nand U4756 (N_4756,In_640,In_1499);
or U4757 (N_4757,In_1494,In_1396);
and U4758 (N_4758,In_445,In_1161);
xnor U4759 (N_4759,In_506,In_1007);
nor U4760 (N_4760,In_1346,In_65);
nand U4761 (N_4761,In_575,In_373);
and U4762 (N_4762,In_669,In_925);
nand U4763 (N_4763,In_1015,In_901);
xor U4764 (N_4764,In_400,In_64);
nor U4765 (N_4765,In_297,In_939);
nand U4766 (N_4766,In_1109,In_1351);
and U4767 (N_4767,In_259,In_25);
and U4768 (N_4768,In_1255,In_99);
xnor U4769 (N_4769,In_90,In_1358);
and U4770 (N_4770,In_1320,In_1073);
nor U4771 (N_4771,In_689,In_1376);
nand U4772 (N_4772,In_556,In_580);
nor U4773 (N_4773,In_438,In_208);
nand U4774 (N_4774,In_346,In_1314);
and U4775 (N_4775,In_747,In_1491);
and U4776 (N_4776,In_88,In_883);
xor U4777 (N_4777,In_13,In_750);
nor U4778 (N_4778,In_717,In_742);
and U4779 (N_4779,In_48,In_709);
nor U4780 (N_4780,In_1089,In_1463);
nand U4781 (N_4781,In_908,In_466);
nand U4782 (N_4782,In_44,In_994);
nor U4783 (N_4783,In_960,In_1441);
and U4784 (N_4784,In_643,In_969);
nand U4785 (N_4785,In_651,In_1392);
xor U4786 (N_4786,In_1083,In_914);
nor U4787 (N_4787,In_1253,In_809);
nor U4788 (N_4788,In_694,In_1353);
nor U4789 (N_4789,In_392,In_1082);
xnor U4790 (N_4790,In_713,In_79);
xnor U4791 (N_4791,In_1279,In_1274);
and U4792 (N_4792,In_518,In_725);
nor U4793 (N_4793,In_1115,In_1208);
xnor U4794 (N_4794,In_558,In_1247);
nand U4795 (N_4795,In_1250,In_284);
and U4796 (N_4796,In_1062,In_334);
nand U4797 (N_4797,In_281,In_432);
nor U4798 (N_4798,In_1480,In_818);
nor U4799 (N_4799,In_1052,In_1406);
and U4800 (N_4800,In_985,In_495);
and U4801 (N_4801,In_942,In_986);
nand U4802 (N_4802,In_295,In_479);
nand U4803 (N_4803,In_890,In_687);
and U4804 (N_4804,In_580,In_996);
nand U4805 (N_4805,In_1232,In_749);
nor U4806 (N_4806,In_955,In_50);
nor U4807 (N_4807,In_1228,In_1171);
nor U4808 (N_4808,In_848,In_1053);
nand U4809 (N_4809,In_1217,In_1083);
and U4810 (N_4810,In_1130,In_270);
and U4811 (N_4811,In_70,In_29);
and U4812 (N_4812,In_1080,In_1194);
nand U4813 (N_4813,In_162,In_943);
or U4814 (N_4814,In_702,In_1306);
or U4815 (N_4815,In_1110,In_409);
nor U4816 (N_4816,In_73,In_506);
nor U4817 (N_4817,In_1012,In_26);
nor U4818 (N_4818,In_978,In_747);
nor U4819 (N_4819,In_811,In_1279);
and U4820 (N_4820,In_1014,In_1056);
nand U4821 (N_4821,In_1253,In_69);
or U4822 (N_4822,In_1039,In_1380);
nand U4823 (N_4823,In_130,In_1300);
nand U4824 (N_4824,In_806,In_1111);
nor U4825 (N_4825,In_792,In_1235);
or U4826 (N_4826,In_439,In_669);
and U4827 (N_4827,In_304,In_431);
nor U4828 (N_4828,In_1334,In_442);
nor U4829 (N_4829,In_1057,In_548);
nor U4830 (N_4830,In_1058,In_50);
and U4831 (N_4831,In_667,In_302);
nand U4832 (N_4832,In_648,In_413);
or U4833 (N_4833,In_139,In_364);
or U4834 (N_4834,In_1177,In_785);
and U4835 (N_4835,In_474,In_735);
or U4836 (N_4836,In_1484,In_637);
and U4837 (N_4837,In_1451,In_994);
nand U4838 (N_4838,In_1488,In_727);
or U4839 (N_4839,In_1399,In_1484);
xor U4840 (N_4840,In_871,In_1027);
and U4841 (N_4841,In_374,In_793);
nand U4842 (N_4842,In_1492,In_959);
nor U4843 (N_4843,In_1110,In_945);
xor U4844 (N_4844,In_398,In_201);
or U4845 (N_4845,In_1082,In_13);
and U4846 (N_4846,In_1453,In_744);
xor U4847 (N_4847,In_637,In_168);
nand U4848 (N_4848,In_629,In_236);
xor U4849 (N_4849,In_934,In_1167);
or U4850 (N_4850,In_331,In_89);
nor U4851 (N_4851,In_19,In_320);
nand U4852 (N_4852,In_635,In_916);
nor U4853 (N_4853,In_401,In_1136);
and U4854 (N_4854,In_201,In_101);
and U4855 (N_4855,In_896,In_39);
and U4856 (N_4856,In_486,In_1212);
and U4857 (N_4857,In_793,In_486);
nor U4858 (N_4858,In_441,In_517);
nor U4859 (N_4859,In_738,In_659);
or U4860 (N_4860,In_1476,In_1288);
or U4861 (N_4861,In_17,In_571);
xnor U4862 (N_4862,In_1480,In_643);
nor U4863 (N_4863,In_1397,In_171);
and U4864 (N_4864,In_68,In_616);
or U4865 (N_4865,In_568,In_582);
xor U4866 (N_4866,In_457,In_504);
nand U4867 (N_4867,In_485,In_1225);
and U4868 (N_4868,In_1380,In_1047);
or U4869 (N_4869,In_1138,In_489);
nand U4870 (N_4870,In_1136,In_831);
or U4871 (N_4871,In_215,In_1403);
and U4872 (N_4872,In_1352,In_905);
xnor U4873 (N_4873,In_213,In_1187);
nor U4874 (N_4874,In_356,In_695);
or U4875 (N_4875,In_237,In_657);
nand U4876 (N_4876,In_757,In_444);
or U4877 (N_4877,In_1206,In_1189);
xor U4878 (N_4878,In_632,In_374);
nand U4879 (N_4879,In_922,In_562);
nor U4880 (N_4880,In_1427,In_885);
nor U4881 (N_4881,In_493,In_328);
xnor U4882 (N_4882,In_112,In_719);
and U4883 (N_4883,In_864,In_1174);
or U4884 (N_4884,In_109,In_1374);
or U4885 (N_4885,In_592,In_761);
nand U4886 (N_4886,In_1194,In_501);
nand U4887 (N_4887,In_439,In_1127);
nor U4888 (N_4888,In_285,In_1339);
and U4889 (N_4889,In_221,In_1464);
nand U4890 (N_4890,In_125,In_820);
nor U4891 (N_4891,In_1293,In_685);
nand U4892 (N_4892,In_1045,In_456);
or U4893 (N_4893,In_968,In_474);
nand U4894 (N_4894,In_806,In_754);
nand U4895 (N_4895,In_481,In_803);
and U4896 (N_4896,In_524,In_961);
nand U4897 (N_4897,In_967,In_85);
or U4898 (N_4898,In_445,In_477);
and U4899 (N_4899,In_1005,In_586);
and U4900 (N_4900,In_1037,In_1498);
nor U4901 (N_4901,In_188,In_141);
and U4902 (N_4902,In_688,In_576);
or U4903 (N_4903,In_1282,In_132);
nand U4904 (N_4904,In_1128,In_740);
xor U4905 (N_4905,In_72,In_906);
xor U4906 (N_4906,In_348,In_1124);
xnor U4907 (N_4907,In_1376,In_21);
nand U4908 (N_4908,In_115,In_765);
or U4909 (N_4909,In_562,In_1372);
nand U4910 (N_4910,In_1488,In_90);
or U4911 (N_4911,In_772,In_1385);
and U4912 (N_4912,In_286,In_253);
or U4913 (N_4913,In_1012,In_884);
xor U4914 (N_4914,In_289,In_874);
nand U4915 (N_4915,In_856,In_198);
nand U4916 (N_4916,In_340,In_1439);
or U4917 (N_4917,In_682,In_249);
and U4918 (N_4918,In_1228,In_682);
and U4919 (N_4919,In_995,In_353);
nand U4920 (N_4920,In_218,In_1055);
or U4921 (N_4921,In_94,In_154);
nand U4922 (N_4922,In_1089,In_550);
and U4923 (N_4923,In_1041,In_1305);
nand U4924 (N_4924,In_1287,In_189);
or U4925 (N_4925,In_984,In_878);
nor U4926 (N_4926,In_1221,In_898);
nand U4927 (N_4927,In_902,In_1087);
xor U4928 (N_4928,In_155,In_1301);
nor U4929 (N_4929,In_1259,In_1028);
nand U4930 (N_4930,In_435,In_1080);
nand U4931 (N_4931,In_1008,In_1233);
or U4932 (N_4932,In_1350,In_1274);
and U4933 (N_4933,In_242,In_73);
and U4934 (N_4934,In_1342,In_795);
and U4935 (N_4935,In_1462,In_51);
or U4936 (N_4936,In_1451,In_44);
and U4937 (N_4937,In_1057,In_581);
nor U4938 (N_4938,In_1439,In_1255);
nor U4939 (N_4939,In_1128,In_2);
nand U4940 (N_4940,In_1306,In_1337);
nand U4941 (N_4941,In_1440,In_438);
or U4942 (N_4942,In_321,In_995);
nand U4943 (N_4943,In_212,In_489);
nand U4944 (N_4944,In_616,In_899);
nor U4945 (N_4945,In_129,In_563);
and U4946 (N_4946,In_654,In_357);
nor U4947 (N_4947,In_421,In_286);
nand U4948 (N_4948,In_29,In_1308);
nor U4949 (N_4949,In_1472,In_1116);
nand U4950 (N_4950,In_365,In_541);
xnor U4951 (N_4951,In_945,In_651);
or U4952 (N_4952,In_1086,In_1185);
xor U4953 (N_4953,In_152,In_1415);
and U4954 (N_4954,In_1216,In_936);
nor U4955 (N_4955,In_956,In_864);
xor U4956 (N_4956,In_1247,In_378);
nand U4957 (N_4957,In_545,In_1063);
or U4958 (N_4958,In_605,In_198);
xor U4959 (N_4959,In_735,In_191);
or U4960 (N_4960,In_1430,In_643);
nor U4961 (N_4961,In_1154,In_304);
and U4962 (N_4962,In_717,In_782);
nor U4963 (N_4963,In_1072,In_1266);
nand U4964 (N_4964,In_1035,In_1385);
nand U4965 (N_4965,In_942,In_240);
nor U4966 (N_4966,In_771,In_63);
nor U4967 (N_4967,In_99,In_1071);
nor U4968 (N_4968,In_396,In_253);
nand U4969 (N_4969,In_630,In_260);
and U4970 (N_4970,In_286,In_342);
and U4971 (N_4971,In_261,In_581);
xnor U4972 (N_4972,In_521,In_1328);
xor U4973 (N_4973,In_214,In_957);
nand U4974 (N_4974,In_495,In_949);
nor U4975 (N_4975,In_1274,In_211);
xnor U4976 (N_4976,In_67,In_1213);
xor U4977 (N_4977,In_691,In_71);
and U4978 (N_4978,In_1392,In_1042);
xor U4979 (N_4979,In_595,In_201);
xnor U4980 (N_4980,In_91,In_168);
nor U4981 (N_4981,In_1308,In_58);
and U4982 (N_4982,In_1144,In_618);
and U4983 (N_4983,In_678,In_46);
nand U4984 (N_4984,In_256,In_436);
or U4985 (N_4985,In_985,In_416);
and U4986 (N_4986,In_1179,In_1047);
or U4987 (N_4987,In_1031,In_480);
nor U4988 (N_4988,In_942,In_139);
xor U4989 (N_4989,In_139,In_446);
and U4990 (N_4990,In_371,In_919);
and U4991 (N_4991,In_23,In_1316);
and U4992 (N_4992,In_851,In_1436);
xor U4993 (N_4993,In_1012,In_854);
nand U4994 (N_4994,In_828,In_1328);
xnor U4995 (N_4995,In_77,In_565);
or U4996 (N_4996,In_125,In_627);
nor U4997 (N_4997,In_188,In_1259);
nand U4998 (N_4998,In_1243,In_1153);
or U4999 (N_4999,In_76,In_1227);
or U5000 (N_5000,N_3710,N_1123);
nor U5001 (N_5001,N_4450,N_1633);
xor U5002 (N_5002,N_3952,N_1189);
or U5003 (N_5003,N_4971,N_3503);
nand U5004 (N_5004,N_1545,N_4186);
nand U5005 (N_5005,N_417,N_4061);
nor U5006 (N_5006,N_3273,N_376);
nand U5007 (N_5007,N_4734,N_1745);
and U5008 (N_5008,N_4042,N_4726);
nor U5009 (N_5009,N_2172,N_3468);
or U5010 (N_5010,N_2995,N_3287);
nand U5011 (N_5011,N_3105,N_3762);
nand U5012 (N_5012,N_4083,N_1072);
nor U5013 (N_5013,N_2876,N_4232);
or U5014 (N_5014,N_1630,N_3110);
nor U5015 (N_5015,N_2889,N_3256);
nor U5016 (N_5016,N_4085,N_1378);
nor U5017 (N_5017,N_2549,N_208);
nand U5018 (N_5018,N_3043,N_1910);
xor U5019 (N_5019,N_1644,N_781);
or U5020 (N_5020,N_3310,N_1220);
nand U5021 (N_5021,N_2632,N_3158);
and U5022 (N_5022,N_4228,N_4922);
nand U5023 (N_5023,N_76,N_4419);
nand U5024 (N_5024,N_4503,N_485);
xnor U5025 (N_5025,N_3062,N_2798);
nand U5026 (N_5026,N_4849,N_1201);
nor U5027 (N_5027,N_4076,N_32);
and U5028 (N_5028,N_4770,N_2036);
or U5029 (N_5029,N_1578,N_2212);
nor U5030 (N_5030,N_3545,N_514);
nand U5031 (N_5031,N_2825,N_799);
xnor U5032 (N_5032,N_1754,N_487);
and U5033 (N_5033,N_3897,N_3599);
nor U5034 (N_5034,N_381,N_4828);
xnor U5035 (N_5035,N_1396,N_4156);
nand U5036 (N_5036,N_1140,N_1520);
or U5037 (N_5037,N_3367,N_232);
xor U5038 (N_5038,N_1181,N_2411);
or U5039 (N_5039,N_3865,N_103);
nand U5040 (N_5040,N_2158,N_111);
nor U5041 (N_5041,N_861,N_2298);
nand U5042 (N_5042,N_3773,N_3239);
and U5043 (N_5043,N_1266,N_2551);
and U5044 (N_5044,N_697,N_3212);
xor U5045 (N_5045,N_4929,N_4401);
and U5046 (N_5046,N_1058,N_2908);
nand U5047 (N_5047,N_4759,N_2260);
nand U5048 (N_5048,N_1525,N_390);
nor U5049 (N_5049,N_808,N_435);
nor U5050 (N_5050,N_1638,N_206);
nor U5051 (N_5051,N_4250,N_4729);
and U5052 (N_5052,N_167,N_4140);
or U5053 (N_5053,N_1255,N_35);
or U5054 (N_5054,N_481,N_2533);
or U5055 (N_5055,N_4622,N_4062);
xor U5056 (N_5056,N_267,N_682);
nand U5057 (N_5057,N_3648,N_4511);
and U5058 (N_5058,N_2858,N_408);
xnor U5059 (N_5059,N_4843,N_1900);
nand U5060 (N_5060,N_3617,N_601);
nor U5061 (N_5061,N_4275,N_681);
xnor U5062 (N_5062,N_934,N_4593);
or U5063 (N_5063,N_1671,N_983);
nor U5064 (N_5064,N_2885,N_794);
nor U5065 (N_5065,N_3511,N_732);
and U5066 (N_5066,N_512,N_3391);
xor U5067 (N_5067,N_4309,N_2199);
xor U5068 (N_5068,N_280,N_3676);
xor U5069 (N_5069,N_4386,N_2396);
or U5070 (N_5070,N_1766,N_4028);
or U5071 (N_5071,N_652,N_4857);
xor U5072 (N_5072,N_3417,N_4404);
xnor U5073 (N_5073,N_1905,N_2224);
nand U5074 (N_5074,N_870,N_4817);
and U5075 (N_5075,N_1293,N_622);
or U5076 (N_5076,N_3284,N_607);
xnor U5077 (N_5077,N_1041,N_2903);
and U5078 (N_5078,N_1818,N_2347);
nor U5079 (N_5079,N_2477,N_827);
or U5080 (N_5080,N_2911,N_4153);
nand U5081 (N_5081,N_3778,N_4168);
nand U5082 (N_5082,N_3642,N_1546);
nand U5083 (N_5083,N_595,N_386);
nor U5084 (N_5084,N_1888,N_142);
or U5085 (N_5085,N_2735,N_3592);
xor U5086 (N_5086,N_1105,N_1261);
nor U5087 (N_5087,N_1403,N_70);
xor U5088 (N_5088,N_3161,N_2796);
nand U5089 (N_5089,N_2540,N_3266);
nor U5090 (N_5090,N_3661,N_4582);
nor U5091 (N_5091,N_177,N_1436);
or U5092 (N_5092,N_3340,N_3974);
and U5093 (N_5093,N_3060,N_3735);
or U5094 (N_5094,N_4072,N_4449);
nor U5095 (N_5095,N_1681,N_3825);
xnor U5096 (N_5096,N_4241,N_2446);
nor U5097 (N_5097,N_4302,N_4767);
xor U5098 (N_5098,N_2425,N_122);
and U5099 (N_5099,N_2469,N_1907);
or U5100 (N_5100,N_698,N_571);
or U5101 (N_5101,N_2936,N_4304);
and U5102 (N_5102,N_4732,N_775);
nor U5103 (N_5103,N_226,N_1314);
xor U5104 (N_5104,N_3615,N_1849);
nand U5105 (N_5105,N_4056,N_4485);
or U5106 (N_5106,N_3264,N_3831);
nor U5107 (N_5107,N_4771,N_3032);
nor U5108 (N_5108,N_847,N_4384);
xor U5109 (N_5109,N_1399,N_4754);
nor U5110 (N_5110,N_1194,N_4390);
and U5111 (N_5111,N_1010,N_258);
nand U5112 (N_5112,N_815,N_3942);
or U5113 (N_5113,N_1457,N_4262);
nor U5114 (N_5114,N_262,N_169);
and U5115 (N_5115,N_1282,N_1137);
or U5116 (N_5116,N_2807,N_3382);
nor U5117 (N_5117,N_686,N_4783);
nand U5118 (N_5118,N_1296,N_1601);
or U5119 (N_5119,N_2358,N_3484);
nor U5120 (N_5120,N_2294,N_3221);
nor U5121 (N_5121,N_1388,N_4336);
nor U5122 (N_5122,N_1066,N_4878);
and U5123 (N_5123,N_3659,N_449);
and U5124 (N_5124,N_53,N_416);
or U5125 (N_5125,N_3554,N_4442);
nor U5126 (N_5126,N_3780,N_4159);
nand U5127 (N_5127,N_138,N_1191);
xnor U5128 (N_5128,N_4043,N_4893);
nor U5129 (N_5129,N_3163,N_4287);
xnor U5130 (N_5130,N_821,N_3818);
nand U5131 (N_5131,N_729,N_39);
or U5132 (N_5132,N_286,N_1004);
or U5133 (N_5133,N_3725,N_3137);
xnor U5134 (N_5134,N_2699,N_26);
or U5135 (N_5135,N_3028,N_303);
xnor U5136 (N_5136,N_3720,N_1940);
nand U5137 (N_5137,N_2081,N_2553);
nand U5138 (N_5138,N_1460,N_1412);
nand U5139 (N_5139,N_4761,N_909);
and U5140 (N_5140,N_3774,N_4632);
nor U5141 (N_5141,N_2314,N_269);
xnor U5142 (N_5142,N_2772,N_920);
nand U5143 (N_5143,N_896,N_3680);
and U5144 (N_5144,N_2990,N_300);
nor U5145 (N_5145,N_4804,N_4999);
xnor U5146 (N_5146,N_4266,N_2855);
and U5147 (N_5147,N_945,N_3875);
xnor U5148 (N_5148,N_971,N_2616);
xor U5149 (N_5149,N_1362,N_4865);
nor U5150 (N_5150,N_3996,N_1980);
nand U5151 (N_5151,N_3874,N_2615);
nor U5152 (N_5152,N_3112,N_3707);
and U5153 (N_5153,N_2386,N_4669);
nand U5154 (N_5154,N_2783,N_1823);
and U5155 (N_5155,N_1283,N_2763);
or U5156 (N_5156,N_4847,N_4306);
nand U5157 (N_5157,N_1530,N_3535);
nand U5158 (N_5158,N_2609,N_766);
nand U5159 (N_5159,N_2297,N_670);
and U5160 (N_5160,N_1312,N_1876);
xnor U5161 (N_5161,N_4092,N_1405);
nor U5162 (N_5162,N_4698,N_4481);
or U5163 (N_5163,N_579,N_2221);
or U5164 (N_5164,N_289,N_1742);
and U5165 (N_5165,N_546,N_2291);
or U5166 (N_5166,N_4594,N_1989);
or U5167 (N_5167,N_1901,N_201);
nand U5168 (N_5168,N_4510,N_3842);
or U5169 (N_5169,N_944,N_2215);
nand U5170 (N_5170,N_4801,N_760);
or U5171 (N_5171,N_2253,N_918);
or U5172 (N_5172,N_4052,N_4677);
nor U5173 (N_5173,N_2710,N_4851);
nor U5174 (N_5174,N_987,N_1169);
nand U5175 (N_5175,N_474,N_2045);
nor U5176 (N_5176,N_4626,N_2142);
nand U5177 (N_5177,N_4272,N_3835);
nand U5178 (N_5178,N_4860,N_438);
or U5179 (N_5179,N_1929,N_2661);
and U5180 (N_5180,N_3167,N_3757);
nor U5181 (N_5181,N_733,N_185);
nand U5182 (N_5182,N_3560,N_4123);
nand U5183 (N_5183,N_4996,N_4727);
nand U5184 (N_5184,N_2547,N_3418);
or U5185 (N_5185,N_3957,N_2875);
nand U5186 (N_5186,N_4926,N_1439);
and U5187 (N_5187,N_2865,N_3422);
or U5188 (N_5188,N_707,N_4741);
xor U5189 (N_5189,N_2157,N_887);
or U5190 (N_5190,N_1802,N_2671);
nand U5191 (N_5191,N_4894,N_3206);
and U5192 (N_5192,N_2502,N_4311);
or U5193 (N_5193,N_1591,N_1418);
nor U5194 (N_5194,N_3144,N_305);
nor U5195 (N_5195,N_2792,N_1159);
xor U5196 (N_5196,N_3797,N_2519);
and U5197 (N_5197,N_1752,N_1974);
and U5198 (N_5198,N_3460,N_109);
nor U5199 (N_5199,N_4395,N_2352);
nand U5200 (N_5200,N_139,N_1338);
nand U5201 (N_5201,N_1598,N_4943);
nor U5202 (N_5202,N_2244,N_3139);
xnor U5203 (N_5203,N_3867,N_4839);
nor U5204 (N_5204,N_496,N_2459);
xnor U5205 (N_5205,N_3671,N_4057);
or U5206 (N_5206,N_1052,N_4636);
xor U5207 (N_5207,N_3941,N_2739);
nor U5208 (N_5208,N_1521,N_3748);
nand U5209 (N_5209,N_699,N_3069);
and U5210 (N_5210,N_3922,N_3537);
xnor U5211 (N_5211,N_245,N_389);
nor U5212 (N_5212,N_4522,N_2342);
nand U5213 (N_5213,N_3356,N_1334);
xnor U5214 (N_5214,N_4631,N_1713);
nor U5215 (N_5215,N_9,N_4885);
xnor U5216 (N_5216,N_1002,N_4921);
or U5217 (N_5217,N_1760,N_4138);
and U5218 (N_5218,N_1080,N_3644);
and U5219 (N_5219,N_4564,N_1902);
xor U5220 (N_5220,N_3132,N_1839);
nor U5221 (N_5221,N_1544,N_54);
nor U5222 (N_5222,N_3734,N_1554);
and U5223 (N_5223,N_3873,N_1136);
nand U5224 (N_5224,N_23,N_2578);
nor U5225 (N_5225,N_3699,N_3243);
and U5226 (N_5226,N_2110,N_217);
and U5227 (N_5227,N_771,N_3740);
nand U5228 (N_5228,N_4339,N_1877);
or U5229 (N_5229,N_4534,N_2429);
or U5230 (N_5230,N_2543,N_691);
nor U5231 (N_5231,N_1350,N_270);
and U5232 (N_5232,N_3806,N_4952);
nand U5233 (N_5233,N_2176,N_3597);
nor U5234 (N_5234,N_2466,N_4116);
nand U5235 (N_5235,N_715,N_4523);
and U5236 (N_5236,N_4528,N_4914);
xnor U5237 (N_5237,N_4239,N_3236);
nand U5238 (N_5238,N_3811,N_2503);
nand U5239 (N_5239,N_2276,N_30);
nand U5240 (N_5240,N_898,N_4301);
and U5241 (N_5241,N_1318,N_4343);
xnor U5242 (N_5242,N_3898,N_3883);
nand U5243 (N_5243,N_3343,N_1112);
nand U5244 (N_5244,N_3843,N_4723);
nor U5245 (N_5245,N_3324,N_6);
nand U5246 (N_5246,N_4044,N_2899);
and U5247 (N_5247,N_4491,N_4928);
and U5248 (N_5248,N_1321,N_3716);
nor U5249 (N_5249,N_2070,N_3001);
and U5250 (N_5250,N_2130,N_4992);
nand U5251 (N_5251,N_2846,N_3697);
xor U5252 (N_5252,N_4171,N_1245);
xor U5253 (N_5253,N_4901,N_3765);
or U5254 (N_5254,N_1696,N_3135);
nand U5255 (N_5255,N_4008,N_1658);
nor U5256 (N_5256,N_410,N_935);
nand U5257 (N_5257,N_3044,N_1934);
or U5258 (N_5258,N_3189,N_450);
nand U5259 (N_5259,N_2853,N_211);
nor U5260 (N_5260,N_1685,N_3403);
nor U5261 (N_5261,N_3142,N_2083);
and U5262 (N_5262,N_1485,N_4397);
and U5263 (N_5263,N_608,N_3904);
and U5264 (N_5264,N_3398,N_3892);
or U5265 (N_5265,N_841,N_3116);
nor U5266 (N_5266,N_4988,N_3050);
nand U5267 (N_5267,N_665,N_3285);
nor U5268 (N_5268,N_3949,N_2815);
xnor U5269 (N_5269,N_4000,N_1132);
or U5270 (N_5270,N_4875,N_403);
xnor U5271 (N_5271,N_2684,N_3448);
and U5272 (N_5272,N_4420,N_4342);
and U5273 (N_5273,N_112,N_930);
nand U5274 (N_5274,N_3886,N_4643);
xnor U5275 (N_5275,N_437,N_4144);
nand U5276 (N_5276,N_1087,N_1593);
or U5277 (N_5277,N_3241,N_4586);
xor U5278 (N_5278,N_3688,N_928);
xnor U5279 (N_5279,N_4270,N_4696);
nor U5280 (N_5280,N_1855,N_4640);
xnor U5281 (N_5281,N_1796,N_4392);
and U5282 (N_5282,N_1674,N_4652);
and U5283 (N_5283,N_295,N_3862);
nor U5284 (N_5284,N_1364,N_516);
and U5285 (N_5285,N_2436,N_876);
xnor U5286 (N_5286,N_2030,N_4105);
nand U5287 (N_5287,N_1107,N_1597);
or U5288 (N_5288,N_1264,N_1677);
or U5289 (N_5289,N_64,N_2056);
xnor U5290 (N_5290,N_2842,N_4149);
and U5291 (N_5291,N_3976,N_1097);
or U5292 (N_5292,N_3690,N_3746);
xnor U5293 (N_5293,N_1056,N_3406);
or U5294 (N_5294,N_3960,N_1883);
nand U5295 (N_5295,N_832,N_2760);
xnor U5296 (N_5296,N_593,N_3254);
nor U5297 (N_5297,N_1919,N_395);
and U5298 (N_5298,N_3294,N_2333);
nor U5299 (N_5299,N_4040,N_311);
nand U5300 (N_5300,N_2415,N_513);
or U5301 (N_5301,N_4748,N_4666);
nand U5302 (N_5302,N_1351,N_2651);
xor U5303 (N_5303,N_2731,N_4280);
and U5304 (N_5304,N_4082,N_4612);
xnor U5305 (N_5305,N_2323,N_308);
xnor U5306 (N_5306,N_1178,N_2574);
nor U5307 (N_5307,N_3117,N_3558);
nand U5308 (N_5308,N_2816,N_3731);
xnor U5309 (N_5309,N_2357,N_0);
and U5310 (N_5310,N_3194,N_2879);
or U5311 (N_5311,N_2658,N_2389);
or U5312 (N_5312,N_3581,N_3758);
or U5313 (N_5313,N_4627,N_1503);
nor U5314 (N_5314,N_2258,N_3430);
and U5315 (N_5315,N_1400,N_241);
and U5316 (N_5316,N_3742,N_1821);
xnor U5317 (N_5317,N_3571,N_4704);
xor U5318 (N_5318,N_421,N_4346);
xnor U5319 (N_5319,N_4601,N_1816);
nand U5320 (N_5320,N_57,N_3967);
and U5321 (N_5321,N_4494,N_2591);
and U5322 (N_5322,N_798,N_3882);
nand U5323 (N_5323,N_2229,N_1853);
xnor U5324 (N_5324,N_2420,N_1489);
nand U5325 (N_5325,N_276,N_4654);
or U5326 (N_5326,N_3351,N_1117);
nand U5327 (N_5327,N_1285,N_3667);
xor U5328 (N_5328,N_3946,N_83);
and U5329 (N_5329,N_2049,N_2385);
nor U5330 (N_5330,N_2487,N_2458);
and U5331 (N_5331,N_1535,N_3990);
nor U5332 (N_5332,N_3788,N_4247);
nor U5333 (N_5333,N_4963,N_4258);
xnor U5334 (N_5334,N_746,N_1561);
xnor U5335 (N_5335,N_116,N_2934);
or U5336 (N_5336,N_1799,N_81);
or U5337 (N_5337,N_3663,N_4620);
or U5338 (N_5338,N_825,N_879);
nand U5339 (N_5339,N_1146,N_647);
xnor U5340 (N_5340,N_230,N_2968);
or U5341 (N_5341,N_1978,N_4284);
nand U5342 (N_5342,N_3864,N_4633);
xnor U5343 (N_5343,N_4530,N_3939);
and U5344 (N_5344,N_4069,N_1676);
nand U5345 (N_5345,N_446,N_183);
or U5346 (N_5346,N_4222,N_1272);
or U5347 (N_5347,N_1789,N_4777);
nor U5348 (N_5348,N_3291,N_3507);
nor U5349 (N_5349,N_1361,N_2098);
xnor U5350 (N_5350,N_1342,N_4840);
xnor U5351 (N_5351,N_924,N_2530);
nand U5352 (N_5352,N_2999,N_176);
and U5353 (N_5353,N_4736,N_3772);
nand U5354 (N_5354,N_1076,N_3975);
nor U5355 (N_5355,N_3523,N_1346);
xnor U5356 (N_5356,N_73,N_4716);
xor U5357 (N_5357,N_368,N_1409);
nand U5358 (N_5358,N_4935,N_1019);
nor U5359 (N_5359,N_108,N_2412);
nor U5360 (N_5360,N_2442,N_2776);
nor U5361 (N_5361,N_846,N_3384);
xor U5362 (N_5362,N_4755,N_3621);
nor U5363 (N_5363,N_3590,N_826);
and U5364 (N_5364,N_4907,N_2734);
nor U5365 (N_5365,N_4165,N_3923);
and U5366 (N_5366,N_980,N_2047);
xor U5367 (N_5367,N_2828,N_1568);
nor U5368 (N_5368,N_3718,N_3878);
and U5369 (N_5369,N_3755,N_4383);
or U5370 (N_5370,N_2507,N_4421);
nand U5371 (N_5371,N_3912,N_598);
or U5372 (N_5372,N_742,N_2374);
or U5373 (N_5373,N_3429,N_1253);
xor U5374 (N_5374,N_4703,N_4439);
xnor U5375 (N_5375,N_537,N_2444);
and U5376 (N_5376,N_3576,N_236);
nand U5377 (N_5377,N_3544,N_2612);
xor U5378 (N_5378,N_4291,N_1805);
and U5379 (N_5379,N_1592,N_2324);
nor U5380 (N_5380,N_2217,N_2062);
or U5381 (N_5381,N_2496,N_1718);
and U5382 (N_5382,N_631,N_1684);
nand U5383 (N_5383,N_4845,N_3346);
or U5384 (N_5384,N_3270,N_1490);
xor U5385 (N_5385,N_1007,N_3006);
or U5386 (N_5386,N_2006,N_3466);
xnor U5387 (N_5387,N_1281,N_2134);
nand U5388 (N_5388,N_2434,N_3414);
xnor U5389 (N_5389,N_1634,N_2315);
nand U5390 (N_5390,N_2698,N_3969);
nand U5391 (N_5391,N_2694,N_1714);
and U5392 (N_5392,N_4548,N_212);
or U5393 (N_5393,N_2541,N_2023);
xnor U5394 (N_5394,N_1099,N_1202);
or U5395 (N_5395,N_4607,N_2539);
nand U5396 (N_5396,N_4024,N_1960);
nand U5397 (N_5397,N_1493,N_520);
nor U5398 (N_5398,N_2219,N_3606);
nor U5399 (N_5399,N_2339,N_2648);
xor U5400 (N_5400,N_1125,N_982);
nor U5401 (N_5401,N_3173,N_1831);
or U5402 (N_5402,N_646,N_2151);
nor U5403 (N_5403,N_162,N_348);
and U5404 (N_5404,N_1455,N_1775);
or U5405 (N_5405,N_3015,N_113);
nand U5406 (N_5406,N_2011,N_1026);
or U5407 (N_5407,N_260,N_4221);
or U5408 (N_5408,N_4685,N_3760);
nand U5409 (N_5409,N_3627,N_2946);
or U5410 (N_5410,N_2237,N_301);
nor U5411 (N_5411,N_3753,N_1657);
or U5412 (N_5412,N_1724,N_3605);
and U5413 (N_5413,N_4424,N_4973);
and U5414 (N_5414,N_360,N_1769);
or U5415 (N_5415,N_1596,N_3980);
or U5416 (N_5416,N_1590,N_2768);
nand U5417 (N_5417,N_706,N_2447);
xnor U5418 (N_5418,N_2280,N_806);
and U5419 (N_5419,N_2129,N_3345);
and U5420 (N_5420,N_3987,N_2849);
or U5421 (N_5421,N_4599,N_3279);
nor U5422 (N_5422,N_779,N_4193);
nand U5423 (N_5423,N_690,N_673);
nor U5424 (N_5424,N_1707,N_2810);
xnor U5425 (N_5425,N_2992,N_602);
nand U5426 (N_5426,N_1499,N_4200);
or U5427 (N_5427,N_1540,N_4359);
and U5428 (N_5428,N_809,N_3233);
xnor U5429 (N_5429,N_3404,N_4223);
and U5430 (N_5430,N_718,N_1549);
or U5431 (N_5431,N_5,N_2190);
nand U5432 (N_5432,N_4163,N_3077);
or U5433 (N_5433,N_2003,N_4715);
nor U5434 (N_5434,N_2965,N_4531);
and U5435 (N_5435,N_3293,N_2432);
nand U5436 (N_5436,N_3223,N_2750);
xnor U5437 (N_5437,N_18,N_4235);
xor U5438 (N_5438,N_2265,N_235);
nand U5439 (N_5439,N_1459,N_638);
and U5440 (N_5440,N_2209,N_1917);
and U5441 (N_5441,N_2398,N_359);
nand U5442 (N_5442,N_2644,N_2405);
and U5443 (N_5443,N_2941,N_1992);
nor U5444 (N_5444,N_2499,N_288);
and U5445 (N_5445,N_3528,N_3073);
nor U5446 (N_5446,N_3107,N_3195);
and U5447 (N_5447,N_1642,N_1149);
and U5448 (N_5448,N_3424,N_2054);
nand U5449 (N_5449,N_4890,N_4217);
nand U5450 (N_5450,N_748,N_1241);
nand U5451 (N_5451,N_20,N_2243);
nand U5452 (N_5452,N_2910,N_1973);
or U5453 (N_5453,N_29,N_4078);
nor U5454 (N_5454,N_1395,N_282);
xor U5455 (N_5455,N_2200,N_4525);
nand U5456 (N_5456,N_318,N_1273);
nor U5457 (N_5457,N_3472,N_1652);
and U5458 (N_5458,N_3930,N_4323);
or U5459 (N_5459,N_1697,N_4189);
nand U5460 (N_5460,N_1310,N_1983);
nor U5461 (N_5461,N_2532,N_2840);
nor U5462 (N_5462,N_4154,N_4286);
nor U5463 (N_5463,N_2144,N_2878);
nor U5464 (N_5464,N_1110,N_3386);
nand U5465 (N_5465,N_3092,N_4130);
nor U5466 (N_5466,N_1476,N_3111);
nor U5467 (N_5467,N_1028,N_4581);
and U5468 (N_5468,N_3623,N_4859);
or U5469 (N_5469,N_40,N_755);
and U5470 (N_5470,N_3113,N_4689);
xor U5471 (N_5471,N_4898,N_2175);
nand U5472 (N_5472,N_999,N_3196);
or U5473 (N_5473,N_1344,N_3657);
nand U5474 (N_5474,N_548,N_4210);
xnor U5475 (N_5475,N_2079,N_3479);
or U5476 (N_5476,N_3958,N_2301);
nor U5477 (N_5477,N_12,N_3443);
xor U5478 (N_5478,N_1031,N_2994);
xor U5479 (N_5479,N_128,N_1967);
xor U5480 (N_5480,N_3869,N_319);
nor U5481 (N_5481,N_1694,N_2978);
or U5482 (N_5482,N_1108,N_358);
nand U5483 (N_5483,N_1847,N_3896);
or U5484 (N_5484,N_2309,N_4546);
or U5485 (N_5485,N_4001,N_4459);
nor U5486 (N_5486,N_1963,N_2950);
or U5487 (N_5487,N_3686,N_553);
nand U5488 (N_5488,N_199,N_44);
or U5489 (N_5489,N_4226,N_2663);
xor U5490 (N_5490,N_1605,N_4051);
and U5491 (N_5491,N_1764,N_1416);
nand U5492 (N_5492,N_4155,N_1508);
nand U5493 (N_5493,N_2617,N_816);
nand U5494 (N_5494,N_3518,N_489);
nor U5495 (N_5495,N_4989,N_3562);
nand U5496 (N_5496,N_3754,N_1180);
xor U5497 (N_5497,N_3464,N_3607);
nor U5498 (N_5498,N_1392,N_1176);
nor U5499 (N_5499,N_2743,N_2747);
and U5500 (N_5500,N_3849,N_2092);
nand U5501 (N_5501,N_317,N_259);
and U5502 (N_5502,N_323,N_1739);
nand U5503 (N_5503,N_3190,N_1472);
xnor U5504 (N_5504,N_1025,N_2489);
or U5505 (N_5505,N_16,N_4709);
or U5506 (N_5506,N_4606,N_4553);
and U5507 (N_5507,N_1687,N_265);
or U5508 (N_5508,N_662,N_4444);
xor U5509 (N_5509,N_885,N_285);
nand U5510 (N_5510,N_3009,N_4166);
nor U5511 (N_5511,N_1154,N_4536);
nand U5512 (N_5512,N_731,N_1570);
and U5513 (N_5513,N_4889,N_3988);
nor U5514 (N_5514,N_429,N_2974);
xor U5515 (N_5515,N_1085,N_4719);
nor U5516 (N_5516,N_1723,N_4431);
xnor U5517 (N_5517,N_1628,N_2657);
nand U5518 (N_5518,N_859,N_4947);
or U5519 (N_5519,N_4782,N_3826);
nor U5520 (N_5520,N_669,N_4969);
or U5521 (N_5521,N_2014,N_3300);
and U5522 (N_5522,N_2834,N_1168);
or U5523 (N_5523,N_1486,N_3297);
nand U5524 (N_5524,N_1864,N_3329);
and U5525 (N_5525,N_3039,N_627);
nor U5526 (N_5526,N_3836,N_574);
nand U5527 (N_5527,N_1933,N_3249);
xnor U5528 (N_5528,N_3079,N_4268);
nand U5529 (N_5529,N_2573,N_36);
nand U5530 (N_5530,N_693,N_2987);
nor U5531 (N_5531,N_1854,N_4816);
or U5532 (N_5532,N_363,N_3594);
or U5533 (N_5533,N_2327,N_1518);
and U5534 (N_5534,N_963,N_28);
nand U5535 (N_5535,N_3660,N_4509);
xor U5536 (N_5536,N_1401,N_554);
xnor U5537 (N_5537,N_1809,N_3280);
xor U5538 (N_5538,N_901,N_2607);
nand U5539 (N_5539,N_1324,N_2559);
and U5540 (N_5540,N_91,N_2234);
nand U5541 (N_5541,N_224,N_2468);
or U5542 (N_5542,N_375,N_1969);
and U5543 (N_5543,N_4364,N_4744);
nand U5544 (N_5544,N_3807,N_2915);
xnor U5545 (N_5545,N_469,N_2206);
or U5546 (N_5546,N_2355,N_1157);
and U5547 (N_5547,N_2714,N_290);
and U5548 (N_5548,N_3210,N_157);
nor U5549 (N_5549,N_2226,N_4029);
and U5550 (N_5550,N_1160,N_3467);
and U5551 (N_5551,N_1613,N_379);
and U5552 (N_5552,N_3260,N_1706);
or U5553 (N_5553,N_564,N_306);
and U5554 (N_5554,N_2645,N_2631);
nor U5555 (N_5555,N_908,N_2299);
nor U5556 (N_5556,N_1461,N_2096);
xnor U5557 (N_5557,N_1984,N_4418);
nor U5558 (N_5558,N_2101,N_4483);
nand U5559 (N_5559,N_4143,N_3940);
or U5560 (N_5560,N_2373,N_154);
nor U5561 (N_5561,N_1820,N_1639);
and U5562 (N_5562,N_2594,N_626);
xnor U5563 (N_5563,N_3870,N_2722);
xor U5564 (N_5564,N_1012,N_4435);
nand U5565 (N_5565,N_1481,N_4285);
xor U5566 (N_5566,N_4470,N_2282);
nand U5567 (N_5567,N_3695,N_4313);
and U5568 (N_5568,N_65,N_321);
xnor U5569 (N_5569,N_1111,N_831);
xnor U5570 (N_5570,N_3454,N_2316);
nor U5571 (N_5571,N_2392,N_52);
xnor U5572 (N_5572,N_3432,N_984);
xor U5573 (N_5573,N_3213,N_2614);
xnor U5574 (N_5574,N_3611,N_182);
xnor U5575 (N_5575,N_4998,N_3548);
and U5576 (N_5576,N_274,N_3595);
and U5577 (N_5577,N_4271,N_4463);
nor U5578 (N_5578,N_2996,N_1061);
and U5579 (N_5579,N_3025,N_1991);
or U5580 (N_5580,N_4399,N_2705);
xor U5581 (N_5581,N_1196,N_1976);
or U5582 (N_5582,N_2837,N_1552);
or U5583 (N_5583,N_674,N_3812);
xor U5584 (N_5584,N_1911,N_1621);
and U5585 (N_5585,N_2225,N_700);
xor U5586 (N_5586,N_790,N_2077);
and U5587 (N_5587,N_3172,N_1523);
nand U5588 (N_5588,N_2848,N_1887);
and U5589 (N_5589,N_2400,N_4263);
nand U5590 (N_5590,N_1243,N_1016);
xnor U5591 (N_5591,N_1550,N_2476);
and U5592 (N_5592,N_4229,N_4571);
and U5593 (N_5593,N_331,N_803);
nor U5594 (N_5594,N_4423,N_2164);
nand U5595 (N_5595,N_4550,N_4682);
nor U5596 (N_5596,N_1637,N_255);
nor U5597 (N_5597,N_3552,N_3331);
or U5598 (N_5598,N_1131,N_4403);
nand U5599 (N_5599,N_1226,N_1040);
nand U5600 (N_5600,N_149,N_2336);
and U5601 (N_5601,N_156,N_467);
and U5602 (N_5602,N_3935,N_38);
or U5603 (N_5603,N_3624,N_1480);
xnor U5604 (N_5604,N_2065,N_1124);
and U5605 (N_5605,N_959,N_4577);
xnor U5606 (N_5606,N_575,N_427);
or U5607 (N_5607,N_4948,N_1914);
xor U5608 (N_5608,N_2369,N_3901);
nand U5609 (N_5609,N_2277,N_3508);
or U5610 (N_5610,N_1725,N_4802);
nor U5611 (N_5611,N_3641,N_68);
nor U5612 (N_5612,N_3540,N_1434);
or U5613 (N_5613,N_1433,N_4412);
nand U5614 (N_5614,N_1083,N_1957);
xor U5615 (N_5615,N_3497,N_371);
and U5616 (N_5616,N_1335,N_2259);
xor U5617 (N_5617,N_4278,N_4327);
and U5618 (N_5618,N_2311,N_2867);
nand U5619 (N_5619,N_293,N_764);
xnor U5620 (N_5620,N_3244,N_937);
nand U5621 (N_5621,N_82,N_2115);
nor U5622 (N_5622,N_3409,N_4913);
or U5623 (N_5623,N_888,N_2544);
xor U5624 (N_5624,N_3240,N_10);
or U5625 (N_5625,N_2111,N_811);
xnor U5626 (N_5626,N_490,N_4101);
nand U5627 (N_5627,N_4429,N_1997);
or U5628 (N_5628,N_3970,N_2882);
and U5629 (N_5629,N_2809,N_3833);
xnor U5630 (N_5630,N_462,N_1257);
xnor U5631 (N_5631,N_3353,N_2080);
nand U5632 (N_5632,N_1404,N_1532);
xnor U5633 (N_5633,N_1701,N_2139);
nor U5634 (N_5634,N_4,N_4780);
and U5635 (N_5635,N_740,N_2856);
and U5636 (N_5636,N_4097,N_1599);
or U5637 (N_5637,N_966,N_1470);
or U5638 (N_5638,N_1408,N_994);
and U5639 (N_5639,N_1954,N_2270);
nor U5640 (N_5640,N_4468,N_2494);
or U5641 (N_5641,N_1574,N_314);
nand U5642 (N_5642,N_3857,N_4858);
or U5643 (N_5643,N_2240,N_502);
nor U5644 (N_5644,N_4374,N_4679);
or U5645 (N_5645,N_71,N_4484);
or U5646 (N_5646,N_1479,N_3415);
xnor U5647 (N_5647,N_525,N_4045);
xnor U5648 (N_5648,N_346,N_2287);
nor U5649 (N_5649,N_4388,N_985);
nand U5650 (N_5650,N_50,N_1235);
and U5651 (N_5651,N_2582,N_4113);
nor U5652 (N_5652,N_3251,N_1013);
and U5653 (N_5653,N_1289,N_3854);
or U5654 (N_5654,N_1187,N_4670);
xor U5655 (N_5655,N_2264,N_974);
nor U5656 (N_5656,N_1719,N_4946);
xnor U5657 (N_5657,N_1130,N_1673);
xor U5658 (N_5658,N_4133,N_858);
nand U5659 (N_5659,N_451,N_2976);
and U5660 (N_5660,N_2500,N_589);
xnor U5661 (N_5661,N_87,N_3764);
xor U5662 (N_5662,N_1729,N_2133);
xor U5663 (N_5663,N_3168,N_342);
nand U5664 (N_5664,N_2531,N_843);
or U5665 (N_5665,N_4888,N_2089);
or U5666 (N_5666,N_4356,N_412);
and U5667 (N_5667,N_4150,N_3492);
nor U5668 (N_5668,N_3822,N_3181);
and U5669 (N_5669,N_4864,N_1541);
xor U5670 (N_5670,N_1495,N_2956);
xor U5671 (N_5671,N_3645,N_3086);
nand U5672 (N_5672,N_1082,N_2896);
nor U5673 (N_5673,N_2775,N_4345);
and U5674 (N_5674,N_3066,N_3792);
and U5675 (N_5675,N_4430,N_3171);
xor U5676 (N_5676,N_3433,N_4778);
xor U5677 (N_5677,N_248,N_98);
nor U5678 (N_5678,N_4683,N_422);
xor U5679 (N_5679,N_2780,N_1075);
nor U5680 (N_5680,N_3379,N_3821);
nor U5681 (N_5681,N_4347,N_3387);
nand U5682 (N_5682,N_1845,N_1113);
and U5683 (N_5683,N_3123,N_2471);
and U5684 (N_5684,N_2185,N_3038);
nor U5685 (N_5685,N_3485,N_2318);
nand U5686 (N_5686,N_1429,N_2831);
nor U5687 (N_5687,N_651,N_2939);
and U5688 (N_5688,N_2569,N_3924);
xor U5689 (N_5689,N_4486,N_4411);
and U5690 (N_5690,N_3744,N_4702);
or U5691 (N_5691,N_1659,N_1055);
and U5692 (N_5692,N_4445,N_906);
or U5693 (N_5693,N_1305,N_249);
and U5694 (N_5694,N_882,N_335);
nand U5695 (N_5695,N_1393,N_2071);
nand U5696 (N_5696,N_3296,N_1144);
and U5697 (N_5697,N_4259,N_1008);
and U5698 (N_5698,N_227,N_805);
nand U5699 (N_5699,N_1450,N_1916);
or U5700 (N_5700,N_1415,N_2382);
xor U5701 (N_5701,N_1512,N_3463);
and U5702 (N_5702,N_2127,N_1100);
nand U5703 (N_5703,N_4371,N_3012);
xnor U5704 (N_5704,N_829,N_1874);
xnor U5705 (N_5705,N_3944,N_777);
and U5706 (N_5706,N_2486,N_4005);
xnor U5707 (N_5707,N_1150,N_414);
xnor U5708 (N_5708,N_3017,N_3231);
or U5709 (N_5709,N_148,N_2247);
nand U5710 (N_5710,N_179,N_1250);
or U5711 (N_5711,N_3736,N_4688);
xnor U5712 (N_5712,N_441,N_2754);
xor U5713 (N_5713,N_4659,N_2504);
xor U5714 (N_5714,N_4274,N_1619);
nor U5715 (N_5715,N_221,N_120);
or U5716 (N_5716,N_3521,N_3119);
nor U5717 (N_5717,N_3947,N_329);
and U5718 (N_5718,N_3400,N_2072);
nor U5719 (N_5719,N_2957,N_1079);
nand U5720 (N_5720,N_3931,N_2482);
and U5721 (N_5721,N_973,N_517);
and U5722 (N_5722,N_948,N_3180);
nand U5723 (N_5723,N_3320,N_763);
nor U5724 (N_5724,N_713,N_1203);
xnor U5725 (N_5725,N_2317,N_1522);
and U5726 (N_5726,N_2975,N_1966);
nor U5727 (N_5727,N_2193,N_3669);
xor U5728 (N_5728,N_4294,N_263);
nor U5729 (N_5729,N_623,N_4282);
nor U5730 (N_5730,N_504,N_711);
or U5731 (N_5731,N_2652,N_445);
and U5732 (N_5732,N_1923,N_4638);
and U5733 (N_5733,N_2741,N_4256);
and U5734 (N_5734,N_3118,N_4657);
nor U5735 (N_5735,N_1941,N_696);
nor U5736 (N_5736,N_3441,N_4330);
and U5737 (N_5737,N_147,N_3965);
and U5738 (N_5738,N_1819,N_1560);
and U5739 (N_5739,N_1580,N_4648);
nand U5740 (N_5740,N_3475,N_1835);
or U5741 (N_5741,N_3968,N_3222);
and U5742 (N_5742,N_630,N_1276);
or U5743 (N_5743,N_605,N_2550);
and U5744 (N_5744,N_4151,N_4198);
or U5745 (N_5745,N_3786,N_3705);
nand U5746 (N_5746,N_256,N_135);
nand U5747 (N_5747,N_577,N_4578);
and U5748 (N_5748,N_3410,N_84);
nand U5749 (N_5749,N_3654,N_3253);
nand U5750 (N_5750,N_765,N_1841);
and U5751 (N_5751,N_3307,N_1611);
nor U5752 (N_5752,N_4554,N_2778);
nor U5753 (N_5753,N_2638,N_4498);
and U5754 (N_5754,N_500,N_557);
nand U5755 (N_5755,N_3525,N_4753);
or U5756 (N_5756,N_4264,N_3911);
or U5757 (N_5757,N_3737,N_524);
nand U5758 (N_5758,N_4324,N_992);
nand U5759 (N_5759,N_1501,N_3261);
nor U5760 (N_5760,N_4749,N_1889);
nand U5761 (N_5761,N_257,N_566);
and U5762 (N_5762,N_2086,N_3616);
and U5763 (N_5763,N_4357,N_3312);
nand U5764 (N_5764,N_4796,N_3588);
nor U5765 (N_5765,N_4714,N_1365);
nand U5766 (N_5766,N_2984,N_2675);
xor U5767 (N_5767,N_2951,N_1224);
or U5768 (N_5768,N_3815,N_845);
or U5769 (N_5769,N_477,N_972);
nand U5770 (N_5770,N_2610,N_3677);
nor U5771 (N_5771,N_2556,N_62);
nor U5772 (N_5772,N_4559,N_978);
or U5773 (N_5773,N_2762,N_1465);
nor U5774 (N_5774,N_4739,N_3613);
nand U5775 (N_5775,N_404,N_3771);
nor U5776 (N_5776,N_2918,N_1937);
nand U5777 (N_5777,N_4708,N_4896);
xnor U5778 (N_5778,N_1035,N_701);
and U5779 (N_5779,N_2337,N_1767);
and U5780 (N_5780,N_1994,N_3421);
xor U5781 (N_5781,N_4184,N_4966);
and U5782 (N_5782,N_2805,N_4317);
nand U5783 (N_5783,N_1683,N_4653);
xnor U5784 (N_5784,N_4733,N_1303);
or U5785 (N_5785,N_2626,N_3250);
nand U5786 (N_5786,N_2283,N_582);
or U5787 (N_5787,N_4765,N_3656);
or U5788 (N_5788,N_3917,N_4788);
xor U5789 (N_5789,N_2155,N_2852);
or U5790 (N_5790,N_1791,N_1093);
or U5791 (N_5791,N_4621,N_4099);
xnor U5792 (N_5792,N_1199,N_2041);
nor U5793 (N_5793,N_2046,N_4844);
or U5794 (N_5794,N_2948,N_1956);
and U5795 (N_5795,N_3573,N_1573);
and U5796 (N_5796,N_2683,N_4792);
or U5797 (N_5797,N_3868,N_2255);
nor U5798 (N_5798,N_3209,N_3153);
nor U5799 (N_5799,N_4982,N_4786);
nand U5800 (N_5800,N_45,N_1060);
and U5801 (N_5801,N_4822,N_96);
xor U5802 (N_5802,N_2207,N_106);
and U5803 (N_5803,N_830,N_3693);
nor U5804 (N_5804,N_1198,N_2456);
nand U5805 (N_5805,N_4147,N_2970);
xnor U5806 (N_5806,N_4505,N_3991);
nand U5807 (N_5807,N_3956,N_1506);
nand U5808 (N_5808,N_1391,N_1368);
or U5809 (N_5809,N_4611,N_4350);
nand U5810 (N_5810,N_2838,N_2345);
nand U5811 (N_5811,N_3768,N_1840);
nand U5812 (N_5812,N_4257,N_3377);
xnor U5813 (N_5813,N_1794,N_1632);
or U5814 (N_5814,N_4533,N_1749);
or U5815 (N_5815,N_3473,N_3520);
nor U5816 (N_5816,N_2426,N_3838);
nor U5817 (N_5817,N_419,N_1565);
nor U5818 (N_5818,N_4096,N_4819);
or U5819 (N_5819,N_1737,N_2938);
and U5820 (N_5820,N_2060,N_4672);
nand U5821 (N_5821,N_1233,N_2565);
nor U5822 (N_5822,N_2929,N_955);
nor U5823 (N_5823,N_220,N_239);
and U5824 (N_5824,N_3738,N_3008);
xor U5825 (N_5825,N_4965,N_2728);
or U5826 (N_5826,N_436,N_2480);
and U5827 (N_5827,N_604,N_717);
nand U5828 (N_5828,N_1297,N_1343);
and U5829 (N_5829,N_4589,N_749);
nor U5830 (N_5830,N_1231,N_494);
nand U5831 (N_5831,N_4967,N_296);
nor U5832 (N_5832,N_277,N_1531);
and U5833 (N_5833,N_361,N_2124);
xor U5834 (N_5834,N_819,N_1374);
or U5835 (N_5835,N_4249,N_2774);
or U5836 (N_5836,N_4465,N_2535);
nor U5837 (N_5837,N_2916,N_720);
nor U5838 (N_5838,N_2795,N_1373);
or U5839 (N_5839,N_3872,N_1548);
nor U5840 (N_5840,N_3850,N_2319);
xor U5841 (N_5841,N_4764,N_1133);
xor U5842 (N_5842,N_1129,N_1141);
or U5843 (N_5843,N_2196,N_88);
and U5844 (N_5844,N_1727,N_1478);
and U5845 (N_5845,N_374,N_1046);
xor U5846 (N_5846,N_1355,N_4089);
nor U5847 (N_5847,N_1833,N_4990);
xor U5848 (N_5848,N_4962,N_2606);
and U5849 (N_5849,N_4959,N_4743);
nor U5850 (N_5850,N_43,N_1912);
xor U5851 (N_5851,N_3381,N_721);
or U5852 (N_5852,N_1543,N_3501);
or U5853 (N_5853,N_339,N_2687);
nor U5854 (N_5854,N_2153,N_3619);
or U5855 (N_5855,N_4245,N_1069);
xor U5856 (N_5856,N_3199,N_714);
nor U5857 (N_5857,N_1120,N_4939);
xor U5858 (N_5858,N_4867,N_3480);
nand U5859 (N_5859,N_923,N_722);
and U5860 (N_5860,N_1449,N_383);
nor U5861 (N_5861,N_1152,N_2841);
nand U5862 (N_5862,N_597,N_1098);
nor U5863 (N_5863,N_1762,N_1139);
nor U5864 (N_5864,N_778,N_1759);
xor U5865 (N_5865,N_1758,N_1249);
nand U5866 (N_5866,N_2346,N_2002);
nand U5867 (N_5867,N_4220,N_3169);
and U5868 (N_5868,N_828,N_773);
and U5869 (N_5869,N_3801,N_2693);
xor U5870 (N_5870,N_2431,N_67);
or U5871 (N_5871,N_677,N_2904);
xor U5872 (N_5872,N_2168,N_3502);
or U5873 (N_5873,N_3729,N_1);
and U5874 (N_5874,N_689,N_3349);
or U5875 (N_5875,N_4160,N_2008);
nor U5876 (N_5876,N_2019,N_1003);
nand U5877 (N_5877,N_860,N_4757);
nand U5878 (N_5878,N_3330,N_931);
and U5879 (N_5879,N_1424,N_4598);
nor U5880 (N_5880,N_442,N_3810);
nor U5881 (N_5881,N_3579,N_1751);
nand U5882 (N_5882,N_1239,N_3512);
xnor U5883 (N_5883,N_2902,N_2917);
nand U5884 (N_5884,N_990,N_4799);
or U5885 (N_5885,N_3547,N_4779);
xor U5886 (N_5886,N_2654,N_74);
and U5887 (N_5887,N_844,N_2395);
xnor U5888 (N_5888,N_181,N_4880);
and U5889 (N_5889,N_1326,N_2082);
or U5890 (N_5890,N_2971,N_4060);
nand U5891 (N_5891,N_4265,N_4674);
or U5892 (N_5892,N_1795,N_2679);
and U5893 (N_5893,N_365,N_976);
xnor U5894 (N_5894,N_2602,N_4167);
nand U5895 (N_5895,N_1053,N_4813);
xnor U5896 (N_5896,N_1074,N_3795);
nand U5897 (N_5897,N_370,N_1741);
xnor U5898 (N_5898,N_2808,N_4396);
nor U5899 (N_5899,N_2653,N_2860);
xnor U5900 (N_5900,N_998,N_4787);
and U5901 (N_5901,N_3666,N_3706);
or U5902 (N_5902,N_1377,N_2379);
or U5903 (N_5903,N_1987,N_2678);
or U5904 (N_5904,N_4118,N_1356);
or U5905 (N_5905,N_527,N_3830);
nand U5906 (N_5906,N_200,N_3428);
or U5907 (N_5907,N_613,N_3321);
nor U5908 (N_5908,N_4541,N_4655);
nand U5909 (N_5909,N_3383,N_4471);
and U5910 (N_5910,N_922,N_2597);
nand U5911 (N_5911,N_1846,N_4862);
and U5912 (N_5912,N_1557,N_4838);
nand U5913 (N_5913,N_1256,N_2370);
and U5914 (N_5914,N_2979,N_1906);
or U5915 (N_5915,N_1627,N_2220);
xnor U5916 (N_5916,N_2779,N_4721);
nand U5917 (N_5917,N_1790,N_180);
nand U5918 (N_5918,N_3517,N_767);
nor U5919 (N_5919,N_4731,N_975);
nand U5920 (N_5920,N_2542,N_3890);
nand U5921 (N_5921,N_823,N_3504);
nand U5922 (N_5922,N_452,N_3625);
nor U5923 (N_5923,N_2292,N_4026);
or U5924 (N_5924,N_2721,N_3691);
nand U5925 (N_5925,N_4663,N_4866);
or U5926 (N_5926,N_1213,N_964);
or U5927 (N_5927,N_298,N_866);
or U5928 (N_5928,N_1229,N_4558);
and U5929 (N_5929,N_4015,N_3395);
nand U5930 (N_5930,N_1765,N_2401);
nor U5931 (N_5931,N_3652,N_1698);
or U5932 (N_5932,N_891,N_3823);
nor U5933 (N_5933,N_3085,N_1274);
and U5934 (N_5934,N_2029,N_1868);
xnor U5935 (N_5935,N_2986,N_1993);
and U5936 (N_5936,N_1363,N_4855);
nand U5937 (N_5937,N_338,N_4318);
xor U5938 (N_5938,N_4916,N_4797);
nand U5939 (N_5939,N_4798,N_3971);
and U5940 (N_5940,N_4331,N_4504);
and U5941 (N_5941,N_505,N_962);
nor U5942 (N_5942,N_4915,N_4818);
nand U5943 (N_5943,N_2312,N_1643);
and U5944 (N_5944,N_3698,N_455);
or U5945 (N_5945,N_4148,N_1468);
xor U5946 (N_5946,N_580,N_344);
nand U5947 (N_5947,N_1519,N_4984);
nand U5948 (N_5948,N_3796,N_2512);
or U5949 (N_5949,N_2862,N_661);
nand U5950 (N_5950,N_4176,N_3003);
and U5951 (N_5951,N_1947,N_3218);
xnor U5952 (N_5952,N_4182,N_1584);
nand U5953 (N_5953,N_1555,N_4567);
nor U5954 (N_5954,N_2921,N_1237);
or U5955 (N_5955,N_3130,N_3866);
nor U5956 (N_5956,N_307,N_357);
nor U5957 (N_5957,N_741,N_2410);
or U5958 (N_5958,N_3574,N_2131);
nor U5959 (N_5959,N_3871,N_3704);
xnor U5960 (N_5960,N_4856,N_1615);
nand U5961 (N_5961,N_3301,N_895);
nand U5962 (N_5962,N_3230,N_1336);
xor U5963 (N_5963,N_1704,N_1190);
nor U5964 (N_5964,N_340,N_592);
nor U5965 (N_5965,N_3121,N_369);
nand U5966 (N_5966,N_1118,N_2749);
xor U5967 (N_5967,N_2173,N_4253);
and U5968 (N_5968,N_3098,N_1448);
xnor U5969 (N_5969,N_1771,N_3457);
nor U5970 (N_5970,N_3805,N_3129);
nand U5971 (N_5971,N_2407,N_2042);
nor U5972 (N_5972,N_1930,N_3136);
xnor U5973 (N_5973,N_2063,N_635);
nor U5974 (N_5974,N_565,N_2349);
and U5975 (N_5975,N_4361,N_3684);
or U5976 (N_5976,N_1953,N_4063);
nand U5977 (N_5977,N_3054,N_216);
nand U5978 (N_5978,N_4203,N_2894);
nand U5979 (N_5979,N_362,N_3775);
nand U5980 (N_5980,N_1755,N_636);
nor U5981 (N_5981,N_3730,N_2959);
and U5982 (N_5982,N_874,N_4179);
nor U5983 (N_5983,N_560,N_2286);
and U5984 (N_5984,N_2109,N_3668);
or U5985 (N_5985,N_4185,N_2608);
nor U5986 (N_5986,N_2981,N_4919);
xor U5987 (N_5987,N_3919,N_3721);
nand U5988 (N_5988,N_1945,N_1184);
nor U5989 (N_5989,N_3268,N_1268);
nor U5990 (N_5990,N_1836,N_3728);
nor U5991 (N_5991,N_4139,N_2634);
nor U5992 (N_5992,N_3055,N_1054);
nor U5993 (N_5993,N_3769,N_2692);
or U5994 (N_5994,N_3238,N_4473);
or U5995 (N_5995,N_2704,N_1774);
nand U5996 (N_5996,N_1828,N_532);
xnor U5997 (N_5997,N_3989,N_2364);
xor U5998 (N_5998,N_2268,N_396);
or U5999 (N_5999,N_309,N_356);
nor U6000 (N_6000,N_761,N_657);
xnor U6001 (N_6001,N_3352,N_299);
or U6002 (N_6002,N_2236,N_1497);
nand U6003 (N_6003,N_3101,N_1979);
nor U6004 (N_6004,N_2724,N_4010);
or U6005 (N_6005,N_1037,N_2621);
nand U6006 (N_6006,N_1167,N_3851);
or U6007 (N_6007,N_4248,N_4861);
or U6008 (N_6008,N_1936,N_2061);
xor U6009 (N_6009,N_1045,N_3078);
and U6010 (N_6010,N_2870,N_3030);
and U6011 (N_6011,N_2884,N_2713);
nor U6012 (N_6012,N_4701,N_330);
nand U6013 (N_6013,N_2348,N_349);
xnor U6014 (N_6014,N_3665,N_1398);
or U6015 (N_6015,N_1660,N_1909);
xnor U6016 (N_6016,N_4126,N_2383);
xor U6017 (N_6017,N_4949,N_3739);
xnor U6018 (N_6018,N_1496,N_1510);
or U6019 (N_6019,N_2149,N_1147);
nand U6020 (N_6020,N_254,N_1104);
or U6021 (N_6021,N_852,N_3143);
xnor U6022 (N_6022,N_1875,N_1536);
nand U6023 (N_6023,N_1843,N_782);
xnor U6024 (N_6024,N_503,N_3814);
xor U6025 (N_6025,N_4665,N_585);
and U6026 (N_6026,N_3819,N_2811);
xnor U6027 (N_6027,N_2361,N_391);
and U6028 (N_6028,N_4178,N_2983);
or U6029 (N_6029,N_4319,N_1693);
nor U6030 (N_6030,N_4529,N_2719);
xor U6031 (N_6031,N_2440,N_3998);
nor U6032 (N_6032,N_4136,N_4124);
nor U6033 (N_6033,N_2898,N_4705);
nand U6034 (N_6034,N_3179,N_683);
nor U6035 (N_6035,N_476,N_877);
nand U6036 (N_6036,N_559,N_1962);
nor U6037 (N_6037,N_1721,N_2690);
nor U6038 (N_6038,N_3577,N_2854);
nor U6039 (N_6039,N_915,N_27);
nand U6040 (N_6040,N_1931,N_1043);
or U6041 (N_6041,N_900,N_1309);
xnor U6042 (N_6042,N_491,N_4563);
xor U6043 (N_6043,N_1217,N_839);
nand U6044 (N_6044,N_4379,N_4337);
and U6045 (N_6045,N_4009,N_234);
nor U6046 (N_6046,N_8,N_378);
and U6047 (N_6047,N_59,N_2021);
and U6048 (N_6048,N_4791,N_3311);
and U6049 (N_6049,N_1651,N_4634);
xnor U6050 (N_6050,N_2015,N_1475);
xor U6051 (N_6051,N_3018,N_1576);
xnor U6052 (N_6052,N_2388,N_2414);
and U6053 (N_6053,N_1667,N_1881);
xor U6054 (N_6054,N_4169,N_2667);
nand U6055 (N_6055,N_4795,N_3147);
nand U6056 (N_6056,N_366,N_237);
nor U6057 (N_6057,N_3363,N_2);
or U6058 (N_6058,N_2707,N_2892);
nor U6059 (N_6059,N_2629,N_3486);
nor U6060 (N_6060,N_2886,N_4054);
or U6061 (N_6061,N_4752,N_2845);
xnor U6062 (N_6062,N_4609,N_3272);
nand U6063 (N_6063,N_171,N_2590);
and U6064 (N_6064,N_3578,N_875);
and U6065 (N_6065,N_1511,N_2833);
or U6066 (N_6066,N_3986,N_1894);
xor U6067 (N_6067,N_4196,N_4829);
and U6068 (N_6068,N_2674,N_1070);
nor U6069 (N_6069,N_401,N_2218);
xnor U6070 (N_6070,N_3088,N_60);
nor U6071 (N_6071,N_1583,N_1610);
nor U6072 (N_6072,N_243,N_1307);
or U6073 (N_6073,N_726,N_659);
xnor U6074 (N_6074,N_4895,N_1731);
and U6075 (N_6075,N_3827,N_2027);
and U6076 (N_6076,N_2010,N_3694);
or U6077 (N_6077,N_1708,N_1328);
and U6078 (N_6078,N_1438,N_2880);
nand U6079 (N_6079,N_4281,N_4521);
or U6080 (N_6080,N_2820,N_2433);
or U6081 (N_6081,N_3255,N_3541);
nor U6082 (N_6082,N_4591,N_3855);
nand U6083 (N_6083,N_1271,N_3099);
nand U6084 (N_6084,N_4881,N_4114);
and U6085 (N_6085,N_1369,N_3647);
xor U6086 (N_6086,N_1063,N_3534);
nor U6087 (N_6087,N_4846,N_2587);
nand U6088 (N_6088,N_3978,N_2285);
xnor U6089 (N_6089,N_4717,N_728);
and U6090 (N_6090,N_4119,N_2998);
nor U6091 (N_6091,N_354,N_19);
and U6092 (N_6092,N_4884,N_1126);
or U6093 (N_6093,N_3041,N_434);
or U6094 (N_6094,N_2488,N_3907);
nor U6095 (N_6095,N_1750,N_2094);
nand U6096 (N_6096,N_151,N_2655);
nor U6097 (N_6097,N_1631,N_2623);
xnor U6098 (N_6098,N_3148,N_4671);
nand U6099 (N_6099,N_4707,N_238);
nor U6100 (N_6100,N_4728,N_1258);
or U6101 (N_6101,N_1228,N_785);
nand U6102 (N_6102,N_1127,N_4848);
or U6103 (N_6103,N_1571,N_1379);
xor U6104 (N_6104,N_2744,N_2166);
xor U6105 (N_6105,N_4830,N_4437);
nor U6106 (N_6106,N_1488,N_1482);
nand U6107 (N_6107,N_4496,N_4462);
and U6108 (N_6108,N_475,N_921);
or U6109 (N_6109,N_2521,N_4053);
and U6110 (N_6110,N_3618,N_1852);
nand U6111 (N_6111,N_2969,N_2394);
nand U6112 (N_6112,N_4506,N_2670);
and U6113 (N_6113,N_1302,N_747);
and U6114 (N_6114,N_460,N_2844);
and U6115 (N_6115,N_3154,N_3664);
or U6116 (N_6116,N_1182,N_2137);
nor U6117 (N_6117,N_2073,N_1949);
nand U6118 (N_6118,N_3093,N_521);
and U6119 (N_6119,N_2963,N_3445);
or U6120 (N_6120,N_4737,N_1792);
or U6121 (N_6121,N_2738,N_904);
nand U6122 (N_6122,N_563,N_4991);
nor U6123 (N_6123,N_1437,N_1640);
xor U6124 (N_6124,N_555,N_223);
or U6125 (N_6125,N_3791,N_195);
or U6126 (N_6126,N_3359,N_2362);
and U6127 (N_6127,N_610,N_79);
nor U6128 (N_6128,N_4580,N_957);
or U6129 (N_6129,N_456,N_2340);
and U6130 (N_6130,N_802,N_886);
or U6131 (N_6131,N_3820,N_4162);
and U6132 (N_6132,N_2302,N_4805);
and U6133 (N_6133,N_4746,N_2620);
nand U6134 (N_6134,N_1101,N_3984);
nand U6135 (N_6135,N_4850,N_562);
xor U6136 (N_6136,N_2589,N_812);
nor U6137 (N_6137,N_77,N_2435);
nor U6138 (N_6138,N_3879,N_4768);
nand U6139 (N_6139,N_4524,N_4252);
or U6140 (N_6140,N_158,N_2740);
nor U6141 (N_6141,N_1062,N_4793);
and U6142 (N_6142,N_4775,N_2701);
xnor U6143 (N_6143,N_2402,N_1279);
nand U6144 (N_6144,N_3702,N_508);
and U6145 (N_6145,N_1023,N_2107);
nor U6146 (N_6146,N_4387,N_2930);
nand U6147 (N_6147,N_3335,N_1230);
or U6148 (N_6148,N_4476,N_2424);
or U6149 (N_6149,N_960,N_4751);
nand U6150 (N_6150,N_1539,N_4540);
nand U6151 (N_6151,N_3399,N_3779);
and U6152 (N_6152,N_1114,N_2169);
xor U6153 (N_6153,N_3104,N_3224);
xnor U6154 (N_6154,N_4583,N_2493);
xor U6155 (N_6155,N_3649,N_4909);
and U6156 (N_6156,N_634,N_3622);
or U6157 (N_6157,N_1959,N_1682);
nand U6158 (N_6158,N_1011,N_1138);
nand U6159 (N_6159,N_3799,N_2350);
nand U6160 (N_6160,N_4644,N_1466);
nor U6161 (N_6161,N_3298,N_2513);
or U6162 (N_6162,N_1515,N_2387);
xor U6163 (N_6163,N_1067,N_759);
nor U6164 (N_6164,N_4320,N_666);
nor U6165 (N_6165,N_3103,N_4814);
nor U6166 (N_6166,N_3549,N_4012);
xor U6167 (N_6167,N_3570,N_17);
nor U6168 (N_6168,N_3175,N_1081);
xnor U6169 (N_6169,N_4441,N_3964);
nor U6170 (N_6170,N_7,N_4276);
nand U6171 (N_6171,N_1387,N_4956);
nor U6172 (N_6172,N_2857,N_2050);
nor U6173 (N_6173,N_1505,N_4300);
nor U6174 (N_6174,N_628,N_275);
nand U6175 (N_6175,N_468,N_4238);
or U6176 (N_6176,N_4006,N_3232);
and U6177 (N_6177,N_4448,N_4628);
xnor U6178 (N_6178,N_1589,N_3832);
nand U6179 (N_6179,N_3114,N_2126);
nand U6180 (N_6180,N_3483,N_4469);
or U6181 (N_6181,N_878,N_3126);
xnor U6182 (N_6182,N_430,N_2472);
xnor U6183 (N_6183,N_1756,N_2891);
and U6184 (N_6184,N_3462,N_1148);
or U6185 (N_6185,N_4870,N_4900);
and U6186 (N_6186,N_836,N_3839);
and U6187 (N_6187,N_3288,N_1920);
nor U6188 (N_6188,N_4934,N_1996);
xor U6189 (N_6189,N_4405,N_2520);
nand U6190 (N_6190,N_3207,N_1380);
nor U6191 (N_6191,N_2443,N_4697);
xnor U6192 (N_6192,N_704,N_3027);
nand U6193 (N_6193,N_4664,N_2603);
or U6194 (N_6194,N_242,N_1918);
nand U6195 (N_6195,N_3242,N_3789);
or U6196 (N_6196,N_3628,N_1193);
xnor U6197 (N_6197,N_1716,N_2007);
and U6198 (N_6198,N_2659,N_1815);
xor U6199 (N_6199,N_1333,N_1430);
or U6200 (N_6200,N_2649,N_995);
or U6201 (N_6201,N_4108,N_202);
xor U6202 (N_6202,N_3732,N_240);
nand U6203 (N_6203,N_3000,N_4516);
or U6204 (N_6204,N_2727,N_568);
and U6205 (N_6205,N_150,N_3784);
nand U6206 (N_6206,N_1017,N_758);
or U6207 (N_6207,N_4658,N_2836);
and U6208 (N_6208,N_1786,N_394);
nand U6209 (N_6209,N_4467,N_130);
nor U6210 (N_6210,N_3211,N_1345);
nand U6211 (N_6211,N_328,N_632);
or U6212 (N_6212,N_117,N_3115);
nor U6213 (N_6213,N_4785,N_2148);
and U6214 (N_6214,N_1366,N_1675);
nor U6215 (N_6215,N_4588,N_3314);
nor U6216 (N_6216,N_3596,N_892);
nor U6217 (N_6217,N_501,N_2864);
and U6218 (N_6218,N_2004,N_1477);
and U6219 (N_6219,N_3900,N_4519);
xnor U6220 (N_6220,N_4373,N_56);
and U6221 (N_6221,N_1664,N_4641);
or U6222 (N_6222,N_2919,N_4100);
and U6223 (N_6223,N_1210,N_3672);
xnor U6224 (N_6224,N_334,N_2506);
nand U6225 (N_6225,N_2203,N_3863);
xor U6226 (N_6226,N_2706,N_2341);
xor U6227 (N_6227,N_1185,N_4508);
nor U6228 (N_6228,N_1581,N_2751);
xnor U6229 (N_6229,N_734,N_1746);
and U6230 (N_6230,N_4093,N_3701);
xnor U6231 (N_6231,N_4417,N_3313);
nor U6232 (N_6232,N_4555,N_3348);
and U6233 (N_6233,N_170,N_578);
and U6234 (N_6234,N_4394,N_4112);
or U6235 (N_6235,N_1872,N_4527);
or U6236 (N_6236,N_4115,N_1402);
xor U6237 (N_6237,N_2514,N_326);
xor U6238 (N_6238,N_4986,N_166);
nor U6239 (N_6239,N_587,N_3629);
or U6240 (N_6240,N_4565,N_4587);
nor U6241 (N_6241,N_1295,N_1850);
nand U6242 (N_6242,N_4098,N_3182);
or U6243 (N_6243,N_2829,N_2457);
and U6244 (N_6244,N_2325,N_3997);
xnor U6245 (N_6245,N_1730,N_1782);
xnor U6246 (N_6246,N_3490,N_3317);
xnor U6247 (N_6247,N_3493,N_925);
or U6248 (N_6248,N_3282,N_2423);
and U6249 (N_6249,N_3380,N_3675);
nand U6250 (N_6250,N_2723,N_4191);
nor U6251 (N_6251,N_3061,N_4211);
nor U6252 (N_6252,N_4547,N_4905);
or U6253 (N_6253,N_4596,N_2248);
xor U6254 (N_6254,N_4526,N_3563);
nor U6255 (N_6255,N_3687,N_3950);
nand U6256 (N_6256,N_1865,N_444);
or U6257 (N_6257,N_4678,N_4906);
or U6258 (N_6258,N_712,N_1078);
or U6259 (N_6259,N_2604,N_1837);
nor U6260 (N_6260,N_2090,N_506);
nor U6261 (N_6261,N_1440,N_544);
nand U6262 (N_6262,N_4202,N_1575);
and U6263 (N_6263,N_2636,N_1626);
or U6264 (N_6264,N_3650,N_4756);
or U6265 (N_6265,N_4623,N_2933);
nand U6266 (N_6266,N_4050,N_3510);
xnor U6267 (N_6267,N_3469,N_3080);
nor U6268 (N_6268,N_2686,N_1320);
and U6269 (N_6269,N_2232,N_3040);
xor U6270 (N_6270,N_4815,N_968);
nor U6271 (N_6271,N_1614,N_4625);
and U6272 (N_6272,N_2806,N_2409);
or U6273 (N_6273,N_1988,N_2843);
xnor U6274 (N_6274,N_1119,N_2084);
and U6275 (N_6275,N_4650,N_482);
and U6276 (N_6276,N_3347,N_3215);
and U6277 (N_6277,N_1800,N_4088);
nor U6278 (N_6278,N_947,N_1188);
nor U6279 (N_6279,N_4910,N_2159);
nand U6280 (N_6280,N_2035,N_4398);
nor U6281 (N_6281,N_3176,N_540);
or U6282 (N_6282,N_4461,N_4329);
nand U6283 (N_6283,N_3376,N_1441);
and U6284 (N_6284,N_1022,N_3390);
or U6285 (N_6285,N_576,N_1990);
or U6286 (N_6286,N_2338,N_1514);
xnor U6287 (N_6287,N_4314,N_2639);
or U6288 (N_6288,N_3572,N_1232);
nand U6289 (N_6289,N_4458,N_2211);
or U6290 (N_6290,N_3198,N_2235);
nor U6291 (N_6291,N_3536,N_2666);
nor U6292 (N_6292,N_2427,N_297);
or U6293 (N_6293,N_4762,N_2676);
and U6294 (N_6294,N_940,N_3292);
nand U6295 (N_6295,N_392,N_668);
nor U6296 (N_6296,N_268,N_127);
and U6297 (N_6297,N_4172,N_988);
nand U6298 (N_6298,N_2097,N_2377);
nand U6299 (N_6299,N_1616,N_3829);
nand U6300 (N_6300,N_752,N_2368);
xor U6301 (N_6301,N_1533,N_3245);
or U6302 (N_6302,N_1301,N_2227);
or U6303 (N_6303,N_97,N_3717);
and U6304 (N_6304,N_4924,N_4974);
or U6305 (N_6305,N_2925,N_4004);
or U6306 (N_6306,N_710,N_2099);
nor U6307 (N_6307,N_2125,N_3802);
and U6308 (N_6308,N_2580,N_3600);
nand U6309 (N_6309,N_4518,N_2977);
or U6310 (N_6310,N_4003,N_4615);
xor U6311 (N_6311,N_4706,N_1009);
xnor U6312 (N_6312,N_2121,N_2628);
xnor U6313 (N_6313,N_2881,N_675);
nand U6314 (N_6314,N_3084,N_2871);
nand U6315 (N_6315,N_708,N_653);
or U6316 (N_6316,N_709,N_1094);
nand U6317 (N_6317,N_1151,N_4560);
nor U6318 (N_6318,N_4480,N_1238);
xnor U6319 (N_6319,N_2822,N_4940);
and U6320 (N_6320,N_4047,N_3064);
nand U6321 (N_6321,N_2057,N_2284);
xor U6322 (N_6322,N_3921,N_3426);
nor U6323 (N_6323,N_680,N_1347);
xor U6324 (N_6324,N_2184,N_3138);
nand U6325 (N_6325,N_48,N_2637);
xnor U6326 (N_6326,N_2306,N_1030);
nor U6327 (N_6327,N_723,N_2461);
and U6328 (N_6328,N_2501,N_4886);
or U6329 (N_6329,N_3326,N_428);
nand U6330 (N_6330,N_3048,N_4645);
or U6331 (N_6331,N_4722,N_2245);
nor U6332 (N_6332,N_643,N_4071);
or U6333 (N_6333,N_2231,N_2020);
and U6334 (N_6334,N_4740,N_2026);
or U6335 (N_6335,N_4360,N_93);
xnor U6336 (N_6336,N_2376,N_3726);
nand U6337 (N_6337,N_4213,N_2406);
and U6338 (N_6338,N_569,N_80);
xnor U6339 (N_6339,N_2784,N_184);
or U6340 (N_6340,N_1927,N_4432);
or U6341 (N_6341,N_1021,N_4590);
or U6342 (N_6342,N_3435,N_61);
or U6343 (N_6343,N_1537,N_4605);
or U6344 (N_6344,N_3178,N_192);
nor U6345 (N_6345,N_2572,N_2961);
nand U6346 (N_6346,N_4987,N_1200);
xor U6347 (N_6347,N_3177,N_1049);
nand U6348 (N_6348,N_2791,N_1585);
nand U6349 (N_6349,N_2418,N_210);
or U6350 (N_6350,N_4941,N_2261);
and U6351 (N_6351,N_4135,N_4573);
or U6352 (N_6352,N_1175,N_3887);
xor U6353 (N_6353,N_1015,N_4556);
and U6354 (N_6354,N_3962,N_3894);
and U6355 (N_6355,N_4013,N_316);
nor U6356 (N_6356,N_4501,N_2770);
xor U6357 (N_6357,N_3580,N_1038);
nand U6358 (N_6358,N_3087,N_913);
nand U6359 (N_6359,N_2566,N_4566);
nor U6360 (N_6360,N_2479,N_2367);
nor U6361 (N_6361,N_163,N_3516);
nand U6362 (N_6362,N_3411,N_3542);
and U6363 (N_6363,N_3653,N_4039);
xor U6364 (N_6364,N_4958,N_4927);
and U6365 (N_6365,N_1375,N_283);
xor U6366 (N_6366,N_4873,N_3834);
nand U6367 (N_6367,N_2522,N_2877);
xor U6368 (N_6368,N_3575,N_2523);
xor U6369 (N_6369,N_1209,N_4686);
and U6370 (N_6370,N_2403,N_2717);
and U6371 (N_6371,N_2818,N_590);
or U6372 (N_6372,N_883,N_3959);
nor U6373 (N_6373,N_2210,N_3122);
nand U6374 (N_6374,N_3816,N_345);
or U6375 (N_6375,N_4206,N_2069);
nand U6376 (N_6376,N_1044,N_4874);
nand U6377 (N_6377,N_2546,N_3229);
and U6378 (N_6378,N_155,N_3470);
nor U6379 (N_6379,N_1084,N_1981);
and U6380 (N_6380,N_2786,N_2037);
nand U6381 (N_6381,N_4372,N_2087);
or U6382 (N_6382,N_2044,N_214);
nor U6383 (N_6383,N_2132,N_4490);
nand U6384 (N_6384,N_853,N_3506);
nand U6385 (N_6385,N_818,N_1109);
nor U6386 (N_6386,N_3566,N_2596);
nand U6387 (N_6387,N_4032,N_833);
nor U6388 (N_6388,N_4340,N_22);
nor U6389 (N_6389,N_2422,N_981);
xnor U6390 (N_6390,N_3569,N_3438);
or U6391 (N_6391,N_3495,N_2570);
or U6392 (N_6392,N_1942,N_2353);
xnor U6393 (N_6393,N_2924,N_2451);
or U6394 (N_6394,N_3374,N_3847);
nor U6395 (N_6395,N_4381,N_3275);
and U6396 (N_6396,N_3083,N_3237);
or U6397 (N_6397,N_3794,N_3828);
or U6398 (N_6398,N_353,N_409);
and U6399 (N_6399,N_3185,N_1036);
nand U6400 (N_6400,N_2033,N_3164);
and U6401 (N_6401,N_4173,N_2515);
and U6402 (N_6402,N_4380,N_3567);
nand U6403 (N_6403,N_1135,N_4216);
nor U6404 (N_6404,N_2528,N_4326);
xor U6405 (N_6405,N_4367,N_1240);
or U6406 (N_6406,N_2181,N_3388);
nor U6407 (N_6407,N_4700,N_1371);
or U6408 (N_6408,N_2538,N_3635);
nand U6409 (N_6409,N_131,N_3709);
nand U6410 (N_6410,N_854,N_4349);
nor U6411 (N_6411,N_3793,N_2688);
nor U6412 (N_6412,N_3909,N_3067);
nor U6413 (N_6413,N_2812,N_281);
nor U6414 (N_6414,N_69,N_2163);
nand U6415 (N_6415,N_402,N_2955);
nand U6416 (N_6416,N_4868,N_4836);
nand U6417 (N_6417,N_198,N_3368);
or U6418 (N_6418,N_2823,N_3727);
xnor U6419 (N_6419,N_1622,N_118);
nand U6420 (N_6420,N_4930,N_3220);
xnor U6421 (N_6421,N_969,N_584);
or U6422 (N_6422,N_1029,N_989);
nor U6423 (N_6423,N_2932,N_4122);
and U6424 (N_6424,N_1498,N_2078);
and U6425 (N_6425,N_3170,N_4413);
and U6426 (N_6426,N_4075,N_24);
nand U6427 (N_6427,N_140,N_1422);
nor U6428 (N_6428,N_1926,N_932);
and U6429 (N_6429,N_49,N_304);
nand U6430 (N_6430,N_4207,N_2561);
and U6431 (N_6431,N_1857,N_3333);
nor U6432 (N_6432,N_1776,N_2510);
or U6433 (N_6433,N_2058,N_961);
and U6434 (N_6434,N_3557,N_2195);
xnor U6435 (N_6435,N_3478,N_2962);
nor U6436 (N_6436,N_3712,N_3166);
nor U6437 (N_6437,N_4234,N_1896);
nand U6438 (N_6438,N_1620,N_1686);
or U6439 (N_6439,N_4613,N_2912);
nor U6440 (N_6440,N_3074,N_2180);
and U6441 (N_6441,N_4592,N_905);
xor U6442 (N_6442,N_3197,N_218);
nand U6443 (N_6443,N_4036,N_1732);
nand U6444 (N_6444,N_768,N_739);
nand U6445 (N_6445,N_4102,N_2378);
nor U6446 (N_6446,N_1891,N_541);
and U6447 (N_6447,N_4497,N_4735);
xnor U6448 (N_6448,N_1327,N_3658);
nor U6449 (N_6449,N_3405,N_507);
nand U6450 (N_6450,N_4892,N_3809);
nor U6451 (N_6451,N_2188,N_3910);
or U6452 (N_6452,N_3953,N_3546);
or U6453 (N_6453,N_3082,N_4219);
xor U6454 (N_6454,N_4920,N_4869);
or U6455 (N_6455,N_2179,N_2380);
nor U6456 (N_6456,N_917,N_2189);
and U6457 (N_6457,N_2304,N_347);
or U6458 (N_6458,N_233,N_2562);
and U6459 (N_6459,N_284,N_2769);
nand U6460 (N_6460,N_3355,N_2966);
xor U6461 (N_6461,N_2117,N_3124);
nor U6462 (N_6462,N_4837,N_2819);
or U6463 (N_6463,N_889,N_2552);
or U6464 (N_6464,N_2307,N_1856);
nor U6465 (N_6465,N_4454,N_425);
xor U6466 (N_6466,N_3174,N_55);
nor U6467 (N_6467,N_3920,N_3026);
nand U6468 (N_6468,N_110,N_4240);
nor U6469 (N_6469,N_4478,N_3278);
and U6470 (N_6470,N_2985,N_4447);
or U6471 (N_6471,N_336,N_3315);
and U6472 (N_6472,N_3994,N_1948);
xnor U6473 (N_6473,N_2205,N_3339);
xnor U6474 (N_6474,N_1740,N_3408);
or U6475 (N_6475,N_4254,N_4389);
and U6476 (N_6476,N_663,N_2720);
and U6477 (N_6477,N_3804,N_4277);
and U6478 (N_6478,N_941,N_1425);
nand U6479 (N_6479,N_4021,N_3992);
and U6480 (N_6480,N_4750,N_2246);
nor U6481 (N_6481,N_1504,N_786);
and U6482 (N_6482,N_1650,N_3674);
nand U6483 (N_6483,N_523,N_2773);
xnor U6484 (N_6484,N_3259,N_3759);
and U6485 (N_6485,N_757,N_3267);
and U6486 (N_6486,N_3914,N_1526);
nand U6487 (N_6487,N_3058,N_3274);
nand U6488 (N_6488,N_310,N_751);
xor U6489 (N_6489,N_3670,N_4086);
nand U6490 (N_6490,N_4290,N_4760);
nor U6491 (N_6491,N_3803,N_499);
or U6492 (N_6492,N_4781,N_2689);
nor U6493 (N_6493,N_2119,N_2764);
xor U6494 (N_6494,N_2085,N_3336);
xor U6495 (N_6495,N_3782,N_1444);
nand U6496 (N_6496,N_4575,N_3915);
nand U6497 (N_6497,N_2588,N_3461);
and U6498 (N_6498,N_4647,N_4789);
and U6499 (N_6499,N_2518,N_2271);
nand U6500 (N_6500,N_2290,N_4763);
nor U6501 (N_6501,N_2761,N_793);
or U6502 (N_6502,N_1288,N_774);
or U6503 (N_6503,N_124,N_856);
nand U6504 (N_6504,N_509,N_1162);
nand U6505 (N_6505,N_1115,N_1382);
xor U6506 (N_6506,N_4452,N_3316);
xor U6507 (N_6507,N_4246,N_4899);
nor U6508 (N_6508,N_4543,N_4842);
xnor U6509 (N_6509,N_1602,N_3004);
nand U6510 (N_6510,N_3402,N_2497);
nand U6511 (N_6511,N_3053,N_397);
nor U6512 (N_6512,N_471,N_1763);
and U6513 (N_6513,N_3561,N_2491);
nor U6514 (N_6514,N_3477,N_466);
nand U6515 (N_6515,N_2753,N_1884);
xor U6516 (N_6516,N_893,N_1892);
nor U6517 (N_6517,N_3476,N_4146);
and U6518 (N_6518,N_993,N_2732);
and U6519 (N_6519,N_3983,N_3305);
nand U6520 (N_6520,N_2601,N_159);
or U6521 (N_6521,N_4852,N_4500);
xor U6522 (N_6522,N_114,N_1502);
or U6523 (N_6523,N_2147,N_15);
and U6524 (N_6524,N_4790,N_1778);
nor U6525 (N_6525,N_1890,N_3063);
and U6526 (N_6526,N_1587,N_4298);
and U6527 (N_6527,N_1838,N_3420);
nand U6528 (N_6528,N_1691,N_672);
and U6529 (N_6529,N_3465,N_2646);
and U6530 (N_6530,N_2906,N_2430);
or U6531 (N_6531,N_3918,N_2863);
and U6532 (N_6532,N_1964,N_2112);
and U6533 (N_6533,N_2759,N_996);
xnor U6534 (N_6534,N_2991,N_4177);
xor U6535 (N_6535,N_3304,N_1316);
xor U6536 (N_6536,N_1091,N_2454);
nand U6537 (N_6537,N_2558,N_543);
xor U6538 (N_6538,N_1880,N_1170);
nand U6539 (N_6539,N_1825,N_3926);
or U6540 (N_6540,N_479,N_2108);
nand U6541 (N_6541,N_1970,N_4237);
and U6542 (N_6542,N_2618,N_2575);
xor U6543 (N_6543,N_3761,N_3837);
nand U6544 (N_6544,N_4980,N_3853);
nand U6545 (N_6545,N_4691,N_1735);
nand U6546 (N_6546,N_4807,N_1869);
and U6547 (N_6547,N_3515,N_4058);
nand U6548 (N_6548,N_3593,N_3002);
and U6549 (N_6549,N_1005,N_4351);
nor U6550 (N_6550,N_1915,N_4810);
and U6551 (N_6551,N_4964,N_1986);
and U6552 (N_6552,N_1965,N_3498);
or U6553 (N_6553,N_2194,N_2954);
and U6554 (N_6554,N_3056,N_4887);
nand U6555 (N_6555,N_2527,N_3308);
nand U6556 (N_6556,N_4711,N_1269);
and U6557 (N_6557,N_2038,N_545);
nand U6558 (N_6558,N_776,N_3662);
and U6559 (N_6559,N_4950,N_385);
nand U6560 (N_6560,N_2758,N_641);
nand U6561 (N_6561,N_2508,N_129);
or U6562 (N_6562,N_2303,N_535);
nor U6563 (N_6563,N_3999,N_4668);
or U6564 (N_6564,N_1783,N_3075);
xor U6565 (N_6565,N_1051,N_1197);
xor U6566 (N_6566,N_2673,N_4635);
nor U6567 (N_6567,N_4835,N_2178);
or U6568 (N_6568,N_2662,N_3733);
xor U6569 (N_6569,N_3609,N_2372);
or U6570 (N_6570,N_938,N_727);
nor U6571 (N_6571,N_186,N_4562);
nor U6572 (N_6572,N_2214,N_4738);
or U6573 (N_6573,N_4758,N_1317);
nand U6574 (N_6574,N_94,N_133);
xor U6575 (N_6575,N_393,N_1690);
or U6576 (N_6576,N_3375,N_4128);
or U6577 (N_6577,N_3425,N_4068);
and U6578 (N_6578,N_4161,N_1895);
or U6579 (N_6579,N_2120,N_1952);
and U6580 (N_6580,N_4876,N_1218);
and U6581 (N_6581,N_2641,N_4046);
and U6582 (N_6582,N_4283,N_291);
or U6583 (N_6583,N_3019,N_1695);
xor U6584 (N_6584,N_1474,N_2222);
nand U6585 (N_6585,N_1715,N_3052);
xor U6586 (N_6586,N_2766,N_1156);
or U6587 (N_6587,N_664,N_745);
and U6588 (N_6588,N_1376,N_848);
and U6589 (N_6589,N_2413,N_3453);
xnor U6590 (N_6590,N_1921,N_3059);
nor U6591 (N_6591,N_530,N_89);
or U6592 (N_6592,N_3246,N_4455);
xor U6593 (N_6593,N_187,N_522);
xor U6594 (N_6594,N_312,N_2474);
or U6595 (N_6595,N_4955,N_958);
nand U6596 (N_6596,N_4197,N_862);
nand U6597 (N_6597,N_4251,N_4199);
xor U6598 (N_6598,N_3614,N_1206);
or U6599 (N_6599,N_1768,N_2835);
nand U6600 (N_6600,N_3047,N_3586);
xnor U6601 (N_6601,N_2100,N_3033);
nand U6602 (N_6602,N_222,N_3423);
nor U6603 (N_6603,N_4684,N_954);
xor U6604 (N_6604,N_1367,N_2254);
nor U6605 (N_6605,N_1827,N_3620);
and U6606 (N_6606,N_4067,N_1042);
or U6607 (N_6607,N_4942,N_178);
and U6608 (N_6608,N_2279,N_857);
nand U6609 (N_6609,N_2242,N_2893);
nor U6610 (N_6610,N_1236,N_1817);
and U6611 (N_6611,N_4863,N_4279);
xor U6612 (N_6612,N_1623,N_2009);
nand U6613 (N_6613,N_3925,N_572);
or U6614 (N_6614,N_3258,N_1858);
xor U6615 (N_6615,N_3108,N_3354);
or U6616 (N_6616,N_1678,N_639);
xor U6617 (N_6617,N_2861,N_41);
nand U6618 (N_6618,N_3927,N_4079);
or U6619 (N_6619,N_2075,N_3529);
nand U6620 (N_6620,N_1975,N_1757);
and U6621 (N_6621,N_929,N_2647);
nor U6622 (N_6622,N_762,N_2525);
and U6623 (N_6623,N_1020,N_1579);
nor U6624 (N_6624,N_1862,N_1473);
or U6625 (N_6625,N_2696,N_320);
nand U6626 (N_6626,N_3152,N_3482);
and U6627 (N_6627,N_1491,N_3509);
or U6628 (N_6628,N_3487,N_3637);
xor U6629 (N_6629,N_3880,N_3936);
and U6630 (N_6630,N_4415,N_1646);
and U6631 (N_6631,N_2922,N_3514);
and U6632 (N_6632,N_3046,N_4175);
nand U6633 (N_6633,N_1517,N_458);
and U6634 (N_6634,N_3800,N_4475);
or U6635 (N_6635,N_1655,N_104);
and U6636 (N_6636,N_3519,N_1617);
nand U6637 (N_6637,N_837,N_705);
nor U6638 (N_6638,N_730,N_3848);
nor U6639 (N_6639,N_1594,N_2793);
xor U6640 (N_6640,N_3982,N_3385);
xnor U6641 (N_6641,N_4624,N_4539);
nand U6642 (N_6642,N_2942,N_1788);
nor U6643 (N_6643,N_1645,N_3630);
nor U6644 (N_6644,N_1903,N_2665);
or U6645 (N_6645,N_4103,N_4224);
nor U6646 (N_6646,N_4656,N_4602);
and U6647 (N_6647,N_4131,N_1027);
nand U6648 (N_6648,N_3133,N_1665);
xor U6649 (N_6649,N_1322,N_2711);
xor U6650 (N_6650,N_3995,N_2952);
nand U6651 (N_6651,N_367,N_1577);
nand U6652 (N_6652,N_2313,N_4692);
nand U6653 (N_6653,N_4585,N_667);
or U6654 (N_6654,N_1609,N_4479);
nand U6655 (N_6655,N_1566,N_2868);
or U6656 (N_6656,N_2028,N_4188);
nand U6657 (N_6657,N_936,N_3434);
nand U6658 (N_6658,N_1542,N_4022);
or U6659 (N_6659,N_599,N_4931);
xor U6660 (N_6660,N_3248,N_3934);
and U6661 (N_6661,N_380,N_1262);
xnor U6662 (N_6662,N_2262,N_1456);
or U6663 (N_6663,N_2895,N_3269);
and U6664 (N_6664,N_2485,N_4299);
nand U6665 (N_6665,N_4877,N_2481);
and U6666 (N_6666,N_3076,N_1246);
nor U6667 (N_6667,N_4164,N_1647);
nand U6668 (N_6668,N_3005,N_679);
or U6669 (N_6669,N_970,N_126);
xor U6670 (N_6670,N_3513,N_2695);
xnor U6671 (N_6671,N_3651,N_1033);
and U6672 (N_6672,N_2331,N_4353);
and U6673 (N_6673,N_2940,N_1121);
or U6674 (N_6674,N_4597,N_3954);
nor U6675 (N_6675,N_3081,N_355);
nor U6676 (N_6676,N_835,N_2736);
xor U6677 (N_6677,N_4158,N_789);
nand U6678 (N_6678,N_1842,N_4363);
and U6679 (N_6679,N_1968,N_1370);
or U6680 (N_6680,N_4194,N_1801);
nand U6681 (N_6681,N_1873,N_405);
nand U6682 (N_6682,N_4409,N_228);
and U6683 (N_6683,N_1341,N_1904);
nor U6684 (N_6684,N_2681,N_3100);
nand U6685 (N_6685,N_2872,N_1319);
and U6686 (N_6686,N_497,N_2972);
nor U6687 (N_6687,N_4017,N_4260);
nor U6688 (N_6688,N_902,N_3715);
nand U6689 (N_6689,N_549,N_4132);
or U6690 (N_6690,N_615,N_3151);
or U6691 (N_6691,N_1972,N_3451);
and U6692 (N_6692,N_253,N_4121);
xnor U6693 (N_6693,N_1492,N_3813);
and U6694 (N_6694,N_121,N_1863);
xor U6695 (N_6695,N_2756,N_4080);
or U6696 (N_6696,N_1166,N_1810);
nor U6697 (N_6697,N_2483,N_4834);
nand U6698 (N_6698,N_287,N_4134);
xnor U6699 (N_6699,N_4978,N_1692);
xnor U6700 (N_6700,N_1442,N_2156);
nor U6701 (N_6701,N_1564,N_2826);
xor U6702 (N_6702,N_2605,N_4853);
xnor U6703 (N_6703,N_3906,N_1689);
or U6704 (N_6704,N_2154,N_750);
xor U6705 (N_6705,N_4091,N_2883);
nand U6706 (N_6706,N_382,N_1808);
xnor U6707 (N_6707,N_3202,N_2554);
xnor U6708 (N_6708,N_2018,N_2567);
and U6709 (N_6709,N_3442,N_2160);
xor U6710 (N_6710,N_2197,N_1607);
nand U6711 (N_6711,N_1225,N_2923);
xnor U6712 (N_6712,N_136,N_418);
xor U6713 (N_6713,N_979,N_2183);
xor U6714 (N_6714,N_4428,N_4917);
nor U6715 (N_6715,N_2718,N_4517);
nor U6716 (N_6716,N_2408,N_373);
nand U6717 (N_6717,N_528,N_4493);
or U6718 (N_6718,N_1995,N_14);
xor U6719 (N_6719,N_1861,N_2737);
nand U6720 (N_6720,N_3322,N_3749);
nor U6721 (N_6721,N_493,N_4094);
or U6722 (N_6722,N_4055,N_3929);
and U6723 (N_6723,N_1360,N_788);
or U6724 (N_6724,N_2599,N_3632);
and U6725 (N_6725,N_4376,N_271);
nor U6726 (N_6726,N_4464,N_2031);
xor U6727 (N_6727,N_4125,N_3750);
or U6728 (N_6728,N_2642,N_1065);
xnor U6729 (N_6729,N_1734,N_2252);
and U6730 (N_6730,N_2122,N_1726);
xnor U6731 (N_6731,N_4303,N_2755);
nor U6732 (N_6732,N_2505,N_3283);
nor U6733 (N_6733,N_1211,N_3361);
nand U6734 (N_6734,N_2672,N_292);
nor U6735 (N_6735,N_3200,N_2660);
xor U6736 (N_6736,N_2146,N_3344);
or U6737 (N_6737,N_194,N_2305);
nand U6738 (N_6738,N_648,N_927);
xnor U6739 (N_6739,N_2726,N_1089);
nand U6740 (N_6740,N_2250,N_1419);
nand U6741 (N_6741,N_2438,N_483);
nor U6742 (N_6742,N_1943,N_1803);
xnor U6743 (N_6743,N_1885,N_3205);
and U6744 (N_6744,N_1781,N_4872);
or U6745 (N_6745,N_2887,N_4106);
and U6746 (N_6746,N_4322,N_4584);
or U6747 (N_6747,N_85,N_459);
nor U6748 (N_6748,N_3840,N_2548);
or U6749 (N_6749,N_2913,N_3049);
or U6750 (N_6750,N_420,N_2495);
nor U6751 (N_6751,N_1722,N_2335);
xnor U6752 (N_6752,N_3214,N_332);
xnor U6753 (N_6753,N_1998,N_2909);
or U6754 (N_6754,N_2790,N_4806);
nand U6755 (N_6755,N_3723,N_197);
xnor U6756 (N_6756,N_3638,N_1844);
nor U6757 (N_6757,N_1462,N_2509);
xnor U6758 (N_6758,N_2295,N_1348);
or U6759 (N_6759,N_107,N_612);
nor U6760 (N_6760,N_2613,N_2989);
or U6761 (N_6761,N_4676,N_2363);
nor U6762 (N_6762,N_1860,N_3394);
nor U6763 (N_6763,N_2360,N_4766);
nand U6764 (N_6764,N_2839,N_2874);
or U6765 (N_6765,N_3678,N_2581);
xor U6766 (N_6766,N_1787,N_687);
nand U6767 (N_6767,N_4713,N_1242);
nor U6768 (N_6768,N_2274,N_518);
or U6769 (N_6769,N_4025,N_1736);
and U6770 (N_6770,N_2016,N_2118);
nor U6771 (N_6771,N_1710,N_2584);
and U6772 (N_6772,N_1384,N_2536);
or U6773 (N_6773,N_484,N_871);
and U6774 (N_6774,N_3446,N_2715);
xnor U6775 (N_6775,N_3945,N_1946);
nand U6776 (N_6776,N_624,N_3844);
or U6777 (N_6777,N_4545,N_1928);
nor U6778 (N_6778,N_495,N_3228);
nand U6779 (N_6779,N_2076,N_4477);
nand U6780 (N_6780,N_914,N_1977);
and U6781 (N_6781,N_3601,N_4608);
and U6782 (N_6782,N_2170,N_1908);
and U6783 (N_6783,N_3016,N_1702);
and U6784 (N_6784,N_3057,N_3626);
xnor U6785 (N_6785,N_1534,N_1709);
and U6786 (N_6786,N_2463,N_4976);
nand U6787 (N_6787,N_3696,N_188);
nor U6788 (N_6788,N_1516,N_4117);
or U6789 (N_6789,N_21,N_2964);
xor U6790 (N_6790,N_1559,N_4416);
nor U6791 (N_6791,N_4375,N_550);
and U6792 (N_6792,N_650,N_350);
and U6793 (N_6793,N_4803,N_3543);
nand U6794 (N_6794,N_911,N_3587);
or U6795 (N_6795,N_4014,N_3555);
or U6796 (N_6796,N_1227,N_4953);
or U6797 (N_6797,N_173,N_3856);
nor U6798 (N_6798,N_2366,N_4059);
or U6799 (N_6799,N_2571,N_4557);
nor U6800 (N_6800,N_1656,N_3373);
xor U6801 (N_6801,N_4328,N_2937);
nand U6802 (N_6802,N_2267,N_100);
and U6803 (N_6803,N_1733,N_2517);
xor U6804 (N_6804,N_3790,N_4825);
or U6805 (N_6805,N_1780,N_633);
xor U6806 (N_6806,N_2511,N_2140);
or U6807 (N_6807,N_967,N_2622);
and U6808 (N_6808,N_510,N_3646);
nand U6809 (N_6809,N_1944,N_145);
nor U6810 (N_6810,N_4808,N_2452);
and U6811 (N_6811,N_4141,N_3889);
or U6812 (N_6812,N_4410,N_4997);
and U6813 (N_6813,N_3150,N_1068);
nand U6814 (N_6814,N_1047,N_4474);
and U6815 (N_6815,N_2460,N_3505);
xor U6816 (N_6816,N_1174,N_4385);
and U6817 (N_6817,N_2730,N_526);
nor U6818 (N_6818,N_795,N_1955);
nor U6819 (N_6819,N_3564,N_4230);
nand U6820 (N_6820,N_3281,N_273);
or U6821 (N_6821,N_1669,N_3903);
and U6822 (N_6822,N_645,N_3337);
nor U6823 (N_6823,N_2040,N_125);
nor U6824 (N_6824,N_3943,N_3095);
or U6825 (N_6825,N_1582,N_3187);
nor U6826 (N_6826,N_547,N_4438);
nor U6827 (N_6827,N_3096,N_534);
nor U6828 (N_6828,N_3751,N_423);
and U6829 (N_6829,N_3603,N_1090);
nand U6830 (N_6830,N_1982,N_2152);
and U6831 (N_6831,N_3413,N_2421);
or U6832 (N_6832,N_2428,N_1411);
and U6833 (N_6833,N_3973,N_3364);
nor U6834 (N_6834,N_95,N_2960);
nor U6835 (N_6835,N_616,N_2059);
nand U6836 (N_6836,N_2150,N_2685);
nand U6837 (N_6837,N_3770,N_1340);
and U6838 (N_6838,N_2419,N_1985);
nor U6839 (N_6839,N_1951,N_90);
xor U6840 (N_6840,N_141,N_3156);
or U6841 (N_6841,N_1527,N_4552);
nand U6842 (N_6842,N_3527,N_2088);
xor U6843 (N_6843,N_2365,N_4630);
nor U6844 (N_6844,N_4205,N_1406);
and U6845 (N_6845,N_3481,N_3397);
nand U6846 (N_6846,N_2814,N_2017);
xnor U6847 (N_6847,N_2708,N_2733);
nor U6848 (N_6848,N_817,N_4572);
nor U6849 (N_6849,N_4341,N_2993);
nor U6850 (N_6850,N_4642,N_1662);
xnor U6851 (N_6851,N_4081,N_637);
nor U6852 (N_6852,N_609,N_3928);
nand U6853 (N_6853,N_4660,N_3884);
and U6854 (N_6854,N_1753,N_865);
and U6855 (N_6855,N_2824,N_4352);
xor U6856 (N_6856,N_1672,N_2484);
nand U6857 (N_6857,N_685,N_3371);
and U6858 (N_6858,N_3604,N_3881);
and U6859 (N_6859,N_480,N_1700);
nor U6860 (N_6860,N_3102,N_4037);
and U6861 (N_6861,N_1867,N_1173);
and U6862 (N_6862,N_4370,N_3766);
nand U6863 (N_6863,N_1001,N_1417);
nor U6864 (N_6864,N_2300,N_161);
nand U6865 (N_6865,N_4269,N_3370);
nand U6866 (N_6866,N_431,N_3341);
or U6867 (N_6867,N_4174,N_946);
nor U6868 (N_6868,N_2467,N_2656);
nor U6869 (N_6869,N_3208,N_1811);
xor U6870 (N_6870,N_863,N_2564);
and U6871 (N_6871,N_3252,N_3319);
or U6872 (N_6872,N_2850,N_3783);
and U6873 (N_6873,N_1509,N_654);
and U6874 (N_6874,N_411,N_1260);
xor U6875 (N_6875,N_3841,N_4065);
and U6876 (N_6876,N_849,N_2709);
nor U6877 (N_6877,N_3798,N_1254);
and U6878 (N_6878,N_2289,N_1711);
xnor U6879 (N_6879,N_4936,N_1164);
and U6880 (N_6880,N_3072,N_3401);
nand U6881 (N_6881,N_3217,N_1077);
nand U6882 (N_6882,N_1588,N_486);
and U6883 (N_6883,N_2186,N_2680);
nand U6884 (N_6884,N_34,N_3450);
xor U6885 (N_6885,N_642,N_2165);
xnor U6886 (N_6886,N_2105,N_956);
nand U6887 (N_6887,N_649,N_4273);
xnor U6888 (N_6888,N_4574,N_2391);
and U6889 (N_6889,N_1922,N_855);
or U6890 (N_6890,N_1432,N_2982);
and U6891 (N_6891,N_949,N_1443);
nand U6892 (N_6892,N_123,N_3673);
nor U6893 (N_6893,N_1699,N_1871);
and U6894 (N_6894,N_1421,N_824);
xnor U6895 (N_6895,N_4111,N_1034);
or U6896 (N_6896,N_511,N_4354);
xor U6897 (N_6897,N_1390,N_2310);
nand U6898 (N_6898,N_1524,N_3763);
nand U6899 (N_6899,N_2859,N_3938);
xor U6900 (N_6900,N_1247,N_4776);
xnor U6901 (N_6901,N_4406,N_4882);
nor U6902 (N_6902,N_1935,N_1299);
nor U6903 (N_6903,N_251,N_3358);
nand U6904 (N_6904,N_2278,N_3532);
and U6905 (N_6905,N_1397,N_591);
and U6906 (N_6906,N_337,N_4568);
and U6907 (N_6907,N_1600,N_620);
xnor U6908 (N_6908,N_413,N_4225);
xnor U6909 (N_6909,N_2093,N_1569);
or U6910 (N_6910,N_203,N_4107);
xor U6911 (N_6911,N_3011,N_3683);
nor U6912 (N_6912,N_3530,N_951);
nand U6913 (N_6913,N_252,N_3334);
xor U6914 (N_6914,N_4233,N_2943);
xnor U6915 (N_6915,N_4561,N_3531);
or U6916 (N_6916,N_3745,N_787);
and U6917 (N_6917,N_1259,N_4981);
nand U6918 (N_6918,N_3787,N_3585);
nand U6919 (N_6919,N_2583,N_78);
nor U6920 (N_6920,N_1308,N_2052);
nor U6921 (N_6921,N_3338,N_754);
nand U6922 (N_6922,N_4064,N_1122);
xor U6923 (N_6923,N_3160,N_1306);
and U6924 (N_6924,N_4932,N_851);
nand U6925 (N_6925,N_1292,N_3494);
and U6926 (N_6926,N_4495,N_1032);
nor U6927 (N_6927,N_3357,N_4215);
nor U6928 (N_6928,N_1747,N_464);
nand U6929 (N_6929,N_4030,N_4651);
xor U6930 (N_6930,N_2113,N_1595);
and U6931 (N_6931,N_611,N_671);
nand U6932 (N_6932,N_13,N_3824);
xnor U6933 (N_6933,N_1431,N_4002);
xnor U6934 (N_6934,N_4305,N_2025);
xor U6935 (N_6935,N_1961,N_2102);
nor U6936 (N_6936,N_2114,N_1128);
or U6937 (N_6937,N_2534,N_2752);
xnor U6938 (N_6938,N_4335,N_3204);
nand U6939 (N_6939,N_884,N_4488);
nand U6940 (N_6940,N_1323,N_1352);
and U6941 (N_6941,N_66,N_457);
nand U6942 (N_6942,N_325,N_2356);
and U6943 (N_6943,N_2393,N_470);
nand U6944 (N_6944,N_3631,N_4617);
and U6945 (N_6945,N_3106,N_3556);
and U6946 (N_6946,N_63,N_4695);
and U6947 (N_6947,N_4244,N_3713);
xor U6948 (N_6948,N_4774,N_3120);
nor U6949 (N_6949,N_3188,N_190);
or U6950 (N_6950,N_2167,N_880);
and U6951 (N_6951,N_3184,N_3412);
nor U6952 (N_6952,N_153,N_4297);
nand U6953 (N_6953,N_1284,N_519);
or U6954 (N_6954,N_4512,N_3440);
and U6955 (N_6955,N_4854,N_2890);
xnor U6956 (N_6956,N_3149,N_37);
nor U6957 (N_6957,N_384,N_174);
nor U6958 (N_6958,N_372,N_2794);
xnor U6959 (N_6959,N_3612,N_4983);
xnor U6960 (N_6960,N_2799,N_2455);
xnor U6961 (N_6961,N_3437,N_807);
or U6962 (N_6962,N_1603,N_753);
nor U6963 (N_6963,N_4614,N_1538);
nand U6964 (N_6964,N_4681,N_4841);
and U6965 (N_6965,N_1414,N_1471);
nor U6966 (N_6966,N_2953,N_244);
nand U6967 (N_6967,N_3309,N_539);
nor U6968 (N_6968,N_3365,N_3290);
and U6969 (N_6969,N_2781,N_2914);
xor U6970 (N_6970,N_1567,N_4724);
or U6971 (N_6971,N_867,N_2334);
nand U6972 (N_6972,N_529,N_3444);
and U6973 (N_6973,N_4035,N_4489);
nor U6974 (N_6974,N_189,N_196);
nor U6975 (N_6975,N_536,N_172);
xnor U6976 (N_6976,N_2034,N_4218);
nor U6977 (N_6977,N_4296,N_1427);
xor U6978 (N_6978,N_558,N_4576);
and U6979 (N_6979,N_264,N_4487);
nor U6980 (N_6980,N_1562,N_2703);
xnor U6981 (N_6981,N_2788,N_4579);
and U6982 (N_6982,N_1586,N_86);
and U6983 (N_6983,N_3846,N_1666);
nor U6984 (N_6984,N_2198,N_99);
or U6985 (N_6985,N_1899,N_3407);
or U6986 (N_6986,N_4451,N_2789);
xnor U6987 (N_6987,N_2344,N_3439);
nor U6988 (N_6988,N_215,N_4492);
xnor U6989 (N_6989,N_881,N_2470);
nand U6990 (N_6990,N_3491,N_4639);
xnor U6991 (N_6991,N_2785,N_3681);
and U6992 (N_6992,N_72,N_2945);
nor U6993 (N_6993,N_4446,N_1372);
xor U6994 (N_6994,N_4730,N_4904);
nor U6995 (N_6995,N_2453,N_1186);
or U6996 (N_6996,N_2216,N_4453);
xor U6997 (N_6997,N_2223,N_4569);
nand U6998 (N_6998,N_143,N_3533);
nand U6999 (N_6999,N_47,N_3031);
nand U7000 (N_7000,N_3785,N_2359);
or U7001 (N_7001,N_3908,N_465);
xor U7002 (N_7002,N_724,N_4460);
and U7003 (N_7003,N_4393,N_1950);
nand U7004 (N_7004,N_890,N_3591);
or U7005 (N_7005,N_2208,N_1797);
nand U7006 (N_7006,N_2263,N_4242);
nor U7007 (N_7007,N_1381,N_2563);
nand U7008 (N_7008,N_2238,N_3286);
xnor U7009 (N_7009,N_2043,N_1556);
or U7010 (N_7010,N_872,N_658);
xnor U7011 (N_7011,N_165,N_3203);
xor U7012 (N_7012,N_2241,N_3071);
nor U7013 (N_7013,N_2116,N_4542);
and U7014 (N_7014,N_498,N_2288);
nor U7015 (N_7015,N_2343,N_1394);
xnor U7016 (N_7016,N_2746,N_4619);
nand U7017 (N_7017,N_2066,N_351);
nor U7018 (N_7018,N_3162,N_2630);
nand U7019 (N_7019,N_1143,N_4823);
nand U7020 (N_7020,N_552,N_4961);
nor U7021 (N_7021,N_3902,N_1924);
xnor U7022 (N_7022,N_3584,N_903);
or U7023 (N_7023,N_1629,N_986);
nand U7024 (N_7024,N_1165,N_2627);
or U7025 (N_7025,N_2928,N_1267);
nor U7026 (N_7026,N_2682,N_2767);
or U7027 (N_7027,N_2351,N_3302);
or U7028 (N_7028,N_3895,N_2765);
nor U7029 (N_7029,N_2851,N_2888);
nor U7030 (N_7030,N_743,N_618);
and U7031 (N_7031,N_4308,N_820);
and U7032 (N_7032,N_231,N_1383);
xnor U7033 (N_7033,N_3299,N_2417);
and U7034 (N_7034,N_432,N_2053);
nor U7035 (N_7035,N_1204,N_1329);
or U7036 (N_7036,N_2439,N_1932);
nand U7037 (N_7037,N_4181,N_1793);
nor U7038 (N_7038,N_4972,N_3756);
nand U7039 (N_7039,N_4769,N_4316);
or U7040 (N_7040,N_3234,N_4600);
nor U7041 (N_7041,N_1636,N_1494);
xnor U7042 (N_7042,N_3155,N_3125);
and U7043 (N_7043,N_4434,N_4968);
nor U7044 (N_7044,N_1423,N_822);
and U7045 (N_7045,N_2329,N_1879);
and U7046 (N_7046,N_716,N_864);
and U7047 (N_7047,N_3679,N_2330);
and U7048 (N_7048,N_3235,N_3455);
xnor U7049 (N_7049,N_1300,N_343);
nand U7050 (N_7050,N_4718,N_756);
or U7051 (N_7051,N_453,N_4826);
nand U7052 (N_7052,N_4440,N_3325);
or U7053 (N_7053,N_4095,N_1248);
and U7054 (N_7054,N_1680,N_4538);
or U7055 (N_7055,N_1898,N_1064);
xor U7056 (N_7056,N_939,N_1814);
or U7057 (N_7057,N_1712,N_3010);
xor U7058 (N_7058,N_1158,N_4120);
and U7059 (N_7059,N_2490,N_3227);
and U7060 (N_7060,N_656,N_838);
nor U7061 (N_7061,N_1183,N_152);
nor U7062 (N_7062,N_3328,N_3682);
xnor U7063 (N_7063,N_1435,N_950);
nor U7064 (N_7064,N_2777,N_4532);
or U7065 (N_7065,N_1103,N_2586);
nand U7066 (N_7066,N_3034,N_4772);
or U7067 (N_7067,N_814,N_261);
and U7068 (N_7068,N_1703,N_2308);
and U7069 (N_7069,N_478,N_2272);
nor U7070 (N_7070,N_463,N_4187);
nor U7071 (N_7071,N_1624,N_2051);
and U7072 (N_7072,N_4673,N_3416);
nand U7073 (N_7073,N_4499,N_783);
and U7074 (N_7074,N_4891,N_399);
nand U7075 (N_7075,N_2557,N_3876);
or U7076 (N_7076,N_3036,N_4049);
or U7077 (N_7077,N_1859,N_4382);
nor U7078 (N_7078,N_1547,N_1337);
or U7079 (N_7079,N_4938,N_3961);
xor U7080 (N_7080,N_2106,N_4693);
nor U7081 (N_7081,N_4720,N_3489);
nand U7082 (N_7082,N_213,N_160);
nor U7083 (N_7083,N_426,N_324);
nor U7084 (N_7084,N_3131,N_573);
and U7085 (N_7085,N_3295,N_1812);
nor U7086 (N_7086,N_4831,N_3752);
xor U7087 (N_7087,N_1463,N_2771);
nor U7088 (N_7088,N_3452,N_2847);
nor U7089 (N_7089,N_2204,N_868);
nor U7090 (N_7090,N_1177,N_2944);
nor U7091 (N_7091,N_341,N_977);
xnor U7092 (N_7092,N_2064,N_533);
or U7093 (N_7093,N_31,N_4333);
nand U7094 (N_7094,N_2091,N_3201);
and U7095 (N_7095,N_1163,N_1265);
nor U7096 (N_7096,N_897,N_2635);
nor U7097 (N_7097,N_1743,N_596);
nor U7098 (N_7098,N_4293,N_4204);
nor U7099 (N_7099,N_3134,N_2182);
or U7100 (N_7100,N_1641,N_1939);
nand U7101 (N_7101,N_2516,N_640);
and U7102 (N_7102,N_4712,N_3937);
or U7103 (N_7103,N_4031,N_570);
nand U7104 (N_7104,N_3979,N_3303);
and U7105 (N_7105,N_4201,N_603);
nor U7106 (N_7106,N_3845,N_4077);
xor U7107 (N_7107,N_791,N_3045);
or U7108 (N_7108,N_2104,N_2700);
nor U7109 (N_7109,N_1263,N_46);
xor U7110 (N_7110,N_2492,N_2598);
nor U7111 (N_7111,N_1145,N_4157);
nor U7112 (N_7112,N_1834,N_1653);
and U7113 (N_7113,N_3350,N_4090);
or U7114 (N_7114,N_1096,N_800);
or U7115 (N_7115,N_2900,N_2619);
nor U7116 (N_7116,N_4104,N_144);
nor U7117 (N_7117,N_3247,N_1215);
nand U7118 (N_7118,N_1006,N_2326);
nor U7119 (N_7119,N_4007,N_2537);
and U7120 (N_7120,N_2162,N_1604);
and U7121 (N_7121,N_810,N_3396);
xnor U7122 (N_7122,N_33,N_1106);
nor U7123 (N_7123,N_2830,N_1116);
and U7124 (N_7124,N_3639,N_943);
or U7125 (N_7125,N_209,N_1452);
and U7126 (N_7126,N_4391,N_219);
nand U7127 (N_7127,N_4667,N_1315);
nor U7128 (N_7128,N_4362,N_1728);
nand U7129 (N_7129,N_415,N_3885);
nor U7130 (N_7130,N_4535,N_1018);
nand U7131 (N_7131,N_1717,N_3389);
nand U7132 (N_7132,N_1048,N_4694);
and U7133 (N_7133,N_4414,N_2600);
xor U7134 (N_7134,N_1913,N_3598);
xor U7135 (N_7135,N_4321,N_1386);
nor U7136 (N_7136,N_4824,N_4466);
nand U7137 (N_7137,N_1886,N_1207);
and U7138 (N_7138,N_3191,N_1095);
xnor U7139 (N_7139,N_991,N_4190);
nor U7140 (N_7140,N_2821,N_725);
nor U7141 (N_7141,N_4066,N_3262);
xor U7142 (N_7142,N_3042,N_1086);
xor U7143 (N_7143,N_3013,N_2478);
or U7144 (N_7144,N_1290,N_1500);
xor U7145 (N_7145,N_3193,N_3808);
and U7146 (N_7146,N_2817,N_2192);
and U7147 (N_7147,N_1102,N_1529);
xor U7148 (N_7148,N_2449,N_1280);
or U7149 (N_7149,N_4977,N_4690);
nand U7150 (N_7150,N_4355,N_352);
or U7151 (N_7151,N_614,N_1882);
and U7152 (N_7152,N_3068,N_3157);
or U7153 (N_7153,N_1720,N_2022);
or U7154 (N_7154,N_1212,N_850);
xor U7155 (N_7155,N_387,N_322);
nor U7156 (N_7156,N_4502,N_2577);
or U7157 (N_7157,N_600,N_3459);
nor U7158 (N_7158,N_3007,N_443);
nand U7159 (N_7159,N_4208,N_2239);
xnor U7160 (N_7160,N_3972,N_1275);
and U7161 (N_7161,N_4933,N_1648);
xnor U7162 (N_7162,N_1208,N_1784);
and U7163 (N_7163,N_2611,N_910);
nand U7164 (N_7164,N_769,N_1453);
nor U7165 (N_7165,N_4209,N_2593);
xor U7166 (N_7166,N_2729,N_3724);
xnor U7167 (N_7167,N_3263,N_1244);
or U7168 (N_7168,N_3966,N_4979);
or U7169 (N_7169,N_1830,N_3722);
or U7170 (N_7170,N_2171,N_75);
nor U7171 (N_7171,N_4456,N_3932);
nor U7172 (N_7172,N_134,N_2005);
or U7173 (N_7173,N_3456,N_3955);
nand U7174 (N_7174,N_2560,N_4699);
or U7175 (N_7175,N_551,N_302);
nand U7176 (N_7176,N_792,N_3685);
or U7177 (N_7177,N_4742,N_2328);
nand U7178 (N_7178,N_2813,N_1428);
xor U7179 (N_7179,N_4985,N_1761);
nor U7180 (N_7180,N_629,N_3090);
nand U7181 (N_7181,N_3431,N_1214);
and U7182 (N_7182,N_4070,N_4649);
nand U7183 (N_7183,N_2450,N_191);
xor U7184 (N_7184,N_2643,N_2748);
nand U7185 (N_7185,N_2702,N_965);
and U7186 (N_7186,N_676,N_4433);
and U7187 (N_7187,N_1670,N_684);
nor U7188 (N_7188,N_4231,N_3145);
and U7189 (N_7189,N_3602,N_842);
nor U7190 (N_7190,N_175,N_4918);
nor U7191 (N_7191,N_4960,N_3714);
xor U7192 (N_7192,N_736,N_1171);
nand U7193 (N_7193,N_916,N_4348);
or U7194 (N_7194,N_2935,N_1777);
nor U7195 (N_7195,N_2332,N_3225);
xnor U7196 (N_7196,N_2068,N_3933);
nand U7197 (N_7197,N_266,N_4255);
nor U7198 (N_7198,N_2251,N_926);
or U7199 (N_7199,N_3700,N_2920);
and U7200 (N_7200,N_3035,N_804);
nand U7201 (N_7201,N_447,N_4687);
or U7202 (N_7202,N_772,N_4315);
nand U7203 (N_7203,N_1454,N_2462);
nor U7204 (N_7204,N_621,N_137);
xor U7205 (N_7205,N_3981,N_688);
and U7206 (N_7206,N_3369,N_4680);
nand U7207 (N_7207,N_1216,N_2448);
nor U7208 (N_7208,N_4292,N_2625);
nor U7209 (N_7209,N_1358,N_168);
or U7210 (N_7210,N_4180,N_2568);
nor U7211 (N_7211,N_2725,N_531);
or U7212 (N_7212,N_813,N_1088);
nand U7213 (N_7213,N_678,N_1304);
nand U7214 (N_7214,N_1410,N_1205);
and U7215 (N_7215,N_3,N_2691);
nor U7216 (N_7216,N_4170,N_3366);
nor U7217 (N_7217,N_3360,N_4011);
nand U7218 (N_7218,N_1357,N_567);
and U7219 (N_7219,N_3094,N_692);
and U7220 (N_7220,N_3318,N_3993);
nor U7221 (N_7221,N_3265,N_2273);
nand U7222 (N_7222,N_3128,N_3767);
or U7223 (N_7223,N_694,N_4145);
and U7224 (N_7224,N_2074,N_784);
and U7225 (N_7225,N_4310,N_1779);
or U7226 (N_7226,N_3692,N_4227);
nand U7227 (N_7227,N_3553,N_2322);
or U7228 (N_7228,N_3568,N_4925);
and U7229 (N_7229,N_1359,N_4288);
nand U7230 (N_7230,N_4809,N_4261);
xor U7231 (N_7231,N_3522,N_2545);
nor U7232 (N_7232,N_625,N_2177);
nor U7233 (N_7233,N_3165,N_3372);
nand U7234 (N_7234,N_3608,N_2640);
xor U7235 (N_7235,N_1222,N_4018);
and U7236 (N_7236,N_1339,N_4443);
or U7237 (N_7237,N_1039,N_3781);
nand U7238 (N_7238,N_2524,N_1451);
and U7239 (N_7239,N_4408,N_488);
nand U7240 (N_7240,N_4970,N_4595);
nand U7241 (N_7241,N_1483,N_2000);
nand U7242 (N_7242,N_2191,N_2873);
or U7243 (N_7243,N_1153,N_4137);
nor U7244 (N_7244,N_3817,N_1354);
nand U7245 (N_7245,N_4537,N_1563);
nor U7246 (N_7246,N_3020,N_4993);
nor U7247 (N_7247,N_1999,N_2973);
xnor U7248 (N_7248,N_400,N_3458);
nor U7249 (N_7249,N_3891,N_454);
and U7250 (N_7250,N_2095,N_4289);
or U7251 (N_7251,N_4214,N_247);
and U7252 (N_7252,N_3127,N_2416);
xnor U7253 (N_7253,N_1134,N_4745);
nor U7254 (N_7254,N_3860,N_4048);
or U7255 (N_7255,N_4425,N_2742);
and U7256 (N_7256,N_2013,N_3743);
or U7257 (N_7257,N_2529,N_4883);
xor U7258 (N_7258,N_4358,N_894);
or U7259 (N_7259,N_737,N_2048);
xnor U7260 (N_7260,N_3636,N_364);
nand U7261 (N_7261,N_3192,N_1155);
and U7262 (N_7262,N_1551,N_1661);
and U7263 (N_7263,N_2404,N_3565);
nand U7264 (N_7264,N_4127,N_3392);
nor U7265 (N_7265,N_4368,N_1420);
and U7266 (N_7266,N_2039,N_1688);
xnor U7267 (N_7267,N_907,N_4832);
and U7268 (N_7268,N_2804,N_4784);
xnor U7269 (N_7269,N_4725,N_3219);
nand U7270 (N_7270,N_4610,N_2321);
or U7271 (N_7271,N_588,N_3905);
xnor U7272 (N_7272,N_4457,N_4183);
xor U7273 (N_7273,N_2980,N_4267);
or U7274 (N_7274,N_3089,N_2797);
xnor U7275 (N_7275,N_4912,N_4334);
or U7276 (N_7276,N_1447,N_3051);
or U7277 (N_7277,N_1866,N_1464);
xnor U7278 (N_7278,N_492,N_3589);
nor U7279 (N_7279,N_4616,N_942);
and U7280 (N_7280,N_2174,N_1057);
nor U7281 (N_7281,N_25,N_4084);
or U7282 (N_7282,N_2161,N_1807);
and U7283 (N_7283,N_2473,N_797);
nand U7284 (N_7284,N_2958,N_583);
nor U7285 (N_7285,N_1770,N_11);
nand U7286 (N_7286,N_3913,N_407);
nor U7287 (N_7287,N_3022,N_1446);
nor U7288 (N_7288,N_2143,N_4325);
nand U7289 (N_7289,N_4827,N_2866);
nor U7290 (N_7290,N_952,N_278);
nand U7291 (N_7291,N_1000,N_2354);
xnor U7292 (N_7292,N_2664,N_2233);
xor U7293 (N_7293,N_796,N_4407);
or U7294 (N_7294,N_4794,N_515);
or U7295 (N_7295,N_4908,N_3065);
and U7296 (N_7296,N_1848,N_2624);
nor U7297 (N_7297,N_4427,N_912);
nand U7298 (N_7298,N_2213,N_2901);
xor U7299 (N_7299,N_115,N_1161);
or U7300 (N_7300,N_3963,N_4074);
nand U7301 (N_7301,N_3526,N_2123);
and U7302 (N_7302,N_1223,N_3070);
or U7303 (N_7303,N_873,N_4800);
nor U7304 (N_7304,N_3559,N_3141);
nand U7305 (N_7305,N_2498,N_2381);
and U7306 (N_7306,N_2907,N_3610);
nand U7307 (N_7307,N_4911,N_3146);
xnor U7308 (N_7308,N_997,N_2256);
or U7309 (N_7309,N_1195,N_2592);
and U7310 (N_7310,N_4637,N_1806);
and U7311 (N_7311,N_2576,N_3582);
or U7312 (N_7312,N_4019,N_1705);
or U7313 (N_7313,N_899,N_3277);
nand U7314 (N_7314,N_1349,N_4195);
nand U7315 (N_7315,N_2375,N_542);
xor U7316 (N_7316,N_4811,N_461);
nand U7317 (N_7317,N_1192,N_3888);
or U7318 (N_7318,N_586,N_2650);
nor U7319 (N_7319,N_4618,N_4402);
nor U7320 (N_7320,N_3109,N_3183);
nor U7321 (N_7321,N_2897,N_2464);
nor U7322 (N_7322,N_780,N_4923);
or U7323 (N_7323,N_1277,N_4020);
or U7324 (N_7324,N_1221,N_702);
and U7325 (N_7325,N_538,N_2668);
xor U7326 (N_7326,N_102,N_4902);
xnor U7327 (N_7327,N_4661,N_2201);
nand U7328 (N_7328,N_1772,N_2905);
nor U7329 (N_7329,N_2787,N_3488);
xnor U7330 (N_7330,N_51,N_2782);
or U7331 (N_7331,N_1612,N_1773);
nand U7332 (N_7332,N_2997,N_1738);
and U7333 (N_7333,N_4603,N_1407);
and U7334 (N_7334,N_3893,N_4142);
nor U7335 (N_7335,N_246,N_2202);
and U7336 (N_7336,N_3323,N_2371);
nand U7337 (N_7337,N_2988,N_3327);
or U7338 (N_7338,N_4027,N_1893);
and U7339 (N_7339,N_3342,N_4034);
xnor U7340 (N_7340,N_1822,N_4152);
and U7341 (N_7341,N_1050,N_4426);
xnor U7342 (N_7342,N_2757,N_556);
nand U7343 (N_7343,N_398,N_205);
xnor U7344 (N_7344,N_204,N_561);
nand U7345 (N_7345,N_3091,N_3640);
nand U7346 (N_7346,N_132,N_770);
xnor U7347 (N_7347,N_1325,N_1445);
and U7348 (N_7348,N_2293,N_4338);
and U7349 (N_7349,N_3471,N_4570);
or U7350 (N_7350,N_3029,N_4369);
xnor U7351 (N_7351,N_2135,N_439);
or U7352 (N_7352,N_4365,N_2296);
nand U7353 (N_7353,N_1798,N_3289);
or U7354 (N_7354,N_4549,N_2926);
nor U7355 (N_7355,N_2633,N_3747);
nand U7356 (N_7356,N_3216,N_4332);
nor U7357 (N_7357,N_193,N_3378);
or U7358 (N_7358,N_333,N_1654);
and U7359 (N_7359,N_279,N_4366);
nor U7360 (N_7360,N_4192,N_4087);
and U7361 (N_7361,N_3186,N_2716);
or U7362 (N_7362,N_250,N_2032);
nor U7363 (N_7363,N_1270,N_225);
and U7364 (N_7364,N_1172,N_272);
xnor U7365 (N_7365,N_1878,N_2475);
or U7366 (N_7366,N_1553,N_2399);
and U7367 (N_7367,N_3436,N_4975);
xor U7368 (N_7368,N_2384,N_4897);
nand U7369 (N_7369,N_4773,N_801);
or U7370 (N_7370,N_4662,N_4378);
or U7371 (N_7371,N_4675,N_655);
nand U7372 (N_7372,N_3539,N_4937);
xor U7373 (N_7373,N_2585,N_4604);
nor U7374 (N_7374,N_738,N_2001);
nand U7375 (N_7375,N_1572,N_3899);
nand U7376 (N_7376,N_4710,N_2595);
xnor U7377 (N_7377,N_1804,N_2136);
and U7378 (N_7378,N_4422,N_101);
nor U7379 (N_7379,N_1679,N_92);
nand U7380 (N_7380,N_3550,N_1331);
nand U7381 (N_7381,N_3499,N_229);
nor U7382 (N_7382,N_4436,N_1851);
and U7383 (N_7383,N_4520,N_1059);
nand U7384 (N_7384,N_1484,N_1829);
or U7385 (N_7385,N_2103,N_3021);
nor U7386 (N_7386,N_1092,N_3719);
or U7387 (N_7387,N_1286,N_2526);
or U7388 (N_7388,N_1251,N_1635);
xor U7389 (N_7389,N_840,N_448);
nor U7390 (N_7390,N_619,N_3703);
xnor U7391 (N_7391,N_719,N_4994);
or U7392 (N_7392,N_2275,N_4307);
and U7393 (N_7393,N_3159,N_3271);
and U7394 (N_7394,N_1313,N_3977);
nand U7395 (N_7395,N_1971,N_315);
or U7396 (N_7396,N_3877,N_2927);
and U7397 (N_7397,N_4212,N_1649);
nand U7398 (N_7398,N_3861,N_4236);
and U7399 (N_7399,N_2390,N_2801);
or U7400 (N_7400,N_3985,N_1294);
nand U7401 (N_7401,N_2745,N_1353);
nor U7402 (N_7402,N_3419,N_4954);
or U7403 (N_7403,N_1558,N_1870);
xor U7404 (N_7404,N_1606,N_4109);
nand U7405 (N_7405,N_4295,N_4821);
nand U7406 (N_7406,N_3427,N_2437);
nor U7407 (N_7407,N_433,N_2465);
nand U7408 (N_7408,N_4957,N_3226);
xnor U7409 (N_7409,N_3037,N_4038);
or U7410 (N_7410,N_606,N_1413);
or U7411 (N_7411,N_3689,N_4023);
or U7412 (N_7412,N_473,N_4544);
and U7413 (N_7413,N_3500,N_2397);
xor U7414 (N_7414,N_3524,N_744);
or U7415 (N_7415,N_3306,N_869);
or U7416 (N_7416,N_1608,N_1925);
nand U7417 (N_7417,N_164,N_3449);
and U7418 (N_7418,N_1744,N_2947);
xnor U7419 (N_7419,N_1014,N_2555);
nand U7420 (N_7420,N_1298,N_4551);
xnor U7421 (N_7421,N_1528,N_58);
xnor U7422 (N_7422,N_2669,N_2677);
nand U7423 (N_7423,N_4945,N_581);
xor U7424 (N_7424,N_2187,N_703);
and U7425 (N_7425,N_2967,N_1748);
or U7426 (N_7426,N_406,N_2445);
or U7427 (N_7427,N_1389,N_3097);
nor U7428 (N_7428,N_4243,N_4515);
or U7429 (N_7429,N_1507,N_4472);
and U7430 (N_7430,N_3634,N_3858);
nor U7431 (N_7431,N_313,N_594);
and U7432 (N_7432,N_1234,N_4629);
and U7433 (N_7433,N_4041,N_105);
nor U7434 (N_7434,N_207,N_3447);
and U7435 (N_7435,N_4344,N_3023);
xor U7436 (N_7436,N_1469,N_3496);
nor U7437 (N_7437,N_3711,N_3257);
nand U7438 (N_7438,N_2067,N_2055);
and U7439 (N_7439,N_2712,N_1179);
xor U7440 (N_7440,N_3643,N_4747);
xnor U7441 (N_7441,N_2269,N_1385);
nor U7442 (N_7442,N_2230,N_2832);
or U7443 (N_7443,N_377,N_1252);
and U7444 (N_7444,N_3583,N_4820);
nand U7445 (N_7445,N_4513,N_3474);
xnor U7446 (N_7446,N_4951,N_4129);
and U7447 (N_7447,N_4903,N_1668);
and U7448 (N_7448,N_1832,N_2266);
or U7449 (N_7449,N_1824,N_3332);
xnor U7450 (N_7450,N_1663,N_2803);
or U7451 (N_7451,N_1330,N_146);
nand U7452 (N_7452,N_695,N_3551);
xnor U7453 (N_7453,N_1311,N_2931);
nor U7454 (N_7454,N_2949,N_4033);
or U7455 (N_7455,N_2141,N_1332);
or U7456 (N_7456,N_2579,N_2697);
nand U7457 (N_7457,N_4377,N_4507);
nand U7458 (N_7458,N_3951,N_2802);
xnor U7459 (N_7459,N_1291,N_1071);
nor U7460 (N_7460,N_1458,N_1897);
and U7461 (N_7461,N_660,N_3140);
xor U7462 (N_7462,N_4646,N_1278);
xnor U7463 (N_7463,N_3776,N_42);
nor U7464 (N_7464,N_3633,N_1938);
nand U7465 (N_7465,N_294,N_1785);
xnor U7466 (N_7466,N_2138,N_4944);
or U7467 (N_7467,N_3655,N_1487);
nor U7468 (N_7468,N_1426,N_1826);
nor U7469 (N_7469,N_3024,N_327);
nand U7470 (N_7470,N_1625,N_2249);
and U7471 (N_7471,N_3916,N_4400);
nand U7472 (N_7472,N_3741,N_424);
nor U7473 (N_7473,N_440,N_4482);
nor U7474 (N_7474,N_3852,N_3393);
and U7475 (N_7475,N_4879,N_472);
or U7476 (N_7476,N_4871,N_4833);
nor U7477 (N_7477,N_3276,N_1287);
nand U7478 (N_7478,N_919,N_4514);
nand U7479 (N_7479,N_3948,N_2869);
nand U7480 (N_7480,N_2441,N_1073);
nand U7481 (N_7481,N_4995,N_1958);
or U7482 (N_7482,N_4812,N_735);
and U7483 (N_7483,N_3708,N_4110);
nand U7484 (N_7484,N_1142,N_3014);
xnor U7485 (N_7485,N_2024,N_3362);
nor U7486 (N_7486,N_1467,N_388);
xor U7487 (N_7487,N_617,N_3538);
or U7488 (N_7488,N_1513,N_1024);
or U7489 (N_7489,N_2827,N_3777);
and U7490 (N_7490,N_119,N_4073);
or U7491 (N_7491,N_2012,N_4016);
xor U7492 (N_7492,N_2320,N_644);
xnor U7493 (N_7493,N_4312,N_1618);
nand U7494 (N_7494,N_2228,N_2145);
or U7495 (N_7495,N_834,N_953);
nor U7496 (N_7496,N_1813,N_1219);
nand U7497 (N_7497,N_2128,N_2281);
nand U7498 (N_7498,N_933,N_2800);
xnor U7499 (N_7499,N_3859,N_2257);
or U7500 (N_7500,N_718,N_2790);
or U7501 (N_7501,N_1750,N_416);
nor U7502 (N_7502,N_1654,N_4441);
nor U7503 (N_7503,N_3069,N_3551);
nor U7504 (N_7504,N_4595,N_2522);
and U7505 (N_7505,N_4241,N_2918);
or U7506 (N_7506,N_404,N_200);
and U7507 (N_7507,N_1150,N_4063);
xor U7508 (N_7508,N_1164,N_4144);
and U7509 (N_7509,N_3547,N_2157);
xnor U7510 (N_7510,N_534,N_1465);
xor U7511 (N_7511,N_4874,N_712);
xor U7512 (N_7512,N_1091,N_806);
nor U7513 (N_7513,N_2062,N_2632);
nand U7514 (N_7514,N_1322,N_2031);
nand U7515 (N_7515,N_3352,N_3058);
nor U7516 (N_7516,N_425,N_2413);
or U7517 (N_7517,N_4226,N_1689);
nor U7518 (N_7518,N_2470,N_3829);
nand U7519 (N_7519,N_3229,N_1243);
xnor U7520 (N_7520,N_889,N_1777);
nand U7521 (N_7521,N_2781,N_1280);
nand U7522 (N_7522,N_4166,N_2385);
or U7523 (N_7523,N_4012,N_466);
nand U7524 (N_7524,N_1372,N_827);
and U7525 (N_7525,N_1900,N_4253);
xor U7526 (N_7526,N_1214,N_2443);
xor U7527 (N_7527,N_1560,N_4437);
and U7528 (N_7528,N_3024,N_1902);
or U7529 (N_7529,N_2912,N_390);
and U7530 (N_7530,N_2718,N_1046);
nor U7531 (N_7531,N_2258,N_2329);
or U7532 (N_7532,N_2005,N_766);
nor U7533 (N_7533,N_2437,N_4343);
nor U7534 (N_7534,N_399,N_564);
nor U7535 (N_7535,N_2744,N_0);
nand U7536 (N_7536,N_3660,N_3452);
nand U7537 (N_7537,N_372,N_3860);
nand U7538 (N_7538,N_3539,N_826);
nand U7539 (N_7539,N_4797,N_1089);
and U7540 (N_7540,N_3001,N_492);
nand U7541 (N_7541,N_2764,N_380);
and U7542 (N_7542,N_2616,N_610);
xor U7543 (N_7543,N_3601,N_4615);
or U7544 (N_7544,N_2070,N_4402);
nand U7545 (N_7545,N_4306,N_3150);
xor U7546 (N_7546,N_3490,N_3071);
nor U7547 (N_7547,N_2680,N_321);
xnor U7548 (N_7548,N_580,N_3198);
xnor U7549 (N_7549,N_3397,N_2464);
and U7550 (N_7550,N_1779,N_3822);
and U7551 (N_7551,N_3745,N_631);
and U7552 (N_7552,N_3023,N_2625);
xnor U7553 (N_7553,N_3576,N_2912);
xnor U7554 (N_7554,N_4149,N_3077);
nor U7555 (N_7555,N_955,N_3360);
or U7556 (N_7556,N_434,N_1690);
or U7557 (N_7557,N_4161,N_4365);
xnor U7558 (N_7558,N_385,N_3649);
xor U7559 (N_7559,N_1651,N_1293);
xor U7560 (N_7560,N_1584,N_4397);
nor U7561 (N_7561,N_2665,N_4743);
nand U7562 (N_7562,N_2329,N_3263);
xnor U7563 (N_7563,N_3120,N_1525);
nand U7564 (N_7564,N_2952,N_4655);
xor U7565 (N_7565,N_4154,N_768);
nand U7566 (N_7566,N_2978,N_3216);
or U7567 (N_7567,N_2707,N_4998);
nand U7568 (N_7568,N_233,N_3);
nand U7569 (N_7569,N_3225,N_4215);
nand U7570 (N_7570,N_4704,N_4940);
nand U7571 (N_7571,N_2497,N_99);
nand U7572 (N_7572,N_1017,N_3886);
nand U7573 (N_7573,N_277,N_1403);
or U7574 (N_7574,N_2134,N_2599);
nand U7575 (N_7575,N_587,N_1373);
and U7576 (N_7576,N_4298,N_3183);
and U7577 (N_7577,N_3376,N_4472);
or U7578 (N_7578,N_1176,N_3713);
or U7579 (N_7579,N_302,N_4774);
nand U7580 (N_7580,N_4533,N_170);
nand U7581 (N_7581,N_3249,N_2141);
nand U7582 (N_7582,N_2994,N_4592);
xor U7583 (N_7583,N_307,N_726);
nand U7584 (N_7584,N_3795,N_1533);
nor U7585 (N_7585,N_129,N_629);
nand U7586 (N_7586,N_2210,N_1785);
and U7587 (N_7587,N_4156,N_1648);
or U7588 (N_7588,N_690,N_4387);
nor U7589 (N_7589,N_4889,N_4396);
or U7590 (N_7590,N_447,N_39);
or U7591 (N_7591,N_4801,N_2125);
xor U7592 (N_7592,N_2308,N_4286);
nor U7593 (N_7593,N_13,N_995);
and U7594 (N_7594,N_1722,N_950);
or U7595 (N_7595,N_2468,N_3330);
and U7596 (N_7596,N_2789,N_4078);
nand U7597 (N_7597,N_1160,N_1890);
or U7598 (N_7598,N_1305,N_3359);
or U7599 (N_7599,N_2644,N_4402);
xnor U7600 (N_7600,N_4761,N_4095);
nand U7601 (N_7601,N_4081,N_1259);
nor U7602 (N_7602,N_4469,N_1884);
nor U7603 (N_7603,N_1251,N_775);
nand U7604 (N_7604,N_2104,N_2353);
xor U7605 (N_7605,N_3341,N_461);
or U7606 (N_7606,N_877,N_4961);
nor U7607 (N_7607,N_2750,N_868);
nor U7608 (N_7608,N_2937,N_550);
xor U7609 (N_7609,N_1670,N_2827);
and U7610 (N_7610,N_1999,N_1808);
nor U7611 (N_7611,N_2835,N_2159);
nor U7612 (N_7612,N_1250,N_4759);
or U7613 (N_7613,N_1510,N_1350);
xnor U7614 (N_7614,N_3574,N_2552);
nand U7615 (N_7615,N_2548,N_3122);
and U7616 (N_7616,N_4200,N_667);
or U7617 (N_7617,N_138,N_4207);
nor U7618 (N_7618,N_3013,N_3467);
nor U7619 (N_7619,N_1494,N_2055);
nand U7620 (N_7620,N_2769,N_4898);
or U7621 (N_7621,N_2408,N_1487);
or U7622 (N_7622,N_2966,N_4430);
nor U7623 (N_7623,N_932,N_4350);
or U7624 (N_7624,N_4837,N_4295);
nor U7625 (N_7625,N_3179,N_1008);
or U7626 (N_7626,N_2453,N_1492);
nor U7627 (N_7627,N_3748,N_1580);
nor U7628 (N_7628,N_3865,N_3875);
and U7629 (N_7629,N_2156,N_4861);
or U7630 (N_7630,N_183,N_459);
nand U7631 (N_7631,N_3242,N_4307);
or U7632 (N_7632,N_1741,N_291);
nor U7633 (N_7633,N_1089,N_555);
or U7634 (N_7634,N_4454,N_3617);
xnor U7635 (N_7635,N_3878,N_4083);
nor U7636 (N_7636,N_3091,N_4260);
nand U7637 (N_7637,N_3381,N_4844);
nor U7638 (N_7638,N_2019,N_1977);
nand U7639 (N_7639,N_1956,N_4341);
and U7640 (N_7640,N_1248,N_3063);
or U7641 (N_7641,N_337,N_1236);
nor U7642 (N_7642,N_1679,N_870);
or U7643 (N_7643,N_1913,N_3017);
and U7644 (N_7644,N_2528,N_3015);
and U7645 (N_7645,N_4736,N_1394);
or U7646 (N_7646,N_3162,N_1598);
xnor U7647 (N_7647,N_4540,N_1789);
xnor U7648 (N_7648,N_369,N_2902);
xnor U7649 (N_7649,N_3704,N_1438);
nand U7650 (N_7650,N_589,N_2299);
xnor U7651 (N_7651,N_257,N_3650);
or U7652 (N_7652,N_2155,N_709);
nor U7653 (N_7653,N_3392,N_727);
nor U7654 (N_7654,N_4596,N_3217);
and U7655 (N_7655,N_4045,N_2141);
xnor U7656 (N_7656,N_3917,N_486);
xor U7657 (N_7657,N_3272,N_812);
nand U7658 (N_7658,N_749,N_4125);
xnor U7659 (N_7659,N_1639,N_1933);
nand U7660 (N_7660,N_4390,N_4102);
nand U7661 (N_7661,N_403,N_2944);
xnor U7662 (N_7662,N_4203,N_632);
and U7663 (N_7663,N_4550,N_3161);
nand U7664 (N_7664,N_4079,N_4375);
or U7665 (N_7665,N_2326,N_3214);
or U7666 (N_7666,N_3140,N_1716);
nand U7667 (N_7667,N_4456,N_939);
nor U7668 (N_7668,N_4202,N_4193);
nand U7669 (N_7669,N_1251,N_2663);
and U7670 (N_7670,N_911,N_4500);
and U7671 (N_7671,N_2065,N_4280);
xor U7672 (N_7672,N_4528,N_120);
nor U7673 (N_7673,N_4244,N_2913);
xnor U7674 (N_7674,N_1927,N_4138);
or U7675 (N_7675,N_3533,N_4253);
xnor U7676 (N_7676,N_2588,N_632);
and U7677 (N_7677,N_3820,N_1039);
xnor U7678 (N_7678,N_3947,N_1676);
and U7679 (N_7679,N_4978,N_244);
xnor U7680 (N_7680,N_1918,N_4907);
nand U7681 (N_7681,N_1098,N_574);
and U7682 (N_7682,N_4523,N_3230);
nor U7683 (N_7683,N_1035,N_510);
and U7684 (N_7684,N_3992,N_1555);
or U7685 (N_7685,N_662,N_32);
nand U7686 (N_7686,N_412,N_4288);
and U7687 (N_7687,N_2245,N_594);
nand U7688 (N_7688,N_4994,N_4506);
xor U7689 (N_7689,N_490,N_52);
nor U7690 (N_7690,N_3531,N_120);
nor U7691 (N_7691,N_1231,N_688);
and U7692 (N_7692,N_3204,N_2426);
nor U7693 (N_7693,N_2957,N_1946);
nor U7694 (N_7694,N_520,N_970);
nor U7695 (N_7695,N_3979,N_972);
xor U7696 (N_7696,N_3755,N_4751);
and U7697 (N_7697,N_3548,N_4486);
xor U7698 (N_7698,N_1770,N_699);
nand U7699 (N_7699,N_943,N_1111);
or U7700 (N_7700,N_4952,N_3950);
and U7701 (N_7701,N_2877,N_1088);
and U7702 (N_7702,N_3761,N_2758);
nand U7703 (N_7703,N_3488,N_1340);
and U7704 (N_7704,N_3447,N_4647);
nor U7705 (N_7705,N_577,N_4328);
xnor U7706 (N_7706,N_4825,N_4401);
nor U7707 (N_7707,N_3795,N_4570);
and U7708 (N_7708,N_4578,N_1952);
nor U7709 (N_7709,N_3894,N_2456);
or U7710 (N_7710,N_3323,N_4258);
nand U7711 (N_7711,N_1843,N_3170);
nor U7712 (N_7712,N_4657,N_4082);
and U7713 (N_7713,N_2145,N_4617);
or U7714 (N_7714,N_3414,N_4365);
nand U7715 (N_7715,N_4926,N_3960);
xor U7716 (N_7716,N_2635,N_3213);
and U7717 (N_7717,N_2091,N_1305);
xor U7718 (N_7718,N_3000,N_4741);
xnor U7719 (N_7719,N_4936,N_1147);
and U7720 (N_7720,N_4692,N_1467);
and U7721 (N_7721,N_2442,N_1947);
and U7722 (N_7722,N_857,N_682);
or U7723 (N_7723,N_438,N_3342);
nand U7724 (N_7724,N_3989,N_1350);
nor U7725 (N_7725,N_3234,N_2806);
nor U7726 (N_7726,N_4648,N_3735);
and U7727 (N_7727,N_2669,N_3534);
nand U7728 (N_7728,N_4372,N_2707);
xnor U7729 (N_7729,N_4480,N_1225);
nor U7730 (N_7730,N_1407,N_3510);
xnor U7731 (N_7731,N_160,N_3230);
or U7732 (N_7732,N_4512,N_340);
and U7733 (N_7733,N_4512,N_3099);
nand U7734 (N_7734,N_1531,N_4790);
or U7735 (N_7735,N_4779,N_3856);
or U7736 (N_7736,N_1014,N_504);
xnor U7737 (N_7737,N_164,N_423);
nand U7738 (N_7738,N_3472,N_2122);
and U7739 (N_7739,N_1899,N_4671);
nor U7740 (N_7740,N_1037,N_1407);
or U7741 (N_7741,N_4636,N_3397);
and U7742 (N_7742,N_4193,N_4431);
or U7743 (N_7743,N_2182,N_3287);
or U7744 (N_7744,N_2759,N_1065);
nor U7745 (N_7745,N_167,N_1866);
or U7746 (N_7746,N_2942,N_2755);
xnor U7747 (N_7747,N_366,N_2311);
nor U7748 (N_7748,N_1022,N_3535);
nand U7749 (N_7749,N_4617,N_4108);
nor U7750 (N_7750,N_3726,N_2222);
nor U7751 (N_7751,N_4140,N_3137);
or U7752 (N_7752,N_841,N_1063);
nor U7753 (N_7753,N_2356,N_3170);
xor U7754 (N_7754,N_4508,N_2992);
or U7755 (N_7755,N_830,N_2946);
xnor U7756 (N_7756,N_3721,N_1460);
and U7757 (N_7757,N_1782,N_1674);
nor U7758 (N_7758,N_4023,N_1372);
and U7759 (N_7759,N_1306,N_3498);
nor U7760 (N_7760,N_3114,N_356);
nor U7761 (N_7761,N_1552,N_4);
xor U7762 (N_7762,N_1977,N_1031);
xor U7763 (N_7763,N_4666,N_3107);
and U7764 (N_7764,N_3881,N_1149);
xnor U7765 (N_7765,N_676,N_1067);
and U7766 (N_7766,N_2413,N_2592);
nand U7767 (N_7767,N_4042,N_3814);
or U7768 (N_7768,N_2546,N_1227);
xnor U7769 (N_7769,N_375,N_4398);
nand U7770 (N_7770,N_3561,N_1663);
and U7771 (N_7771,N_1004,N_1303);
and U7772 (N_7772,N_4871,N_1755);
nor U7773 (N_7773,N_364,N_455);
nor U7774 (N_7774,N_4556,N_2419);
or U7775 (N_7775,N_3603,N_1450);
and U7776 (N_7776,N_1185,N_2322);
nand U7777 (N_7777,N_314,N_2218);
nor U7778 (N_7778,N_225,N_4464);
nand U7779 (N_7779,N_1386,N_4189);
or U7780 (N_7780,N_811,N_2914);
nor U7781 (N_7781,N_364,N_4148);
or U7782 (N_7782,N_3924,N_4468);
nor U7783 (N_7783,N_1574,N_1379);
nand U7784 (N_7784,N_2796,N_3727);
nor U7785 (N_7785,N_3332,N_1979);
or U7786 (N_7786,N_2072,N_4963);
nand U7787 (N_7787,N_1920,N_1647);
and U7788 (N_7788,N_4969,N_2805);
nor U7789 (N_7789,N_1707,N_1946);
and U7790 (N_7790,N_4654,N_1966);
and U7791 (N_7791,N_2186,N_1317);
nand U7792 (N_7792,N_4363,N_772);
nand U7793 (N_7793,N_800,N_550);
nor U7794 (N_7794,N_1331,N_653);
nand U7795 (N_7795,N_3131,N_3552);
and U7796 (N_7796,N_1438,N_1584);
nand U7797 (N_7797,N_238,N_1983);
nor U7798 (N_7798,N_3092,N_2903);
or U7799 (N_7799,N_2700,N_3042);
xnor U7800 (N_7800,N_3081,N_2593);
xor U7801 (N_7801,N_1474,N_862);
nor U7802 (N_7802,N_2131,N_1110);
nand U7803 (N_7803,N_4037,N_4033);
and U7804 (N_7804,N_4135,N_4217);
and U7805 (N_7805,N_4488,N_4507);
or U7806 (N_7806,N_3153,N_1702);
nor U7807 (N_7807,N_332,N_2398);
or U7808 (N_7808,N_4715,N_4899);
xnor U7809 (N_7809,N_2722,N_1246);
nor U7810 (N_7810,N_1295,N_3214);
xnor U7811 (N_7811,N_3823,N_1280);
nor U7812 (N_7812,N_1604,N_3687);
xor U7813 (N_7813,N_441,N_1321);
nor U7814 (N_7814,N_2204,N_1398);
and U7815 (N_7815,N_712,N_3199);
and U7816 (N_7816,N_2602,N_4322);
nand U7817 (N_7817,N_784,N_4916);
xor U7818 (N_7818,N_915,N_608);
or U7819 (N_7819,N_4643,N_1902);
nor U7820 (N_7820,N_2523,N_1282);
xnor U7821 (N_7821,N_1887,N_173);
and U7822 (N_7822,N_271,N_2870);
xnor U7823 (N_7823,N_3334,N_2593);
or U7824 (N_7824,N_1210,N_1756);
nor U7825 (N_7825,N_622,N_4284);
or U7826 (N_7826,N_3895,N_2330);
nor U7827 (N_7827,N_412,N_260);
or U7828 (N_7828,N_1316,N_124);
or U7829 (N_7829,N_2366,N_2170);
nor U7830 (N_7830,N_2703,N_789);
nand U7831 (N_7831,N_1918,N_3307);
or U7832 (N_7832,N_3680,N_1170);
xor U7833 (N_7833,N_155,N_1218);
or U7834 (N_7834,N_1189,N_621);
and U7835 (N_7835,N_362,N_631);
and U7836 (N_7836,N_1257,N_257);
nand U7837 (N_7837,N_350,N_1341);
nor U7838 (N_7838,N_3787,N_1409);
or U7839 (N_7839,N_1498,N_4094);
xnor U7840 (N_7840,N_4781,N_2407);
nand U7841 (N_7841,N_1019,N_3434);
or U7842 (N_7842,N_2577,N_547);
nor U7843 (N_7843,N_4039,N_2476);
nand U7844 (N_7844,N_2898,N_2025);
nor U7845 (N_7845,N_4894,N_2534);
nand U7846 (N_7846,N_4540,N_2987);
and U7847 (N_7847,N_1611,N_4693);
xor U7848 (N_7848,N_3928,N_1819);
or U7849 (N_7849,N_3576,N_813);
xnor U7850 (N_7850,N_1463,N_4830);
or U7851 (N_7851,N_808,N_1993);
xor U7852 (N_7852,N_4995,N_3771);
and U7853 (N_7853,N_3120,N_906);
nor U7854 (N_7854,N_3063,N_4788);
xor U7855 (N_7855,N_2749,N_3252);
nand U7856 (N_7856,N_4050,N_4414);
nor U7857 (N_7857,N_1693,N_1341);
xor U7858 (N_7858,N_428,N_3614);
nor U7859 (N_7859,N_1211,N_654);
and U7860 (N_7860,N_1901,N_3631);
xnor U7861 (N_7861,N_2765,N_353);
xnor U7862 (N_7862,N_4232,N_3341);
nand U7863 (N_7863,N_3230,N_2320);
nand U7864 (N_7864,N_1590,N_3386);
nand U7865 (N_7865,N_763,N_970);
xnor U7866 (N_7866,N_2525,N_1478);
and U7867 (N_7867,N_868,N_3681);
or U7868 (N_7868,N_1592,N_3066);
nand U7869 (N_7869,N_3864,N_4166);
or U7870 (N_7870,N_4780,N_2198);
nor U7871 (N_7871,N_1689,N_1656);
and U7872 (N_7872,N_2308,N_3282);
or U7873 (N_7873,N_282,N_4881);
nand U7874 (N_7874,N_2014,N_1351);
nand U7875 (N_7875,N_657,N_4177);
xnor U7876 (N_7876,N_3789,N_3303);
xnor U7877 (N_7877,N_2885,N_1901);
xnor U7878 (N_7878,N_2359,N_4551);
xnor U7879 (N_7879,N_2877,N_1141);
xor U7880 (N_7880,N_1721,N_4585);
nor U7881 (N_7881,N_1973,N_698);
nand U7882 (N_7882,N_3037,N_3797);
or U7883 (N_7883,N_2165,N_3254);
and U7884 (N_7884,N_3941,N_3770);
nor U7885 (N_7885,N_2005,N_1521);
xor U7886 (N_7886,N_1416,N_1016);
xnor U7887 (N_7887,N_2238,N_2593);
xnor U7888 (N_7888,N_4005,N_4681);
nand U7889 (N_7889,N_2503,N_2405);
and U7890 (N_7890,N_1866,N_908);
xnor U7891 (N_7891,N_3267,N_4227);
and U7892 (N_7892,N_2241,N_4394);
nand U7893 (N_7893,N_3258,N_2168);
nand U7894 (N_7894,N_730,N_2453);
and U7895 (N_7895,N_2244,N_2251);
nand U7896 (N_7896,N_1702,N_3734);
or U7897 (N_7897,N_758,N_252);
or U7898 (N_7898,N_2730,N_3680);
or U7899 (N_7899,N_1959,N_2039);
nand U7900 (N_7900,N_4888,N_2323);
and U7901 (N_7901,N_1360,N_3988);
or U7902 (N_7902,N_1005,N_4786);
nor U7903 (N_7903,N_3561,N_2560);
xnor U7904 (N_7904,N_113,N_1247);
and U7905 (N_7905,N_4717,N_3851);
nor U7906 (N_7906,N_4247,N_4410);
xor U7907 (N_7907,N_1137,N_3343);
xnor U7908 (N_7908,N_192,N_1255);
and U7909 (N_7909,N_365,N_2009);
xnor U7910 (N_7910,N_3799,N_2125);
and U7911 (N_7911,N_3046,N_4050);
xnor U7912 (N_7912,N_2316,N_2357);
xor U7913 (N_7913,N_1303,N_4382);
nor U7914 (N_7914,N_70,N_2970);
or U7915 (N_7915,N_3026,N_3482);
nand U7916 (N_7916,N_3092,N_1734);
and U7917 (N_7917,N_3476,N_2551);
or U7918 (N_7918,N_3200,N_3096);
xnor U7919 (N_7919,N_4304,N_178);
nand U7920 (N_7920,N_2806,N_4150);
and U7921 (N_7921,N_4987,N_3798);
xnor U7922 (N_7922,N_190,N_2951);
or U7923 (N_7923,N_3623,N_2969);
xor U7924 (N_7924,N_3440,N_1389);
and U7925 (N_7925,N_2992,N_2368);
nor U7926 (N_7926,N_4542,N_3578);
or U7927 (N_7927,N_4034,N_4400);
nand U7928 (N_7928,N_1466,N_4440);
xnor U7929 (N_7929,N_3632,N_3110);
nand U7930 (N_7930,N_2578,N_3301);
and U7931 (N_7931,N_726,N_934);
nand U7932 (N_7932,N_1176,N_3573);
xnor U7933 (N_7933,N_1306,N_620);
nand U7934 (N_7934,N_261,N_474);
or U7935 (N_7935,N_1851,N_2377);
xor U7936 (N_7936,N_760,N_4902);
nand U7937 (N_7937,N_3714,N_1906);
and U7938 (N_7938,N_1386,N_4756);
nor U7939 (N_7939,N_1275,N_2816);
nand U7940 (N_7940,N_129,N_3220);
xor U7941 (N_7941,N_811,N_4412);
and U7942 (N_7942,N_3349,N_1735);
nand U7943 (N_7943,N_3236,N_640);
and U7944 (N_7944,N_1517,N_316);
or U7945 (N_7945,N_3334,N_1722);
or U7946 (N_7946,N_2011,N_3289);
or U7947 (N_7947,N_3430,N_3435);
and U7948 (N_7948,N_2046,N_263);
or U7949 (N_7949,N_1466,N_1182);
xnor U7950 (N_7950,N_1281,N_2995);
or U7951 (N_7951,N_1098,N_536);
or U7952 (N_7952,N_3636,N_3477);
xor U7953 (N_7953,N_4578,N_4312);
nand U7954 (N_7954,N_1279,N_1965);
nor U7955 (N_7955,N_4434,N_3566);
nor U7956 (N_7956,N_4253,N_1266);
or U7957 (N_7957,N_1995,N_409);
xor U7958 (N_7958,N_4637,N_16);
xnor U7959 (N_7959,N_3752,N_354);
xor U7960 (N_7960,N_3629,N_515);
and U7961 (N_7961,N_2106,N_484);
nand U7962 (N_7962,N_3580,N_877);
and U7963 (N_7963,N_1825,N_2169);
xor U7964 (N_7964,N_203,N_3135);
or U7965 (N_7965,N_1118,N_4315);
nor U7966 (N_7966,N_393,N_539);
or U7967 (N_7967,N_1134,N_609);
and U7968 (N_7968,N_3632,N_3962);
nand U7969 (N_7969,N_1913,N_2731);
and U7970 (N_7970,N_540,N_4463);
nor U7971 (N_7971,N_1342,N_4968);
and U7972 (N_7972,N_4844,N_246);
or U7973 (N_7973,N_2033,N_813);
nand U7974 (N_7974,N_3054,N_3454);
and U7975 (N_7975,N_3937,N_381);
nor U7976 (N_7976,N_3511,N_3568);
and U7977 (N_7977,N_3106,N_3575);
or U7978 (N_7978,N_2080,N_257);
nand U7979 (N_7979,N_2236,N_607);
nor U7980 (N_7980,N_718,N_2675);
nand U7981 (N_7981,N_1384,N_1770);
xnor U7982 (N_7982,N_3792,N_4616);
nand U7983 (N_7983,N_4,N_2807);
nand U7984 (N_7984,N_3526,N_2565);
nor U7985 (N_7985,N_4014,N_338);
xnor U7986 (N_7986,N_4299,N_2608);
xnor U7987 (N_7987,N_2744,N_1024);
nor U7988 (N_7988,N_2262,N_2521);
nand U7989 (N_7989,N_1661,N_1328);
nand U7990 (N_7990,N_4646,N_497);
nand U7991 (N_7991,N_4018,N_2297);
or U7992 (N_7992,N_2622,N_846);
or U7993 (N_7993,N_1941,N_3130);
nand U7994 (N_7994,N_3586,N_1820);
nand U7995 (N_7995,N_4062,N_3997);
nand U7996 (N_7996,N_4335,N_4630);
nand U7997 (N_7997,N_1835,N_356);
and U7998 (N_7998,N_2421,N_14);
or U7999 (N_7999,N_1681,N_195);
xnor U8000 (N_8000,N_2700,N_1438);
nand U8001 (N_8001,N_2602,N_2661);
xnor U8002 (N_8002,N_2290,N_1865);
xnor U8003 (N_8003,N_1147,N_3762);
or U8004 (N_8004,N_4972,N_3444);
nand U8005 (N_8005,N_591,N_2504);
xnor U8006 (N_8006,N_3360,N_830);
nand U8007 (N_8007,N_2327,N_88);
xnor U8008 (N_8008,N_1506,N_1590);
nand U8009 (N_8009,N_1463,N_2637);
nand U8010 (N_8010,N_1802,N_3447);
nand U8011 (N_8011,N_4432,N_3322);
xor U8012 (N_8012,N_3225,N_3953);
nand U8013 (N_8013,N_3944,N_4792);
xnor U8014 (N_8014,N_2013,N_4666);
nand U8015 (N_8015,N_3415,N_1662);
nand U8016 (N_8016,N_3715,N_3221);
nor U8017 (N_8017,N_3311,N_706);
nor U8018 (N_8018,N_2730,N_1234);
and U8019 (N_8019,N_3162,N_4423);
or U8020 (N_8020,N_3532,N_4889);
and U8021 (N_8021,N_1020,N_4971);
xor U8022 (N_8022,N_3250,N_1901);
and U8023 (N_8023,N_2789,N_2117);
and U8024 (N_8024,N_3826,N_1808);
nand U8025 (N_8025,N_309,N_1738);
nand U8026 (N_8026,N_3148,N_1820);
or U8027 (N_8027,N_379,N_2242);
nor U8028 (N_8028,N_3448,N_3428);
nor U8029 (N_8029,N_3523,N_4013);
or U8030 (N_8030,N_4097,N_3639);
nor U8031 (N_8031,N_2255,N_4038);
nor U8032 (N_8032,N_6,N_2812);
and U8033 (N_8033,N_1636,N_4282);
nand U8034 (N_8034,N_1744,N_803);
nand U8035 (N_8035,N_4429,N_4257);
nand U8036 (N_8036,N_2598,N_134);
and U8037 (N_8037,N_230,N_2218);
xnor U8038 (N_8038,N_4925,N_2202);
nor U8039 (N_8039,N_1931,N_197);
xnor U8040 (N_8040,N_73,N_2473);
or U8041 (N_8041,N_3878,N_3843);
xnor U8042 (N_8042,N_2219,N_3220);
and U8043 (N_8043,N_4599,N_4922);
xnor U8044 (N_8044,N_1888,N_917);
xor U8045 (N_8045,N_2447,N_2861);
nand U8046 (N_8046,N_2544,N_3520);
and U8047 (N_8047,N_3325,N_4715);
nor U8048 (N_8048,N_3047,N_2601);
xnor U8049 (N_8049,N_1565,N_3192);
xnor U8050 (N_8050,N_278,N_2947);
nand U8051 (N_8051,N_2876,N_3308);
nor U8052 (N_8052,N_2172,N_77);
or U8053 (N_8053,N_602,N_4351);
and U8054 (N_8054,N_3173,N_487);
xnor U8055 (N_8055,N_4935,N_3598);
or U8056 (N_8056,N_3423,N_2697);
nor U8057 (N_8057,N_2207,N_3104);
xor U8058 (N_8058,N_2429,N_912);
nand U8059 (N_8059,N_4941,N_3327);
nor U8060 (N_8060,N_4209,N_59);
xnor U8061 (N_8061,N_510,N_1154);
nor U8062 (N_8062,N_1349,N_1958);
and U8063 (N_8063,N_4660,N_20);
nor U8064 (N_8064,N_968,N_4646);
nand U8065 (N_8065,N_2486,N_1789);
and U8066 (N_8066,N_1862,N_948);
or U8067 (N_8067,N_613,N_850);
xnor U8068 (N_8068,N_3370,N_1700);
nand U8069 (N_8069,N_1431,N_225);
and U8070 (N_8070,N_321,N_2855);
or U8071 (N_8071,N_3494,N_3389);
nor U8072 (N_8072,N_3011,N_1568);
or U8073 (N_8073,N_2253,N_3970);
nor U8074 (N_8074,N_699,N_3919);
xnor U8075 (N_8075,N_159,N_325);
nand U8076 (N_8076,N_1399,N_2841);
xnor U8077 (N_8077,N_2004,N_1961);
nand U8078 (N_8078,N_2833,N_532);
nor U8079 (N_8079,N_4473,N_819);
or U8080 (N_8080,N_1501,N_2087);
or U8081 (N_8081,N_3647,N_3662);
nand U8082 (N_8082,N_3666,N_2725);
nand U8083 (N_8083,N_2912,N_4723);
xnor U8084 (N_8084,N_2154,N_2592);
nor U8085 (N_8085,N_1079,N_4954);
nand U8086 (N_8086,N_1720,N_3902);
nor U8087 (N_8087,N_1691,N_2970);
or U8088 (N_8088,N_4446,N_2940);
and U8089 (N_8089,N_1187,N_4789);
nor U8090 (N_8090,N_4325,N_3147);
nor U8091 (N_8091,N_2819,N_1766);
nand U8092 (N_8092,N_2911,N_3621);
nand U8093 (N_8093,N_3090,N_3874);
xor U8094 (N_8094,N_776,N_1194);
or U8095 (N_8095,N_1913,N_425);
and U8096 (N_8096,N_4253,N_2283);
and U8097 (N_8097,N_3266,N_907);
and U8098 (N_8098,N_3964,N_489);
xnor U8099 (N_8099,N_484,N_1352);
nor U8100 (N_8100,N_3433,N_3507);
xor U8101 (N_8101,N_3970,N_4392);
or U8102 (N_8102,N_1397,N_839);
xnor U8103 (N_8103,N_2418,N_2039);
or U8104 (N_8104,N_794,N_3383);
xnor U8105 (N_8105,N_2024,N_4482);
or U8106 (N_8106,N_439,N_3154);
nand U8107 (N_8107,N_1128,N_2893);
nor U8108 (N_8108,N_2140,N_686);
nand U8109 (N_8109,N_3226,N_3093);
nor U8110 (N_8110,N_432,N_295);
or U8111 (N_8111,N_2497,N_4565);
xor U8112 (N_8112,N_3975,N_677);
or U8113 (N_8113,N_1693,N_2893);
xor U8114 (N_8114,N_3910,N_3432);
nand U8115 (N_8115,N_3985,N_3104);
nor U8116 (N_8116,N_1731,N_417);
nor U8117 (N_8117,N_4973,N_1557);
nor U8118 (N_8118,N_2477,N_3706);
xnor U8119 (N_8119,N_1269,N_1963);
nand U8120 (N_8120,N_3949,N_3801);
nor U8121 (N_8121,N_2252,N_341);
and U8122 (N_8122,N_3563,N_1021);
xnor U8123 (N_8123,N_2320,N_4750);
or U8124 (N_8124,N_51,N_584);
or U8125 (N_8125,N_1297,N_2117);
xor U8126 (N_8126,N_4219,N_2398);
and U8127 (N_8127,N_2208,N_4927);
nand U8128 (N_8128,N_663,N_1385);
and U8129 (N_8129,N_14,N_412);
and U8130 (N_8130,N_4232,N_3978);
nor U8131 (N_8131,N_4589,N_2585);
xor U8132 (N_8132,N_3980,N_3141);
and U8133 (N_8133,N_4912,N_4848);
and U8134 (N_8134,N_1954,N_778);
nor U8135 (N_8135,N_3733,N_116);
and U8136 (N_8136,N_215,N_358);
nand U8137 (N_8137,N_3293,N_1685);
nand U8138 (N_8138,N_2528,N_3276);
xor U8139 (N_8139,N_3449,N_3898);
xor U8140 (N_8140,N_3760,N_4444);
and U8141 (N_8141,N_939,N_533);
nand U8142 (N_8142,N_2416,N_1475);
and U8143 (N_8143,N_1841,N_3798);
nor U8144 (N_8144,N_1223,N_4777);
or U8145 (N_8145,N_2878,N_24);
and U8146 (N_8146,N_4030,N_1725);
or U8147 (N_8147,N_4690,N_2473);
or U8148 (N_8148,N_4417,N_570);
nand U8149 (N_8149,N_4638,N_656);
nor U8150 (N_8150,N_4476,N_4243);
and U8151 (N_8151,N_2904,N_473);
and U8152 (N_8152,N_1881,N_1312);
xnor U8153 (N_8153,N_3675,N_147);
or U8154 (N_8154,N_3779,N_2323);
or U8155 (N_8155,N_690,N_359);
nand U8156 (N_8156,N_530,N_547);
and U8157 (N_8157,N_1984,N_1348);
nand U8158 (N_8158,N_3956,N_1990);
nor U8159 (N_8159,N_4813,N_444);
nand U8160 (N_8160,N_4324,N_4669);
xnor U8161 (N_8161,N_1829,N_4297);
nand U8162 (N_8162,N_2406,N_3362);
and U8163 (N_8163,N_1504,N_1073);
nor U8164 (N_8164,N_4387,N_2602);
xnor U8165 (N_8165,N_410,N_2871);
nor U8166 (N_8166,N_42,N_3341);
xor U8167 (N_8167,N_1185,N_3432);
xor U8168 (N_8168,N_31,N_283);
xnor U8169 (N_8169,N_2709,N_2693);
nor U8170 (N_8170,N_1634,N_4580);
xnor U8171 (N_8171,N_4724,N_4354);
nand U8172 (N_8172,N_525,N_3376);
or U8173 (N_8173,N_1631,N_2874);
xor U8174 (N_8174,N_1954,N_1345);
nor U8175 (N_8175,N_2968,N_1279);
nor U8176 (N_8176,N_1932,N_230);
nand U8177 (N_8177,N_3134,N_397);
xnor U8178 (N_8178,N_3143,N_645);
or U8179 (N_8179,N_1741,N_2193);
nor U8180 (N_8180,N_3627,N_2001);
xnor U8181 (N_8181,N_4430,N_4976);
and U8182 (N_8182,N_2015,N_402);
nor U8183 (N_8183,N_4095,N_3237);
and U8184 (N_8184,N_1556,N_3691);
and U8185 (N_8185,N_1752,N_3622);
nand U8186 (N_8186,N_1965,N_981);
and U8187 (N_8187,N_455,N_4160);
and U8188 (N_8188,N_224,N_1743);
or U8189 (N_8189,N_3308,N_2860);
or U8190 (N_8190,N_3034,N_3258);
or U8191 (N_8191,N_3399,N_3884);
nand U8192 (N_8192,N_1771,N_891);
nand U8193 (N_8193,N_1212,N_2275);
and U8194 (N_8194,N_2219,N_1033);
nand U8195 (N_8195,N_1413,N_1987);
or U8196 (N_8196,N_447,N_3835);
or U8197 (N_8197,N_1819,N_2386);
nor U8198 (N_8198,N_517,N_1189);
nand U8199 (N_8199,N_3969,N_2217);
nor U8200 (N_8200,N_4960,N_4001);
xor U8201 (N_8201,N_424,N_2951);
nand U8202 (N_8202,N_2626,N_3028);
nand U8203 (N_8203,N_2063,N_1865);
nor U8204 (N_8204,N_1029,N_2117);
nor U8205 (N_8205,N_1479,N_3313);
xor U8206 (N_8206,N_2644,N_4622);
nor U8207 (N_8207,N_4023,N_4680);
nand U8208 (N_8208,N_3961,N_2239);
and U8209 (N_8209,N_4845,N_33);
and U8210 (N_8210,N_886,N_4710);
xnor U8211 (N_8211,N_2619,N_2046);
and U8212 (N_8212,N_1817,N_4595);
nand U8213 (N_8213,N_1173,N_1774);
and U8214 (N_8214,N_1267,N_4143);
nor U8215 (N_8215,N_1757,N_1410);
and U8216 (N_8216,N_1647,N_2413);
nand U8217 (N_8217,N_2715,N_2936);
and U8218 (N_8218,N_2727,N_284);
nor U8219 (N_8219,N_2223,N_4643);
and U8220 (N_8220,N_2344,N_1332);
xnor U8221 (N_8221,N_458,N_1589);
nand U8222 (N_8222,N_448,N_4173);
nor U8223 (N_8223,N_4500,N_3975);
and U8224 (N_8224,N_400,N_1038);
nand U8225 (N_8225,N_2606,N_2417);
nand U8226 (N_8226,N_3708,N_4875);
and U8227 (N_8227,N_4612,N_1086);
nand U8228 (N_8228,N_4626,N_4992);
nor U8229 (N_8229,N_2233,N_4421);
xor U8230 (N_8230,N_300,N_3668);
xnor U8231 (N_8231,N_4440,N_2696);
or U8232 (N_8232,N_3074,N_1374);
and U8233 (N_8233,N_546,N_752);
xnor U8234 (N_8234,N_829,N_3659);
nor U8235 (N_8235,N_3721,N_2239);
xnor U8236 (N_8236,N_1915,N_308);
nand U8237 (N_8237,N_519,N_1456);
nor U8238 (N_8238,N_4771,N_2969);
or U8239 (N_8239,N_965,N_324);
nor U8240 (N_8240,N_2542,N_3481);
and U8241 (N_8241,N_858,N_3333);
or U8242 (N_8242,N_2303,N_907);
and U8243 (N_8243,N_201,N_190);
or U8244 (N_8244,N_2444,N_81);
xor U8245 (N_8245,N_2530,N_1306);
nor U8246 (N_8246,N_968,N_3148);
nand U8247 (N_8247,N_4055,N_2253);
or U8248 (N_8248,N_2911,N_534);
or U8249 (N_8249,N_2608,N_909);
nand U8250 (N_8250,N_3716,N_1135);
nor U8251 (N_8251,N_3567,N_2374);
or U8252 (N_8252,N_2850,N_885);
nand U8253 (N_8253,N_974,N_3485);
nand U8254 (N_8254,N_4592,N_1569);
nor U8255 (N_8255,N_3159,N_1596);
nor U8256 (N_8256,N_3691,N_3271);
xor U8257 (N_8257,N_680,N_1572);
nand U8258 (N_8258,N_4841,N_1673);
nand U8259 (N_8259,N_2572,N_2965);
and U8260 (N_8260,N_3191,N_4886);
or U8261 (N_8261,N_4023,N_408);
or U8262 (N_8262,N_2455,N_2955);
nor U8263 (N_8263,N_755,N_2279);
and U8264 (N_8264,N_924,N_1675);
nand U8265 (N_8265,N_1394,N_3630);
nor U8266 (N_8266,N_3600,N_1983);
or U8267 (N_8267,N_4265,N_1853);
nor U8268 (N_8268,N_3861,N_1687);
nor U8269 (N_8269,N_4984,N_4185);
xor U8270 (N_8270,N_3050,N_2010);
or U8271 (N_8271,N_853,N_4942);
xnor U8272 (N_8272,N_2093,N_872);
xnor U8273 (N_8273,N_2312,N_3409);
and U8274 (N_8274,N_4689,N_819);
or U8275 (N_8275,N_4771,N_3813);
or U8276 (N_8276,N_3797,N_4746);
or U8277 (N_8277,N_639,N_4003);
nand U8278 (N_8278,N_1456,N_138);
xor U8279 (N_8279,N_2534,N_290);
or U8280 (N_8280,N_4596,N_1168);
and U8281 (N_8281,N_807,N_2861);
or U8282 (N_8282,N_2539,N_765);
or U8283 (N_8283,N_1739,N_4753);
and U8284 (N_8284,N_2105,N_1225);
xor U8285 (N_8285,N_2800,N_4858);
or U8286 (N_8286,N_1762,N_829);
nor U8287 (N_8287,N_4653,N_1568);
nand U8288 (N_8288,N_995,N_2678);
nand U8289 (N_8289,N_1328,N_2586);
nor U8290 (N_8290,N_1199,N_563);
or U8291 (N_8291,N_1172,N_4800);
nor U8292 (N_8292,N_4981,N_4284);
xor U8293 (N_8293,N_4613,N_4537);
xor U8294 (N_8294,N_1532,N_4963);
nor U8295 (N_8295,N_2028,N_3046);
xor U8296 (N_8296,N_818,N_3970);
nor U8297 (N_8297,N_42,N_175);
or U8298 (N_8298,N_1439,N_3600);
nor U8299 (N_8299,N_3740,N_2422);
or U8300 (N_8300,N_4064,N_2810);
nor U8301 (N_8301,N_2251,N_4976);
and U8302 (N_8302,N_1182,N_62);
nand U8303 (N_8303,N_1745,N_4045);
nor U8304 (N_8304,N_2779,N_2822);
or U8305 (N_8305,N_2478,N_1959);
nor U8306 (N_8306,N_4326,N_4452);
and U8307 (N_8307,N_824,N_1728);
nand U8308 (N_8308,N_1566,N_4921);
xor U8309 (N_8309,N_1648,N_3669);
or U8310 (N_8310,N_3181,N_4820);
xnor U8311 (N_8311,N_997,N_2179);
or U8312 (N_8312,N_1264,N_4504);
and U8313 (N_8313,N_78,N_2712);
nor U8314 (N_8314,N_2929,N_2187);
xnor U8315 (N_8315,N_4674,N_2059);
and U8316 (N_8316,N_4266,N_4455);
xnor U8317 (N_8317,N_1295,N_1716);
nor U8318 (N_8318,N_2855,N_4325);
nand U8319 (N_8319,N_1573,N_3312);
and U8320 (N_8320,N_474,N_1605);
and U8321 (N_8321,N_2509,N_1771);
xnor U8322 (N_8322,N_1102,N_269);
nor U8323 (N_8323,N_1592,N_3584);
xor U8324 (N_8324,N_2618,N_4988);
xor U8325 (N_8325,N_2430,N_2207);
nor U8326 (N_8326,N_384,N_3259);
or U8327 (N_8327,N_3981,N_2132);
or U8328 (N_8328,N_1573,N_1981);
nor U8329 (N_8329,N_434,N_1622);
and U8330 (N_8330,N_2374,N_1291);
and U8331 (N_8331,N_881,N_1865);
or U8332 (N_8332,N_1025,N_4320);
xnor U8333 (N_8333,N_1950,N_4013);
xnor U8334 (N_8334,N_425,N_4740);
and U8335 (N_8335,N_4570,N_3568);
or U8336 (N_8336,N_3657,N_3397);
nand U8337 (N_8337,N_571,N_452);
nor U8338 (N_8338,N_1316,N_2968);
nor U8339 (N_8339,N_4909,N_4261);
xor U8340 (N_8340,N_1036,N_3385);
and U8341 (N_8341,N_2883,N_3585);
nor U8342 (N_8342,N_508,N_2092);
nand U8343 (N_8343,N_4974,N_2090);
and U8344 (N_8344,N_173,N_1462);
xor U8345 (N_8345,N_1722,N_2737);
nor U8346 (N_8346,N_1652,N_1768);
nor U8347 (N_8347,N_514,N_2823);
xnor U8348 (N_8348,N_4906,N_1622);
and U8349 (N_8349,N_3404,N_3343);
and U8350 (N_8350,N_729,N_1797);
or U8351 (N_8351,N_1043,N_1008);
or U8352 (N_8352,N_3775,N_3880);
and U8353 (N_8353,N_4661,N_488);
nand U8354 (N_8354,N_1850,N_2128);
or U8355 (N_8355,N_2750,N_971);
or U8356 (N_8356,N_4886,N_42);
xor U8357 (N_8357,N_1738,N_2848);
or U8358 (N_8358,N_4123,N_3309);
nand U8359 (N_8359,N_335,N_340);
and U8360 (N_8360,N_3919,N_513);
and U8361 (N_8361,N_4399,N_3168);
and U8362 (N_8362,N_389,N_2804);
xnor U8363 (N_8363,N_3649,N_3494);
or U8364 (N_8364,N_1025,N_4139);
nor U8365 (N_8365,N_1477,N_3220);
nand U8366 (N_8366,N_3535,N_2790);
nand U8367 (N_8367,N_1451,N_3412);
xor U8368 (N_8368,N_40,N_4599);
nand U8369 (N_8369,N_3838,N_2561);
or U8370 (N_8370,N_758,N_228);
or U8371 (N_8371,N_755,N_2445);
xor U8372 (N_8372,N_1783,N_67);
and U8373 (N_8373,N_2751,N_4625);
nor U8374 (N_8374,N_3027,N_3800);
nand U8375 (N_8375,N_2697,N_2991);
or U8376 (N_8376,N_4424,N_1974);
xor U8377 (N_8377,N_2493,N_4555);
xnor U8378 (N_8378,N_661,N_4835);
or U8379 (N_8379,N_3602,N_1569);
or U8380 (N_8380,N_1026,N_3555);
nor U8381 (N_8381,N_25,N_4346);
nor U8382 (N_8382,N_2561,N_3382);
or U8383 (N_8383,N_4299,N_1467);
nor U8384 (N_8384,N_59,N_75);
nand U8385 (N_8385,N_1560,N_2049);
and U8386 (N_8386,N_4601,N_1282);
or U8387 (N_8387,N_4448,N_2936);
nor U8388 (N_8388,N_3704,N_174);
or U8389 (N_8389,N_3032,N_1444);
nor U8390 (N_8390,N_3649,N_2339);
nand U8391 (N_8391,N_2340,N_1013);
or U8392 (N_8392,N_328,N_4203);
or U8393 (N_8393,N_715,N_3912);
and U8394 (N_8394,N_1448,N_1549);
nand U8395 (N_8395,N_2113,N_2926);
xor U8396 (N_8396,N_4366,N_4409);
xnor U8397 (N_8397,N_2561,N_3347);
nor U8398 (N_8398,N_928,N_2596);
nor U8399 (N_8399,N_837,N_2849);
or U8400 (N_8400,N_3646,N_1086);
or U8401 (N_8401,N_13,N_2053);
xor U8402 (N_8402,N_1466,N_1872);
nor U8403 (N_8403,N_964,N_2296);
nand U8404 (N_8404,N_968,N_2921);
xor U8405 (N_8405,N_2940,N_1012);
or U8406 (N_8406,N_3455,N_4127);
and U8407 (N_8407,N_3385,N_1297);
or U8408 (N_8408,N_728,N_4503);
nand U8409 (N_8409,N_429,N_4678);
nor U8410 (N_8410,N_4580,N_2432);
nor U8411 (N_8411,N_4015,N_2659);
and U8412 (N_8412,N_4706,N_201);
or U8413 (N_8413,N_762,N_4205);
xnor U8414 (N_8414,N_4197,N_1698);
nor U8415 (N_8415,N_2866,N_3811);
or U8416 (N_8416,N_2837,N_2328);
xor U8417 (N_8417,N_1671,N_226);
nand U8418 (N_8418,N_675,N_2937);
nand U8419 (N_8419,N_741,N_2331);
xnor U8420 (N_8420,N_1765,N_866);
nand U8421 (N_8421,N_750,N_1157);
xor U8422 (N_8422,N_1112,N_2616);
or U8423 (N_8423,N_4977,N_3611);
nand U8424 (N_8424,N_3915,N_3754);
or U8425 (N_8425,N_2431,N_1853);
nand U8426 (N_8426,N_1051,N_1213);
nor U8427 (N_8427,N_2103,N_1271);
nand U8428 (N_8428,N_3825,N_2885);
or U8429 (N_8429,N_877,N_422);
nor U8430 (N_8430,N_1679,N_4912);
nor U8431 (N_8431,N_4219,N_2519);
nor U8432 (N_8432,N_3124,N_3640);
nor U8433 (N_8433,N_3092,N_3026);
xnor U8434 (N_8434,N_3777,N_895);
nor U8435 (N_8435,N_4038,N_4604);
nand U8436 (N_8436,N_2258,N_604);
or U8437 (N_8437,N_3546,N_1278);
nand U8438 (N_8438,N_1445,N_3184);
and U8439 (N_8439,N_4718,N_390);
xor U8440 (N_8440,N_378,N_3196);
or U8441 (N_8441,N_1283,N_2962);
and U8442 (N_8442,N_2375,N_1287);
nor U8443 (N_8443,N_1369,N_4968);
and U8444 (N_8444,N_2922,N_1765);
or U8445 (N_8445,N_3650,N_1411);
or U8446 (N_8446,N_4913,N_4164);
xnor U8447 (N_8447,N_1287,N_4543);
nor U8448 (N_8448,N_3056,N_2326);
xnor U8449 (N_8449,N_3875,N_1486);
nand U8450 (N_8450,N_4493,N_4096);
nand U8451 (N_8451,N_4032,N_327);
nand U8452 (N_8452,N_1268,N_3531);
nor U8453 (N_8453,N_2527,N_1947);
and U8454 (N_8454,N_1064,N_2062);
nor U8455 (N_8455,N_15,N_2096);
and U8456 (N_8456,N_881,N_272);
nand U8457 (N_8457,N_3581,N_4370);
nor U8458 (N_8458,N_1664,N_2894);
nand U8459 (N_8459,N_2581,N_3803);
xor U8460 (N_8460,N_2232,N_1039);
nand U8461 (N_8461,N_3355,N_2737);
nor U8462 (N_8462,N_1625,N_1090);
or U8463 (N_8463,N_1992,N_856);
or U8464 (N_8464,N_4251,N_2364);
xnor U8465 (N_8465,N_3511,N_4453);
nor U8466 (N_8466,N_1182,N_1355);
nor U8467 (N_8467,N_4408,N_4364);
and U8468 (N_8468,N_2922,N_2853);
nor U8469 (N_8469,N_4689,N_1395);
and U8470 (N_8470,N_228,N_3642);
and U8471 (N_8471,N_4467,N_3030);
nor U8472 (N_8472,N_2526,N_3153);
nand U8473 (N_8473,N_2391,N_4121);
xnor U8474 (N_8474,N_915,N_3395);
nor U8475 (N_8475,N_1469,N_3573);
or U8476 (N_8476,N_3843,N_1559);
or U8477 (N_8477,N_1759,N_4922);
nor U8478 (N_8478,N_751,N_3545);
nand U8479 (N_8479,N_2415,N_2522);
nand U8480 (N_8480,N_4653,N_3023);
xnor U8481 (N_8481,N_1040,N_4583);
and U8482 (N_8482,N_2205,N_205);
nand U8483 (N_8483,N_3305,N_2786);
xor U8484 (N_8484,N_362,N_506);
and U8485 (N_8485,N_1874,N_4493);
xnor U8486 (N_8486,N_737,N_2496);
xnor U8487 (N_8487,N_2706,N_3704);
nand U8488 (N_8488,N_3590,N_2025);
nand U8489 (N_8489,N_3403,N_1546);
and U8490 (N_8490,N_4679,N_2110);
nor U8491 (N_8491,N_200,N_1973);
or U8492 (N_8492,N_545,N_1635);
nor U8493 (N_8493,N_509,N_2875);
xnor U8494 (N_8494,N_2738,N_220);
nor U8495 (N_8495,N_1112,N_1937);
nand U8496 (N_8496,N_3725,N_3294);
nor U8497 (N_8497,N_2977,N_4378);
xor U8498 (N_8498,N_942,N_102);
nand U8499 (N_8499,N_2923,N_4766);
and U8500 (N_8500,N_182,N_3594);
xnor U8501 (N_8501,N_2058,N_1751);
nor U8502 (N_8502,N_1290,N_4383);
xnor U8503 (N_8503,N_4165,N_3388);
nand U8504 (N_8504,N_2840,N_2038);
xor U8505 (N_8505,N_4770,N_3219);
nand U8506 (N_8506,N_2275,N_2101);
nor U8507 (N_8507,N_4635,N_4782);
and U8508 (N_8508,N_5,N_4221);
and U8509 (N_8509,N_1946,N_1968);
nor U8510 (N_8510,N_3858,N_1592);
or U8511 (N_8511,N_4739,N_2770);
nand U8512 (N_8512,N_717,N_1097);
or U8513 (N_8513,N_3548,N_64);
xor U8514 (N_8514,N_72,N_3944);
nor U8515 (N_8515,N_2466,N_3919);
and U8516 (N_8516,N_3574,N_4645);
and U8517 (N_8517,N_1479,N_2645);
nand U8518 (N_8518,N_4059,N_2164);
nand U8519 (N_8519,N_3647,N_4490);
or U8520 (N_8520,N_3486,N_2386);
or U8521 (N_8521,N_1004,N_3278);
nor U8522 (N_8522,N_589,N_4089);
nand U8523 (N_8523,N_2369,N_4067);
xnor U8524 (N_8524,N_3553,N_257);
nand U8525 (N_8525,N_1984,N_3615);
and U8526 (N_8526,N_2432,N_4729);
nor U8527 (N_8527,N_236,N_4111);
and U8528 (N_8528,N_3279,N_3920);
or U8529 (N_8529,N_287,N_1512);
or U8530 (N_8530,N_2538,N_4230);
nand U8531 (N_8531,N_3072,N_2043);
xor U8532 (N_8532,N_3915,N_1899);
or U8533 (N_8533,N_815,N_819);
or U8534 (N_8534,N_1300,N_3525);
nand U8535 (N_8535,N_1390,N_671);
or U8536 (N_8536,N_2964,N_2015);
or U8537 (N_8537,N_164,N_1352);
and U8538 (N_8538,N_3839,N_4861);
nor U8539 (N_8539,N_3707,N_3993);
nor U8540 (N_8540,N_728,N_1222);
xor U8541 (N_8541,N_2438,N_677);
or U8542 (N_8542,N_118,N_3658);
and U8543 (N_8543,N_4593,N_3290);
and U8544 (N_8544,N_2911,N_4597);
or U8545 (N_8545,N_3434,N_1841);
nor U8546 (N_8546,N_564,N_2966);
or U8547 (N_8547,N_980,N_3631);
nand U8548 (N_8548,N_2527,N_889);
and U8549 (N_8549,N_1603,N_4766);
and U8550 (N_8550,N_737,N_960);
or U8551 (N_8551,N_2638,N_4918);
xnor U8552 (N_8552,N_4625,N_1001);
or U8553 (N_8553,N_893,N_4821);
xnor U8554 (N_8554,N_4760,N_4705);
or U8555 (N_8555,N_3876,N_817);
or U8556 (N_8556,N_2709,N_4079);
nor U8557 (N_8557,N_4730,N_4135);
xor U8558 (N_8558,N_2249,N_4908);
nor U8559 (N_8559,N_2266,N_539);
xor U8560 (N_8560,N_3941,N_3140);
and U8561 (N_8561,N_1446,N_572);
or U8562 (N_8562,N_2405,N_2573);
or U8563 (N_8563,N_1806,N_1654);
nand U8564 (N_8564,N_1053,N_908);
nand U8565 (N_8565,N_1453,N_4223);
or U8566 (N_8566,N_2301,N_1128);
and U8567 (N_8567,N_1681,N_1230);
nand U8568 (N_8568,N_2590,N_4073);
xnor U8569 (N_8569,N_3181,N_3497);
and U8570 (N_8570,N_1292,N_2408);
and U8571 (N_8571,N_3694,N_1299);
and U8572 (N_8572,N_3002,N_2271);
and U8573 (N_8573,N_2628,N_4128);
nor U8574 (N_8574,N_458,N_3154);
and U8575 (N_8575,N_4177,N_1476);
xor U8576 (N_8576,N_1933,N_1697);
xnor U8577 (N_8577,N_3500,N_4107);
or U8578 (N_8578,N_3506,N_3402);
nor U8579 (N_8579,N_4785,N_3176);
xnor U8580 (N_8580,N_4301,N_1810);
and U8581 (N_8581,N_3184,N_4133);
and U8582 (N_8582,N_3535,N_1280);
nand U8583 (N_8583,N_112,N_55);
or U8584 (N_8584,N_3848,N_3880);
or U8585 (N_8585,N_2234,N_2982);
xor U8586 (N_8586,N_869,N_466);
xor U8587 (N_8587,N_4567,N_3169);
or U8588 (N_8588,N_3076,N_3736);
and U8589 (N_8589,N_1470,N_1995);
nor U8590 (N_8590,N_4596,N_3618);
xnor U8591 (N_8591,N_605,N_2675);
nand U8592 (N_8592,N_4570,N_2868);
nor U8593 (N_8593,N_1723,N_2739);
and U8594 (N_8594,N_796,N_2355);
and U8595 (N_8595,N_4512,N_3185);
or U8596 (N_8596,N_4162,N_4936);
nor U8597 (N_8597,N_3252,N_4661);
xnor U8598 (N_8598,N_3452,N_4299);
xnor U8599 (N_8599,N_3289,N_4478);
nand U8600 (N_8600,N_3518,N_2787);
xor U8601 (N_8601,N_1789,N_2413);
xor U8602 (N_8602,N_2271,N_1665);
and U8603 (N_8603,N_1805,N_4565);
and U8604 (N_8604,N_2163,N_1801);
xor U8605 (N_8605,N_1947,N_4858);
and U8606 (N_8606,N_1546,N_818);
and U8607 (N_8607,N_264,N_4737);
nor U8608 (N_8608,N_857,N_902);
nor U8609 (N_8609,N_3712,N_1734);
xnor U8610 (N_8610,N_371,N_1713);
or U8611 (N_8611,N_4890,N_3986);
xor U8612 (N_8612,N_2271,N_1568);
nor U8613 (N_8613,N_2471,N_1538);
xnor U8614 (N_8614,N_2611,N_3384);
nor U8615 (N_8615,N_1629,N_2768);
nor U8616 (N_8616,N_4703,N_818);
or U8617 (N_8617,N_3551,N_3888);
nand U8618 (N_8618,N_2786,N_4870);
nor U8619 (N_8619,N_414,N_996);
and U8620 (N_8620,N_91,N_256);
nor U8621 (N_8621,N_4712,N_171);
or U8622 (N_8622,N_4040,N_223);
nand U8623 (N_8623,N_676,N_4214);
and U8624 (N_8624,N_3348,N_4733);
and U8625 (N_8625,N_3125,N_2688);
or U8626 (N_8626,N_3145,N_4847);
or U8627 (N_8627,N_3420,N_2060);
nand U8628 (N_8628,N_626,N_2641);
nand U8629 (N_8629,N_3613,N_4764);
or U8630 (N_8630,N_2532,N_1742);
or U8631 (N_8631,N_1464,N_1732);
xor U8632 (N_8632,N_657,N_2662);
and U8633 (N_8633,N_592,N_4742);
nand U8634 (N_8634,N_324,N_4599);
and U8635 (N_8635,N_599,N_3478);
or U8636 (N_8636,N_1454,N_778);
nand U8637 (N_8637,N_64,N_1661);
and U8638 (N_8638,N_532,N_1778);
and U8639 (N_8639,N_1725,N_712);
and U8640 (N_8640,N_4772,N_4610);
nor U8641 (N_8641,N_917,N_1761);
nor U8642 (N_8642,N_4519,N_4650);
or U8643 (N_8643,N_4303,N_3422);
and U8644 (N_8644,N_337,N_3565);
or U8645 (N_8645,N_1655,N_3440);
xor U8646 (N_8646,N_130,N_1063);
nor U8647 (N_8647,N_2545,N_2504);
and U8648 (N_8648,N_4704,N_261);
and U8649 (N_8649,N_4378,N_1013);
xor U8650 (N_8650,N_2348,N_203);
nor U8651 (N_8651,N_4404,N_3918);
nor U8652 (N_8652,N_4618,N_1122);
nand U8653 (N_8653,N_4184,N_2483);
nor U8654 (N_8654,N_4665,N_1634);
nor U8655 (N_8655,N_704,N_4311);
nand U8656 (N_8656,N_3824,N_3762);
nand U8657 (N_8657,N_1394,N_1403);
and U8658 (N_8658,N_2994,N_1699);
xnor U8659 (N_8659,N_1220,N_4817);
nand U8660 (N_8660,N_4071,N_29);
xnor U8661 (N_8661,N_3424,N_2978);
nor U8662 (N_8662,N_2023,N_502);
and U8663 (N_8663,N_2250,N_1583);
and U8664 (N_8664,N_4312,N_1915);
nand U8665 (N_8665,N_3065,N_861);
or U8666 (N_8666,N_2673,N_3353);
and U8667 (N_8667,N_4425,N_733);
xor U8668 (N_8668,N_2095,N_3674);
xor U8669 (N_8669,N_2071,N_2317);
or U8670 (N_8670,N_4680,N_3412);
nand U8671 (N_8671,N_4107,N_703);
nand U8672 (N_8672,N_1173,N_4846);
nand U8673 (N_8673,N_1634,N_2673);
nand U8674 (N_8674,N_2069,N_3176);
or U8675 (N_8675,N_1865,N_3029);
or U8676 (N_8676,N_4519,N_2645);
and U8677 (N_8677,N_359,N_3410);
xnor U8678 (N_8678,N_205,N_4021);
nor U8679 (N_8679,N_1873,N_4587);
and U8680 (N_8680,N_1417,N_970);
or U8681 (N_8681,N_1269,N_2121);
or U8682 (N_8682,N_279,N_4701);
nor U8683 (N_8683,N_737,N_2015);
nor U8684 (N_8684,N_1405,N_1327);
nor U8685 (N_8685,N_3416,N_2074);
nor U8686 (N_8686,N_2113,N_2136);
and U8687 (N_8687,N_3269,N_1404);
or U8688 (N_8688,N_4868,N_3202);
and U8689 (N_8689,N_3100,N_2985);
or U8690 (N_8690,N_2626,N_3690);
or U8691 (N_8691,N_490,N_3556);
or U8692 (N_8692,N_4555,N_3855);
nand U8693 (N_8693,N_2269,N_2254);
nor U8694 (N_8694,N_455,N_2244);
or U8695 (N_8695,N_2423,N_4000);
and U8696 (N_8696,N_2464,N_402);
nand U8697 (N_8697,N_3383,N_4675);
xor U8698 (N_8698,N_2684,N_4811);
and U8699 (N_8699,N_2842,N_4549);
and U8700 (N_8700,N_3054,N_41);
or U8701 (N_8701,N_4464,N_351);
nor U8702 (N_8702,N_1173,N_2951);
nand U8703 (N_8703,N_920,N_2143);
nand U8704 (N_8704,N_3058,N_1929);
nand U8705 (N_8705,N_927,N_2250);
or U8706 (N_8706,N_831,N_2759);
nor U8707 (N_8707,N_4334,N_3442);
or U8708 (N_8708,N_2606,N_2377);
nand U8709 (N_8709,N_187,N_3442);
and U8710 (N_8710,N_211,N_3284);
and U8711 (N_8711,N_3103,N_2380);
xnor U8712 (N_8712,N_4404,N_1631);
nand U8713 (N_8713,N_3163,N_858);
and U8714 (N_8714,N_975,N_4481);
xor U8715 (N_8715,N_3466,N_362);
or U8716 (N_8716,N_1808,N_480);
nor U8717 (N_8717,N_2329,N_2446);
and U8718 (N_8718,N_3762,N_752);
xnor U8719 (N_8719,N_4508,N_4056);
or U8720 (N_8720,N_4119,N_2735);
or U8721 (N_8721,N_2450,N_4509);
nor U8722 (N_8722,N_4031,N_3454);
or U8723 (N_8723,N_487,N_1566);
nor U8724 (N_8724,N_948,N_2155);
nand U8725 (N_8725,N_2584,N_1814);
nor U8726 (N_8726,N_4702,N_1477);
or U8727 (N_8727,N_1529,N_4830);
nor U8728 (N_8728,N_2347,N_4246);
and U8729 (N_8729,N_1878,N_2730);
nor U8730 (N_8730,N_3384,N_4694);
or U8731 (N_8731,N_1447,N_1889);
and U8732 (N_8732,N_2485,N_2403);
nand U8733 (N_8733,N_4056,N_3759);
xor U8734 (N_8734,N_3543,N_2750);
and U8735 (N_8735,N_4737,N_4481);
and U8736 (N_8736,N_2390,N_2566);
xor U8737 (N_8737,N_2685,N_1183);
or U8738 (N_8738,N_2284,N_3628);
or U8739 (N_8739,N_1221,N_3540);
xor U8740 (N_8740,N_4558,N_265);
and U8741 (N_8741,N_4486,N_3980);
xor U8742 (N_8742,N_359,N_869);
xnor U8743 (N_8743,N_775,N_757);
nand U8744 (N_8744,N_283,N_3194);
nand U8745 (N_8745,N_876,N_2758);
or U8746 (N_8746,N_2643,N_1508);
and U8747 (N_8747,N_4397,N_1483);
and U8748 (N_8748,N_2786,N_3520);
or U8749 (N_8749,N_590,N_1185);
and U8750 (N_8750,N_2329,N_615);
xnor U8751 (N_8751,N_2873,N_3782);
or U8752 (N_8752,N_4340,N_782);
nand U8753 (N_8753,N_3955,N_3685);
nor U8754 (N_8754,N_399,N_4381);
xor U8755 (N_8755,N_3494,N_748);
and U8756 (N_8756,N_62,N_2432);
or U8757 (N_8757,N_2188,N_925);
xnor U8758 (N_8758,N_2472,N_4392);
xnor U8759 (N_8759,N_2429,N_147);
nor U8760 (N_8760,N_25,N_4956);
or U8761 (N_8761,N_1832,N_3575);
nand U8762 (N_8762,N_2528,N_2658);
nor U8763 (N_8763,N_3764,N_2482);
nand U8764 (N_8764,N_3063,N_1085);
and U8765 (N_8765,N_1750,N_1046);
or U8766 (N_8766,N_3504,N_4704);
and U8767 (N_8767,N_2492,N_4252);
xor U8768 (N_8768,N_1310,N_2840);
xor U8769 (N_8769,N_2342,N_4026);
and U8770 (N_8770,N_3492,N_2956);
nor U8771 (N_8771,N_860,N_410);
nand U8772 (N_8772,N_350,N_2932);
nand U8773 (N_8773,N_2159,N_4212);
or U8774 (N_8774,N_496,N_1453);
or U8775 (N_8775,N_893,N_1108);
nand U8776 (N_8776,N_4843,N_4281);
xor U8777 (N_8777,N_4112,N_3726);
nand U8778 (N_8778,N_1156,N_65);
xnor U8779 (N_8779,N_195,N_4871);
and U8780 (N_8780,N_3145,N_2098);
and U8781 (N_8781,N_4768,N_227);
or U8782 (N_8782,N_2658,N_3096);
or U8783 (N_8783,N_4749,N_3349);
xor U8784 (N_8784,N_4205,N_2986);
or U8785 (N_8785,N_689,N_1004);
and U8786 (N_8786,N_1975,N_834);
nand U8787 (N_8787,N_4283,N_4197);
nand U8788 (N_8788,N_1193,N_3207);
nor U8789 (N_8789,N_2850,N_4538);
and U8790 (N_8790,N_1985,N_892);
or U8791 (N_8791,N_2121,N_3882);
or U8792 (N_8792,N_506,N_4011);
and U8793 (N_8793,N_142,N_3013);
or U8794 (N_8794,N_412,N_1682);
nor U8795 (N_8795,N_945,N_4193);
nand U8796 (N_8796,N_3180,N_3149);
xnor U8797 (N_8797,N_930,N_1229);
xnor U8798 (N_8798,N_529,N_1317);
xor U8799 (N_8799,N_2087,N_2056);
xnor U8800 (N_8800,N_1352,N_3824);
or U8801 (N_8801,N_2123,N_2762);
nor U8802 (N_8802,N_1156,N_3601);
nand U8803 (N_8803,N_1569,N_678);
nand U8804 (N_8804,N_4116,N_955);
and U8805 (N_8805,N_732,N_3456);
and U8806 (N_8806,N_4687,N_2236);
and U8807 (N_8807,N_488,N_3936);
nand U8808 (N_8808,N_3303,N_1852);
or U8809 (N_8809,N_4900,N_1789);
or U8810 (N_8810,N_1144,N_3058);
nand U8811 (N_8811,N_1735,N_3804);
nand U8812 (N_8812,N_3422,N_869);
and U8813 (N_8813,N_3619,N_4606);
or U8814 (N_8814,N_4484,N_960);
xnor U8815 (N_8815,N_4869,N_2792);
or U8816 (N_8816,N_1199,N_657);
and U8817 (N_8817,N_2289,N_4026);
or U8818 (N_8818,N_472,N_2543);
and U8819 (N_8819,N_4540,N_312);
nor U8820 (N_8820,N_3851,N_1696);
and U8821 (N_8821,N_2101,N_3890);
and U8822 (N_8822,N_56,N_2144);
nor U8823 (N_8823,N_823,N_2078);
or U8824 (N_8824,N_4472,N_3555);
xor U8825 (N_8825,N_2447,N_1556);
xnor U8826 (N_8826,N_4266,N_3542);
nor U8827 (N_8827,N_432,N_554);
nand U8828 (N_8828,N_2059,N_4299);
xnor U8829 (N_8829,N_4967,N_420);
or U8830 (N_8830,N_4222,N_4445);
xor U8831 (N_8831,N_4541,N_3120);
xnor U8832 (N_8832,N_1848,N_4044);
and U8833 (N_8833,N_2768,N_3654);
xor U8834 (N_8834,N_2424,N_1441);
nand U8835 (N_8835,N_4794,N_681);
nand U8836 (N_8836,N_330,N_1836);
nand U8837 (N_8837,N_3944,N_4950);
nand U8838 (N_8838,N_3858,N_2419);
or U8839 (N_8839,N_1406,N_4056);
nand U8840 (N_8840,N_1306,N_3558);
nand U8841 (N_8841,N_171,N_2697);
and U8842 (N_8842,N_486,N_3808);
and U8843 (N_8843,N_3232,N_682);
or U8844 (N_8844,N_1324,N_2965);
nor U8845 (N_8845,N_3232,N_3541);
and U8846 (N_8846,N_498,N_1397);
xor U8847 (N_8847,N_4733,N_1638);
xnor U8848 (N_8848,N_4667,N_3351);
and U8849 (N_8849,N_845,N_3774);
xnor U8850 (N_8850,N_3091,N_328);
nor U8851 (N_8851,N_2399,N_4586);
nand U8852 (N_8852,N_3055,N_2181);
and U8853 (N_8853,N_1026,N_3362);
xnor U8854 (N_8854,N_3364,N_2271);
nand U8855 (N_8855,N_4295,N_3056);
and U8856 (N_8856,N_2624,N_2603);
nand U8857 (N_8857,N_2944,N_2734);
and U8858 (N_8858,N_39,N_1518);
nor U8859 (N_8859,N_3594,N_3909);
nor U8860 (N_8860,N_2805,N_3225);
or U8861 (N_8861,N_3234,N_608);
nand U8862 (N_8862,N_37,N_3106);
nor U8863 (N_8863,N_2216,N_4983);
nand U8864 (N_8864,N_4919,N_4746);
and U8865 (N_8865,N_468,N_1305);
and U8866 (N_8866,N_699,N_1608);
nor U8867 (N_8867,N_2218,N_217);
or U8868 (N_8868,N_3484,N_3957);
or U8869 (N_8869,N_399,N_595);
or U8870 (N_8870,N_510,N_3696);
or U8871 (N_8871,N_2779,N_4756);
nand U8872 (N_8872,N_4253,N_355);
xnor U8873 (N_8873,N_185,N_1402);
xor U8874 (N_8874,N_3793,N_1774);
or U8875 (N_8875,N_3751,N_4862);
nand U8876 (N_8876,N_549,N_4374);
or U8877 (N_8877,N_2242,N_361);
and U8878 (N_8878,N_4594,N_992);
nand U8879 (N_8879,N_4334,N_3578);
xor U8880 (N_8880,N_2364,N_4656);
xnor U8881 (N_8881,N_463,N_2483);
nor U8882 (N_8882,N_4854,N_3883);
nor U8883 (N_8883,N_161,N_4492);
nand U8884 (N_8884,N_3931,N_3596);
nand U8885 (N_8885,N_1453,N_3214);
nor U8886 (N_8886,N_129,N_2144);
xor U8887 (N_8887,N_24,N_2416);
nand U8888 (N_8888,N_3416,N_3365);
and U8889 (N_8889,N_2235,N_4637);
or U8890 (N_8890,N_2939,N_4109);
and U8891 (N_8891,N_352,N_4153);
or U8892 (N_8892,N_3448,N_3507);
or U8893 (N_8893,N_588,N_4198);
or U8894 (N_8894,N_612,N_2917);
xnor U8895 (N_8895,N_2437,N_2081);
nand U8896 (N_8896,N_2226,N_2796);
nand U8897 (N_8897,N_3033,N_725);
and U8898 (N_8898,N_2175,N_3653);
nor U8899 (N_8899,N_1373,N_449);
and U8900 (N_8900,N_1140,N_2849);
nand U8901 (N_8901,N_615,N_2356);
and U8902 (N_8902,N_4792,N_1519);
or U8903 (N_8903,N_1509,N_2250);
nor U8904 (N_8904,N_2348,N_1803);
xor U8905 (N_8905,N_1807,N_376);
nor U8906 (N_8906,N_4984,N_4670);
or U8907 (N_8907,N_1885,N_813);
nor U8908 (N_8908,N_496,N_2762);
xor U8909 (N_8909,N_4199,N_2244);
nand U8910 (N_8910,N_2062,N_1215);
or U8911 (N_8911,N_2498,N_965);
nor U8912 (N_8912,N_4835,N_1853);
xnor U8913 (N_8913,N_3492,N_4583);
nor U8914 (N_8914,N_4828,N_2435);
and U8915 (N_8915,N_3224,N_4985);
xor U8916 (N_8916,N_3209,N_667);
nand U8917 (N_8917,N_1754,N_2445);
xor U8918 (N_8918,N_2631,N_2766);
nor U8919 (N_8919,N_3513,N_3982);
nand U8920 (N_8920,N_4924,N_3077);
xor U8921 (N_8921,N_3663,N_1787);
xnor U8922 (N_8922,N_4197,N_4589);
nor U8923 (N_8923,N_1349,N_4793);
or U8924 (N_8924,N_1796,N_451);
and U8925 (N_8925,N_3186,N_4448);
xnor U8926 (N_8926,N_3843,N_1348);
xnor U8927 (N_8927,N_1546,N_4461);
nor U8928 (N_8928,N_1719,N_4461);
nor U8929 (N_8929,N_4989,N_3465);
xnor U8930 (N_8930,N_4759,N_4998);
xor U8931 (N_8931,N_47,N_2073);
xor U8932 (N_8932,N_188,N_1489);
or U8933 (N_8933,N_2586,N_4546);
xor U8934 (N_8934,N_4171,N_97);
and U8935 (N_8935,N_4447,N_4939);
nand U8936 (N_8936,N_757,N_3661);
and U8937 (N_8937,N_2686,N_2716);
or U8938 (N_8938,N_2754,N_4628);
nand U8939 (N_8939,N_4760,N_3527);
nand U8940 (N_8940,N_785,N_200);
or U8941 (N_8941,N_3668,N_4647);
nand U8942 (N_8942,N_2971,N_3506);
nor U8943 (N_8943,N_2042,N_2220);
and U8944 (N_8944,N_2592,N_564);
or U8945 (N_8945,N_612,N_3707);
or U8946 (N_8946,N_193,N_937);
nor U8947 (N_8947,N_4069,N_3433);
xor U8948 (N_8948,N_292,N_712);
and U8949 (N_8949,N_3654,N_522);
or U8950 (N_8950,N_511,N_1880);
nor U8951 (N_8951,N_2417,N_1003);
nand U8952 (N_8952,N_1775,N_1949);
and U8953 (N_8953,N_2213,N_4761);
xor U8954 (N_8954,N_3264,N_2858);
nand U8955 (N_8955,N_2143,N_2001);
xor U8956 (N_8956,N_3529,N_3221);
or U8957 (N_8957,N_4528,N_1368);
xnor U8958 (N_8958,N_3502,N_1240);
nor U8959 (N_8959,N_278,N_1997);
xor U8960 (N_8960,N_2274,N_4574);
and U8961 (N_8961,N_130,N_1435);
or U8962 (N_8962,N_3092,N_2617);
and U8963 (N_8963,N_448,N_3361);
or U8964 (N_8964,N_3132,N_4640);
xor U8965 (N_8965,N_4164,N_3398);
nand U8966 (N_8966,N_2038,N_3747);
or U8967 (N_8967,N_1881,N_3283);
xnor U8968 (N_8968,N_701,N_3526);
and U8969 (N_8969,N_3124,N_1552);
xor U8970 (N_8970,N_4506,N_3716);
and U8971 (N_8971,N_3580,N_167);
or U8972 (N_8972,N_2618,N_3166);
xor U8973 (N_8973,N_3096,N_1563);
nand U8974 (N_8974,N_3007,N_204);
and U8975 (N_8975,N_1283,N_2608);
and U8976 (N_8976,N_4782,N_4528);
or U8977 (N_8977,N_4743,N_3440);
xor U8978 (N_8978,N_2070,N_420);
nand U8979 (N_8979,N_2813,N_3692);
and U8980 (N_8980,N_1565,N_2642);
nor U8981 (N_8981,N_1338,N_4981);
nor U8982 (N_8982,N_4857,N_1097);
nor U8983 (N_8983,N_995,N_2504);
nand U8984 (N_8984,N_1887,N_4026);
or U8985 (N_8985,N_1830,N_3565);
and U8986 (N_8986,N_1474,N_3744);
nor U8987 (N_8987,N_1199,N_2293);
xor U8988 (N_8988,N_2479,N_2879);
nor U8989 (N_8989,N_2055,N_2068);
nand U8990 (N_8990,N_1993,N_3918);
nor U8991 (N_8991,N_531,N_3615);
or U8992 (N_8992,N_897,N_2286);
and U8993 (N_8993,N_2629,N_2326);
nor U8994 (N_8994,N_3437,N_562);
and U8995 (N_8995,N_1036,N_176);
nor U8996 (N_8996,N_3337,N_4834);
and U8997 (N_8997,N_859,N_3201);
or U8998 (N_8998,N_4438,N_363);
nor U8999 (N_8999,N_2856,N_3329);
xor U9000 (N_9000,N_3459,N_970);
nor U9001 (N_9001,N_4124,N_4927);
nand U9002 (N_9002,N_4781,N_3286);
or U9003 (N_9003,N_3726,N_635);
nand U9004 (N_9004,N_3002,N_1102);
or U9005 (N_9005,N_114,N_341);
or U9006 (N_9006,N_2137,N_3087);
nand U9007 (N_9007,N_2730,N_2010);
and U9008 (N_9008,N_2345,N_4380);
and U9009 (N_9009,N_3313,N_1673);
nor U9010 (N_9010,N_2139,N_482);
xor U9011 (N_9011,N_547,N_2887);
or U9012 (N_9012,N_2451,N_4094);
nor U9013 (N_9013,N_488,N_2911);
xor U9014 (N_9014,N_4884,N_144);
nor U9015 (N_9015,N_1423,N_420);
xnor U9016 (N_9016,N_1494,N_2984);
xnor U9017 (N_9017,N_487,N_3231);
nand U9018 (N_9018,N_3562,N_1077);
xor U9019 (N_9019,N_1229,N_986);
or U9020 (N_9020,N_3710,N_1584);
nand U9021 (N_9021,N_236,N_3680);
and U9022 (N_9022,N_1229,N_4432);
nand U9023 (N_9023,N_4830,N_1153);
xnor U9024 (N_9024,N_3182,N_3120);
xor U9025 (N_9025,N_769,N_248);
or U9026 (N_9026,N_149,N_76);
xor U9027 (N_9027,N_1317,N_2994);
and U9028 (N_9028,N_2755,N_2027);
xnor U9029 (N_9029,N_3599,N_3275);
xor U9030 (N_9030,N_4998,N_3498);
nor U9031 (N_9031,N_2859,N_1727);
nor U9032 (N_9032,N_1728,N_4265);
nand U9033 (N_9033,N_1122,N_4213);
nor U9034 (N_9034,N_1085,N_4928);
and U9035 (N_9035,N_4358,N_229);
nor U9036 (N_9036,N_2420,N_4257);
nand U9037 (N_9037,N_2461,N_991);
and U9038 (N_9038,N_3529,N_4732);
nor U9039 (N_9039,N_4224,N_4914);
nor U9040 (N_9040,N_1271,N_1506);
xnor U9041 (N_9041,N_1595,N_4901);
nor U9042 (N_9042,N_2628,N_1493);
and U9043 (N_9043,N_4194,N_2077);
xor U9044 (N_9044,N_427,N_3388);
and U9045 (N_9045,N_1997,N_655);
or U9046 (N_9046,N_3788,N_375);
and U9047 (N_9047,N_3595,N_4029);
nor U9048 (N_9048,N_3458,N_862);
nor U9049 (N_9049,N_2259,N_3180);
or U9050 (N_9050,N_1407,N_2491);
or U9051 (N_9051,N_2839,N_3732);
and U9052 (N_9052,N_3210,N_1975);
and U9053 (N_9053,N_3492,N_4351);
nor U9054 (N_9054,N_1761,N_2676);
or U9055 (N_9055,N_1987,N_1164);
or U9056 (N_9056,N_1303,N_3990);
and U9057 (N_9057,N_3407,N_4479);
and U9058 (N_9058,N_1187,N_525);
and U9059 (N_9059,N_4149,N_3505);
nand U9060 (N_9060,N_4178,N_1474);
and U9061 (N_9061,N_1497,N_636);
nand U9062 (N_9062,N_1643,N_1112);
nand U9063 (N_9063,N_2525,N_4157);
xor U9064 (N_9064,N_3926,N_4213);
nand U9065 (N_9065,N_4578,N_3810);
or U9066 (N_9066,N_2698,N_772);
or U9067 (N_9067,N_2344,N_1498);
xnor U9068 (N_9068,N_4813,N_3937);
and U9069 (N_9069,N_1079,N_1097);
or U9070 (N_9070,N_2226,N_778);
xnor U9071 (N_9071,N_550,N_1633);
nor U9072 (N_9072,N_4382,N_1484);
nor U9073 (N_9073,N_4631,N_1497);
nand U9074 (N_9074,N_477,N_1826);
nand U9075 (N_9075,N_2195,N_110);
xnor U9076 (N_9076,N_3403,N_579);
or U9077 (N_9077,N_2599,N_3647);
nor U9078 (N_9078,N_112,N_2193);
nor U9079 (N_9079,N_1078,N_333);
or U9080 (N_9080,N_4916,N_4661);
nand U9081 (N_9081,N_303,N_1259);
nand U9082 (N_9082,N_3579,N_987);
xor U9083 (N_9083,N_2849,N_3292);
or U9084 (N_9084,N_2156,N_1717);
nor U9085 (N_9085,N_4744,N_1743);
xor U9086 (N_9086,N_3514,N_3838);
nor U9087 (N_9087,N_849,N_1558);
or U9088 (N_9088,N_289,N_397);
and U9089 (N_9089,N_1858,N_4186);
or U9090 (N_9090,N_360,N_1816);
nand U9091 (N_9091,N_2609,N_950);
and U9092 (N_9092,N_596,N_2213);
nand U9093 (N_9093,N_2116,N_2978);
or U9094 (N_9094,N_4940,N_448);
nand U9095 (N_9095,N_3787,N_4774);
nand U9096 (N_9096,N_1235,N_1370);
nand U9097 (N_9097,N_2517,N_1826);
nand U9098 (N_9098,N_4842,N_4321);
xnor U9099 (N_9099,N_4344,N_2059);
and U9100 (N_9100,N_1393,N_1253);
or U9101 (N_9101,N_4517,N_4073);
nor U9102 (N_9102,N_3857,N_2682);
nor U9103 (N_9103,N_126,N_972);
nand U9104 (N_9104,N_4149,N_149);
xnor U9105 (N_9105,N_711,N_172);
xnor U9106 (N_9106,N_3166,N_3554);
nor U9107 (N_9107,N_35,N_2653);
and U9108 (N_9108,N_4210,N_3109);
nor U9109 (N_9109,N_3641,N_2705);
xnor U9110 (N_9110,N_979,N_4018);
or U9111 (N_9111,N_3261,N_4114);
and U9112 (N_9112,N_1138,N_2365);
and U9113 (N_9113,N_715,N_937);
or U9114 (N_9114,N_627,N_315);
and U9115 (N_9115,N_905,N_2583);
and U9116 (N_9116,N_2674,N_3041);
nand U9117 (N_9117,N_2359,N_2155);
nor U9118 (N_9118,N_4896,N_104);
nor U9119 (N_9119,N_3517,N_775);
nand U9120 (N_9120,N_2520,N_3816);
xor U9121 (N_9121,N_2470,N_3141);
or U9122 (N_9122,N_868,N_4903);
nor U9123 (N_9123,N_3984,N_2814);
or U9124 (N_9124,N_303,N_177);
or U9125 (N_9125,N_1917,N_1707);
or U9126 (N_9126,N_1150,N_4011);
nand U9127 (N_9127,N_570,N_3154);
and U9128 (N_9128,N_2719,N_3522);
and U9129 (N_9129,N_2392,N_3744);
xor U9130 (N_9130,N_423,N_2480);
xor U9131 (N_9131,N_4378,N_1028);
xor U9132 (N_9132,N_1646,N_2210);
and U9133 (N_9133,N_1609,N_4867);
and U9134 (N_9134,N_1657,N_3338);
xor U9135 (N_9135,N_2149,N_3499);
or U9136 (N_9136,N_1863,N_4470);
or U9137 (N_9137,N_2931,N_2258);
xor U9138 (N_9138,N_1499,N_2055);
nor U9139 (N_9139,N_1095,N_4517);
and U9140 (N_9140,N_1637,N_3639);
xor U9141 (N_9141,N_3950,N_2588);
and U9142 (N_9142,N_234,N_2645);
xnor U9143 (N_9143,N_3509,N_3991);
and U9144 (N_9144,N_1391,N_2372);
nand U9145 (N_9145,N_3100,N_2544);
and U9146 (N_9146,N_3015,N_3001);
nor U9147 (N_9147,N_1156,N_2752);
nand U9148 (N_9148,N_695,N_4563);
nor U9149 (N_9149,N_715,N_4232);
nand U9150 (N_9150,N_2697,N_4619);
nor U9151 (N_9151,N_392,N_4314);
and U9152 (N_9152,N_2452,N_2461);
nor U9153 (N_9153,N_444,N_4396);
nor U9154 (N_9154,N_2055,N_72);
and U9155 (N_9155,N_3758,N_1507);
or U9156 (N_9156,N_1507,N_1519);
or U9157 (N_9157,N_1237,N_4994);
nor U9158 (N_9158,N_2103,N_1966);
or U9159 (N_9159,N_3482,N_2399);
xnor U9160 (N_9160,N_580,N_3859);
xnor U9161 (N_9161,N_4772,N_3463);
or U9162 (N_9162,N_1320,N_4580);
xor U9163 (N_9163,N_4623,N_2031);
and U9164 (N_9164,N_193,N_1295);
nand U9165 (N_9165,N_3970,N_2718);
xor U9166 (N_9166,N_4597,N_2625);
xnor U9167 (N_9167,N_1132,N_4237);
or U9168 (N_9168,N_1623,N_79);
and U9169 (N_9169,N_629,N_3263);
xor U9170 (N_9170,N_3352,N_1068);
nand U9171 (N_9171,N_712,N_3578);
nand U9172 (N_9172,N_3945,N_2195);
xor U9173 (N_9173,N_996,N_1676);
xnor U9174 (N_9174,N_3536,N_3741);
xnor U9175 (N_9175,N_2652,N_1797);
and U9176 (N_9176,N_211,N_4654);
or U9177 (N_9177,N_891,N_1515);
and U9178 (N_9178,N_96,N_1522);
and U9179 (N_9179,N_1630,N_1032);
or U9180 (N_9180,N_3713,N_4740);
and U9181 (N_9181,N_540,N_118);
nand U9182 (N_9182,N_4622,N_3521);
nor U9183 (N_9183,N_700,N_4215);
nand U9184 (N_9184,N_801,N_3478);
or U9185 (N_9185,N_2345,N_862);
nand U9186 (N_9186,N_2191,N_191);
and U9187 (N_9187,N_595,N_2734);
and U9188 (N_9188,N_2073,N_2380);
nor U9189 (N_9189,N_3274,N_1936);
nand U9190 (N_9190,N_4337,N_3961);
nor U9191 (N_9191,N_4441,N_335);
nor U9192 (N_9192,N_1856,N_2308);
nor U9193 (N_9193,N_1378,N_2934);
nor U9194 (N_9194,N_2079,N_4735);
and U9195 (N_9195,N_3886,N_2765);
and U9196 (N_9196,N_1869,N_4564);
or U9197 (N_9197,N_4314,N_620);
nor U9198 (N_9198,N_4660,N_2487);
or U9199 (N_9199,N_1985,N_1846);
nand U9200 (N_9200,N_2338,N_3476);
and U9201 (N_9201,N_2699,N_3063);
nor U9202 (N_9202,N_4349,N_1605);
nor U9203 (N_9203,N_3520,N_2329);
and U9204 (N_9204,N_3094,N_1828);
or U9205 (N_9205,N_1535,N_3355);
xnor U9206 (N_9206,N_2265,N_2303);
nand U9207 (N_9207,N_3859,N_3520);
or U9208 (N_9208,N_4903,N_2540);
nand U9209 (N_9209,N_886,N_2931);
xnor U9210 (N_9210,N_1298,N_2644);
xor U9211 (N_9211,N_1136,N_480);
or U9212 (N_9212,N_1779,N_2910);
nand U9213 (N_9213,N_3109,N_1704);
nor U9214 (N_9214,N_1148,N_3237);
nor U9215 (N_9215,N_1351,N_3030);
or U9216 (N_9216,N_836,N_550);
or U9217 (N_9217,N_919,N_627);
or U9218 (N_9218,N_3640,N_2498);
or U9219 (N_9219,N_202,N_337);
or U9220 (N_9220,N_3626,N_3647);
or U9221 (N_9221,N_3090,N_3206);
or U9222 (N_9222,N_1692,N_4644);
xnor U9223 (N_9223,N_1549,N_3598);
xnor U9224 (N_9224,N_3547,N_3132);
xor U9225 (N_9225,N_1901,N_3666);
or U9226 (N_9226,N_253,N_3907);
nand U9227 (N_9227,N_2244,N_892);
and U9228 (N_9228,N_345,N_3954);
nor U9229 (N_9229,N_3263,N_3365);
nand U9230 (N_9230,N_1842,N_2990);
or U9231 (N_9231,N_689,N_1901);
or U9232 (N_9232,N_334,N_3373);
nand U9233 (N_9233,N_4769,N_2677);
xor U9234 (N_9234,N_4218,N_1014);
nor U9235 (N_9235,N_1200,N_4766);
xnor U9236 (N_9236,N_462,N_1640);
or U9237 (N_9237,N_3307,N_2143);
xor U9238 (N_9238,N_1966,N_3368);
nor U9239 (N_9239,N_3681,N_2395);
nand U9240 (N_9240,N_4003,N_1226);
nor U9241 (N_9241,N_1631,N_1156);
or U9242 (N_9242,N_4000,N_2748);
and U9243 (N_9243,N_4462,N_384);
xor U9244 (N_9244,N_3139,N_283);
nand U9245 (N_9245,N_419,N_3114);
xnor U9246 (N_9246,N_2569,N_633);
nand U9247 (N_9247,N_1911,N_2477);
nor U9248 (N_9248,N_537,N_1339);
or U9249 (N_9249,N_1632,N_2856);
and U9250 (N_9250,N_40,N_231);
nand U9251 (N_9251,N_1164,N_1547);
nor U9252 (N_9252,N_2716,N_637);
or U9253 (N_9253,N_2312,N_1445);
nor U9254 (N_9254,N_1421,N_2734);
and U9255 (N_9255,N_86,N_1734);
nor U9256 (N_9256,N_1350,N_2734);
nor U9257 (N_9257,N_1977,N_811);
or U9258 (N_9258,N_1573,N_2054);
and U9259 (N_9259,N_1202,N_1538);
nor U9260 (N_9260,N_2297,N_3052);
nor U9261 (N_9261,N_1911,N_4535);
xnor U9262 (N_9262,N_2708,N_2728);
xnor U9263 (N_9263,N_495,N_1401);
xnor U9264 (N_9264,N_415,N_480);
xnor U9265 (N_9265,N_4703,N_1062);
or U9266 (N_9266,N_4658,N_820);
nor U9267 (N_9267,N_1673,N_1200);
nand U9268 (N_9268,N_255,N_3760);
nor U9269 (N_9269,N_755,N_3359);
nor U9270 (N_9270,N_2820,N_1295);
nor U9271 (N_9271,N_2686,N_4098);
nand U9272 (N_9272,N_1179,N_866);
nor U9273 (N_9273,N_3255,N_1372);
xnor U9274 (N_9274,N_2718,N_996);
and U9275 (N_9275,N_1684,N_2629);
xnor U9276 (N_9276,N_2842,N_2136);
nand U9277 (N_9277,N_243,N_2937);
nor U9278 (N_9278,N_582,N_1563);
nand U9279 (N_9279,N_3910,N_4763);
and U9280 (N_9280,N_2307,N_1204);
xor U9281 (N_9281,N_3004,N_3138);
xnor U9282 (N_9282,N_4360,N_1549);
xnor U9283 (N_9283,N_3156,N_4403);
nand U9284 (N_9284,N_35,N_3357);
nor U9285 (N_9285,N_1870,N_3095);
nand U9286 (N_9286,N_427,N_4143);
or U9287 (N_9287,N_2208,N_2032);
nand U9288 (N_9288,N_3637,N_4658);
and U9289 (N_9289,N_1685,N_4867);
nand U9290 (N_9290,N_3302,N_1703);
or U9291 (N_9291,N_1240,N_2041);
nor U9292 (N_9292,N_3727,N_4420);
xor U9293 (N_9293,N_4268,N_2550);
and U9294 (N_9294,N_4819,N_2525);
xor U9295 (N_9295,N_819,N_209);
nand U9296 (N_9296,N_4810,N_990);
and U9297 (N_9297,N_2576,N_1805);
and U9298 (N_9298,N_2802,N_3255);
and U9299 (N_9299,N_718,N_2832);
nor U9300 (N_9300,N_1332,N_4307);
xnor U9301 (N_9301,N_1426,N_3649);
nand U9302 (N_9302,N_1753,N_56);
nand U9303 (N_9303,N_1928,N_1696);
or U9304 (N_9304,N_3511,N_2081);
or U9305 (N_9305,N_4647,N_3840);
and U9306 (N_9306,N_3542,N_4822);
nand U9307 (N_9307,N_3379,N_4585);
and U9308 (N_9308,N_1673,N_788);
nor U9309 (N_9309,N_4106,N_2356);
or U9310 (N_9310,N_3496,N_4866);
or U9311 (N_9311,N_2187,N_2900);
nor U9312 (N_9312,N_89,N_1651);
xor U9313 (N_9313,N_4323,N_1513);
or U9314 (N_9314,N_3502,N_933);
xor U9315 (N_9315,N_954,N_4147);
nor U9316 (N_9316,N_937,N_3751);
nand U9317 (N_9317,N_4382,N_3254);
or U9318 (N_9318,N_3864,N_3260);
xor U9319 (N_9319,N_4554,N_1493);
and U9320 (N_9320,N_3975,N_2583);
nand U9321 (N_9321,N_1755,N_2930);
nand U9322 (N_9322,N_4480,N_1346);
nand U9323 (N_9323,N_3475,N_2180);
nor U9324 (N_9324,N_352,N_1782);
xnor U9325 (N_9325,N_2319,N_3069);
or U9326 (N_9326,N_3598,N_1842);
nand U9327 (N_9327,N_961,N_1969);
or U9328 (N_9328,N_629,N_4499);
and U9329 (N_9329,N_2320,N_1932);
and U9330 (N_9330,N_1064,N_412);
and U9331 (N_9331,N_890,N_4619);
and U9332 (N_9332,N_1150,N_2929);
nor U9333 (N_9333,N_3278,N_118);
or U9334 (N_9334,N_2574,N_4737);
nand U9335 (N_9335,N_3499,N_3534);
nand U9336 (N_9336,N_213,N_3613);
nand U9337 (N_9337,N_1403,N_3867);
or U9338 (N_9338,N_2039,N_1787);
nor U9339 (N_9339,N_2525,N_3507);
nor U9340 (N_9340,N_831,N_2082);
or U9341 (N_9341,N_2208,N_4325);
or U9342 (N_9342,N_3911,N_237);
or U9343 (N_9343,N_221,N_2692);
xnor U9344 (N_9344,N_4775,N_1653);
nor U9345 (N_9345,N_3103,N_3576);
or U9346 (N_9346,N_1746,N_360);
or U9347 (N_9347,N_2942,N_1902);
nand U9348 (N_9348,N_1681,N_1125);
and U9349 (N_9349,N_753,N_1461);
nor U9350 (N_9350,N_925,N_61);
nor U9351 (N_9351,N_2044,N_4618);
nand U9352 (N_9352,N_732,N_1831);
or U9353 (N_9353,N_2583,N_3937);
and U9354 (N_9354,N_3513,N_2438);
xor U9355 (N_9355,N_2267,N_4257);
xor U9356 (N_9356,N_1354,N_940);
nor U9357 (N_9357,N_916,N_3313);
or U9358 (N_9358,N_3472,N_1700);
nor U9359 (N_9359,N_4480,N_263);
and U9360 (N_9360,N_4266,N_3201);
or U9361 (N_9361,N_3022,N_322);
or U9362 (N_9362,N_338,N_3604);
xor U9363 (N_9363,N_1067,N_258);
xnor U9364 (N_9364,N_3453,N_3952);
nor U9365 (N_9365,N_3334,N_4661);
xnor U9366 (N_9366,N_557,N_3100);
or U9367 (N_9367,N_1737,N_3731);
nor U9368 (N_9368,N_294,N_3125);
or U9369 (N_9369,N_1992,N_4478);
and U9370 (N_9370,N_704,N_1263);
xor U9371 (N_9371,N_1847,N_4319);
and U9372 (N_9372,N_4045,N_2509);
or U9373 (N_9373,N_965,N_1730);
and U9374 (N_9374,N_3579,N_2788);
nor U9375 (N_9375,N_258,N_225);
or U9376 (N_9376,N_4546,N_249);
or U9377 (N_9377,N_1656,N_4946);
nor U9378 (N_9378,N_2503,N_4105);
xnor U9379 (N_9379,N_2990,N_3622);
xor U9380 (N_9380,N_2728,N_1984);
nand U9381 (N_9381,N_2636,N_1644);
nand U9382 (N_9382,N_3621,N_2208);
or U9383 (N_9383,N_1893,N_4859);
nor U9384 (N_9384,N_3052,N_635);
nor U9385 (N_9385,N_4699,N_4787);
xnor U9386 (N_9386,N_2548,N_4720);
nor U9387 (N_9387,N_4390,N_1451);
and U9388 (N_9388,N_894,N_1086);
or U9389 (N_9389,N_3876,N_2967);
xnor U9390 (N_9390,N_1064,N_1954);
xor U9391 (N_9391,N_1730,N_1182);
nor U9392 (N_9392,N_1734,N_4470);
nor U9393 (N_9393,N_3508,N_3505);
nor U9394 (N_9394,N_3807,N_4057);
xnor U9395 (N_9395,N_3451,N_4284);
nor U9396 (N_9396,N_3056,N_100);
and U9397 (N_9397,N_1708,N_108);
xor U9398 (N_9398,N_2953,N_4797);
xor U9399 (N_9399,N_3649,N_3206);
nor U9400 (N_9400,N_2075,N_4432);
xor U9401 (N_9401,N_1611,N_3516);
or U9402 (N_9402,N_3575,N_742);
nand U9403 (N_9403,N_4733,N_3821);
or U9404 (N_9404,N_814,N_3109);
and U9405 (N_9405,N_3330,N_1364);
and U9406 (N_9406,N_2848,N_1858);
nor U9407 (N_9407,N_4752,N_1411);
or U9408 (N_9408,N_1309,N_647);
nand U9409 (N_9409,N_2353,N_2287);
or U9410 (N_9410,N_1657,N_3637);
or U9411 (N_9411,N_2043,N_1397);
nor U9412 (N_9412,N_148,N_179);
nand U9413 (N_9413,N_20,N_1578);
nor U9414 (N_9414,N_4920,N_2659);
nand U9415 (N_9415,N_1470,N_784);
xnor U9416 (N_9416,N_4189,N_2932);
xor U9417 (N_9417,N_1933,N_1873);
nor U9418 (N_9418,N_4735,N_75);
and U9419 (N_9419,N_430,N_4400);
nand U9420 (N_9420,N_981,N_255);
or U9421 (N_9421,N_3859,N_3561);
nand U9422 (N_9422,N_2397,N_4537);
and U9423 (N_9423,N_4997,N_4223);
nand U9424 (N_9424,N_1043,N_3446);
nand U9425 (N_9425,N_1707,N_4533);
and U9426 (N_9426,N_3830,N_651);
or U9427 (N_9427,N_3353,N_3670);
or U9428 (N_9428,N_4365,N_420);
and U9429 (N_9429,N_1706,N_1462);
nor U9430 (N_9430,N_3635,N_1506);
or U9431 (N_9431,N_3563,N_3310);
and U9432 (N_9432,N_4082,N_1867);
or U9433 (N_9433,N_1091,N_2686);
nor U9434 (N_9434,N_4871,N_3891);
xnor U9435 (N_9435,N_1277,N_4705);
and U9436 (N_9436,N_4275,N_2227);
and U9437 (N_9437,N_449,N_461);
xnor U9438 (N_9438,N_2265,N_4659);
or U9439 (N_9439,N_1289,N_1410);
or U9440 (N_9440,N_2681,N_1748);
nor U9441 (N_9441,N_642,N_3202);
xnor U9442 (N_9442,N_3050,N_1708);
or U9443 (N_9443,N_2795,N_3848);
nand U9444 (N_9444,N_2539,N_1117);
and U9445 (N_9445,N_2602,N_2523);
or U9446 (N_9446,N_2477,N_2379);
nor U9447 (N_9447,N_495,N_3355);
nand U9448 (N_9448,N_3387,N_2955);
or U9449 (N_9449,N_4247,N_748);
or U9450 (N_9450,N_3497,N_904);
and U9451 (N_9451,N_4367,N_1546);
and U9452 (N_9452,N_948,N_4480);
or U9453 (N_9453,N_2803,N_2057);
xnor U9454 (N_9454,N_4480,N_1189);
and U9455 (N_9455,N_2182,N_4653);
and U9456 (N_9456,N_4519,N_475);
or U9457 (N_9457,N_4748,N_2690);
nor U9458 (N_9458,N_2938,N_4576);
xnor U9459 (N_9459,N_127,N_1001);
or U9460 (N_9460,N_4162,N_4934);
and U9461 (N_9461,N_4901,N_2514);
nor U9462 (N_9462,N_509,N_4854);
xor U9463 (N_9463,N_648,N_2945);
nand U9464 (N_9464,N_1319,N_2859);
xor U9465 (N_9465,N_1833,N_4654);
xor U9466 (N_9466,N_1061,N_1590);
nand U9467 (N_9467,N_4958,N_483);
nand U9468 (N_9468,N_1604,N_2115);
xor U9469 (N_9469,N_3515,N_2247);
and U9470 (N_9470,N_511,N_704);
nor U9471 (N_9471,N_3130,N_824);
nor U9472 (N_9472,N_1990,N_4213);
nand U9473 (N_9473,N_2694,N_3164);
or U9474 (N_9474,N_4241,N_2822);
and U9475 (N_9475,N_623,N_4936);
nand U9476 (N_9476,N_387,N_909);
or U9477 (N_9477,N_2709,N_3588);
or U9478 (N_9478,N_4399,N_4161);
xor U9479 (N_9479,N_3813,N_1369);
xnor U9480 (N_9480,N_1503,N_611);
nor U9481 (N_9481,N_2850,N_2834);
and U9482 (N_9482,N_50,N_2607);
nor U9483 (N_9483,N_4379,N_3815);
or U9484 (N_9484,N_2112,N_2710);
xor U9485 (N_9485,N_2678,N_1949);
nor U9486 (N_9486,N_3899,N_4062);
xor U9487 (N_9487,N_519,N_2987);
nor U9488 (N_9488,N_1723,N_1373);
nor U9489 (N_9489,N_2869,N_46);
nand U9490 (N_9490,N_2067,N_3673);
xnor U9491 (N_9491,N_2397,N_2322);
nor U9492 (N_9492,N_1476,N_1001);
or U9493 (N_9493,N_3097,N_4056);
nor U9494 (N_9494,N_602,N_3041);
and U9495 (N_9495,N_2599,N_2174);
and U9496 (N_9496,N_3886,N_4655);
nor U9497 (N_9497,N_4184,N_304);
nand U9498 (N_9498,N_3203,N_1348);
or U9499 (N_9499,N_2206,N_1850);
and U9500 (N_9500,N_4414,N_4821);
or U9501 (N_9501,N_1916,N_496);
or U9502 (N_9502,N_4547,N_1524);
nand U9503 (N_9503,N_4660,N_207);
or U9504 (N_9504,N_2154,N_4956);
nor U9505 (N_9505,N_2163,N_3336);
or U9506 (N_9506,N_1167,N_263);
nor U9507 (N_9507,N_4307,N_946);
or U9508 (N_9508,N_116,N_3925);
nor U9509 (N_9509,N_2793,N_314);
nor U9510 (N_9510,N_942,N_4748);
and U9511 (N_9511,N_2264,N_3341);
nand U9512 (N_9512,N_717,N_2767);
xnor U9513 (N_9513,N_494,N_3401);
xor U9514 (N_9514,N_2541,N_218);
or U9515 (N_9515,N_4863,N_2768);
nand U9516 (N_9516,N_447,N_109);
xnor U9517 (N_9517,N_1734,N_4762);
nor U9518 (N_9518,N_827,N_3651);
xor U9519 (N_9519,N_3065,N_4167);
or U9520 (N_9520,N_2868,N_1393);
nor U9521 (N_9521,N_4451,N_2664);
xnor U9522 (N_9522,N_4395,N_4024);
or U9523 (N_9523,N_4892,N_2343);
xnor U9524 (N_9524,N_3998,N_4311);
or U9525 (N_9525,N_4202,N_167);
or U9526 (N_9526,N_3398,N_994);
nor U9527 (N_9527,N_62,N_1021);
or U9528 (N_9528,N_2734,N_1614);
or U9529 (N_9529,N_4339,N_1182);
xor U9530 (N_9530,N_2535,N_2221);
nor U9531 (N_9531,N_1527,N_972);
nand U9532 (N_9532,N_83,N_376);
nor U9533 (N_9533,N_1844,N_146);
xor U9534 (N_9534,N_3240,N_4728);
or U9535 (N_9535,N_1973,N_3112);
and U9536 (N_9536,N_3013,N_4887);
xnor U9537 (N_9537,N_1050,N_2512);
nor U9538 (N_9538,N_754,N_1258);
xnor U9539 (N_9539,N_3488,N_2500);
xor U9540 (N_9540,N_2659,N_3959);
or U9541 (N_9541,N_2337,N_1576);
xnor U9542 (N_9542,N_3678,N_2030);
xnor U9543 (N_9543,N_4116,N_1170);
xnor U9544 (N_9544,N_2049,N_4460);
nand U9545 (N_9545,N_975,N_1717);
or U9546 (N_9546,N_3087,N_3929);
and U9547 (N_9547,N_4001,N_2968);
xnor U9548 (N_9548,N_4733,N_1647);
nor U9549 (N_9549,N_4924,N_4158);
and U9550 (N_9550,N_2427,N_2374);
and U9551 (N_9551,N_334,N_533);
or U9552 (N_9552,N_2703,N_1714);
and U9553 (N_9553,N_2535,N_891);
and U9554 (N_9554,N_392,N_3856);
and U9555 (N_9555,N_3035,N_3499);
nand U9556 (N_9556,N_1678,N_3732);
nand U9557 (N_9557,N_4247,N_4158);
or U9558 (N_9558,N_4582,N_994);
nor U9559 (N_9559,N_1070,N_1355);
nor U9560 (N_9560,N_4274,N_1233);
nor U9561 (N_9561,N_2964,N_3533);
nor U9562 (N_9562,N_3459,N_4350);
or U9563 (N_9563,N_4285,N_132);
nor U9564 (N_9564,N_1283,N_1387);
and U9565 (N_9565,N_4509,N_2940);
and U9566 (N_9566,N_4618,N_4990);
and U9567 (N_9567,N_2140,N_3320);
and U9568 (N_9568,N_3980,N_57);
and U9569 (N_9569,N_1064,N_36);
nor U9570 (N_9570,N_2902,N_865);
xor U9571 (N_9571,N_2324,N_2502);
nand U9572 (N_9572,N_4173,N_2788);
nor U9573 (N_9573,N_673,N_2499);
nor U9574 (N_9574,N_3361,N_977);
nor U9575 (N_9575,N_2825,N_2515);
nor U9576 (N_9576,N_3977,N_933);
nand U9577 (N_9577,N_4730,N_2123);
nor U9578 (N_9578,N_4813,N_3834);
nand U9579 (N_9579,N_4117,N_1390);
nand U9580 (N_9580,N_1820,N_1351);
xnor U9581 (N_9581,N_4980,N_3814);
or U9582 (N_9582,N_2935,N_121);
and U9583 (N_9583,N_135,N_965);
xor U9584 (N_9584,N_2814,N_2141);
nor U9585 (N_9585,N_4385,N_541);
nand U9586 (N_9586,N_1546,N_3070);
or U9587 (N_9587,N_2493,N_889);
xor U9588 (N_9588,N_4178,N_791);
and U9589 (N_9589,N_1015,N_171);
xnor U9590 (N_9590,N_1869,N_4662);
and U9591 (N_9591,N_11,N_1979);
and U9592 (N_9592,N_4889,N_807);
and U9593 (N_9593,N_1810,N_746);
xnor U9594 (N_9594,N_1588,N_4617);
or U9595 (N_9595,N_3154,N_4058);
nand U9596 (N_9596,N_4608,N_938);
and U9597 (N_9597,N_2214,N_3183);
and U9598 (N_9598,N_4888,N_4129);
or U9599 (N_9599,N_3257,N_517);
or U9600 (N_9600,N_468,N_2222);
or U9601 (N_9601,N_483,N_3113);
or U9602 (N_9602,N_3790,N_1082);
and U9603 (N_9603,N_492,N_241);
or U9604 (N_9604,N_4691,N_1322);
nand U9605 (N_9605,N_2319,N_2189);
nand U9606 (N_9606,N_4495,N_1143);
or U9607 (N_9607,N_4023,N_4885);
xnor U9608 (N_9608,N_1973,N_71);
and U9609 (N_9609,N_2708,N_3650);
nor U9610 (N_9610,N_2309,N_1059);
and U9611 (N_9611,N_4610,N_4961);
and U9612 (N_9612,N_4313,N_1232);
nor U9613 (N_9613,N_2867,N_3305);
nand U9614 (N_9614,N_820,N_4757);
or U9615 (N_9615,N_4058,N_4858);
or U9616 (N_9616,N_641,N_3679);
or U9617 (N_9617,N_2817,N_4987);
or U9618 (N_9618,N_4381,N_2619);
nor U9619 (N_9619,N_1264,N_1017);
and U9620 (N_9620,N_290,N_2878);
xnor U9621 (N_9621,N_3117,N_799);
or U9622 (N_9622,N_1777,N_3556);
and U9623 (N_9623,N_1522,N_666);
xnor U9624 (N_9624,N_2787,N_1885);
and U9625 (N_9625,N_1420,N_1768);
or U9626 (N_9626,N_2616,N_3577);
or U9627 (N_9627,N_3288,N_3506);
and U9628 (N_9628,N_2113,N_351);
and U9629 (N_9629,N_1573,N_204);
xnor U9630 (N_9630,N_4544,N_765);
nand U9631 (N_9631,N_3054,N_1670);
xor U9632 (N_9632,N_4834,N_329);
xor U9633 (N_9633,N_2294,N_4677);
xnor U9634 (N_9634,N_922,N_1772);
and U9635 (N_9635,N_3807,N_660);
nand U9636 (N_9636,N_4978,N_3210);
and U9637 (N_9637,N_4557,N_4661);
nand U9638 (N_9638,N_3832,N_1881);
or U9639 (N_9639,N_178,N_354);
or U9640 (N_9640,N_3921,N_3095);
nand U9641 (N_9641,N_4084,N_126);
and U9642 (N_9642,N_693,N_1045);
and U9643 (N_9643,N_1566,N_1529);
or U9644 (N_9644,N_1486,N_4448);
xnor U9645 (N_9645,N_4651,N_3286);
nand U9646 (N_9646,N_2151,N_2596);
xor U9647 (N_9647,N_4989,N_1689);
and U9648 (N_9648,N_89,N_1268);
and U9649 (N_9649,N_1772,N_4850);
or U9650 (N_9650,N_2994,N_2251);
and U9651 (N_9651,N_4161,N_3238);
nor U9652 (N_9652,N_2014,N_3086);
nor U9653 (N_9653,N_928,N_2527);
xor U9654 (N_9654,N_1647,N_992);
and U9655 (N_9655,N_672,N_4731);
and U9656 (N_9656,N_4714,N_246);
or U9657 (N_9657,N_546,N_2456);
and U9658 (N_9658,N_4765,N_3117);
and U9659 (N_9659,N_4444,N_1899);
nor U9660 (N_9660,N_3444,N_3993);
nand U9661 (N_9661,N_2732,N_4284);
nor U9662 (N_9662,N_1027,N_297);
nor U9663 (N_9663,N_4589,N_4264);
and U9664 (N_9664,N_3297,N_4297);
nor U9665 (N_9665,N_1312,N_4884);
xnor U9666 (N_9666,N_842,N_2669);
or U9667 (N_9667,N_1798,N_4979);
nor U9668 (N_9668,N_4733,N_484);
or U9669 (N_9669,N_2111,N_1286);
xor U9670 (N_9670,N_1491,N_3468);
and U9671 (N_9671,N_1651,N_937);
xnor U9672 (N_9672,N_1120,N_519);
xnor U9673 (N_9673,N_278,N_3259);
xnor U9674 (N_9674,N_75,N_275);
and U9675 (N_9675,N_3823,N_4041);
and U9676 (N_9676,N_1119,N_3030);
nand U9677 (N_9677,N_73,N_676);
nand U9678 (N_9678,N_4755,N_4507);
nor U9679 (N_9679,N_1941,N_3338);
xnor U9680 (N_9680,N_517,N_2501);
nand U9681 (N_9681,N_3598,N_3891);
xnor U9682 (N_9682,N_3705,N_3228);
and U9683 (N_9683,N_2410,N_803);
xnor U9684 (N_9684,N_3473,N_1434);
nand U9685 (N_9685,N_4198,N_4191);
and U9686 (N_9686,N_3471,N_1570);
nor U9687 (N_9687,N_2303,N_3631);
or U9688 (N_9688,N_518,N_3699);
and U9689 (N_9689,N_3524,N_4449);
nor U9690 (N_9690,N_2528,N_324);
or U9691 (N_9691,N_1888,N_1781);
nand U9692 (N_9692,N_690,N_128);
nand U9693 (N_9693,N_3307,N_4298);
nand U9694 (N_9694,N_3937,N_1045);
nand U9695 (N_9695,N_3986,N_2776);
nor U9696 (N_9696,N_2611,N_2198);
nand U9697 (N_9697,N_647,N_2835);
nand U9698 (N_9698,N_201,N_4833);
or U9699 (N_9699,N_1770,N_563);
or U9700 (N_9700,N_3113,N_4601);
nand U9701 (N_9701,N_4727,N_3292);
and U9702 (N_9702,N_2238,N_1493);
nand U9703 (N_9703,N_1986,N_2818);
and U9704 (N_9704,N_731,N_927);
or U9705 (N_9705,N_2273,N_2633);
and U9706 (N_9706,N_220,N_3618);
nand U9707 (N_9707,N_2777,N_424);
nand U9708 (N_9708,N_4426,N_273);
and U9709 (N_9709,N_1956,N_369);
nor U9710 (N_9710,N_1338,N_3227);
nand U9711 (N_9711,N_3084,N_1232);
nor U9712 (N_9712,N_4775,N_2597);
nand U9713 (N_9713,N_4144,N_1420);
or U9714 (N_9714,N_4006,N_1737);
nor U9715 (N_9715,N_3631,N_2991);
nand U9716 (N_9716,N_1286,N_675);
xnor U9717 (N_9717,N_1438,N_2540);
nor U9718 (N_9718,N_1506,N_3021);
or U9719 (N_9719,N_4644,N_125);
xor U9720 (N_9720,N_3959,N_2829);
xor U9721 (N_9721,N_2764,N_1181);
or U9722 (N_9722,N_609,N_4668);
or U9723 (N_9723,N_36,N_2701);
and U9724 (N_9724,N_2009,N_1070);
or U9725 (N_9725,N_2882,N_3836);
xor U9726 (N_9726,N_3544,N_4304);
or U9727 (N_9727,N_1936,N_4808);
nand U9728 (N_9728,N_2271,N_4633);
and U9729 (N_9729,N_2490,N_4590);
nor U9730 (N_9730,N_2012,N_3087);
and U9731 (N_9731,N_536,N_1846);
or U9732 (N_9732,N_1272,N_2871);
and U9733 (N_9733,N_3818,N_1566);
xnor U9734 (N_9734,N_4119,N_3052);
nor U9735 (N_9735,N_3020,N_3911);
nand U9736 (N_9736,N_27,N_3115);
nand U9737 (N_9737,N_545,N_3398);
xnor U9738 (N_9738,N_1861,N_263);
nor U9739 (N_9739,N_1114,N_2519);
nor U9740 (N_9740,N_1929,N_4879);
nor U9741 (N_9741,N_4122,N_4239);
nor U9742 (N_9742,N_4388,N_2032);
xor U9743 (N_9743,N_2453,N_1474);
nor U9744 (N_9744,N_344,N_4416);
or U9745 (N_9745,N_859,N_4441);
xor U9746 (N_9746,N_4929,N_2131);
xor U9747 (N_9747,N_4469,N_4094);
nor U9748 (N_9748,N_3830,N_800);
nor U9749 (N_9749,N_35,N_1715);
and U9750 (N_9750,N_4218,N_2426);
and U9751 (N_9751,N_3057,N_2563);
or U9752 (N_9752,N_887,N_321);
and U9753 (N_9753,N_270,N_255);
nand U9754 (N_9754,N_4333,N_1370);
or U9755 (N_9755,N_3574,N_1166);
or U9756 (N_9756,N_4271,N_4007);
and U9757 (N_9757,N_1281,N_2920);
or U9758 (N_9758,N_692,N_194);
xor U9759 (N_9759,N_4634,N_3996);
nand U9760 (N_9760,N_4252,N_4074);
nor U9761 (N_9761,N_3646,N_4288);
nand U9762 (N_9762,N_4131,N_1300);
or U9763 (N_9763,N_1960,N_3423);
xnor U9764 (N_9764,N_1233,N_2662);
or U9765 (N_9765,N_348,N_4208);
nor U9766 (N_9766,N_3337,N_2374);
nand U9767 (N_9767,N_3002,N_2465);
xor U9768 (N_9768,N_2806,N_2528);
or U9769 (N_9769,N_4009,N_1759);
or U9770 (N_9770,N_2520,N_3882);
nor U9771 (N_9771,N_546,N_4572);
nor U9772 (N_9772,N_3927,N_3714);
or U9773 (N_9773,N_1558,N_2426);
nor U9774 (N_9774,N_1386,N_4895);
nand U9775 (N_9775,N_1207,N_4373);
and U9776 (N_9776,N_828,N_89);
xor U9777 (N_9777,N_2509,N_3693);
nand U9778 (N_9778,N_3269,N_2759);
and U9779 (N_9779,N_549,N_3678);
or U9780 (N_9780,N_4486,N_1762);
xnor U9781 (N_9781,N_1022,N_3726);
and U9782 (N_9782,N_2054,N_3345);
xor U9783 (N_9783,N_2009,N_2181);
or U9784 (N_9784,N_3297,N_1584);
xor U9785 (N_9785,N_1711,N_4674);
and U9786 (N_9786,N_1032,N_4625);
or U9787 (N_9787,N_1653,N_3458);
nor U9788 (N_9788,N_4246,N_1837);
and U9789 (N_9789,N_3724,N_3556);
nor U9790 (N_9790,N_3047,N_1446);
and U9791 (N_9791,N_3319,N_2934);
and U9792 (N_9792,N_4347,N_1120);
nand U9793 (N_9793,N_540,N_2246);
nand U9794 (N_9794,N_4948,N_4783);
or U9795 (N_9795,N_3101,N_13);
nand U9796 (N_9796,N_1382,N_4270);
xnor U9797 (N_9797,N_4737,N_2757);
nand U9798 (N_9798,N_3871,N_3549);
and U9799 (N_9799,N_2988,N_2052);
nand U9800 (N_9800,N_3272,N_4386);
nand U9801 (N_9801,N_1200,N_1229);
nor U9802 (N_9802,N_1476,N_3740);
or U9803 (N_9803,N_2220,N_4430);
xor U9804 (N_9804,N_3478,N_3961);
or U9805 (N_9805,N_1222,N_373);
and U9806 (N_9806,N_231,N_3584);
and U9807 (N_9807,N_3432,N_1094);
xnor U9808 (N_9808,N_3811,N_1989);
nand U9809 (N_9809,N_138,N_1796);
nor U9810 (N_9810,N_506,N_1831);
nor U9811 (N_9811,N_4633,N_4895);
and U9812 (N_9812,N_823,N_4591);
nor U9813 (N_9813,N_4046,N_3932);
and U9814 (N_9814,N_444,N_3702);
xor U9815 (N_9815,N_2401,N_1524);
xnor U9816 (N_9816,N_3244,N_1081);
or U9817 (N_9817,N_4911,N_3772);
xnor U9818 (N_9818,N_43,N_1287);
and U9819 (N_9819,N_1909,N_3129);
nand U9820 (N_9820,N_3741,N_3090);
xnor U9821 (N_9821,N_1659,N_485);
nand U9822 (N_9822,N_2151,N_2929);
xor U9823 (N_9823,N_3903,N_2164);
nor U9824 (N_9824,N_2397,N_4619);
xor U9825 (N_9825,N_4901,N_2049);
or U9826 (N_9826,N_2037,N_1137);
xnor U9827 (N_9827,N_1709,N_2412);
and U9828 (N_9828,N_1600,N_4999);
and U9829 (N_9829,N_2074,N_319);
or U9830 (N_9830,N_2683,N_1254);
xor U9831 (N_9831,N_584,N_1164);
nor U9832 (N_9832,N_2894,N_1792);
nor U9833 (N_9833,N_2108,N_4730);
or U9834 (N_9834,N_3011,N_4131);
or U9835 (N_9835,N_4241,N_2438);
and U9836 (N_9836,N_746,N_4962);
nand U9837 (N_9837,N_426,N_4601);
xnor U9838 (N_9838,N_3675,N_4592);
nand U9839 (N_9839,N_888,N_305);
or U9840 (N_9840,N_3371,N_2109);
or U9841 (N_9841,N_569,N_4413);
and U9842 (N_9842,N_4897,N_3863);
nor U9843 (N_9843,N_4462,N_1033);
and U9844 (N_9844,N_1540,N_529);
nand U9845 (N_9845,N_4042,N_114);
and U9846 (N_9846,N_2121,N_36);
nand U9847 (N_9847,N_1614,N_281);
nand U9848 (N_9848,N_3944,N_4223);
xor U9849 (N_9849,N_1819,N_4932);
or U9850 (N_9850,N_3494,N_4909);
xor U9851 (N_9851,N_4743,N_2181);
xnor U9852 (N_9852,N_171,N_1227);
nand U9853 (N_9853,N_4087,N_1147);
and U9854 (N_9854,N_4883,N_3289);
nor U9855 (N_9855,N_2699,N_4463);
nand U9856 (N_9856,N_4184,N_4577);
or U9857 (N_9857,N_2657,N_4386);
xor U9858 (N_9858,N_342,N_2786);
nand U9859 (N_9859,N_2064,N_4543);
or U9860 (N_9860,N_36,N_1023);
xnor U9861 (N_9861,N_3222,N_1779);
or U9862 (N_9862,N_1047,N_4988);
and U9863 (N_9863,N_4730,N_4339);
xnor U9864 (N_9864,N_709,N_1278);
xor U9865 (N_9865,N_4373,N_2682);
and U9866 (N_9866,N_4170,N_1401);
xnor U9867 (N_9867,N_2055,N_3442);
xor U9868 (N_9868,N_560,N_2495);
and U9869 (N_9869,N_1412,N_1340);
nor U9870 (N_9870,N_2193,N_4740);
nor U9871 (N_9871,N_2752,N_1972);
or U9872 (N_9872,N_4632,N_4681);
xor U9873 (N_9873,N_4585,N_761);
nor U9874 (N_9874,N_3945,N_1167);
and U9875 (N_9875,N_1528,N_2863);
or U9876 (N_9876,N_1081,N_1929);
xor U9877 (N_9877,N_3363,N_3338);
or U9878 (N_9878,N_2145,N_215);
xnor U9879 (N_9879,N_702,N_3931);
nor U9880 (N_9880,N_2160,N_3950);
or U9881 (N_9881,N_3012,N_4812);
xnor U9882 (N_9882,N_2790,N_3916);
xor U9883 (N_9883,N_4879,N_2920);
and U9884 (N_9884,N_3640,N_1927);
nor U9885 (N_9885,N_4337,N_4533);
or U9886 (N_9886,N_663,N_2114);
xnor U9887 (N_9887,N_1012,N_4181);
xnor U9888 (N_9888,N_972,N_496);
and U9889 (N_9889,N_1828,N_4631);
xnor U9890 (N_9890,N_504,N_4613);
xnor U9891 (N_9891,N_3188,N_3760);
and U9892 (N_9892,N_4711,N_259);
or U9893 (N_9893,N_335,N_1112);
xor U9894 (N_9894,N_3849,N_2133);
nand U9895 (N_9895,N_1905,N_3446);
nor U9896 (N_9896,N_1801,N_111);
nor U9897 (N_9897,N_3012,N_90);
and U9898 (N_9898,N_4521,N_226);
nor U9899 (N_9899,N_4162,N_955);
or U9900 (N_9900,N_4662,N_3922);
xor U9901 (N_9901,N_603,N_2459);
nand U9902 (N_9902,N_4014,N_1528);
nand U9903 (N_9903,N_134,N_3714);
or U9904 (N_9904,N_4077,N_3388);
and U9905 (N_9905,N_3852,N_128);
xor U9906 (N_9906,N_2667,N_3240);
nand U9907 (N_9907,N_2485,N_190);
nor U9908 (N_9908,N_463,N_3311);
nand U9909 (N_9909,N_2632,N_798);
nor U9910 (N_9910,N_2657,N_4091);
or U9911 (N_9911,N_3702,N_4671);
nor U9912 (N_9912,N_1169,N_2182);
nor U9913 (N_9913,N_4991,N_1980);
xnor U9914 (N_9914,N_1187,N_3884);
nor U9915 (N_9915,N_1146,N_2850);
nor U9916 (N_9916,N_824,N_3793);
or U9917 (N_9917,N_2627,N_700);
or U9918 (N_9918,N_3321,N_4364);
and U9919 (N_9919,N_3360,N_1383);
nor U9920 (N_9920,N_1204,N_2713);
nand U9921 (N_9921,N_2514,N_1096);
nor U9922 (N_9922,N_4475,N_4377);
or U9923 (N_9923,N_2487,N_4300);
and U9924 (N_9924,N_2450,N_3552);
and U9925 (N_9925,N_4921,N_4143);
nor U9926 (N_9926,N_446,N_1626);
or U9927 (N_9927,N_3401,N_3139);
or U9928 (N_9928,N_239,N_2448);
xnor U9929 (N_9929,N_4933,N_2195);
and U9930 (N_9930,N_1871,N_4054);
xnor U9931 (N_9931,N_266,N_4294);
or U9932 (N_9932,N_1102,N_3231);
xor U9933 (N_9933,N_1237,N_200);
nand U9934 (N_9934,N_1960,N_763);
nor U9935 (N_9935,N_1108,N_1608);
nor U9936 (N_9936,N_538,N_433);
xnor U9937 (N_9937,N_1232,N_446);
nor U9938 (N_9938,N_2645,N_712);
and U9939 (N_9939,N_4566,N_918);
or U9940 (N_9940,N_77,N_2748);
nand U9941 (N_9941,N_4228,N_356);
nor U9942 (N_9942,N_3864,N_4458);
xnor U9943 (N_9943,N_1392,N_2563);
and U9944 (N_9944,N_3807,N_1712);
and U9945 (N_9945,N_2206,N_639);
and U9946 (N_9946,N_2218,N_785);
nand U9947 (N_9947,N_457,N_2570);
and U9948 (N_9948,N_3468,N_1699);
nand U9949 (N_9949,N_3453,N_4115);
nor U9950 (N_9950,N_48,N_1092);
and U9951 (N_9951,N_3747,N_370);
and U9952 (N_9952,N_1783,N_1749);
nand U9953 (N_9953,N_4607,N_2565);
xnor U9954 (N_9954,N_1935,N_1417);
and U9955 (N_9955,N_3699,N_855);
xor U9956 (N_9956,N_1833,N_3470);
or U9957 (N_9957,N_876,N_2674);
nand U9958 (N_9958,N_2090,N_3362);
and U9959 (N_9959,N_3771,N_2305);
nand U9960 (N_9960,N_1926,N_4269);
nor U9961 (N_9961,N_3920,N_4842);
or U9962 (N_9962,N_3143,N_866);
and U9963 (N_9963,N_265,N_291);
or U9964 (N_9964,N_2418,N_3966);
xnor U9965 (N_9965,N_3975,N_993);
nor U9966 (N_9966,N_2901,N_2352);
xor U9967 (N_9967,N_4821,N_1208);
nor U9968 (N_9968,N_3900,N_170);
or U9969 (N_9969,N_4267,N_4538);
nor U9970 (N_9970,N_2755,N_3278);
or U9971 (N_9971,N_3553,N_1371);
nand U9972 (N_9972,N_370,N_730);
nor U9973 (N_9973,N_616,N_1016);
nand U9974 (N_9974,N_4434,N_1864);
nor U9975 (N_9975,N_2496,N_4706);
and U9976 (N_9976,N_2653,N_2245);
xor U9977 (N_9977,N_3833,N_1087);
nand U9978 (N_9978,N_4528,N_234);
nand U9979 (N_9979,N_588,N_707);
nand U9980 (N_9980,N_211,N_4312);
nor U9981 (N_9981,N_2022,N_743);
nor U9982 (N_9982,N_2833,N_1654);
or U9983 (N_9983,N_1769,N_4323);
and U9984 (N_9984,N_2178,N_424);
xor U9985 (N_9985,N_4763,N_87);
nand U9986 (N_9986,N_39,N_3475);
xnor U9987 (N_9987,N_1237,N_567);
and U9988 (N_9988,N_3660,N_1834);
nor U9989 (N_9989,N_1798,N_3305);
or U9990 (N_9990,N_208,N_4105);
or U9991 (N_9991,N_3682,N_3617);
xnor U9992 (N_9992,N_1699,N_3595);
nand U9993 (N_9993,N_2358,N_4021);
nor U9994 (N_9994,N_4794,N_4716);
nor U9995 (N_9995,N_3566,N_4498);
nor U9996 (N_9996,N_3331,N_4008);
nand U9997 (N_9997,N_2937,N_706);
or U9998 (N_9998,N_4663,N_3400);
or U9999 (N_9999,N_646,N_4856);
nand U10000 (N_10000,N_7864,N_5028);
nand U10001 (N_10001,N_7306,N_6110);
and U10002 (N_10002,N_8128,N_8347);
and U10003 (N_10003,N_9361,N_6221);
and U10004 (N_10004,N_8444,N_6828);
or U10005 (N_10005,N_7050,N_6664);
and U10006 (N_10006,N_8810,N_6674);
nor U10007 (N_10007,N_5496,N_5173);
nor U10008 (N_10008,N_9842,N_5722);
nor U10009 (N_10009,N_9131,N_7532);
and U10010 (N_10010,N_9005,N_8169);
and U10011 (N_10011,N_7068,N_7857);
xnor U10012 (N_10012,N_9996,N_8212);
or U10013 (N_10013,N_6984,N_9899);
xnor U10014 (N_10014,N_7843,N_8164);
or U10015 (N_10015,N_9541,N_9935);
nor U10016 (N_10016,N_5671,N_6764);
nand U10017 (N_10017,N_6797,N_8342);
nand U10018 (N_10018,N_9101,N_7938);
nand U10019 (N_10019,N_7420,N_9794);
nand U10020 (N_10020,N_8176,N_8421);
nand U10021 (N_10021,N_5220,N_8693);
xor U10022 (N_10022,N_8745,N_8251);
or U10023 (N_10023,N_7931,N_8933);
nand U10024 (N_10024,N_9027,N_9446);
nor U10025 (N_10025,N_5253,N_6825);
xor U10026 (N_10026,N_9181,N_5561);
and U10027 (N_10027,N_7492,N_7926);
or U10028 (N_10028,N_6057,N_6934);
or U10029 (N_10029,N_8096,N_5935);
xor U10030 (N_10030,N_7309,N_5506);
nand U10031 (N_10031,N_7890,N_5251);
xor U10032 (N_10032,N_9487,N_9622);
or U10033 (N_10033,N_6077,N_5338);
and U10034 (N_10034,N_9301,N_6465);
or U10035 (N_10035,N_9906,N_6331);
nand U10036 (N_10036,N_8847,N_7371);
xnor U10037 (N_10037,N_5100,N_7599);
nor U10038 (N_10038,N_6337,N_6416);
nand U10039 (N_10039,N_9388,N_7765);
xnor U10040 (N_10040,N_7279,N_5818);
xnor U10041 (N_10041,N_9727,N_5403);
or U10042 (N_10042,N_9734,N_8638);
nand U10043 (N_10043,N_6267,N_7645);
xor U10044 (N_10044,N_8768,N_8833);
or U10045 (N_10045,N_5801,N_5388);
xnor U10046 (N_10046,N_9391,N_6639);
nand U10047 (N_10047,N_5250,N_7159);
xor U10048 (N_10048,N_5924,N_7958);
and U10049 (N_10049,N_5227,N_9843);
and U10050 (N_10050,N_9819,N_9195);
nor U10051 (N_10051,N_8455,N_8433);
nand U10052 (N_10052,N_7125,N_5948);
and U10053 (N_10053,N_8920,N_9854);
xor U10054 (N_10054,N_7283,N_8598);
xor U10055 (N_10055,N_9862,N_7282);
and U10056 (N_10056,N_7084,N_9248);
or U10057 (N_10057,N_6201,N_7587);
nand U10058 (N_10058,N_8182,N_8758);
or U10059 (N_10059,N_6715,N_5115);
nand U10060 (N_10060,N_8245,N_5456);
and U10061 (N_10061,N_9038,N_6495);
or U10062 (N_10062,N_5822,N_6821);
and U10063 (N_10063,N_8230,N_5938);
nand U10064 (N_10064,N_7650,N_7742);
xnor U10065 (N_10065,N_6233,N_7628);
xor U10066 (N_10066,N_5840,N_5476);
xor U10067 (N_10067,N_9406,N_5928);
or U10068 (N_10068,N_5482,N_6161);
and U10069 (N_10069,N_8706,N_8961);
and U10070 (N_10070,N_7034,N_8189);
xor U10071 (N_10071,N_8020,N_6211);
or U10072 (N_10072,N_5753,N_7995);
or U10073 (N_10073,N_5952,N_6017);
nand U10074 (N_10074,N_6444,N_6086);
xnor U10075 (N_10075,N_9865,N_9345);
xor U10076 (N_10076,N_7554,N_7848);
and U10077 (N_10077,N_8405,N_6689);
xor U10078 (N_10078,N_8333,N_5518);
nor U10079 (N_10079,N_7360,N_9158);
and U10080 (N_10080,N_6354,N_5961);
nor U10081 (N_10081,N_9864,N_8701);
or U10082 (N_10082,N_5153,N_9015);
and U10083 (N_10083,N_8938,N_8157);
nor U10084 (N_10084,N_7867,N_9236);
and U10085 (N_10085,N_8793,N_8763);
nor U10086 (N_10086,N_8992,N_8228);
nand U10087 (N_10087,N_7392,N_6502);
and U10088 (N_10088,N_7751,N_8801);
or U10089 (N_10089,N_7953,N_9231);
nor U10090 (N_10090,N_9934,N_8932);
nor U10091 (N_10091,N_8173,N_7838);
nand U10092 (N_10092,N_9871,N_6215);
nor U10093 (N_10093,N_5603,N_8748);
xor U10094 (N_10094,N_7053,N_6670);
and U10095 (N_10095,N_7381,N_9139);
and U10096 (N_10096,N_6072,N_6371);
nor U10097 (N_10097,N_7302,N_5445);
nor U10098 (N_10098,N_6928,N_9562);
and U10099 (N_10099,N_9775,N_9769);
nor U10100 (N_10100,N_9550,N_6148);
and U10101 (N_10101,N_7464,N_5148);
or U10102 (N_10102,N_8741,N_7552);
nor U10103 (N_10103,N_7986,N_7689);
nand U10104 (N_10104,N_9922,N_5014);
or U10105 (N_10105,N_8217,N_7107);
nor U10106 (N_10106,N_9907,N_9490);
nand U10107 (N_10107,N_6711,N_9247);
or U10108 (N_10108,N_8472,N_7969);
nor U10109 (N_10109,N_8561,N_8272);
xnor U10110 (N_10110,N_6508,N_5215);
or U10111 (N_10111,N_8897,N_8734);
and U10112 (N_10112,N_5748,N_8773);
and U10113 (N_10113,N_6969,N_5993);
nor U10114 (N_10114,N_8590,N_8591);
xor U10115 (N_10115,N_7019,N_6183);
nand U10116 (N_10116,N_9923,N_8990);
or U10117 (N_10117,N_6523,N_8718);
or U10118 (N_10118,N_5046,N_7895);
xor U10119 (N_10119,N_9289,N_6656);
nand U10120 (N_10120,N_9477,N_7896);
nand U10121 (N_10121,N_8735,N_6248);
nand U10122 (N_10122,N_5214,N_5971);
nor U10123 (N_10123,N_7688,N_6351);
nor U10124 (N_10124,N_6198,N_9260);
nand U10125 (N_10125,N_7516,N_8923);
nand U10126 (N_10126,N_7951,N_5188);
and U10127 (N_10127,N_8406,N_6587);
nand U10128 (N_10128,N_7517,N_8499);
nand U10129 (N_10129,N_6016,N_5260);
xnor U10130 (N_10130,N_8130,N_8152);
nand U10131 (N_10131,N_9690,N_8142);
xor U10132 (N_10132,N_8686,N_9306);
xnor U10133 (N_10133,N_8330,N_9605);
nor U10134 (N_10134,N_6743,N_5544);
nor U10135 (N_10135,N_5957,N_7183);
nor U10136 (N_10136,N_8034,N_9272);
nor U10137 (N_10137,N_5252,N_5637);
xnor U10138 (N_10138,N_6230,N_7209);
nor U10139 (N_10139,N_8694,N_9692);
nor U10140 (N_10140,N_9489,N_9679);
or U10141 (N_10141,N_5293,N_5198);
or U10142 (N_10142,N_5925,N_6503);
xor U10143 (N_10143,N_5238,N_5084);
and U10144 (N_10144,N_7128,N_6930);
and U10145 (N_10145,N_5313,N_8894);
nor U10146 (N_10146,N_6679,N_7006);
or U10147 (N_10147,N_6339,N_5172);
nor U10148 (N_10148,N_9989,N_9269);
nor U10149 (N_10149,N_9523,N_6784);
and U10150 (N_10150,N_7174,N_6265);
and U10151 (N_10151,N_6202,N_9688);
and U10152 (N_10152,N_6687,N_9790);
xor U10153 (N_10153,N_5768,N_8149);
and U10154 (N_10154,N_5815,N_8458);
and U10155 (N_10155,N_6659,N_9543);
nor U10156 (N_10156,N_8683,N_8380);
nand U10157 (N_10157,N_8231,N_7402);
and U10158 (N_10158,N_9891,N_5047);
xnor U10159 (N_10159,N_7333,N_5093);
nor U10160 (N_10160,N_9175,N_7832);
xor U10161 (N_10161,N_8611,N_6557);
or U10162 (N_10162,N_6063,N_6996);
and U10163 (N_10163,N_9300,N_7262);
nor U10164 (N_10164,N_9048,N_6757);
nand U10165 (N_10165,N_6193,N_5132);
xnor U10166 (N_10166,N_6264,N_8141);
or U10167 (N_10167,N_9662,N_5413);
or U10168 (N_10168,N_6239,N_7403);
xor U10169 (N_10169,N_9009,N_8781);
nor U10170 (N_10170,N_7862,N_5414);
nand U10171 (N_10171,N_5221,N_9024);
nor U10172 (N_10172,N_9396,N_5343);
nand U10173 (N_10173,N_6350,N_9022);
nand U10174 (N_10174,N_6634,N_6652);
nor U10175 (N_10175,N_6088,N_9157);
nor U10176 (N_10176,N_9431,N_8240);
and U10177 (N_10177,N_9916,N_6987);
xnor U10178 (N_10178,N_7796,N_9837);
nor U10179 (N_10179,N_7394,N_8653);
and U10180 (N_10180,N_7244,N_5258);
nand U10181 (N_10181,N_5599,N_6253);
xnor U10182 (N_10182,N_5996,N_8829);
xnor U10183 (N_10183,N_9618,N_9671);
or U10184 (N_10184,N_6991,N_7866);
nand U10185 (N_10185,N_9804,N_8378);
xnor U10186 (N_10186,N_8058,N_7303);
or U10187 (N_10187,N_8014,N_9349);
or U10188 (N_10188,N_6777,N_9963);
and U10189 (N_10189,N_7294,N_9321);
and U10190 (N_10190,N_6599,N_5721);
and U10191 (N_10191,N_6007,N_9820);
nand U10192 (N_10192,N_8370,N_7760);
or U10193 (N_10193,N_5960,N_5479);
nor U10194 (N_10194,N_7920,N_9560);
and U10195 (N_10195,N_7851,N_7583);
nand U10196 (N_10196,N_6864,N_8605);
nor U10197 (N_10197,N_9389,N_7978);
and U10198 (N_10198,N_6677,N_8427);
and U10199 (N_10199,N_7768,N_6517);
and U10200 (N_10200,N_8952,N_8003);
xnor U10201 (N_10201,N_5991,N_9786);
nand U10202 (N_10202,N_7405,N_5713);
nor U10203 (N_10203,N_8418,N_8756);
or U10204 (N_10204,N_6438,N_6542);
and U10205 (N_10205,N_5033,N_8423);
and U10206 (N_10206,N_7500,N_5005);
xor U10207 (N_10207,N_8443,N_6405);
and U10208 (N_10208,N_9990,N_5542);
or U10209 (N_10209,N_6621,N_9378);
xnor U10210 (N_10210,N_5017,N_8644);
nand U10211 (N_10211,N_7005,N_5012);
nor U10212 (N_10212,N_5585,N_9970);
nand U10213 (N_10213,N_7063,N_9567);
xnor U10214 (N_10214,N_7273,N_8247);
nor U10215 (N_10215,N_6190,N_9287);
xor U10216 (N_10216,N_5798,N_8996);
xnor U10217 (N_10217,N_7823,N_7519);
nand U10218 (N_10218,N_9604,N_8885);
xnor U10219 (N_10219,N_6841,N_7376);
and U10220 (N_10220,N_9137,N_8125);
and U10221 (N_10221,N_8634,N_9733);
xor U10222 (N_10222,N_8078,N_6893);
and U10223 (N_10223,N_5695,N_7581);
or U10224 (N_10224,N_8654,N_9316);
nand U10225 (N_10225,N_9075,N_7509);
or U10226 (N_10226,N_8827,N_5568);
and U10227 (N_10227,N_6129,N_9546);
and U10228 (N_10228,N_5369,N_5090);
or U10229 (N_10229,N_8875,N_6464);
nand U10230 (N_10230,N_8165,N_7409);
and U10231 (N_10231,N_6237,N_5291);
and U10232 (N_10232,N_6366,N_9932);
or U10233 (N_10233,N_5076,N_5788);
and U10234 (N_10234,N_8056,N_6716);
nand U10235 (N_10235,N_6628,N_9793);
xnor U10236 (N_10236,N_6657,N_7132);
nor U10237 (N_10237,N_8174,N_8767);
nor U10238 (N_10238,N_6483,N_9817);
and U10239 (N_10239,N_5868,N_5044);
and U10240 (N_10240,N_6873,N_9776);
nor U10241 (N_10241,N_7707,N_6959);
and U10242 (N_10242,N_8011,N_8349);
or U10243 (N_10243,N_8846,N_9186);
nor U10244 (N_10244,N_6736,N_6999);
nor U10245 (N_10245,N_7683,N_9438);
nor U10246 (N_10246,N_6471,N_6281);
nor U10247 (N_10247,N_5177,N_9276);
and U10248 (N_10248,N_6270,N_9405);
nor U10249 (N_10249,N_7661,N_6385);
and U10250 (N_10250,N_7593,N_7865);
nor U10251 (N_10251,N_9191,N_7887);
nor U10252 (N_10252,N_9747,N_7199);
or U10253 (N_10253,N_8604,N_5200);
and U10254 (N_10254,N_9711,N_6972);
xnor U10255 (N_10255,N_6291,N_5997);
nand U10256 (N_10256,N_5643,N_6322);
xor U10257 (N_10257,N_6878,N_6698);
and U10258 (N_10258,N_7348,N_9982);
nor U10259 (N_10259,N_8432,N_6328);
nand U10260 (N_10260,N_6808,N_6593);
nand U10261 (N_10261,N_6831,N_5335);
nand U10262 (N_10262,N_8028,N_6895);
nor U10263 (N_10263,N_5320,N_9224);
nor U10264 (N_10264,N_5789,N_9814);
and U10265 (N_10265,N_5652,N_5239);
xor U10266 (N_10266,N_5183,N_9271);
xor U10267 (N_10267,N_7894,N_9595);
xor U10268 (N_10268,N_9514,N_8752);
and U10269 (N_10269,N_7379,N_5539);
or U10270 (N_10270,N_8185,N_6970);
nor U10271 (N_10271,N_8621,N_5500);
xor U10272 (N_10272,N_7803,N_7215);
and U10273 (N_10273,N_6163,N_9593);
xnor U10274 (N_10274,N_5931,N_6045);
xnor U10275 (N_10275,N_6229,N_6901);
xnor U10276 (N_10276,N_7748,N_5596);
nand U10277 (N_10277,N_6159,N_8656);
and U10278 (N_10278,N_5397,N_7542);
xor U10279 (N_10279,N_9293,N_8184);
or U10280 (N_10280,N_7042,N_7793);
nor U10281 (N_10281,N_7000,N_6436);
and U10282 (N_10282,N_8377,N_7595);
xnor U10283 (N_10283,N_6141,N_6580);
nor U10284 (N_10284,N_9440,N_7233);
or U10285 (N_10285,N_5906,N_7809);
or U10286 (N_10286,N_8613,N_6766);
xnor U10287 (N_10287,N_7845,N_6426);
nor U10288 (N_10288,N_5196,N_5680);
nand U10289 (N_10289,N_9323,N_7237);
nand U10290 (N_10290,N_8966,N_9347);
nand U10291 (N_10291,N_8581,N_7004);
nor U10292 (N_10292,N_7772,N_9423);
nor U10293 (N_10293,N_5186,N_7563);
nor U10294 (N_10294,N_8258,N_6362);
and U10295 (N_10295,N_6536,N_9680);
and U10296 (N_10296,N_6914,N_5999);
xor U10297 (N_10297,N_9374,N_6922);
nand U10298 (N_10298,N_9860,N_9246);
or U10299 (N_10299,N_6983,N_5576);
or U10300 (N_10300,N_5703,N_5303);
or U10301 (N_10301,N_9146,N_8974);
xnor U10302 (N_10302,N_8063,N_6187);
or U10303 (N_10303,N_7469,N_7624);
and U10304 (N_10304,N_7657,N_5669);
nand U10305 (N_10305,N_7750,N_7441);
xnor U10306 (N_10306,N_5591,N_6039);
xor U10307 (N_10307,N_6617,N_9753);
and U10308 (N_10308,N_8595,N_9946);
nand U10309 (N_10309,N_6332,N_9766);
or U10310 (N_10310,N_6848,N_6518);
nor U10311 (N_10311,N_7136,N_6310);
nor U10312 (N_10312,N_9233,N_7726);
nor U10313 (N_10313,N_8337,N_9126);
nand U10314 (N_10314,N_9098,N_5638);
nor U10315 (N_10315,N_6466,N_8401);
xor U10316 (N_10316,N_8809,N_5463);
nand U10317 (N_10317,N_6643,N_6907);
and U10318 (N_10318,N_5490,N_9194);
xor U10319 (N_10319,N_9141,N_6568);
and U10320 (N_10320,N_5472,N_5083);
nor U10321 (N_10321,N_6316,N_8220);
or U10322 (N_10322,N_7586,N_7644);
nor U10323 (N_10323,N_9108,N_9893);
and U10324 (N_10324,N_7961,N_7588);
and U10325 (N_10325,N_8681,N_6528);
nand U10326 (N_10326,N_8042,N_8102);
nor U10327 (N_10327,N_9205,N_8050);
xnor U10328 (N_10328,N_8221,N_7898);
nand U10329 (N_10329,N_8296,N_9756);
and U10330 (N_10330,N_7734,N_6939);
and U10331 (N_10331,N_7269,N_7071);
nand U10332 (N_10332,N_7443,N_7806);
and U10333 (N_10333,N_7470,N_6406);
or U10334 (N_10334,N_5541,N_7841);
nand U10335 (N_10335,N_6131,N_5963);
and U10336 (N_10336,N_8738,N_5056);
and U10337 (N_10337,N_7417,N_7222);
nand U10338 (N_10338,N_5793,N_8105);
or U10339 (N_10339,N_7118,N_9802);
xnor U10340 (N_10340,N_5199,N_8420);
xnor U10341 (N_10341,N_5311,N_9274);
xor U10342 (N_10342,N_7124,N_5147);
nand U10343 (N_10343,N_5074,N_5185);
xnor U10344 (N_10344,N_7701,N_5061);
or U10345 (N_10345,N_7672,N_5441);
xnor U10346 (N_10346,N_7332,N_6205);
and U10347 (N_10347,N_7550,N_5812);
or U10348 (N_10348,N_5455,N_5572);
xnor U10349 (N_10349,N_6725,N_6364);
nand U10350 (N_10350,N_6137,N_8314);
xor U10351 (N_10351,N_7915,N_6737);
nand U10352 (N_10352,N_9770,N_5515);
nor U10353 (N_10353,N_9103,N_9043);
and U10354 (N_10354,N_6635,N_7559);
nor U10355 (N_10355,N_9521,N_5571);
and U10356 (N_10356,N_6619,N_8584);
or U10357 (N_10357,N_9579,N_5091);
and U10358 (N_10358,N_8862,N_7681);
nor U10359 (N_10359,N_8731,N_5597);
or U10360 (N_10360,N_6001,N_8260);
and U10361 (N_10361,N_6411,N_7103);
nor U10362 (N_10362,N_5725,N_5946);
and U10363 (N_10363,N_9386,N_8825);
xnor U10364 (N_10364,N_8859,N_8373);
nand U10365 (N_10365,N_8392,N_8172);
and U10366 (N_10366,N_7069,N_5284);
xnor U10367 (N_10367,N_5848,N_6717);
xnor U10368 (N_10368,N_7411,N_8136);
and U10369 (N_10369,N_6974,N_8188);
nor U10370 (N_10370,N_6839,N_5257);
and U10371 (N_10371,N_8065,N_6038);
nor U10372 (N_10372,N_7266,N_8283);
nor U10373 (N_10373,N_9535,N_8775);
nor U10374 (N_10374,N_7919,N_7081);
nor U10375 (N_10375,N_7208,N_5255);
xnor U10376 (N_10376,N_7461,N_9844);
nor U10377 (N_10377,N_9299,N_8218);
nand U10378 (N_10378,N_5893,N_5867);
and U10379 (N_10379,N_7922,N_5174);
and U10380 (N_10380,N_7206,N_8080);
and U10381 (N_10381,N_5069,N_5022);
xnor U10382 (N_10382,N_5094,N_9668);
xnor U10383 (N_10383,N_6071,N_9956);
nor U10384 (N_10384,N_5319,N_8652);
xor U10385 (N_10385,N_8310,N_7972);
xor U10386 (N_10386,N_5276,N_7076);
nand U10387 (N_10387,N_7690,N_7070);
xor U10388 (N_10388,N_9206,N_5315);
and U10389 (N_10389,N_9150,N_6139);
and U10390 (N_10390,N_7531,N_6434);
nor U10391 (N_10391,N_7160,N_6932);
nand U10392 (N_10392,N_9187,N_7404);
xnor U10393 (N_10393,N_9459,N_8040);
and U10394 (N_10394,N_5088,N_6047);
and U10395 (N_10395,N_9602,N_9852);
xnor U10396 (N_10396,N_5895,N_7501);
nor U10397 (N_10397,N_9429,N_6624);
nand U10398 (N_10398,N_7195,N_5246);
nor U10399 (N_10399,N_9221,N_5570);
and U10400 (N_10400,N_8289,N_7388);
or U10401 (N_10401,N_5334,N_5743);
or U10402 (N_10402,N_8651,N_9913);
nand U10403 (N_10403,N_9288,N_5751);
nor U10404 (N_10404,N_7655,N_7329);
and U10405 (N_10405,N_7180,N_8249);
xor U10406 (N_10406,N_5802,N_6213);
nand U10407 (N_10407,N_5922,N_9828);
or U10408 (N_10408,N_8836,N_8803);
or U10409 (N_10409,N_7236,N_8857);
nand U10410 (N_10410,N_9133,N_7521);
xnor U10411 (N_10411,N_7792,N_8379);
or U10412 (N_10412,N_5179,N_8538);
nor U10413 (N_10413,N_7182,N_8119);
xnor U10414 (N_10414,N_8163,N_5411);
xor U10415 (N_10415,N_6286,N_7369);
xnor U10416 (N_10416,N_7775,N_5181);
nand U10417 (N_10417,N_8144,N_5027);
xnor U10418 (N_10418,N_6767,N_6055);
nand U10419 (N_10419,N_8566,N_5773);
or U10420 (N_10420,N_6319,N_8626);
nand U10421 (N_10421,N_5026,N_7704);
xor U10422 (N_10422,N_5308,N_9132);
nor U10423 (N_10423,N_7770,N_9456);
or U10424 (N_10424,N_5740,N_7495);
or U10425 (N_10425,N_8618,N_9371);
and U10426 (N_10426,N_5341,N_6924);
nand U10427 (N_10427,N_9637,N_6919);
nand U10428 (N_10428,N_6858,N_8623);
nand U10429 (N_10429,N_6299,N_7013);
nor U10430 (N_10430,N_6827,N_6942);
and U10431 (N_10431,N_5964,N_6494);
nor U10432 (N_10432,N_7873,N_5939);
nor U10433 (N_10433,N_7390,N_5594);
and U10434 (N_10434,N_9196,N_6025);
and U10435 (N_10435,N_8229,N_8945);
and U10436 (N_10436,N_7391,N_5365);
and U10437 (N_10437,N_9121,N_5843);
nand U10438 (N_10438,N_5363,N_8697);
xor U10439 (N_10439,N_8387,N_5126);
and U10440 (N_10440,N_6641,N_8121);
nor U10441 (N_10441,N_6285,N_5914);
or U10442 (N_10442,N_9156,N_7105);
nor U10443 (N_10443,N_9969,N_8340);
or U10444 (N_10444,N_6391,N_5771);
or U10445 (N_10445,N_6775,N_9724);
xnor U10446 (N_10446,N_9503,N_5042);
xnor U10447 (N_10447,N_7758,N_5977);
and U10448 (N_10448,N_5078,N_5466);
nor U10449 (N_10449,N_8822,N_7738);
nor U10450 (N_10450,N_5098,N_6029);
and U10451 (N_10451,N_7223,N_5647);
or U10452 (N_10452,N_7842,N_8834);
nand U10453 (N_10453,N_8870,N_6588);
and U10454 (N_10454,N_6257,N_9882);
or U10455 (N_10455,N_9473,N_8344);
and U10456 (N_10456,N_6348,N_8737);
and U10457 (N_10457,N_9011,N_5831);
xor U10458 (N_10458,N_7565,N_7361);
and U10459 (N_10459,N_9443,N_5998);
nand U10460 (N_10460,N_7692,N_7295);
and U10461 (N_10461,N_5543,N_5342);
and U10462 (N_10462,N_7205,N_5399);
xnor U10463 (N_10463,N_5858,N_8343);
nor U10464 (N_10464,N_6747,N_5814);
nand U10465 (N_10465,N_9120,N_9308);
or U10466 (N_10466,N_7307,N_7207);
nand U10467 (N_10467,N_6951,N_7072);
and U10468 (N_10468,N_6565,N_8855);
or U10469 (N_10469,N_7483,N_5218);
nand U10470 (N_10470,N_7663,N_9741);
xnor U10471 (N_10471,N_8509,N_6719);
and U10472 (N_10472,N_7572,N_6718);
xnor U10473 (N_10473,N_9165,N_6463);
and U10474 (N_10474,N_6931,N_8872);
nand U10475 (N_10475,N_5432,N_8410);
or U10476 (N_10476,N_6100,N_6309);
or U10477 (N_10477,N_6756,N_5374);
nand U10478 (N_10478,N_5507,N_7436);
nor U10479 (N_10479,N_6021,N_8197);
and U10480 (N_10480,N_5934,N_7187);
nand U10481 (N_10481,N_8650,N_5982);
and U10482 (N_10482,N_6491,N_5009);
and U10483 (N_10483,N_9557,N_6519);
xor U10484 (N_10484,N_7364,N_9627);
and U10485 (N_10485,N_5888,N_9482);
nand U10486 (N_10486,N_5485,N_8000);
xor U10487 (N_10487,N_7292,N_7714);
xor U10488 (N_10488,N_7173,N_5645);
nand U10489 (N_10489,N_7524,N_8930);
nand U10490 (N_10490,N_9988,N_5471);
or U10491 (N_10491,N_9324,N_9938);
xor U10492 (N_10492,N_5757,N_9207);
nand U10493 (N_10493,N_9949,N_8394);
or U10494 (N_10494,N_9572,N_5623);
or U10495 (N_10495,N_8783,N_7619);
nand U10496 (N_10496,N_7860,N_7030);
nand U10497 (N_10497,N_9588,N_7607);
or U10498 (N_10498,N_8570,N_9597);
xor U10499 (N_10499,N_8278,N_8946);
nor U10500 (N_10500,N_9792,N_9174);
nor U10501 (N_10501,N_8147,N_5166);
xnor U10502 (N_10502,N_6439,N_5692);
nand U10503 (N_10503,N_5567,N_6729);
nand U10504 (N_10504,N_9416,N_7192);
nor U10505 (N_10505,N_8964,N_5011);
and U10506 (N_10506,N_8304,N_7048);
nor U10507 (N_10507,N_8760,N_9905);
or U10508 (N_10508,N_7067,N_5975);
and U10509 (N_10509,N_5156,N_8030);
nor U10510 (N_10510,N_5165,N_6723);
or U10511 (N_10511,N_9409,N_9408);
and U10512 (N_10512,N_6002,N_6345);
and U10513 (N_10513,N_7203,N_7757);
and U10514 (N_10514,N_6184,N_5684);
and U10515 (N_10515,N_8919,N_5241);
nand U10516 (N_10516,N_9166,N_9190);
or U10517 (N_10517,N_7238,N_7749);
or U10518 (N_10518,N_8633,N_5618);
or U10519 (N_10519,N_8057,N_8181);
xor U10520 (N_10520,N_6302,N_7615);
nand U10521 (N_10521,N_5475,N_8442);
or U10522 (N_10522,N_6510,N_6946);
nor U10523 (N_10523,N_5118,N_6611);
and U10524 (N_10524,N_9055,N_7699);
and U10525 (N_10525,N_6167,N_5950);
or U10526 (N_10526,N_9890,N_6780);
xor U10527 (N_10527,N_6115,N_8639);
nor U10528 (N_10528,N_9708,N_9483);
and U10529 (N_10529,N_6091,N_7066);
nor U10530 (N_10530,N_5383,N_7473);
and U10531 (N_10531,N_5862,N_6846);
or U10532 (N_10532,N_7732,N_7086);
and U10533 (N_10533,N_5614,N_5720);
or U10534 (N_10534,N_6855,N_6745);
nor U10535 (N_10535,N_5689,N_7312);
and U10536 (N_10536,N_8944,N_9642);
and U10537 (N_10537,N_5412,N_5106);
xor U10538 (N_10538,N_8098,N_5911);
nor U10539 (N_10539,N_6544,N_6457);
xnor U10540 (N_10540,N_7393,N_6440);
and U10541 (N_10541,N_6709,N_5318);
or U10542 (N_10542,N_9341,N_9313);
and U10543 (N_10543,N_8550,N_9846);
or U10544 (N_10544,N_5244,N_5292);
and U10545 (N_10545,N_8101,N_5393);
and U10546 (N_10546,N_8109,N_9192);
or U10547 (N_10547,N_5916,N_7786);
and U10548 (N_10548,N_8271,N_9360);
nor U10549 (N_10549,N_9807,N_9978);
or U10550 (N_10550,N_7540,N_7600);
or U10551 (N_10551,N_9384,N_9874);
or U10552 (N_10552,N_7646,N_6806);
and U10553 (N_10553,N_9880,N_6106);
and U10554 (N_10554,N_5796,N_9566);
or U10555 (N_10555,N_5514,N_8035);
xnor U10556 (N_10556,N_7543,N_7813);
nand U10557 (N_10557,N_9020,N_7727);
xnor U10558 (N_10558,N_8692,N_9544);
nor U10559 (N_10559,N_6226,N_6520);
xor U10560 (N_10560,N_7406,N_6347);
or U10561 (N_10561,N_5575,N_5873);
xnor U10562 (N_10562,N_6144,N_7909);
nor U10563 (N_10563,N_9617,N_8879);
or U10564 (N_10564,N_7398,N_7598);
nand U10565 (N_10565,N_6866,N_7480);
nor U10566 (N_10566,N_6437,N_6240);
nand U10567 (N_10567,N_8845,N_5065);
or U10568 (N_10568,N_7530,N_7319);
xor U10569 (N_10569,N_6526,N_7226);
and U10570 (N_10570,N_7057,N_8154);
xor U10571 (N_10571,N_5770,N_9109);
and U10572 (N_10572,N_6596,N_8367);
nand U10573 (N_10573,N_6997,N_7161);
nand U10574 (N_10574,N_8309,N_8253);
xor U10575 (N_10575,N_6685,N_9035);
and U10576 (N_10576,N_9461,N_8587);
nand U10577 (N_10577,N_6355,N_8636);
nor U10578 (N_10578,N_6003,N_9314);
or U10579 (N_10579,N_5877,N_9661);
xnor U10580 (N_10580,N_6172,N_9689);
or U10581 (N_10581,N_7077,N_8129);
nand U10582 (N_10582,N_6076,N_5520);
xor U10583 (N_10583,N_9859,N_7037);
and U10584 (N_10584,N_5826,N_6234);
nor U10585 (N_10585,N_8112,N_5937);
nor U10586 (N_10586,N_7177,N_8015);
and U10587 (N_10587,N_5330,N_8562);
nor U10588 (N_10588,N_6238,N_5972);
xor U10589 (N_10589,N_8493,N_7908);
nand U10590 (N_10590,N_8564,N_5470);
xor U10591 (N_10591,N_9755,N_5429);
nor U10592 (N_10592,N_9434,N_8202);
or U10593 (N_10593,N_6393,N_9587);
nor U10594 (N_10594,N_5442,N_9608);
nor U10595 (N_10595,N_8274,N_5333);
and U10596 (N_10596,N_9516,N_7242);
nor U10597 (N_10597,N_8482,N_9478);
and U10598 (N_10598,N_9244,N_9464);
and U10599 (N_10599,N_8876,N_6196);
xor U10600 (N_10600,N_6695,N_5854);
and U10601 (N_10601,N_9309,N_6597);
or U10602 (N_10602,N_5842,N_8089);
xor U10603 (N_10603,N_9315,N_9466);
and U10604 (N_10604,N_5679,N_8012);
or U10605 (N_10605,N_6578,N_5787);
or U10606 (N_10606,N_5786,N_5423);
nand U10607 (N_10607,N_8530,N_8655);
xnor U10608 (N_10608,N_6273,N_5728);
nor U10609 (N_10609,N_8821,N_8353);
or U10610 (N_10610,N_5527,N_6102);
nor U10611 (N_10611,N_6079,N_8287);
nand U10612 (N_10612,N_5712,N_5197);
nand U10613 (N_10613,N_7785,N_9512);
and U10614 (N_10614,N_5841,N_7477);
nor U10615 (N_10615,N_5955,N_8479);
nand U10616 (N_10616,N_5987,N_6852);
or U10617 (N_10617,N_8940,N_5117);
nand U10618 (N_10618,N_5560,N_5744);
xnor U10619 (N_10619,N_5903,N_7023);
or U10620 (N_10620,N_9509,N_8252);
or U10621 (N_10621,N_5593,N_8890);
nor U10622 (N_10622,N_6423,N_7780);
and U10623 (N_10623,N_5875,N_8723);
and U10624 (N_10624,N_9243,N_5817);
or U10625 (N_10625,N_5367,N_9071);
nand U10626 (N_10626,N_8901,N_7625);
nor U10627 (N_10627,N_6814,N_9017);
and U10628 (N_10628,N_6262,N_9006);
xor U10629 (N_10629,N_7837,N_5792);
nand U10630 (N_10630,N_7674,N_8439);
xnor U10631 (N_10631,N_8403,N_7994);
and U10632 (N_10632,N_6921,N_6323);
and U10633 (N_10633,N_5557,N_9284);
xor U10634 (N_10634,N_6646,N_8515);
and U10635 (N_10635,N_5436,N_6053);
or U10636 (N_10636,N_7642,N_8673);
nor U10637 (N_10637,N_7670,N_7795);
and U10638 (N_10638,N_5688,N_9678);
xor U10639 (N_10639,N_9052,N_6485);
or U10640 (N_10640,N_8390,N_6453);
nor U10641 (N_10641,N_8973,N_9220);
or U10642 (N_10642,N_5600,N_6636);
xnor U10643 (N_10643,N_6706,N_7534);
or U10644 (N_10644,N_6208,N_8941);
and U10645 (N_10645,N_8350,N_8660);
and U10646 (N_10646,N_9280,N_7120);
nor U10647 (N_10647,N_5462,N_6573);
nor U10648 (N_10648,N_8994,N_5425);
and U10649 (N_10649,N_7881,N_5702);
or U10650 (N_10650,N_5431,N_8558);
and U10651 (N_10651,N_9983,N_9021);
nor U10652 (N_10652,N_5306,N_5497);
xor U10653 (N_10653,N_7126,N_8934);
nor U10654 (N_10654,N_9827,N_6802);
or U10655 (N_10655,N_5382,N_8610);
xor U10656 (N_10656,N_7110,N_8428);
and U10657 (N_10657,N_7429,N_8688);
xor U10658 (N_10658,N_9665,N_7889);
nor U10659 (N_10659,N_6977,N_9547);
nand U10660 (N_10660,N_9710,N_7367);
nor U10661 (N_10661,N_7141,N_8484);
nor U10662 (N_10662,N_7825,N_9063);
nand U10663 (N_10663,N_8438,N_5970);
or U10664 (N_10664,N_5266,N_7497);
nand U10665 (N_10665,N_8474,N_7580);
or U10666 (N_10666,N_8494,N_8279);
xor U10667 (N_10667,N_8397,N_6069);
xnor U10668 (N_10668,N_5095,N_9718);
nor U10669 (N_10669,N_8594,N_6188);
or U10670 (N_10670,N_5805,N_9059);
or U10671 (N_10671,N_5384,N_6595);
nor U10672 (N_10672,N_6378,N_8327);
xnor U10673 (N_10673,N_5724,N_5628);
or U10674 (N_10674,N_5346,N_5579);
nor U10675 (N_10675,N_9367,N_7505);
xnor U10676 (N_10676,N_5681,N_9823);
and U10677 (N_10677,N_5355,N_9351);
nor U10678 (N_10678,N_9200,N_5336);
xor U10679 (N_10679,N_8667,N_5853);
and U10680 (N_10680,N_5405,N_7941);
nor U10681 (N_10681,N_7353,N_8388);
nor U10682 (N_10682,N_8345,N_8715);
or U10683 (N_10683,N_8580,N_7956);
nand U10684 (N_10684,N_9070,N_7479);
xor U10685 (N_10685,N_9312,N_6662);
nor U10686 (N_10686,N_6417,N_9585);
nand U10687 (N_10687,N_6392,N_9060);
and U10688 (N_10688,N_5504,N_8711);
and U10689 (N_10689,N_6452,N_7687);
and U10690 (N_10690,N_5779,N_6562);
and U10691 (N_10691,N_9686,N_7491);
nand U10692 (N_10692,N_5529,N_7784);
nor U10693 (N_10693,N_7754,N_7088);
or U10694 (N_10694,N_7822,N_8526);
or U10695 (N_10695,N_7073,N_8571);
or U10696 (N_10696,N_9354,N_9803);
nor U10697 (N_10697,N_7043,N_8800);
or U10698 (N_10698,N_8045,N_6530);
nand U10699 (N_10699,N_6293,N_6620);
nor U10700 (N_10700,N_9250,N_5120);
and U10701 (N_10701,N_5344,N_9829);
xor U10702 (N_10702,N_8702,N_6449);
and U10703 (N_10703,N_5985,N_9594);
and U10704 (N_10704,N_8574,N_8004);
and U10705 (N_10705,N_9387,N_8140);
nor U10706 (N_10706,N_9799,N_7389);
or U10707 (N_10707,N_9119,N_9716);
nor U10708 (N_10708,N_5123,N_6896);
nand U10709 (N_10709,N_7817,N_5104);
nand U10710 (N_10710,N_8044,N_8312);
nand U10711 (N_10711,N_7893,N_7286);
xnor U10712 (N_10712,N_9835,N_9981);
nand U10713 (N_10713,N_8362,N_8720);
nor U10714 (N_10714,N_5730,N_8820);
or U10715 (N_10715,N_5886,N_8092);
nand U10716 (N_10716,N_9833,N_8199);
nand U10717 (N_10717,N_9879,N_7408);
nor U10718 (N_10718,N_8915,N_5797);
or U10719 (N_10719,N_8782,N_9222);
and U10720 (N_10720,N_6067,N_9954);
xnor U10721 (N_10721,N_7267,N_8881);
nor U10722 (N_10722,N_9783,N_8346);
nand U10723 (N_10723,N_9528,N_8398);
xor U10724 (N_10724,N_6909,N_8434);
or U10725 (N_10725,N_9178,N_7151);
nand U10726 (N_10726,N_8522,N_8975);
or U10727 (N_10727,N_9674,N_6146);
nand U10728 (N_10728,N_9379,N_5624);
xor U10729 (N_10729,N_8488,N_7239);
and U10730 (N_10730,N_8062,N_5857);
and U10731 (N_10731,N_8424,N_9014);
nand U10732 (N_10732,N_9331,N_5583);
nand U10733 (N_10733,N_7377,N_8452);
and U10734 (N_10734,N_7623,N_7133);
nor U10735 (N_10735,N_9573,N_7422);
or U10736 (N_10736,N_9866,N_6168);
and U10737 (N_10737,N_7009,N_7527);
xor U10738 (N_10738,N_5735,N_7849);
nand U10739 (N_10739,N_9984,N_8518);
nand U10740 (N_10740,N_6157,N_8556);
or U10741 (N_10741,N_7257,N_7324);
nand U10742 (N_10742,N_5799,N_6033);
nand U10743 (N_10743,N_8641,N_6650);
xor U10744 (N_10744,N_9073,N_9366);
nor U10745 (N_10745,N_7759,N_5362);
nor U10746 (N_10746,N_9903,N_7546);
and U10747 (N_10747,N_7627,N_8954);
and U10748 (N_10748,N_8292,N_8959);
nor U10749 (N_10749,N_6360,N_8785);
and U10750 (N_10750,N_5240,N_7248);
xor U10751 (N_10751,N_7117,N_9857);
nor U10752 (N_10752,N_5395,N_8805);
and U10753 (N_10753,N_5556,N_5268);
xor U10754 (N_10754,N_5769,N_6627);
and U10755 (N_10755,N_6898,N_7496);
or U10756 (N_10756,N_6153,N_7346);
xor U10757 (N_10757,N_5347,N_8481);
or U10758 (N_10758,N_8951,N_8840);
xor U10759 (N_10759,N_7153,N_5150);
nor U10760 (N_10760,N_9162,N_6812);
nor U10761 (N_10761,N_5619,N_8884);
nor U10762 (N_10762,N_9397,N_5536);
and U10763 (N_10763,N_9453,N_9717);
nand U10764 (N_10764,N_6049,N_5634);
nor U10765 (N_10765,N_5607,N_7287);
or U10766 (N_10766,N_7033,N_5169);
xor U10767 (N_10767,N_7155,N_6004);
xnor U10768 (N_10768,N_7557,N_5328);
and U10769 (N_10769,N_5114,N_5510);
or U10770 (N_10770,N_9995,N_6971);
nor U10771 (N_10771,N_8678,N_6842);
nand U10772 (N_10772,N_9259,N_7590);
nor U10773 (N_10773,N_5936,N_5190);
nor U10774 (N_10774,N_9558,N_6694);
xor U10775 (N_10775,N_8843,N_6515);
and U10776 (N_10776,N_7090,N_5865);
nand U10777 (N_10777,N_5049,N_7047);
nor U10778 (N_10778,N_8361,N_7440);
or U10779 (N_10779,N_6728,N_8366);
or U10780 (N_10780,N_6222,N_7083);
and U10781 (N_10781,N_5243,N_7566);
xor U10782 (N_10782,N_6258,N_5498);
xor U10783 (N_10783,N_7096,N_5324);
and U10784 (N_10784,N_7603,N_9676);
and U10785 (N_10785,N_6681,N_9917);
and U10786 (N_10786,N_9037,N_8646);
nor U10787 (N_10787,N_7256,N_7163);
and U10788 (N_10788,N_7062,N_7733);
xor U10789 (N_10789,N_8049,N_7721);
nor U10790 (N_10790,N_5981,N_7028);
or U10791 (N_10791,N_5021,N_5844);
or U10792 (N_10792,N_5135,N_5316);
or U10793 (N_10793,N_9053,N_9411);
nand U10794 (N_10794,N_6561,N_7474);
nor U10795 (N_10795,N_9427,N_6622);
or U10796 (N_10796,N_6583,N_8213);
and U10797 (N_10797,N_7297,N_6478);
or U10798 (N_10798,N_6236,N_7745);
xnor U10799 (N_10799,N_6014,N_6394);
xnor U10800 (N_10800,N_9441,N_8575);
nand U10801 (N_10801,N_8717,N_6868);
nor U10802 (N_10802,N_5145,N_8236);
xor U10803 (N_10803,N_7224,N_9278);
nor U10804 (N_10804,N_6567,N_5016);
nor U10805 (N_10805,N_5280,N_8407);
nor U10806 (N_10806,N_8107,N_9135);
nand U10807 (N_10807,N_5503,N_9920);
xnor U10808 (N_10808,N_7675,N_8237);
nand U10809 (N_10809,N_7658,N_5040);
or U10810 (N_10810,N_7917,N_7631);
xnor U10811 (N_10811,N_7696,N_8450);
or U10812 (N_10812,N_8979,N_8175);
or U10813 (N_10813,N_5063,N_9414);
xnor U10814 (N_10814,N_7164,N_8541);
nor U10815 (N_10815,N_9326,N_8334);
nor U10816 (N_10816,N_8313,N_9143);
nand U10817 (N_10817,N_6082,N_5050);
nand U10818 (N_10818,N_5254,N_8922);
or U10819 (N_10819,N_6329,N_7960);
and U10820 (N_10820,N_8208,N_7129);
nor U10821 (N_10821,N_7433,N_6287);
nor U10822 (N_10822,N_6982,N_9470);
or U10823 (N_10823,N_9836,N_6404);
nand U10824 (N_10824,N_9636,N_7574);
and U10825 (N_10825,N_6555,N_9018);
nand U10826 (N_10826,N_8732,N_7575);
or U10827 (N_10827,N_8227,N_7684);
nand U10828 (N_10828,N_7790,N_8275);
xnor U10829 (N_10829,N_8757,N_9067);
nor U10830 (N_10830,N_8740,N_6488);
and U10831 (N_10831,N_6585,N_9508);
nand U10832 (N_10832,N_5180,N_5224);
or U10833 (N_10833,N_9974,N_9270);
or U10834 (N_10834,N_9130,N_7318);
nor U10835 (N_10835,N_9094,N_6135);
xnor U10836 (N_10836,N_6823,N_9959);
nor U10837 (N_10837,N_8023,N_5666);
or U10838 (N_10838,N_5143,N_5926);
nand U10839 (N_10839,N_9425,N_6476);
nand U10840 (N_10840,N_5790,N_8811);
or U10841 (N_10841,N_7833,N_6327);
nor U10842 (N_10842,N_5249,N_9136);
nand U10843 (N_10843,N_8856,N_8095);
and U10844 (N_10844,N_5708,N_8435);
or U10845 (N_10845,N_5785,N_7700);
and U10846 (N_10846,N_8409,N_7445);
nor U10847 (N_10847,N_8013,N_9238);
xor U10848 (N_10848,N_6575,N_7880);
nor U10849 (N_10849,N_6778,N_5125);
or U10850 (N_10850,N_6604,N_6177);
and U10851 (N_10851,N_5247,N_5784);
and U10852 (N_10852,N_5205,N_8848);
nand U10853 (N_10853,N_9979,N_9062);
and U10854 (N_10854,N_5228,N_6145);
and U10855 (N_10855,N_6395,N_7121);
nand U10856 (N_10856,N_6985,N_7476);
nand U10857 (N_10857,N_7413,N_8892);
nand U10858 (N_10858,N_7425,N_8900);
or U10859 (N_10859,N_7997,N_9040);
or U10860 (N_10860,N_8490,N_5766);
nand U10861 (N_10861,N_9448,N_5909);
and U10862 (N_10862,N_6487,N_8828);
nor U10863 (N_10863,N_8480,N_8106);
and U10864 (N_10864,N_7847,N_5731);
xor U10865 (N_10865,N_6845,N_6960);
and U10866 (N_10866,N_6116,N_9796);
nor U10867 (N_10867,N_9003,N_5162);
or U10868 (N_10868,N_8352,N_5706);
nor U10869 (N_10869,N_8725,N_9118);
xor U10870 (N_10870,N_5357,N_7787);
xnor U10871 (N_10871,N_6692,N_6905);
nor U10872 (N_10872,N_7985,N_7697);
nand U10873 (N_10873,N_7525,N_7115);
nor U10874 (N_10874,N_5908,N_7410);
xor U10875 (N_10875,N_8348,N_9311);
or U10876 (N_10876,N_9462,N_8921);
nand U10877 (N_10877,N_7812,N_9265);
xor U10878 (N_10878,N_9941,N_7723);
nor U10879 (N_10879,N_6867,N_9561);
nand U10880 (N_10880,N_6407,N_6397);
xnor U10881 (N_10881,N_9486,N_9177);
nand U10882 (N_10882,N_8709,N_6048);
nand U10883 (N_10883,N_7639,N_9707);
nand U10884 (N_10884,N_7100,N_5435);
xor U10885 (N_10885,N_6467,N_9026);
or U10886 (N_10886,N_8449,N_5749);
and U10887 (N_10887,N_8273,N_7407);
and U10888 (N_10888,N_9390,N_5694);
or U10889 (N_10889,N_7314,N_6853);
xnor U10890 (N_10890,N_8670,N_9320);
nor U10891 (N_10891,N_8277,N_6242);
or U10892 (N_10892,N_5777,N_8573);
nor U10893 (N_10893,N_5929,N_9513);
nor U10894 (N_10894,N_5810,N_5474);
nor U10895 (N_10895,N_5420,N_6294);
or U10896 (N_10896,N_9179,N_9444);
nand U10897 (N_10897,N_8118,N_6796);
and U10898 (N_10898,N_8671,N_5294);
nand U10899 (N_10899,N_6263,N_9418);
xnor U10900 (N_10900,N_5245,N_5872);
or U10901 (N_10901,N_6031,N_9683);
or U10902 (N_10902,N_8592,N_7241);
and U10903 (N_10903,N_8116,N_5437);
or U10904 (N_10904,N_9667,N_8528);
xor U10905 (N_10905,N_9745,N_7899);
nand U10906 (N_10906,N_7736,N_6154);
and U10907 (N_10907,N_9632,N_5163);
and U10908 (N_10908,N_5915,N_6833);
nor U10909 (N_10909,N_7630,N_5043);
xnor U10910 (N_10910,N_8708,N_5923);
and U10911 (N_10911,N_6386,N_7015);
or U10912 (N_10912,N_6305,N_9080);
or U10913 (N_10913,N_7400,N_7189);
nand U10914 (N_10914,N_6647,N_7944);
and U10915 (N_10915,N_8364,N_6344);
xnor U10916 (N_10916,N_9851,N_9184);
nand U10917 (N_10917,N_8315,N_7092);
and U10918 (N_10918,N_5407,N_7570);
nor U10919 (N_10919,N_7840,N_9001);
nor U10920 (N_10920,N_6320,N_7358);
nand U10921 (N_10921,N_9450,N_9237);
and U10922 (N_10922,N_7140,N_5531);
xor U10923 (N_10923,N_9815,N_7891);
nor U10924 (N_10924,N_6968,N_7489);
or U10925 (N_10925,N_6284,N_9555);
or U10926 (N_10926,N_9655,N_7265);
xor U10927 (N_10927,N_7850,N_8835);
xnor U10928 (N_10928,N_8579,N_9554);
nor U10929 (N_10929,N_5781,N_8565);
nor U10930 (N_10930,N_6479,N_5387);
xor U10931 (N_10931,N_6422,N_5677);
or U10932 (N_10932,N_5396,N_9987);
nor U10933 (N_10933,N_7686,N_6164);
or U10934 (N_10934,N_5839,N_6752);
nand U10935 (N_10935,N_7482,N_5661);
nand U10936 (N_10936,N_8815,N_5402);
nor U10937 (N_10937,N_5956,N_6326);
xor U10938 (N_10938,N_6107,N_5765);
and U10939 (N_10939,N_6333,N_9915);
nand U10940 (N_10940,N_5615,N_7870);
xor U10941 (N_10941,N_8916,N_7991);
and U10942 (N_10942,N_7448,N_8032);
nand U10943 (N_10943,N_5538,N_7648);
nand U10944 (N_10944,N_6195,N_7150);
xnor U10945 (N_10945,N_7585,N_8234);
xor U10946 (N_10946,N_6176,N_7487);
nand U10947 (N_10947,N_6926,N_8099);
nor U10948 (N_10948,N_8658,N_5444);
nand U10949 (N_10949,N_8989,N_6251);
nand U10950 (N_10950,N_8371,N_5540);
and U10951 (N_10951,N_8585,N_5272);
nor U10952 (N_10952,N_8318,N_8323);
xnor U10953 (N_10953,N_9977,N_5783);
or U10954 (N_10954,N_5732,N_9318);
xnor U10955 (N_10955,N_6220,N_9629);
xnor U10956 (N_10956,N_6840,N_8661);
or U10957 (N_10957,N_5035,N_9909);
or U10958 (N_10958,N_8259,N_5870);
nor U10959 (N_10959,N_8985,N_8103);
and U10960 (N_10960,N_9589,N_5979);
or U10961 (N_10961,N_7641,N_5427);
nand U10962 (N_10962,N_7737,N_8981);
nand U10963 (N_10963,N_7612,N_8663);
nor U10964 (N_10964,N_9383,N_7194);
or U10965 (N_10965,N_7438,N_6103);
xor U10966 (N_10966,N_7872,N_7229);
nor U10967 (N_10967,N_5409,N_7344);
or U10968 (N_10968,N_7419,N_6203);
nor U10969 (N_10969,N_6368,N_9282);
nor U10970 (N_10970,N_6776,N_8086);
nor U10971 (N_10971,N_9031,N_9404);
xor U10972 (N_10972,N_5102,N_6358);
xnor U10973 (N_10973,N_7345,N_6429);
xnor U10974 (N_10974,N_6829,N_5454);
xor U10975 (N_10975,N_8902,N_6083);
and U10976 (N_10976,N_7387,N_6147);
or U10977 (N_10977,N_6489,N_9600);
nand U10978 (N_10978,N_5986,N_5314);
or U10979 (N_10979,N_9654,N_7826);
or U10980 (N_10980,N_7810,N_9342);
and U10981 (N_10981,N_5234,N_6911);
xor U10982 (N_10982,N_6908,N_6710);
xor U10983 (N_10983,N_7210,N_8917);
or U10984 (N_10984,N_9507,N_9991);
and U10985 (N_10985,N_6384,N_9649);
nor U10986 (N_10986,N_6995,N_7227);
nand U10987 (N_10987,N_5824,N_5562);
nor U10988 (N_10988,N_6420,N_9732);
and U10989 (N_10989,N_9641,N_6124);
and U10990 (N_10990,N_7828,N_9885);
xnor U10991 (N_10991,N_9047,N_7499);
xor U10992 (N_10992,N_8672,N_6486);
and U10993 (N_10993,N_8158,N_6667);
nand U10994 (N_10994,N_9525,N_5670);
and U10995 (N_10995,N_7982,N_8824);
and U10996 (N_10996,N_6459,N_8582);
and U10997 (N_10997,N_9170,N_7412);
nor U10998 (N_10998,N_9578,N_8052);
or U10999 (N_10999,N_9111,N_6274);
nor U11000 (N_11000,N_5532,N_5134);
or U11001 (N_11001,N_9407,N_7171);
xnor U11002 (N_11002,N_9791,N_7056);
and U11003 (N_11003,N_7604,N_9942);
and U11004 (N_11004,N_9840,N_5301);
nand U11005 (N_11005,N_9025,N_5738);
nand U11006 (N_11006,N_9064,N_6292);
nand U11007 (N_11007,N_7041,N_6531);
nor U11008 (N_11008,N_9254,N_7636);
nor U11009 (N_11009,N_5248,N_6762);
xor U11010 (N_11010,N_6272,N_5299);
nor U11011 (N_11011,N_9606,N_6649);
nand U11012 (N_11012,N_9317,N_7220);
and U11013 (N_11013,N_9110,N_5919);
xor U11014 (N_11014,N_8491,N_6010);
or U11015 (N_11015,N_7122,N_9127);
xor U11016 (N_11016,N_6191,N_8774);
xor U11017 (N_11017,N_5690,N_5325);
nor U11018 (N_11018,N_6398,N_5795);
and U11019 (N_11019,N_5918,N_5229);
nor U11020 (N_11020,N_5465,N_7020);
and U11021 (N_11021,N_7616,N_6787);
xnor U11022 (N_11022,N_8151,N_8019);
xor U11023 (N_11023,N_7304,N_9385);
nand U11024 (N_11024,N_7632,N_6614);
xor U11025 (N_11025,N_7962,N_8882);
nor U11026 (N_11026,N_7844,N_5499);
xor U11027 (N_11027,N_7275,N_8301);
and U11028 (N_11028,N_8502,N_9723);
nor U11029 (N_11029,N_9626,N_9861);
xor U11030 (N_11030,N_7720,N_8150);
xor U11031 (N_11031,N_9531,N_5552);
xnor U11032 (N_11032,N_8699,N_7827);
xnor U11033 (N_11033,N_5217,N_7934);
and U11034 (N_11034,N_5417,N_5385);
nor U11035 (N_11035,N_8751,N_7253);
nor U11036 (N_11036,N_9832,N_8754);
nand U11037 (N_11037,N_5309,N_5237);
or U11038 (N_11038,N_5639,N_5855);
nand U11039 (N_11039,N_5332,N_6092);
or U11040 (N_11040,N_6735,N_5426);
nor U11041 (N_11041,N_8700,N_6629);
or U11042 (N_11042,N_5210,N_6906);
nand U11043 (N_11043,N_9010,N_9551);
or U11044 (N_11044,N_8048,N_5509);
nand U11045 (N_11045,N_6181,N_5460);
or U11046 (N_11046,N_7486,N_7715);
nand U11047 (N_11047,N_5945,N_5664);
and U11048 (N_11048,N_6425,N_5778);
nor U11049 (N_11049,N_7526,N_9898);
nand U11050 (N_11050,N_7659,N_8248);
nor U11051 (N_11051,N_9908,N_6862);
xnor U11052 (N_11052,N_9615,N_5847);
nor U11053 (N_11053,N_8545,N_7948);
and U11054 (N_11054,N_8878,N_7541);
xnor U11055 (N_11055,N_8083,N_7446);
xnor U11056 (N_11056,N_7968,N_9943);
nor U11057 (N_11057,N_5060,N_5629);
nand U11058 (N_11058,N_5519,N_5055);
nand U11059 (N_11059,N_7490,N_6020);
and U11060 (N_11060,N_8860,N_7202);
nand U11061 (N_11061,N_9788,N_6482);
nand U11062 (N_11062,N_7080,N_8445);
nand U11063 (N_11063,N_9161,N_8997);
and U11064 (N_11064,N_9930,N_8389);
xor U11065 (N_11065,N_8666,N_5622);
or U11066 (N_11066,N_8517,N_6070);
and U11067 (N_11067,N_7942,N_8643);
and U11068 (N_11068,N_7018,N_9782);
or U11069 (N_11069,N_7717,N_9474);
or U11070 (N_11070,N_6978,N_6490);
xnor U11071 (N_11071,N_7694,N_9310);
xor U11072 (N_11072,N_8363,N_5845);
nand U11073 (N_11073,N_8539,N_5469);
or U11074 (N_11074,N_8467,N_9344);
xor U11075 (N_11075,N_8729,N_7074);
nor U11076 (N_11076,N_8906,N_8295);
xor U11077 (N_11077,N_8139,N_5350);
and U11078 (N_11078,N_9000,N_6539);
nand U11079 (N_11079,N_5947,N_7762);
and U11080 (N_11080,N_5477,N_9424);
nor U11081 (N_11081,N_7051,N_5007);
and U11082 (N_11082,N_7957,N_7556);
nand U11083 (N_11083,N_7638,N_5461);
nor U11084 (N_11084,N_5726,N_8091);
or U11085 (N_11085,N_8413,N_9400);
and U11086 (N_11086,N_8257,N_7913);
and U11087 (N_11087,N_7036,N_9830);
or U11088 (N_11088,N_5904,N_6475);
or U11089 (N_11089,N_9962,N_6805);
and U11090 (N_11090,N_6955,N_9534);
and U11091 (N_11091,N_7888,N_9234);
nor U11092 (N_11092,N_6899,N_7910);
nand U11093 (N_11093,N_9381,N_6799);
and U11094 (N_11094,N_5883,N_6838);
or U11095 (N_11095,N_7829,N_5296);
or U11096 (N_11096,N_6113,N_7232);
and U11097 (N_11097,N_5121,N_6795);
xnor U11098 (N_11098,N_7200,N_5051);
nand U11099 (N_11099,N_8485,N_9332);
xor U11100 (N_11100,N_9787,N_8513);
and U11101 (N_11101,N_7510,N_5714);
and U11102 (N_11102,N_7702,N_9771);
nor U11103 (N_11103,N_8788,N_7235);
nand U11104 (N_11104,N_5380,N_5852);
xnor U11105 (N_11105,N_7251,N_8280);
nand U11106 (N_11106,N_6742,N_7094);
and U11107 (N_11107,N_9709,N_8061);
or U11108 (N_11108,N_5105,N_8395);
nand U11109 (N_11109,N_6295,N_8798);
or U11110 (N_11110,N_5273,N_6558);
nand U11111 (N_11111,N_9058,N_8070);
nand U11112 (N_11112,N_7743,N_9261);
or U11113 (N_11113,N_6543,N_5832);
nand U11114 (N_11114,N_5109,N_9729);
and U11115 (N_11115,N_6616,N_8126);
or U11116 (N_11116,N_7415,N_8615);
or U11117 (N_11117,N_7753,N_5232);
or U11118 (N_11118,N_8470,N_9849);
xnor U11119 (N_11119,N_9818,N_5746);
xor U11120 (N_11120,N_9742,N_5548);
or U11121 (N_11121,N_5816,N_6095);
or U11122 (N_11122,N_6052,N_9215);
and U11123 (N_11123,N_7892,N_9072);
and U11124 (N_11124,N_7401,N_5626);
or U11125 (N_11125,N_6035,N_7537);
and U11126 (N_11126,N_8647,N_8516);
nand U11127 (N_11127,N_8873,N_7098);
xor U11128 (N_11128,N_9697,N_7230);
and U11129 (N_11129,N_8110,N_6089);
xor U11130 (N_11130,N_9881,N_8802);
nand U11131 (N_11131,N_9994,N_9245);
xor U11132 (N_11132,N_5608,N_8786);
xor U11133 (N_11133,N_9936,N_8795);
or U11134 (N_11134,N_8483,N_8852);
nor U11135 (N_11135,N_7976,N_5378);
and U11136 (N_11136,N_9115,N_8950);
and U11137 (N_11137,N_7370,N_9504);
and U11138 (N_11138,N_9012,N_9002);
xnor U11139 (N_11139,N_8400,N_5459);
or U11140 (N_11140,N_6149,N_5484);
nor U11141 (N_11141,N_7052,N_7512);
xnor U11142 (N_11142,N_7589,N_8896);
or U11143 (N_11143,N_7315,N_6945);
or U11144 (N_11144,N_7602,N_9848);
and U11145 (N_11145,N_6625,N_7965);
nor U11146 (N_11146,N_6199,N_9816);
nand U11147 (N_11147,N_5124,N_7284);
and U11148 (N_11148,N_8447,N_5211);
nor U11149 (N_11149,N_6455,N_9552);
and U11150 (N_11150,N_8425,N_8649);
nor U11151 (N_11151,N_6474,N_7139);
xnor U11152 (N_11152,N_7168,N_6356);
xor U11153 (N_11153,N_7363,N_9650);
and U11154 (N_11154,N_5791,N_6441);
nand U11155 (N_11155,N_8662,N_6374);
or U11156 (N_11156,N_7955,N_9451);
nand U11157 (N_11157,N_7945,N_6809);
nor U11158 (N_11158,N_7116,N_9182);
xor U11159 (N_11159,N_5943,N_6606);
nand U11160 (N_11160,N_7426,N_6418);
nor U11161 (N_11161,N_9773,N_5263);
xnor U11162 (N_11162,N_7678,N_6093);
nand U11163 (N_11163,N_6581,N_9730);
and U11164 (N_11164,N_6973,N_7313);
and U11165 (N_11165,N_9795,N_5451);
and U11166 (N_11166,N_6313,N_8778);
nor U11167 (N_11167,N_9210,N_7134);
or U11168 (N_11168,N_8868,N_8791);
and U11169 (N_11169,N_5269,N_6064);
nand U11170 (N_11170,N_7170,N_7162);
and U11171 (N_11171,N_5992,N_7097);
or U11172 (N_11172,N_6713,N_8408);
or U11173 (N_11173,N_7231,N_9492);
nand U11174 (N_11174,N_6612,N_6661);
nand U11175 (N_11175,N_9357,N_6654);
and U11176 (N_11176,N_7093,N_8842);
and U11177 (N_11177,N_9677,N_6245);
xnor U11178 (N_11178,N_8281,N_8664);
nand U11179 (N_11179,N_5602,N_9426);
and U11180 (N_11180,N_5545,N_7017);
nor U11181 (N_11181,N_6005,N_8903);
and U11182 (N_11182,N_6330,N_7298);
nor U11183 (N_11183,N_5297,N_9124);
xor U11184 (N_11184,N_8368,N_8223);
or U11185 (N_11185,N_9069,N_9435);
xor U11186 (N_11186,N_7321,N_5905);
xnor U11187 (N_11187,N_9117,N_6361);
or U11188 (N_11188,N_7740,N_5780);
nor U11189 (N_11189,N_8907,N_5658);
or U11190 (N_11190,N_8351,N_5804);
or U11191 (N_11191,N_6632,N_5450);
or U11192 (N_11192,N_9479,N_9279);
nor U11193 (N_11193,N_6990,N_8018);
xor U11194 (N_11194,N_9319,N_7854);
and U11195 (N_11195,N_8160,N_6150);
xor U11196 (N_11196,N_7853,N_9160);
nand U11197 (N_11197,N_9785,N_8625);
and U11198 (N_11198,N_7640,N_6410);
and U11199 (N_11199,N_7087,N_9392);
nand U11200 (N_11200,N_5128,N_8963);
nand U11201 (N_11201,N_5995,N_6605);
nor U11202 (N_11202,N_9051,N_5096);
xor U11203 (N_11203,N_8739,N_7729);
xnor U11204 (N_11204,N_9433,N_5729);
xnor U11205 (N_11205,N_9948,N_8766);
nor U11206 (N_11206,N_8913,N_6943);
and U11207 (N_11207,N_6727,N_7016);
and U11208 (N_11208,N_6739,N_9968);
and U11209 (N_11209,N_9183,N_7952);
nor U11210 (N_11210,N_9750,N_5351);
nor U11211 (N_11211,N_8514,N_5534);
or U11212 (N_11212,N_8602,N_5067);
or U11213 (N_11213,N_6492,N_5821);
or U11214 (N_11214,N_7779,N_5754);
and U11215 (N_11215,N_5606,N_7713);
nor U11216 (N_11216,N_8713,N_9258);
or U11217 (N_11217,N_8269,N_5565);
or U11218 (N_11218,N_7774,N_5625);
nand U11219 (N_11219,N_9611,N_7988);
nor U11220 (N_11220,N_5398,N_5302);
nor U11221 (N_11221,N_7055,N_9564);
and U11222 (N_11222,N_5361,N_5523);
nand U11223 (N_11223,N_5231,N_9256);
nand U11224 (N_11224,N_9897,N_7883);
and U11225 (N_11225,N_6850,N_6498);
xnor U11226 (N_11226,N_8027,N_9926);
nand U11227 (N_11227,N_6232,N_7112);
nor U11228 (N_11228,N_6904,N_7609);
xor U11229 (N_11229,N_6794,N_5010);
xor U11230 (N_11230,N_6789,N_6648);
nor U11231 (N_11231,N_9394,N_5352);
or U11232 (N_11232,N_7127,N_6963);
nand U11233 (N_11233,N_6682,N_6377);
nand U11234 (N_11234,N_8784,N_5707);
and U11235 (N_11235,N_5535,N_6760);
and U11236 (N_11236,N_8642,N_8721);
and U11237 (N_11237,N_7493,N_6865);
and U11238 (N_11238,N_8716,N_6369);
nand U11239 (N_11239,N_5236,N_9036);
xor U11240 (N_11240,N_9752,N_7234);
and U11241 (N_11241,N_6078,N_8055);
and U11242 (N_11242,N_8054,N_9148);
nor U11243 (N_11243,N_9845,N_6288);
or U11244 (N_11244,N_9945,N_5693);
nand U11245 (N_11245,N_8559,N_9621);
nor U11246 (N_11246,N_7834,N_6480);
xnor U11247 (N_11247,N_6929,N_6925);
xor U11248 (N_11248,N_7964,N_9919);
and U11249 (N_11249,N_6382,N_6250);
nand U11250 (N_11250,N_7341,N_6910);
and U11251 (N_11251,N_7651,N_9497);
nor U11252 (N_11252,N_6882,N_5481);
nor U11253 (N_11253,N_6594,N_6421);
xnor U11254 (N_11254,N_7011,N_9330);
and U11255 (N_11255,N_5920,N_8429);
or U11256 (N_11256,N_9701,N_7350);
and U11257 (N_11257,N_6000,N_7264);
nand U11258 (N_11258,N_8402,N_8426);
or U11259 (N_11259,N_6888,N_6754);
nor U11260 (N_11260,N_8794,N_9878);
and U11261 (N_11261,N_5391,N_8335);
nor U11262 (N_11262,N_6372,N_7947);
xor U11263 (N_11263,N_9253,N_5701);
xnor U11264 (N_11264,N_7999,N_8640);
xnor U11265 (N_11265,N_5133,N_6138);
and U11266 (N_11266,N_5823,N_5809);
nand U11267 (N_11267,N_8026,N_9029);
nor U11268 (N_11268,N_5739,N_6376);
nor U11269 (N_11269,N_7544,N_6755);
or U11270 (N_11270,N_5072,N_6121);
xor U11271 (N_11271,N_8059,N_5965);
nand U11272 (N_11272,N_8512,N_7091);
or U11273 (N_11273,N_5097,N_6704);
or U11274 (N_11274,N_5610,N_5187);
or U11275 (N_11275,N_5676,N_9041);
nor U11276 (N_11276,N_9731,N_7769);
or U11277 (N_11277,N_9154,N_9302);
nor U11278 (N_11278,N_6976,N_9746);
and U11279 (N_11279,N_7989,N_8386);
xnor U11280 (N_11280,N_6998,N_8770);
and U11281 (N_11281,N_5458,N_9653);
nor U11282 (N_11282,N_5742,N_9761);
and U11283 (N_11283,N_9696,N_8858);
nand U11284 (N_11284,N_9475,N_5168);
nor U11285 (N_11285,N_6388,N_9577);
xor U11286 (N_11286,N_8769,N_7529);
xor U11287 (N_11287,N_9298,N_7060);
nand U11288 (N_11288,N_9809,N_7031);
nor U11289 (N_11289,N_5082,N_6607);
nand U11290 (N_11290,N_8451,N_7744);
nor U11291 (N_11291,N_9501,N_7399);
nor U11292 (N_11292,N_8303,N_9092);
nor U11293 (N_11293,N_5674,N_7667);
or U11294 (N_11294,N_6912,N_8060);
nand U11295 (N_11295,N_8461,N_5864);
or U11296 (N_11296,N_7677,N_8064);
nand U11297 (N_11297,N_9872,N_9568);
and U11298 (N_11298,N_6965,N_7970);
or U11299 (N_11299,N_7188,N_7375);
xor U11300 (N_11300,N_7165,N_9624);
nor U11301 (N_11301,N_9412,N_7921);
or U11302 (N_11302,N_8532,N_6570);
and U11303 (N_11303,N_6224,N_5446);
xnor U11304 (N_11304,N_6903,N_6790);
nand U11305 (N_11305,N_6891,N_9125);
and U11306 (N_11306,N_8609,N_9575);
nor U11307 (N_11307,N_5265,N_5657);
and U11308 (N_11308,N_8462,N_6271);
nor U11309 (N_11309,N_8384,N_6036);
xor U11310 (N_11310,N_8216,N_5577);
nor U11311 (N_11311,N_6690,N_8355);
nand U11312 (N_11312,N_7708,N_8986);
and U11313 (N_11313,N_8308,N_9266);
xor U11314 (N_11314,N_6712,N_6056);
xnor U11315 (N_11315,N_7882,N_8736);
or U11316 (N_11316,N_6962,N_9924);
nor U11317 (N_11317,N_7305,N_5449);
and U11318 (N_11318,N_5546,N_8730);
nand U11319 (N_11319,N_7937,N_8883);
nand U11320 (N_11320,N_7289,N_7855);
nand U11321 (N_11321,N_7245,N_9255);
or U11322 (N_11322,N_7261,N_6887);
nand U11323 (N_11323,N_9242,N_9805);
or U11324 (N_11324,N_5158,N_8276);
nand U11325 (N_11325,N_6726,N_7278);
or U11326 (N_11326,N_8282,N_5140);
nand U11327 (N_11327,N_6011,N_8417);
xnor U11328 (N_11328,N_6598,N_6028);
or U11329 (N_11329,N_7561,N_5151);
nand U11330 (N_11330,N_9420,N_8005);
nand U11331 (N_11331,N_9768,N_5803);
and U11332 (N_11332,N_8679,N_9527);
nand U11333 (N_11333,N_7916,N_6750);
nand U11334 (N_11334,N_8839,N_5213);
xnor U11335 (N_11335,N_6927,N_9449);
nand U11336 (N_11336,N_8168,N_7351);
xnor U11337 (N_11337,N_7184,N_7943);
xnor U11338 (N_11338,N_8525,N_7374);
nand U11339 (N_11339,N_5192,N_9609);
nand U11340 (N_11340,N_8473,N_8155);
or U11341 (N_11341,N_5704,N_8544);
xnor U11342 (N_11342,N_9740,N_9153);
and U11343 (N_11343,N_8998,N_5899);
or U11344 (N_11344,N_7874,N_5691);
nor U11345 (N_11345,N_8263,N_9128);
and U11346 (N_11346,N_8039,N_6105);
xnor U11347 (N_11347,N_5175,N_7901);
or U11348 (N_11348,N_9706,N_5127);
and U11349 (N_11349,N_9620,N_9596);
nor U11350 (N_11350,N_7311,N_5846);
nor U11351 (N_11351,N_7794,N_5734);
and U11352 (N_11352,N_5080,N_7191);
and U11353 (N_11353,N_7582,N_7378);
and U11354 (N_11354,N_5772,N_9563);
and U11355 (N_11355,N_9960,N_7453);
nor U11356 (N_11356,N_8543,N_9669);
xnor U11357 (N_11357,N_8844,N_8874);
and U11358 (N_11358,N_9283,N_8689);
or U11359 (N_11359,N_6289,N_8603);
nand U11360 (N_11360,N_6660,N_9410);
nand U11361 (N_11361,N_9066,N_7871);
nor U11362 (N_11362,N_5222,N_9966);
nand U11363 (N_11363,N_5559,N_6500);
or U11364 (N_11364,N_9635,N_8300);
or U11365 (N_11365,N_9413,N_5776);
or U11366 (N_11366,N_8006,N_7781);
xor U11367 (N_11367,N_8123,N_8466);
nand U11368 (N_11368,N_9904,N_5304);
and U11369 (N_11369,N_8419,N_8486);
nand U11370 (N_11370,N_6571,N_6554);
and U11371 (N_11371,N_8967,N_6753);
or U11372 (N_11372,N_5089,N_5212);
nand U11373 (N_11373,N_6915,N_6216);
xor U11374 (N_11374,N_9488,N_7123);
or U11375 (N_11375,N_7725,N_7852);
or U11376 (N_11376,N_7349,N_9362);
nand U11377 (N_11377,N_5161,N_8536);
or U11378 (N_11378,N_9743,N_6816);
and U11379 (N_11379,N_6869,N_6564);
nand U11380 (N_11380,N_7594,N_6080);
and U11381 (N_11381,N_7463,N_9571);
nor U11382 (N_11382,N_6872,N_7861);
or U11383 (N_11383,N_7940,N_7975);
xnor U11384 (N_11384,N_7272,N_5287);
nand U11385 (N_11385,N_5980,N_6683);
or U11386 (N_11386,N_9993,N_6979);
and U11387 (N_11387,N_6023,N_5081);
xnor U11388 (N_11388,N_6297,N_5467);
or U11389 (N_11389,N_7382,N_6306);
or U11390 (N_11390,N_5001,N_6856);
nand U11391 (N_11391,N_5079,N_5551);
nand U11392 (N_11392,N_7260,N_5439);
xnor U11393 (N_11393,N_5041,N_7032);
and U11394 (N_11394,N_7372,N_6259);
xor U11395 (N_11395,N_6408,N_9822);
nor U11396 (N_11396,N_5085,N_5353);
xor U11397 (N_11397,N_7933,N_9658);
or U11398 (N_11398,N_5549,N_6566);
nor U11399 (N_11399,N_7506,N_6084);
nand U11400 (N_11400,N_8524,N_9294);
xnor U11401 (N_11401,N_5573,N_6325);
nand U11402 (N_11402,N_7010,N_9591);
xor U11403 (N_11403,N_9565,N_9875);
xor U11404 (N_11404,N_6935,N_9432);
nor U11405 (N_11405,N_7154,N_6321);
and U11406 (N_11406,N_8132,N_8365);
or U11407 (N_11407,N_5176,N_6046);
or U11408 (N_11408,N_6830,N_5530);
xor U11409 (N_11409,N_6917,N_7148);
or U11410 (N_11410,N_6553,N_5587);
xnor U11411 (N_11411,N_5617,N_8090);
nor U11412 (N_11412,N_7863,N_5611);
and U11413 (N_11413,N_6551,N_9698);
and U11414 (N_11414,N_7735,N_6058);
nor U11415 (N_11415,N_9442,N_9876);
and U11416 (N_11416,N_5331,N_6448);
nand U11417 (N_11417,N_5654,N_7296);
and U11418 (N_11418,N_6913,N_7152);
xnor U11419 (N_11419,N_6860,N_7201);
nor U11420 (N_11420,N_7467,N_5741);
nor U11421 (N_11421,N_7059,N_7930);
nor U11422 (N_11422,N_6847,N_7706);
nand U11423 (N_11423,N_6779,N_7169);
nand U11424 (N_11424,N_9295,N_6277);
nand U11425 (N_11425,N_9239,N_7777);
xor U11426 (N_11426,N_7946,N_7724);
nor U11427 (N_11427,N_8001,N_7167);
xnor U11428 (N_11428,N_8143,N_8733);
nor U11429 (N_11429,N_6550,N_9275);
nor U11430 (N_11430,N_8608,N_9778);
xor U11431 (N_11431,N_7254,N_6505);
nand U11432 (N_11432,N_8861,N_6380);
nand U11433 (N_11433,N_9209,N_6290);
or U11434 (N_11434,N_9764,N_5107);
nor U11435 (N_11435,N_6577,N_8549);
and U11436 (N_11436,N_7515,N_8504);
nand U11437 (N_11437,N_6732,N_7611);
nand U11438 (N_11438,N_5667,N_9639);
nand U11439 (N_11439,N_5434,N_7022);
or U11440 (N_11440,N_7633,N_5505);
or U11441 (N_11441,N_7355,N_8299);
nand U11442 (N_11442,N_5058,N_8816);
or U11443 (N_11443,N_6548,N_7325);
nand U11444 (N_11444,N_9694,N_6210);
nor U11445 (N_11445,N_9748,N_5863);
and U11446 (N_11446,N_5337,N_7886);
or U11447 (N_11447,N_9700,N_8588);
or U11448 (N_11448,N_6579,N_8555);
nor U11449 (N_11449,N_6114,N_6334);
nor U11450 (N_11450,N_9417,N_9095);
nor U11451 (N_11451,N_8134,N_6613);
nand U11452 (N_11452,N_5059,N_7075);
xor U11453 (N_11453,N_7386,N_5764);
nor U11454 (N_11454,N_7507,N_7478);
nand U11455 (N_11455,N_5762,N_9651);
and U11456 (N_11456,N_5526,N_9812);
and U11457 (N_11457,N_7503,N_6545);
nand U11458 (N_11458,N_5370,N_5878);
and U11459 (N_11459,N_6013,N_6462);
xnor U11460 (N_11460,N_7330,N_7746);
nand U11461 (N_11461,N_5015,N_6022);
nand U11462 (N_11462,N_9725,N_6324);
xor U11463 (N_11463,N_8804,N_9877);
nor U11464 (N_11464,N_9359,N_9171);
and U11465 (N_11465,N_8250,N_6916);
or U11466 (N_11466,N_7522,N_9559);
nor U11467 (N_11467,N_5193,N_8317);
nor U11468 (N_11468,N_6162,N_6940);
or U11469 (N_11469,N_9106,N_7214);
or U11470 (N_11470,N_9869,N_8137);
nand U11471 (N_11471,N_6458,N_6094);
and U11472 (N_11472,N_7014,N_6143);
nor U11473 (N_11473,N_8567,N_8936);
or U11474 (N_11474,N_6506,N_9896);
nor U11475 (N_11475,N_7212,N_8108);
and U11476 (N_11476,N_8468,N_7494);
and U11477 (N_11477,N_7824,N_9382);
or U11478 (N_11478,N_6252,N_8156);
and U11479 (N_11479,N_9116,N_7973);
or U11480 (N_11480,N_5678,N_7221);
and U11481 (N_11481,N_9199,N_9918);
xnor U11482 (N_11482,N_7104,N_7029);
nand U11483 (N_11483,N_8261,N_6521);
nand U11484 (N_11484,N_6450,N_8969);
or U11485 (N_11485,N_6206,N_9185);
nor U11486 (N_11486,N_8779,N_5290);
or U11487 (N_11487,N_8657,N_9980);
nand U11488 (N_11488,N_9520,N_9841);
xnor U11489 (N_11489,N_7875,N_8224);
and U11490 (N_11490,N_6428,N_8041);
nor U11491 (N_11491,N_8617,N_6673);
and U11492 (N_11492,N_9039,N_8067);
xor U11493 (N_11493,N_5037,N_7601);
nor U11494 (N_11494,N_5068,N_7731);
nand U11495 (N_11495,N_9738,N_6387);
and U11496 (N_11496,N_7339,N_5967);
nor U11497 (N_11497,N_6524,N_9601);
nand U11498 (N_11498,N_8750,N_7705);
nand U11499 (N_11499,N_9149,N_9947);
or U11500 (N_11500,N_7679,N_9811);
nand U11501 (N_11501,N_6958,N_8456);
nor U11502 (N_11502,N_9403,N_7021);
xnor U11503 (N_11503,N_9322,N_7773);
and U11504 (N_11504,N_6892,N_7712);
or U11505 (N_11505,N_9078,N_9728);
nand U11506 (N_11506,N_6701,N_9032);
nand U11507 (N_11507,N_9496,N_9576);
nor U11508 (N_11508,N_8454,N_8807);
and U11509 (N_11509,N_6516,N_5644);
nand U11510 (N_11510,N_8908,N_7597);
or U11511 (N_11511,N_5808,N_6136);
or U11512 (N_11512,N_5632,N_6774);
xor U11513 (N_11513,N_6721,N_7481);
nor U11514 (N_11514,N_7385,N_8826);
or U11515 (N_11515,N_8325,N_6547);
xnor U11516 (N_11516,N_8510,N_9458);
xor U11517 (N_11517,N_9971,N_5111);
and U11518 (N_11518,N_6431,N_5880);
nand U11519 (N_11519,N_9664,N_7981);
nand U11520 (N_11520,N_6112,N_9140);
xnor U11521 (N_11521,N_6818,N_9142);
and U11522 (N_11522,N_6889,N_7290);
xnor U11523 (N_11523,N_8331,N_8904);
or U11524 (N_11524,N_9495,N_5048);
and U11525 (N_11525,N_8830,N_9720);
nor U11526 (N_11526,N_6043,N_9806);
xnor U11527 (N_11527,N_9607,N_8812);
xnor U11528 (N_11528,N_6375,N_6854);
and U11529 (N_11529,N_7571,N_9113);
and U11530 (N_11530,N_7328,N_5415);
and U11531 (N_11531,N_8912,N_5697);
xor U11532 (N_11532,N_8146,N_7211);
nor U11533 (N_11533,N_5406,N_7811);
xor U11534 (N_11534,N_6389,N_5528);
nor U11535 (N_11535,N_7008,N_5641);
nand U11536 (N_11536,N_5648,N_5604);
or U11537 (N_11537,N_9262,N_7568);
nand U11538 (N_11538,N_9223,N_9625);
and U11539 (N_11539,N_6559,N_5032);
or U11540 (N_11540,N_8557,N_8322);
nand U11541 (N_11541,N_9958,N_8094);
and U11542 (N_11542,N_6473,N_9856);
and U11543 (N_11543,N_5949,N_8396);
nor U11544 (N_11544,N_5881,N_8560);
and U11545 (N_11545,N_6993,N_6365);
or U11546 (N_11546,N_8949,N_7045);
xnor U11547 (N_11547,N_8599,N_5057);
xnor U11548 (N_11548,N_7584,N_7983);
nand U11549 (N_11549,N_9570,N_6875);
xnor U11550 (N_11550,N_5900,N_5774);
or U11551 (N_11551,N_9089,N_6938);
nand U11552 (N_11552,N_7326,N_6837);
or U11553 (N_11553,N_8025,N_9675);
or U11554 (N_11554,N_8422,N_6822);
or U11555 (N_11555,N_9670,N_7316);
nand U11556 (N_11556,N_9638,N_6424);
nor U11557 (N_11557,N_8311,N_6200);
or U11558 (N_11558,N_9813,N_8546);
or U11559 (N_11559,N_8431,N_8256);
and U11560 (N_11560,N_7320,N_9976);
nor U11561 (N_11561,N_9484,N_7243);
or U11562 (N_11562,N_7755,N_8506);
or U11563 (N_11563,N_9044,N_6881);
nor U11564 (N_11564,N_9702,N_5687);
nor U11565 (N_11565,N_6770,N_6655);
nor U11566 (N_11566,N_6773,N_8680);
nor U11567 (N_11567,N_7698,N_6119);
or U11568 (N_11568,N_6920,N_9499);
nand U11569 (N_11569,N_7560,N_7250);
xor U11570 (N_11570,N_5989,N_9076);
and U11571 (N_11571,N_9985,N_9682);
or U11572 (N_11572,N_5348,N_9227);
and U11573 (N_11573,N_6189,N_9065);
nor U11574 (N_11574,N_5242,N_6346);
xnor U11575 (N_11575,N_7247,N_6744);
xnor U11576 (N_11576,N_9164,N_9049);
nor U11577 (N_11577,N_9228,N_6249);
xnor U11578 (N_11578,N_9648,N_5209);
and U11579 (N_11579,N_5208,N_9084);
xnor U11580 (N_11580,N_6412,N_5062);
xor U11581 (N_11581,N_6600,N_9167);
and U11582 (N_11582,N_7293,N_9623);
nor U11583 (N_11583,N_6696,N_9291);
and U11584 (N_11584,N_7808,N_9197);
and U11585 (N_11585,N_6108,N_5555);
and U11586 (N_11586,N_7992,N_6218);
nand U11587 (N_11587,N_7741,N_7783);
nor U11588 (N_11588,N_9735,N_5871);
nand U11589 (N_11589,N_6280,N_6749);
nand U11590 (N_11590,N_6493,N_9693);
xnor U11591 (N_11591,N_5827,N_6484);
or U11592 (N_11592,N_5584,N_9774);
nor U11593 (N_11593,N_9824,N_6890);
and U11594 (N_11594,N_5281,N_7662);
or U11595 (N_11595,N_8093,N_6783);
and U11596 (N_11596,N_8637,N_6247);
xnor U11597 (N_11597,N_7836,N_9998);
nor U11598 (N_11598,N_9176,N_8622);
nor U11599 (N_11599,N_6765,N_7747);
nand U11600 (N_11600,N_8459,N_6741);
or U11601 (N_11601,N_6472,N_9530);
nand U11602 (N_11602,N_8124,N_7869);
xor U11603 (N_11603,N_8628,N_9645);
xor U11604 (N_11604,N_5310,N_6675);
nand U11605 (N_11605,N_6691,N_8232);
and U11606 (N_11606,N_8437,N_9515);
nand U11607 (N_11607,N_7929,N_8226);
or U11608 (N_11608,N_8111,N_6068);
xnor U11609 (N_11609,N_7703,N_6175);
or U11610 (N_11610,N_5747,N_5130);
or U11611 (N_11611,N_5892,N_6403);
nand U11612 (N_11612,N_5282,N_5073);
xnor U11613 (N_11613,N_7001,N_9428);
xnor U11614 (N_11614,N_6849,N_7977);
xor U11615 (N_11615,N_5902,N_9744);
nand U11616 (N_11616,N_9901,N_6260);
nor U11617 (N_11617,N_9365,N_6949);
and U11618 (N_11618,N_8867,N_8326);
nand U11619 (N_11619,N_8947,N_9972);
xnor U11620 (N_11620,N_7835,N_9986);
xor U11621 (N_11621,N_7455,N_7271);
and U11622 (N_11622,N_8358,N_9719);
or U11623 (N_11623,N_5554,N_7610);
and U11624 (N_11624,N_8596,N_9870);
and U11625 (N_11625,N_7252,N_5230);
and U11626 (N_11626,N_7149,N_6885);
xor U11627 (N_11627,N_7805,N_5024);
and U11628 (N_11628,N_5642,N_5326);
nor U11629 (N_11629,N_5660,N_7647);
nand U11630 (N_11630,N_9524,N_7484);
nand U11631 (N_11631,N_8659,N_8255);
nand U11632 (N_11632,N_9801,N_9569);
xor U11633 (N_11633,N_6307,N_7979);
nor U11634 (N_11634,N_5138,N_5053);
or U11635 (N_11635,N_6225,N_9545);
or U11636 (N_11636,N_7596,N_6008);
nor U11637 (N_11637,N_5563,N_9445);
nor U11638 (N_11638,N_8955,N_5286);
xnor U11639 (N_11639,N_8206,N_5894);
and U11640 (N_11640,N_8620,N_8297);
nor U11641 (N_11641,N_5489,N_7468);
xor U11642 (N_11642,N_5204,N_6601);
nand U11643 (N_11643,N_8850,N_6642);
nand U11644 (N_11644,N_9914,N_6414);
and U11645 (N_11645,N_8984,N_9068);
nand U11646 (N_11646,N_8009,N_6844);
xnor U11647 (N_11647,N_8631,N_5891);
xnor U11648 (N_11648,N_9532,N_8081);
nor U11649 (N_11649,N_6894,N_7643);
nand U11650 (N_11650,N_5023,N_8115);
and U11651 (N_11651,N_7936,N_5836);
or U11652 (N_11652,N_7990,N_7911);
xnor U11653 (N_11653,N_7928,N_7288);
nand U11654 (N_11654,N_9057,N_7444);
xnor U11655 (N_11655,N_9713,N_8508);
xor U11656 (N_11656,N_9808,N_7089);
nand U11657 (N_11657,N_5849,N_6062);
and U11658 (N_11658,N_8073,N_5025);
or U11659 (N_11659,N_5170,N_9931);
nand U11660 (N_11660,N_7137,N_8749);
or U11661 (N_11661,N_6874,N_7569);
xnor U11662 (N_11662,N_8266,N_7450);
and U11663 (N_11663,N_6087,N_6156);
nor U11664 (N_11664,N_9086,N_5994);
or U11665 (N_11665,N_7485,N_8787);
nor U11666 (N_11666,N_7605,N_8764);
and U11667 (N_11667,N_5400,N_7514);
or U11668 (N_11668,N_9940,N_8547);
xnor U11669 (N_11669,N_7058,N_5379);
xor U11670 (N_11670,N_5650,N_6209);
nand U11671 (N_11671,N_6301,N_8356);
xnor U11672 (N_11672,N_7181,N_5912);
xnor U11673 (N_11673,N_6379,N_8851);
nor U11674 (N_11674,N_6791,N_8033);
nand U11675 (N_11675,N_9910,N_7498);
or U11676 (N_11676,N_7722,N_8161);
or U11677 (N_11677,N_8970,N_9494);
nor U11678 (N_11678,N_5521,N_6096);
or U11679 (N_11679,N_9230,N_9401);
nand U11680 (N_11680,N_7668,N_9598);
and U11681 (N_11681,N_7025,N_6591);
nor U11682 (N_11682,N_8492,N_9539);
nor U11683 (N_11683,N_9867,N_5207);
nor U11684 (N_11684,N_6688,N_8939);
or U11685 (N_11685,N_7142,N_9212);
nand U11686 (N_11686,N_8294,N_9208);
nand U11687 (N_11687,N_7676,N_6637);
nand U11688 (N_11688,N_8606,N_5984);
xor U11689 (N_11689,N_7434,N_5659);
or U11690 (N_11690,N_6312,N_7459);
or U11691 (N_11691,N_9023,N_7903);
or U11692 (N_11692,N_7323,N_5054);
and U11693 (N_11693,N_7281,N_5835);
or U11694 (N_11694,N_8307,N_7621);
xnor U11695 (N_11695,N_7818,N_9471);
xnor U11696 (N_11696,N_5381,N_7145);
or U11697 (N_11697,N_7912,N_6509);
and U11698 (N_11698,N_5113,N_6269);
xnor U11699 (N_11699,N_6653,N_6461);
and U11700 (N_11700,N_9691,N_8799);
nand U11701 (N_11701,N_6303,N_7186);
nand U11702 (N_11702,N_5942,N_7523);
xor U11703 (N_11703,N_9352,N_7340);
nand U11704 (N_11704,N_6186,N_9647);
xor U11705 (N_11705,N_9281,N_9454);
xor U11706 (N_11706,N_6782,N_7225);
and U11707 (N_11707,N_5616,N_6447);
xnor U11708 (N_11708,N_6142,N_9292);
xnor U11709 (N_11709,N_6178,N_9925);
nor U11710 (N_11710,N_7576,N_8104);
xnor U11711 (N_11711,N_8880,N_7217);
nand U11712 (N_11712,N_5533,N_8576);
nor U11713 (N_11713,N_5340,N_8962);
nand U11714 (N_11714,N_7308,N_5756);
nand U11715 (N_11715,N_6373,N_9542);
and U11716 (N_11716,N_9797,N_9380);
nand U11717 (N_11717,N_8187,N_9422);
or U11718 (N_11718,N_9656,N_6672);
or U11719 (N_11719,N_9145,N_5000);
nand U11720 (N_11720,N_9325,N_8999);
nand U11721 (N_11721,N_7900,N_8899);
nand U11722 (N_11722,N_7143,N_9739);
xnor U11723 (N_11723,N_7331,N_7558);
xor U11724 (N_11724,N_6586,N_6352);
or U11725 (N_11725,N_7423,N_5494);
xnor U11726 (N_11726,N_8219,N_7927);
and U11727 (N_11727,N_6989,N_9395);
and U11728 (N_11728,N_5834,N_8074);
nor U11729 (N_11729,N_8359,N_9114);
nor U11730 (N_11730,N_6219,N_5493);
nand U11731 (N_11731,N_5564,N_8162);
xor U11732 (N_11732,N_8520,N_9343);
or U11733 (N_11733,N_8910,N_8535);
xor U11734 (N_11734,N_5869,N_8953);
and U11735 (N_11735,N_5807,N_9225);
nor U11736 (N_11736,N_5988,N_5673);
nor U11737 (N_11737,N_9217,N_6884);
xnor U11738 (N_11738,N_5711,N_6937);
nor U11739 (N_11739,N_8186,N_9198);
or U11740 (N_11740,N_8977,N_6966);
nand U11741 (N_11741,N_8931,N_7778);
or U11742 (N_11742,N_9975,N_5767);
xor U11743 (N_11743,N_6859,N_5866);
nand U11744 (N_11744,N_7971,N_5004);
nor U11745 (N_11745,N_5194,N_8796);
and U11746 (N_11746,N_5910,N_9173);
xor U11747 (N_11747,N_8235,N_8727);
and U11748 (N_11748,N_7166,N_6630);
nor U11749 (N_11749,N_7669,N_8806);
and U11750 (N_11750,N_9973,N_9083);
nand U11751 (N_11751,N_7277,N_8578);
and U11752 (N_11752,N_9485,N_8987);
and U11753 (N_11753,N_9169,N_7046);
nand U11754 (N_11754,N_7003,N_9714);
and U11755 (N_11755,N_6731,N_5480);
nand U11756 (N_11756,N_9640,N_7213);
or U11757 (N_11757,N_7274,N_8958);
xor U11758 (N_11758,N_6527,N_9900);
xor U11759 (N_11759,N_5859,N_5574);
and U11760 (N_11760,N_6582,N_6574);
and U11761 (N_11761,N_7460,N_6941);
or U11762 (N_11762,N_5092,N_7879);
nor U11763 (N_11763,N_7219,N_8082);
nand U11764 (N_11764,N_8691,N_7618);
and U11765 (N_11765,N_5696,N_6697);
nor U11766 (N_11766,N_9144,N_9377);
and U11767 (N_11767,N_9285,N_5178);
nand U11768 (N_11768,N_6268,N_8037);
and U11769 (N_11769,N_8288,N_8457);
nor U11770 (N_11770,N_7520,N_6603);
and U11771 (N_11771,N_9249,N_9286);
or U11772 (N_11772,N_8238,N_6015);
xnor U11773 (N_11773,N_5146,N_6759);
and U11774 (N_11774,N_5410,N_6876);
nor U11775 (N_11775,N_7673,N_7653);
nor U11776 (N_11776,N_9460,N_5759);
nor U11777 (N_11777,N_9333,N_6227);
and U11778 (N_11778,N_6194,N_8761);
and U11779 (N_11779,N_7276,N_9355);
and U11780 (N_11780,N_8849,N_6836);
xor U11781 (N_11781,N_8819,N_7814);
xor U11782 (N_11782,N_6684,N_5329);
and U11783 (N_11783,N_7752,N_8886);
and U11784 (N_11784,N_5430,N_6512);
nand U11785 (N_11785,N_5825,N_6282);
and U11786 (N_11786,N_9088,N_6552);
nand U11787 (N_11787,N_5203,N_7365);
or U11788 (N_11788,N_6041,N_5665);
nand U11789 (N_11789,N_5019,N_7204);
and U11790 (N_11790,N_8117,N_7397);
nor U11791 (N_11791,N_6496,N_5672);
nand U11792 (N_11792,N_8676,N_6576);
and U11793 (N_11793,N_7336,N_7111);
nand U11794 (N_11794,N_9469,N_9574);
xnor U11795 (N_11795,N_8233,N_9630);
and U11796 (N_11796,N_6800,N_6126);
nor U11797 (N_11797,N_7577,N_8624);
or U11798 (N_11798,N_8262,N_5930);
or U11799 (N_11799,N_9536,N_6788);
or U11800 (N_11800,N_8166,N_7432);
nand U11801 (N_11801,N_9455,N_5149);
nor U11802 (N_11802,N_5216,N_9372);
or U11803 (N_11803,N_7437,N_5278);
and U11804 (N_11804,N_5718,N_9937);
xnor U11805 (N_11805,N_6857,N_8521);
or U11806 (N_11806,N_9888,N_7876);
nand U11807 (N_11807,N_8284,N_9921);
or U11808 (N_11808,N_9831,N_6693);
or U11809 (N_11809,N_9540,N_9226);
nand U11810 (N_11810,N_5131,N_7966);
xnor U11811 (N_11811,N_5763,N_5264);
xor U11812 (N_11812,N_5838,N_8937);
and U11813 (N_11813,N_5160,N_8551);
xor U11814 (N_11814,N_8321,N_7130);
xor U11815 (N_11815,N_9633,N_5375);
xnor U11816 (N_11816,N_6228,N_5419);
or U11817 (N_11817,N_6834,N_6192);
nand U11818 (N_11818,N_8329,N_6130);
xor U11819 (N_11819,N_6026,N_7418);
nor U11820 (N_11820,N_6499,N_8925);
xnor U11821 (N_11821,N_9472,N_7980);
and U11822 (N_11822,N_8135,N_8088);
or U11823 (N_11823,N_5235,N_6870);
nor U11824 (N_11824,N_9421,N_7106);
and U11825 (N_11825,N_5502,N_7820);
nand U11826 (N_11826,N_6390,N_8957);
or U11827 (N_11827,N_8293,N_7144);
xor U11828 (N_11828,N_6758,N_7291);
nor U11829 (N_11829,N_6556,N_8863);
and U11830 (N_11830,N_6584,N_8865);
xor U11831 (N_11831,N_5052,N_5990);
xnor U11832 (N_11832,N_8339,N_6383);
xnor U11833 (N_11833,N_8131,N_8866);
nor U11834 (N_11834,N_9967,N_9202);
nand U11835 (N_11835,N_9491,N_8674);
xnor U11836 (N_11836,N_5525,N_5271);
nand U11837 (N_11837,N_8563,N_5897);
and U11838 (N_11838,N_9335,N_8614);
or U11839 (N_11839,N_7513,N_8891);
or U11840 (N_11840,N_9193,N_6572);
xnor U11841 (N_11841,N_8215,N_7085);
nor U11842 (N_11842,N_9616,N_5323);
nand U11843 (N_11843,N_5478,N_5876);
nand U11844 (N_11844,N_6994,N_9091);
or U11845 (N_11845,N_7285,N_9028);
xnor U11846 (N_11846,N_9229,N_8976);
nor U11847 (N_11847,N_9155,N_9612);
xor U11848 (N_11848,N_6009,N_9699);
and U11849 (N_11849,N_9643,N_5675);
nand U11850 (N_11850,N_8648,N_8475);
and U11851 (N_11851,N_5103,N_9928);
xnor U11852 (N_11852,N_5129,N_6761);
nor U11853 (N_11853,N_8416,N_9364);
nor U11854 (N_11854,N_6032,N_7301);
and U11855 (N_11855,N_7421,N_8122);
or U11856 (N_11856,N_8968,N_9219);
xnor U11857 (N_11857,N_8724,N_7027);
xor U11858 (N_11858,N_8077,N_9850);
xor U11859 (N_11859,N_6430,N_9760);
nor U11860 (N_11860,N_6610,N_8519);
xnor U11861 (N_11861,N_5408,N_9537);
and U11862 (N_11862,N_5295,N_9074);
and U11863 (N_11863,N_7475,N_8719);
nor U11864 (N_11864,N_6396,N_5279);
nor U11865 (N_11865,N_6185,N_9538);
and U11866 (N_11866,N_5723,N_6734);
or U11867 (N_11867,N_9779,N_5070);
xor U11868 (N_11868,N_6442,N_8704);
xor U11869 (N_11869,N_7024,N_9961);
and U11870 (N_11870,N_9415,N_7012);
nand U11871 (N_11871,N_6785,N_9950);
and U11872 (N_11872,N_7799,N_6666);
and U11873 (N_11873,N_9687,N_7716);
and U11874 (N_11874,N_5110,N_5537);
xor U11875 (N_11875,N_5189,N_5416);
xor U11876 (N_11876,N_7442,N_5550);
or U11877 (N_11877,N_6738,N_9398);
and U11878 (N_11878,N_8669,N_5944);
nand U11879 (N_11879,N_5036,N_5418);
nand U11880 (N_11880,N_5951,N_7380);
or U11881 (N_11881,N_5917,N_8864);
xor U11882 (N_11882,N_5453,N_9476);
nand U11883 (N_11883,N_6173,N_8935);
xor U11884 (N_11884,N_6877,N_9765);
and U11885 (N_11885,N_7466,N_6663);
nand U11886 (N_11886,N_8838,N_9781);
xor U11887 (N_11887,N_6879,N_9582);
or U11888 (N_11888,N_8291,N_6132);
nand U11889 (N_11889,N_8066,N_6986);
nor U11890 (N_11890,N_7685,N_6793);
nor U11891 (N_11891,N_6413,N_7830);
nand U11892 (N_11892,N_7562,N_9965);
nor U11893 (N_11893,N_5884,N_6871);
nor U11894 (N_11894,N_5157,N_9439);
xor U11895 (N_11895,N_8742,N_9481);
xor U11896 (N_11896,N_9614,N_7190);
nor U11897 (N_11897,N_9218,N_9348);
or U11898 (N_11898,N_5569,N_5716);
nand U11899 (N_11899,N_5887,N_9203);
nor U11900 (N_11900,N_5404,N_5006);
and U11901 (N_11901,N_9839,N_7342);
and U11902 (N_11902,N_5155,N_5682);
nor U11903 (N_11903,N_9767,N_6956);
and U11904 (N_11904,N_5141,N_5386);
nand U11905 (N_11905,N_6633,N_9363);
or U11906 (N_11906,N_9213,N_9257);
xor U11907 (N_11907,N_7771,N_5003);
xnor U11908 (N_11908,N_9373,N_6151);
or U11909 (N_11909,N_6560,N_7998);
nor U11910 (N_11910,N_7268,N_9685);
xor U11911 (N_11911,N_5099,N_5511);
nor U11912 (N_11912,N_6279,N_9712);
nand U11913 (N_11913,N_9657,N_8430);
and U11914 (N_11914,N_6085,N_5898);
or U11915 (N_11915,N_5116,N_6097);
or U11916 (N_11916,N_8503,N_7310);
xnor U11917 (N_11917,N_9465,N_9556);
and U11918 (N_11918,N_8627,N_8817);
or U11919 (N_11919,N_6343,N_8316);
xor U11920 (N_11920,N_9214,N_5376);
or U11921 (N_11921,N_6254,N_7691);
nor U11922 (N_11922,N_5829,N_5636);
or U11923 (N_11923,N_5851,N_6098);
nor U11924 (N_11924,N_8022,N_7877);
and U11925 (N_11925,N_5039,N_7449);
nand U11926 (N_11926,N_5705,N_6980);
xnor U11927 (N_11927,N_5813,N_7573);
or U11928 (N_11928,N_7907,N_9338);
and U11929 (N_11929,N_5752,N_6090);
nand U11930 (N_11930,N_9082,N_7959);
xor U11931 (N_11931,N_6514,N_9772);
xnor U11932 (N_11932,N_7798,N_9393);
xor U11933 (N_11933,N_7430,N_5277);
nor U11934 (N_11934,N_8712,N_6111);
nor U11935 (N_11935,N_8244,N_9800);
nand U11936 (N_11936,N_6256,N_8500);
nand U11937 (N_11937,N_6296,N_7666);
nand U11938 (N_11938,N_6214,N_7065);
and U11939 (N_11939,N_8703,N_8687);
xor U11940 (N_11940,N_8531,N_7660);
or U11941 (N_11941,N_8707,N_6549);
or U11942 (N_11942,N_8148,N_5358);
or U11943 (N_11943,N_5142,N_5612);
and U11944 (N_11944,N_8841,N_9847);
nand U11945 (N_11945,N_6246,N_8993);
nor U11946 (N_11946,N_9353,N_7454);
or U11947 (N_11947,N_5709,N_8616);
nor U11948 (N_11948,N_5727,N_6128);
nor U11949 (N_11949,N_7819,N_9997);
xnor U11950 (N_11950,N_6686,N_8823);
nor U11951 (N_11951,N_6469,N_7416);
or U11952 (N_11952,N_8607,N_6954);
xor U11953 (N_11953,N_7665,N_6468);
nand U11954 (N_11954,N_7038,N_9754);
nor U11955 (N_11955,N_9789,N_5524);
and U11956 (N_11956,N_8051,N_8391);
and U11957 (N_11957,N_6720,N_8630);
and U11958 (N_11958,N_6623,N_8145);
xor U11959 (N_11959,N_6363,N_9004);
xnor U11960 (N_11960,N_7831,N_5020);
and U11961 (N_11961,N_8927,N_8911);
and U11962 (N_11962,N_5806,N_8290);
xor U11963 (N_11963,N_5976,N_5627);
nand U11964 (N_11964,N_7317,N_6243);
nand U11965 (N_11965,N_7396,N_9356);
or U11966 (N_11966,N_6751,N_9721);
xor U11967 (N_11967,N_9863,N_9873);
xor U11968 (N_11968,N_7119,N_6967);
or U11969 (N_11969,N_9517,N_9519);
and U11970 (N_11970,N_8814,N_8554);
and U11971 (N_11971,N_6820,N_9334);
or U11972 (N_11972,N_8929,N_7904);
nor U11973 (N_11973,N_9297,N_5663);
nand U11974 (N_11974,N_6359,N_9704);
xor U11975 (N_11975,N_7906,N_6099);
and U11976 (N_11976,N_6590,N_7518);
xnor U11977 (N_11977,N_9016,N_5811);
and U11978 (N_11978,N_5775,N_8777);
and U11979 (N_11979,N_5206,N_7384);
and U11980 (N_11980,N_5339,N_8167);
xnor U11981 (N_11981,N_9046,N_8381);
and U11982 (N_11982,N_7539,N_6724);
xor U11983 (N_11983,N_9810,N_5457);
or U11984 (N_11984,N_5907,N_8414);
xor U11985 (N_11985,N_6304,N_9502);
xnor U11986 (N_11986,N_9054,N_6073);
and U11987 (N_11987,N_5640,N_8448);
or U11988 (N_11988,N_9663,N_7327);
xnor U11989 (N_11989,N_8190,N_5698);
nand U11990 (N_11990,N_8320,N_5558);
and U11991 (N_11991,N_9929,N_6123);
nor U11992 (N_11992,N_9102,N_6819);
and U11993 (N_11993,N_9368,N_9522);
and U11994 (N_11994,N_5154,N_9912);
nand U11995 (N_11995,N_7763,N_8178);
and U11996 (N_11996,N_7950,N_7693);
or U11997 (N_11997,N_6644,N_8586);
or U11998 (N_11998,N_7974,N_7026);
or U11999 (N_11999,N_7334,N_9500);
xnor U12000 (N_12000,N_8265,N_5635);
xnor U12001 (N_12001,N_8665,N_7606);
nand U12002 (N_12002,N_8534,N_5077);
and U12003 (N_12003,N_8031,N_5586);
xnor U12004 (N_12004,N_9511,N_6569);
nand U12005 (N_12005,N_9050,N_5087);
or U12006 (N_12006,N_8113,N_8471);
xnor U12007 (N_12007,N_5598,N_8127);
or U12008 (N_12008,N_8179,N_7885);
nand U12009 (N_12009,N_9463,N_6166);
or U12010 (N_12010,N_7528,N_5366);
and U12011 (N_12011,N_7357,N_5298);
nand U12012 (N_12012,N_8960,N_5717);
or U12013 (N_12013,N_8928,N_5262);
nand U12014 (N_12014,N_9467,N_9939);
nor U12015 (N_12015,N_6703,N_8505);
nand U12016 (N_12016,N_5424,N_9447);
nand U12017 (N_12017,N_6975,N_5966);
nand U12018 (N_12018,N_6546,N_7939);
xor U12019 (N_12019,N_5921,N_8374);
and U12020 (N_12020,N_5440,N_5137);
xor U12021 (N_12021,N_7061,N_8682);
or U12022 (N_12022,N_6042,N_8412);
or U12023 (N_12023,N_7424,N_6435);
and U12024 (N_12024,N_9329,N_9715);
nand U12025 (N_12025,N_6540,N_7035);
nand U12026 (N_12026,N_7428,N_6748);
nand U12027 (N_12027,N_6525,N_6059);
nand U12028 (N_12028,N_6537,N_7457);
nor U12029 (N_12029,N_8685,N_8813);
and U12030 (N_12030,N_9437,N_6318);
nor U12031 (N_12031,N_7996,N_5261);
nand U12032 (N_12032,N_6276,N_7347);
or U12033 (N_12033,N_6179,N_5547);
xor U12034 (N_12034,N_6283,N_6456);
or U12035 (N_12035,N_8460,N_8270);
and U12036 (N_12036,N_5761,N_7664);
nor U12037 (N_12037,N_5152,N_9583);
xnor U12038 (N_12038,N_5655,N_7629);
nand U12039 (N_12039,N_5595,N_6900);
xor U12040 (N_12040,N_8487,N_9964);
or U12041 (N_12041,N_9858,N_7649);
nor U12042 (N_12042,N_8024,N_8533);
nor U12043 (N_12043,N_8204,N_7635);
or U12044 (N_12044,N_5968,N_6212);
xnor U12045 (N_12045,N_6504,N_9953);
and U12046 (N_12046,N_6399,N_9533);
nand U12047 (N_12047,N_8047,N_5372);
xor U12048 (N_12048,N_8205,N_8501);
nand U12049 (N_12049,N_9749,N_7131);
or U12050 (N_12050,N_5008,N_8211);
nand U12051 (N_12051,N_7954,N_7654);
and U12052 (N_12052,N_6615,N_7788);
nor U12053 (N_12053,N_5447,N_6060);
xor U12054 (N_12054,N_8114,N_7427);
and U12055 (N_12055,N_6733,N_5580);
nor U12056 (N_12056,N_6125,N_9757);
nor U12057 (N_12057,N_9007,N_8696);
xnor U12058 (N_12058,N_8583,N_8242);
and U12059 (N_12059,N_9304,N_5256);
and U12060 (N_12060,N_8375,N_6065);
and U12061 (N_12061,N_7932,N_9889);
and U12062 (N_12062,N_5860,N_9505);
nand U12063 (N_12063,N_6532,N_7451);
nor U12064 (N_12064,N_6278,N_5275);
nand U12065 (N_12065,N_8120,N_6501);
nor U12066 (N_12066,N_6645,N_8177);
nand U12067 (N_12067,N_7884,N_8888);
xor U12068 (N_12068,N_7095,N_5018);
or U12069 (N_12069,N_5901,N_5322);
or U12070 (N_12070,N_7578,N_8053);
or U12071 (N_12071,N_8017,N_5983);
or U12072 (N_12072,N_7456,N_8207);
and U12073 (N_12073,N_5389,N_8744);
nor U12074 (N_12074,N_9821,N_7504);
or U12075 (N_12075,N_5750,N_7280);
xnor U12076 (N_12076,N_6923,N_9834);
nor U12077 (N_12077,N_5700,N_7452);
xor U12078 (N_12078,N_6353,N_7049);
and U12079 (N_12079,N_5651,N_8780);
or U12080 (N_12080,N_7791,N_7536);
nand U12081 (N_12081,N_5321,N_7176);
and U12082 (N_12082,N_5913,N_7634);
nand U12083 (N_12083,N_8069,N_6522);
nand U12084 (N_12084,N_5613,N_5045);
and U12085 (N_12085,N_5428,N_7591);
and U12086 (N_12086,N_8593,N_7614);
nor U12087 (N_12087,N_7555,N_5492);
xnor U12088 (N_12088,N_9189,N_6535);
nand U12089 (N_12089,N_8357,N_6255);
or U12090 (N_12090,N_8635,N_7993);
or U12091 (N_12091,N_6223,N_8469);
or U12092 (N_12092,N_5223,N_7567);
xor U12093 (N_12093,N_8898,N_9264);
and U12094 (N_12094,N_7099,N_8553);
xor U12095 (N_12095,N_9268,N_5371);
or U12096 (N_12096,N_8203,N_8497);
nor U12097 (N_12097,N_9457,N_7114);
xor U12098 (N_12098,N_7789,N_6180);
nand U12099 (N_12099,N_5553,N_7923);
xnor U12100 (N_12100,N_6300,N_7816);
and U12101 (N_12101,N_9350,N_6217);
nor U12102 (N_12102,N_9290,N_8043);
nor U12103 (N_12103,N_6602,N_6702);
nor U12104 (N_12104,N_6235,N_7193);
xor U12105 (N_12105,N_6231,N_6027);
xnor U12106 (N_12106,N_8972,N_6826);
and U12107 (N_12107,N_6152,N_6275);
and U12108 (N_12108,N_5219,N_8338);
and U12109 (N_12109,N_6804,N_8753);
xnor U12110 (N_12110,N_6075,N_5002);
and U12111 (N_12111,N_9999,N_7511);
and U12112 (N_12112,N_5373,N_8980);
xor U12113 (N_12113,N_8905,N_8246);
nor U12114 (N_12114,N_8909,N_7807);
and U12115 (N_12115,N_6034,N_7007);
and U12116 (N_12116,N_5473,N_9887);
and U12117 (N_12117,N_5136,N_8200);
or U12118 (N_12118,N_9090,N_6961);
and U12119 (N_12119,N_5882,N_9952);
and U12120 (N_12120,N_6311,N_5885);
or U12121 (N_12121,N_6460,N_5259);
nor U12122 (N_12122,N_8589,N_8871);
nand U12123 (N_12123,N_6446,N_9762);
nand U12124 (N_12124,N_9763,N_8399);
or U12125 (N_12125,N_8336,N_6470);
xor U12126 (N_12126,N_9631,N_8789);
xnor U12127 (N_12127,N_5828,N_5890);
or U12128 (N_12128,N_5962,N_8138);
nor U12129 (N_12129,N_8572,N_9868);
xor U12130 (N_12130,N_8552,N_9911);
and U12131 (N_12131,N_9081,N_9251);
nand U12132 (N_12132,N_6786,N_6401);
nand U12133 (N_12133,N_8209,N_6768);
and U12134 (N_12134,N_7249,N_9666);
and U12135 (N_12135,N_9646,N_6824);
nor U12136 (N_12136,N_8214,N_9277);
nand U12137 (N_12137,N_6054,N_9201);
nor U12138 (N_12138,N_7776,N_8404);
or U12139 (N_12139,N_5513,N_6012);
and U12140 (N_12140,N_8914,N_8369);
xor U12141 (N_12141,N_5646,N_6415);
nor U12142 (N_12142,N_8577,N_8016);
and U12143 (N_12143,N_6609,N_5030);
nor U12144 (N_12144,N_5274,N_7255);
nand U12145 (N_12145,N_5668,N_7801);
and U12146 (N_12146,N_5820,N_5830);
nor U12147 (N_12147,N_8192,N_6207);
or U12148 (N_12148,N_7465,N_5195);
xor U12149 (N_12149,N_7258,N_5782);
nor U12150 (N_12150,N_8542,N_5933);
nand U12151 (N_12151,N_5590,N_6513);
or U12152 (N_12152,N_7335,N_9296);
nor U12153 (N_12153,N_6367,N_8759);
and U12154 (N_12154,N_6676,N_9659);
xor U12155 (N_12155,N_7078,N_5377);
xnor U12156 (N_12156,N_9267,N_6477);
and U12157 (N_12157,N_8601,N_9123);
and U12158 (N_12158,N_8097,N_6171);
nand U12159 (N_12159,N_8159,N_7147);
xnor U12160 (N_12160,N_6511,N_7172);
or U12161 (N_12161,N_9163,N_8021);
xnor U12162 (N_12162,N_8991,N_6341);
nor U12163 (N_12163,N_7547,N_6658);
and U12164 (N_12164,N_8965,N_9737);
and U12165 (N_12165,N_6454,N_9825);
nor U12166 (N_12166,N_8877,N_5360);
or U12167 (N_12167,N_7739,N_9105);
and U12168 (N_12168,N_8222,N_5491);
nand U12169 (N_12169,N_8869,N_6044);
nand U12170 (N_12170,N_6669,N_8194);
xnor U12171 (N_12171,N_6953,N_7218);
or U12172 (N_12172,N_7359,N_9327);
or U12173 (N_12173,N_6843,N_6066);
or U12174 (N_12174,N_8818,N_8385);
and U12175 (N_12175,N_5710,N_8453);
nand U12176 (N_12176,N_5448,N_5932);
and U12177 (N_12177,N_9634,N_9673);
or U12178 (N_12178,N_8302,N_8746);
nand U12179 (N_12179,N_9549,N_7859);
xor U12180 (N_12180,N_6618,N_5289);
nor U12181 (N_12181,N_9955,N_8887);
nand U12182 (N_12182,N_6952,N_6722);
nand U12183 (N_12183,N_8029,N_5733);
and U12184 (N_12184,N_5486,N_9506);
nand U12185 (N_12185,N_5182,N_5958);
nand U12186 (N_12186,N_8046,N_9902);
or U12187 (N_12187,N_7711,N_6118);
xor U12188 (N_12188,N_8180,N_8747);
or U12189 (N_12189,N_9430,N_6507);
or U12190 (N_12190,N_9211,N_8726);
and U12191 (N_12191,N_8632,N_9077);
and U12192 (N_12192,N_8286,N_6933);
nor U12193 (N_12193,N_8195,N_5401);
nor U12194 (N_12194,N_7079,N_9097);
or U12195 (N_12195,N_6037,N_6155);
and U12196 (N_12196,N_5394,N_6451);
or U12197 (N_12197,N_8790,N_6671);
nand U12198 (N_12198,N_7839,N_8527);
xnor U12199 (N_12199,N_9328,N_7471);
nand U12200 (N_12200,N_5685,N_7462);
xnor U12201 (N_12201,N_8982,N_7146);
and U12202 (N_12202,N_7502,N_9138);
xor U12203 (N_12203,N_6626,N_8477);
nand U12204 (N_12204,N_9100,N_9510);
or U12205 (N_12205,N_8995,N_8171);
nand U12206 (N_12206,N_9493,N_8415);
nor U12207 (N_12207,N_9726,N_6006);
or U12208 (N_12208,N_9263,N_6024);
nand U12209 (N_12209,N_8010,N_5758);
or U12210 (N_12210,N_7337,N_8677);
nor U12211 (N_12211,N_5288,N_9172);
xor U12212 (N_12212,N_8393,N_7044);
or U12213 (N_12213,N_7538,N_6700);
nor U12214 (N_12214,N_8210,N_7064);
or U12215 (N_12215,N_8978,N_9061);
nand U12216 (N_12216,N_7395,N_8511);
or U12217 (N_12217,N_8268,N_9498);
nand U12218 (N_12218,N_7902,N_5683);
or U12219 (N_12219,N_6445,N_8684);
xnor U12220 (N_12220,N_9099,N_8743);
or U12221 (N_12221,N_9034,N_5508);
and U12222 (N_12222,N_7447,N_6261);
xnor U12223 (N_12223,N_5086,N_5954);
or U12224 (N_12224,N_9358,N_5483);
xor U12225 (N_12225,N_9927,N_6746);
and U12226 (N_12226,N_5270,N_6497);
and U12227 (N_12227,N_7897,N_7300);
xnor U12228 (N_12228,N_6050,N_7362);
xnor U12229 (N_12229,N_8440,N_5940);
nand U12230 (N_12230,N_8170,N_7472);
and U12231 (N_12231,N_7113,N_6680);
nor U12232 (N_12232,N_9705,N_8698);
or U12233 (N_12233,N_8762,N_5959);
or U12234 (N_12234,N_9337,N_8926);
xor U12235 (N_12235,N_5969,N_9336);
or U12236 (N_12236,N_5101,N_7728);
nand U12237 (N_12237,N_8772,N_8446);
nor U12238 (N_12238,N_9652,N_7435);
or U12239 (N_12239,N_9147,N_7259);
nor U12240 (N_12240,N_6019,N_5686);
xor U12241 (N_12241,N_8306,N_7535);
and U12242 (N_12242,N_9660,N_7764);
xnor U12243 (N_12243,N_5108,N_5438);
or U12244 (N_12244,N_8619,N_6699);
and U12245 (N_12245,N_5512,N_7458);
and U12246 (N_12246,N_5588,N_7175);
and U12247 (N_12247,N_7414,N_9603);
nand U12248 (N_12248,N_7709,N_5171);
and U12249 (N_12249,N_6981,N_6563);
or U12250 (N_12250,N_5464,N_5649);
xnor U12251 (N_12251,N_5392,N_8918);
and U12252 (N_12252,N_8198,N_7800);
xor U12253 (N_12253,N_5631,N_7198);
xor U12254 (N_12254,N_6051,N_6081);
xor U12255 (N_12255,N_6170,N_7196);
xor U12256 (N_12256,N_6851,N_7652);
nor U12257 (N_12257,N_8201,N_7671);
xor U12258 (N_12258,N_9644,N_7858);
nand U12259 (N_12259,N_5225,N_5368);
or U12260 (N_12260,N_5433,N_9419);
or U12261 (N_12261,N_6883,N_7216);
nor U12262 (N_12262,N_8971,N_6241);
nor U12263 (N_12263,N_7878,N_9216);
nor U12264 (N_12264,N_7815,N_6120);
nor U12265 (N_12265,N_6342,N_9033);
and U12266 (N_12266,N_6117,N_8372);
and U12267 (N_12267,N_5285,N_7354);
and U12268 (N_12268,N_9798,N_7637);
or U12269 (N_12269,N_7905,N_7197);
or U12270 (N_12270,N_8225,N_9030);
nor U12271 (N_12271,N_9894,N_9376);
nor U12272 (N_12272,N_8776,N_7987);
or U12273 (N_12273,N_6807,N_7608);
xnor U12274 (N_12274,N_5495,N_5038);
xnor U12275 (N_12275,N_8600,N_9590);
nor U12276 (N_12276,N_8007,N_6533);
nor U12277 (N_12277,N_7352,N_5167);
nand U12278 (N_12278,N_5468,N_6947);
nand U12279 (N_12279,N_6165,N_5317);
or U12280 (N_12280,N_8193,N_6801);
or U12281 (N_12281,N_8072,N_9722);
and U12282 (N_12282,N_8071,N_9180);
nor U12283 (N_12283,N_8383,N_8629);
or U12284 (N_12284,N_7366,N_5144);
nor U12285 (N_12285,N_9307,N_6813);
nor U12286 (N_12286,N_7138,N_6109);
nor U12287 (N_12287,N_7821,N_9580);
nand U12288 (N_12288,N_7270,N_9232);
nand U12289 (N_12289,N_6957,N_6592);
nor U12290 (N_12290,N_9305,N_5364);
xnor U12291 (N_12291,N_6772,N_9273);
xor U12292 (N_12292,N_9152,N_6936);
nand U12293 (N_12293,N_5581,N_8068);
or U12294 (N_12294,N_5184,N_7782);
nor U12295 (N_12295,N_6708,N_9045);
or U12296 (N_12296,N_7488,N_6133);
and U12297 (N_12297,N_8714,N_7343);
and U12298 (N_12298,N_9518,N_9303);
and U12299 (N_12299,N_5312,N_7949);
or U12300 (N_12300,N_5201,N_6651);
nor U12301 (N_12301,N_5071,N_6140);
nand U12302 (N_12302,N_7682,N_8895);
and U12303 (N_12303,N_5119,N_6640);
nor U12304 (N_12304,N_7246,N_6160);
nor U12305 (N_12305,N_8441,N_6335);
or U12306 (N_12306,N_5488,N_6918);
xnor U12307 (N_12307,N_6204,N_8319);
xnor U12308 (N_12308,N_6370,N_5953);
and U12309 (N_12309,N_7368,N_8382);
or U12310 (N_12310,N_7761,N_5421);
xor U12311 (N_12311,N_8771,N_9777);
and U12312 (N_12312,N_7549,N_6880);
nand U12313 (N_12313,N_9838,N_7718);
xor U12314 (N_12314,N_9096,N_5013);
nor U12315 (N_12315,N_5879,N_6707);
and U12316 (N_12316,N_9452,N_6964);
nand U12317 (N_12317,N_5927,N_6897);
xnor U12318 (N_12318,N_6538,N_8837);
or U12319 (N_12319,N_9610,N_6357);
nand U12320 (N_12320,N_9375,N_7656);
nor U12321 (N_12321,N_5856,N_9933);
nor U12322 (N_12322,N_8341,N_9951);
or U12323 (N_12323,N_6992,N_8755);
nor U12324 (N_12324,N_5973,N_5159);
xnor U12325 (N_12325,N_8285,N_9188);
and U12326 (N_12326,N_7228,N_6182);
or U12327 (N_12327,N_5359,N_5736);
or U12328 (N_12328,N_7626,N_6811);
or U12329 (N_12329,N_8943,N_5582);
and U12330 (N_12330,N_8264,N_5267);
xnor U12331 (N_12331,N_6781,N_6400);
nand U12332 (N_12332,N_5760,N_9784);
or U12333 (N_12333,N_5452,N_9695);
or U12334 (N_12334,N_5850,N_9122);
nand U12335 (N_12335,N_8710,N_6798);
and U12336 (N_12336,N_8540,N_8085);
nor U12337 (N_12337,N_9736,N_8476);
and U12338 (N_12338,N_8705,N_6608);
or U12339 (N_12339,N_6169,N_9436);
nand U12340 (N_12340,N_5978,N_9892);
nand U12341 (N_12341,N_8889,N_6668);
xor U12342 (N_12342,N_8489,N_8675);
and U12343 (N_12343,N_5974,N_5566);
or U12344 (N_12344,N_6730,N_7719);
nor U12345 (N_12345,N_7158,N_8529);
nor U12346 (N_12346,N_9628,N_8728);
and U12347 (N_12347,N_6817,N_8354);
xnor U12348 (N_12348,N_6317,N_9241);
or U12349 (N_12349,N_5283,N_9529);
and U12350 (N_12350,N_5345,N_6589);
or U12351 (N_12351,N_7383,N_7551);
xor U12352 (N_12352,N_5064,N_8924);
nor U12353 (N_12353,N_9895,N_7178);
and U12354 (N_12354,N_6040,N_6832);
xor U12355 (N_12355,N_6349,N_8465);
or U12356 (N_12356,N_7963,N_6861);
or U12357 (N_12357,N_6988,N_5029);
nand U12358 (N_12358,N_7984,N_6266);
or U12359 (N_12359,N_8792,N_9855);
nor U12360 (N_12360,N_9107,N_9992);
or U12361 (N_12361,N_6944,N_7135);
xor U12362 (N_12362,N_6381,N_5656);
xor U12363 (N_12363,N_7592,N_5589);
nor U12364 (N_12364,N_7553,N_9159);
xnor U12365 (N_12365,N_9134,N_8498);
or U12366 (N_12366,N_7935,N_7924);
and U12367 (N_12367,N_5896,N_7109);
xor U12368 (N_12368,N_5422,N_8239);
or U12369 (N_12369,N_8597,N_8196);
xor U12370 (N_12370,N_8569,N_8956);
nor U12371 (N_12371,N_5517,N_6427);
nand U12372 (N_12372,N_9548,N_5307);
xor U12373 (N_12373,N_8690,N_8079);
nor U12374 (N_12374,N_8076,N_6101);
or U12375 (N_12375,N_6104,N_6134);
xor U12376 (N_12376,N_5833,N_8478);
and U12377 (N_12377,N_8853,N_8568);
and U12378 (N_12378,N_8087,N_7439);
or U12379 (N_12379,N_7856,N_9235);
nand U12380 (N_12380,N_6835,N_5354);
or U12381 (N_12381,N_9240,N_6197);
nand U12382 (N_12382,N_6018,N_8084);
nand U12383 (N_12383,N_9339,N_6174);
and U12384 (N_12384,N_8464,N_7613);
nor U12385 (N_12385,N_5300,N_9526);
xor U12386 (N_12386,N_5164,N_8100);
and U12387 (N_12387,N_7156,N_6792);
or U12388 (N_12388,N_5715,N_7002);
nand U12389 (N_12389,N_6158,N_8983);
or U12390 (N_12390,N_5327,N_9340);
xor U12391 (N_12391,N_7967,N_7622);
nor U12392 (N_12392,N_7579,N_6769);
nand U12393 (N_12393,N_8612,N_6810);
nand U12394 (N_12394,N_8360,N_6409);
nand U12395 (N_12395,N_9703,N_5737);
and U12396 (N_12396,N_5034,N_8243);
nor U12397 (N_12397,N_7338,N_8075);
xnor U12398 (N_12398,N_9093,N_7766);
nor U12399 (N_12399,N_8523,N_6902);
nor U12400 (N_12400,N_9008,N_5226);
and U12401 (N_12401,N_8332,N_5621);
nand U12402 (N_12402,N_7918,N_7564);
or U12403 (N_12403,N_5620,N_8831);
nor U12404 (N_12404,N_9468,N_9584);
xor U12405 (N_12405,N_9853,N_9780);
xor U12406 (N_12406,N_5031,N_5874);
or U12407 (N_12407,N_9751,N_8495);
xnor U12408 (N_12408,N_8765,N_9613);
and U12409 (N_12409,N_6244,N_6950);
xnor U12410 (N_12410,N_6638,N_9553);
xnor U12411 (N_12411,N_9884,N_8436);
or U12412 (N_12412,N_6122,N_6714);
or U12413 (N_12413,N_8808,N_8832);
nor U12414 (N_12414,N_7102,N_5630);
and U12415 (N_12415,N_9586,N_5122);
nor U12416 (N_12416,N_6678,N_7797);
and U12417 (N_12417,N_5653,N_7756);
and U12418 (N_12418,N_5516,N_9480);
nor U12419 (N_12419,N_9087,N_9112);
xor U12420 (N_12420,N_7548,N_6763);
nand U12421 (N_12421,N_5443,N_8645);
or U12422 (N_12422,N_6419,N_5349);
or U12423 (N_12423,N_9085,N_5941);
nand U12424 (N_12424,N_5719,N_5755);
or U12425 (N_12425,N_9957,N_8254);
nor U12426 (N_12426,N_7545,N_7040);
xnor U12427 (N_12427,N_7082,N_9402);
nand U12428 (N_12428,N_9369,N_7356);
xor U12429 (N_12429,N_8153,N_7617);
nand U12430 (N_12430,N_8036,N_9151);
nand U12431 (N_12431,N_6541,N_6127);
or U12432 (N_12432,N_9104,N_7054);
or U12433 (N_12433,N_5075,N_6074);
nand U12434 (N_12434,N_7730,N_6948);
and U12435 (N_12435,N_7263,N_5794);
nand U12436 (N_12436,N_7431,N_9252);
xnor U12437 (N_12437,N_9944,N_8183);
nand U12438 (N_12438,N_7108,N_7868);
and U12439 (N_12439,N_8988,N_9619);
nand U12440 (N_12440,N_5305,N_5112);
and U12441 (N_12441,N_9370,N_7802);
or U12442 (N_12442,N_5800,N_5819);
or U12443 (N_12443,N_8038,N_6665);
and U12444 (N_12444,N_6529,N_8328);
nand U12445 (N_12445,N_8463,N_7767);
nor U12446 (N_12446,N_7695,N_6336);
nand U12447 (N_12447,N_5837,N_5139);
nor U12448 (N_12448,N_5522,N_9599);
and U12449 (N_12449,N_7240,N_5202);
nand U12450 (N_12450,N_5191,N_9592);
nand U12451 (N_12451,N_6338,N_8411);
nor U12452 (N_12452,N_5699,N_5578);
nand U12453 (N_12453,N_9672,N_9346);
nor U12454 (N_12454,N_8241,N_7299);
xnor U12455 (N_12455,N_8298,N_6315);
xnor U12456 (N_12456,N_8797,N_8854);
or U12457 (N_12457,N_8191,N_6340);
or U12458 (N_12458,N_6433,N_9013);
xor U12459 (N_12459,N_8133,N_9883);
xor U12460 (N_12460,N_9042,N_8942);
xnor U12461 (N_12461,N_5066,N_9168);
xnor U12462 (N_12462,N_5601,N_6481);
nand U12463 (N_12463,N_7620,N_9758);
or U12464 (N_12464,N_8893,N_6815);
or U12465 (N_12465,N_7914,N_6030);
nand U12466 (N_12466,N_9079,N_8324);
nor U12467 (N_12467,N_5592,N_8722);
xnor U12468 (N_12468,N_9826,N_7179);
nand U12469 (N_12469,N_6314,N_6740);
or U12470 (N_12470,N_5487,N_8507);
nand U12471 (N_12471,N_9684,N_8537);
and U12472 (N_12472,N_9129,N_8548);
nand U12473 (N_12473,N_7710,N_6886);
and U12474 (N_12474,N_7925,N_6534);
xor U12475 (N_12475,N_8496,N_5605);
nand U12476 (N_12476,N_5390,N_5501);
and U12477 (N_12477,N_5889,N_7101);
xnor U12478 (N_12478,N_9019,N_7373);
xnor U12479 (N_12479,N_7039,N_9204);
xnor U12480 (N_12480,N_6443,N_6705);
nor U12481 (N_12481,N_6771,N_6803);
nand U12482 (N_12482,N_9399,N_6631);
or U12483 (N_12483,N_6061,N_9056);
and U12484 (N_12484,N_6298,N_5356);
and U12485 (N_12485,N_8376,N_5633);
and U12486 (N_12486,N_6308,N_8948);
xnor U12487 (N_12487,N_6432,N_8002);
and U12488 (N_12488,N_8267,N_8305);
xor U12489 (N_12489,N_7846,N_7804);
or U12490 (N_12490,N_5745,N_7680);
nand U12491 (N_12491,N_5662,N_6863);
and U12492 (N_12492,N_9886,N_5233);
or U12493 (N_12493,N_9759,N_7157);
xor U12494 (N_12494,N_8695,N_8668);
nand U12495 (N_12495,N_7185,N_9581);
or U12496 (N_12496,N_5861,N_6402);
or U12497 (N_12497,N_9681,N_8008);
xor U12498 (N_12498,N_7322,N_5609);
or U12499 (N_12499,N_7508,N_7533);
xnor U12500 (N_12500,N_9842,N_9877);
and U12501 (N_12501,N_8809,N_9125);
and U12502 (N_12502,N_8235,N_9378);
xnor U12503 (N_12503,N_7565,N_7626);
nor U12504 (N_12504,N_9508,N_5427);
nor U12505 (N_12505,N_8818,N_7805);
nor U12506 (N_12506,N_5536,N_9959);
nand U12507 (N_12507,N_8953,N_9156);
or U12508 (N_12508,N_6039,N_5408);
nor U12509 (N_12509,N_8153,N_9152);
or U12510 (N_12510,N_9094,N_8933);
xor U12511 (N_12511,N_6420,N_9388);
or U12512 (N_12512,N_6241,N_8859);
and U12513 (N_12513,N_7355,N_6924);
and U12514 (N_12514,N_5606,N_8189);
nor U12515 (N_12515,N_7850,N_8096);
or U12516 (N_12516,N_5550,N_8338);
nand U12517 (N_12517,N_8283,N_8729);
or U12518 (N_12518,N_6701,N_6024);
nor U12519 (N_12519,N_9312,N_9840);
nor U12520 (N_12520,N_5827,N_8738);
nand U12521 (N_12521,N_9439,N_8035);
nand U12522 (N_12522,N_5205,N_6035);
nand U12523 (N_12523,N_8565,N_8306);
nor U12524 (N_12524,N_8853,N_9790);
nand U12525 (N_12525,N_9375,N_8181);
and U12526 (N_12526,N_5359,N_7717);
or U12527 (N_12527,N_8461,N_7391);
nor U12528 (N_12528,N_5111,N_8993);
or U12529 (N_12529,N_6582,N_7854);
or U12530 (N_12530,N_6398,N_8791);
or U12531 (N_12531,N_6632,N_6030);
nor U12532 (N_12532,N_9971,N_5285);
nor U12533 (N_12533,N_6416,N_8738);
xnor U12534 (N_12534,N_6073,N_8954);
xor U12535 (N_12535,N_5123,N_7879);
or U12536 (N_12536,N_9431,N_8770);
xnor U12537 (N_12537,N_9898,N_7389);
nor U12538 (N_12538,N_6857,N_7441);
nand U12539 (N_12539,N_5189,N_6931);
and U12540 (N_12540,N_6101,N_9755);
or U12541 (N_12541,N_5129,N_5426);
nand U12542 (N_12542,N_9282,N_9342);
nand U12543 (N_12543,N_7660,N_7171);
or U12544 (N_12544,N_7094,N_6914);
or U12545 (N_12545,N_6345,N_6715);
and U12546 (N_12546,N_8417,N_9478);
or U12547 (N_12547,N_8144,N_5401);
and U12548 (N_12548,N_6857,N_7626);
or U12549 (N_12549,N_6108,N_9611);
or U12550 (N_12550,N_8842,N_5106);
nand U12551 (N_12551,N_7823,N_8297);
or U12552 (N_12552,N_5163,N_8736);
xnor U12553 (N_12553,N_8449,N_6487);
and U12554 (N_12554,N_5202,N_5861);
nor U12555 (N_12555,N_7358,N_5676);
xor U12556 (N_12556,N_7196,N_7825);
or U12557 (N_12557,N_6291,N_9619);
nor U12558 (N_12558,N_6948,N_6761);
nor U12559 (N_12559,N_8794,N_7597);
and U12560 (N_12560,N_7013,N_9083);
nand U12561 (N_12561,N_8521,N_9640);
xnor U12562 (N_12562,N_7806,N_9610);
xor U12563 (N_12563,N_5210,N_8161);
xor U12564 (N_12564,N_7362,N_5139);
or U12565 (N_12565,N_6114,N_5381);
nor U12566 (N_12566,N_7891,N_7599);
nand U12567 (N_12567,N_9833,N_5334);
xor U12568 (N_12568,N_9029,N_8873);
nand U12569 (N_12569,N_7102,N_5791);
and U12570 (N_12570,N_6134,N_6238);
nand U12571 (N_12571,N_6305,N_9033);
nor U12572 (N_12572,N_9027,N_6969);
nor U12573 (N_12573,N_5805,N_8683);
nor U12574 (N_12574,N_7354,N_7710);
nand U12575 (N_12575,N_5016,N_8873);
or U12576 (N_12576,N_7572,N_8776);
nand U12577 (N_12577,N_5005,N_6979);
and U12578 (N_12578,N_9365,N_8374);
xnor U12579 (N_12579,N_6365,N_8891);
nand U12580 (N_12580,N_9639,N_5657);
xnor U12581 (N_12581,N_5427,N_9703);
or U12582 (N_12582,N_9306,N_6817);
nand U12583 (N_12583,N_7197,N_7598);
or U12584 (N_12584,N_6805,N_8463);
xor U12585 (N_12585,N_7664,N_8511);
and U12586 (N_12586,N_8951,N_6032);
and U12587 (N_12587,N_8457,N_5806);
and U12588 (N_12588,N_9967,N_5189);
nand U12589 (N_12589,N_7358,N_7723);
xor U12590 (N_12590,N_9899,N_6535);
or U12591 (N_12591,N_7104,N_5482);
nand U12592 (N_12592,N_9300,N_6051);
nor U12593 (N_12593,N_8689,N_8706);
nand U12594 (N_12594,N_5772,N_5047);
or U12595 (N_12595,N_5677,N_8047);
or U12596 (N_12596,N_7482,N_9992);
or U12597 (N_12597,N_7883,N_7001);
or U12598 (N_12598,N_6157,N_6122);
nand U12599 (N_12599,N_7416,N_9517);
nor U12600 (N_12600,N_6436,N_6742);
nor U12601 (N_12601,N_7463,N_8005);
and U12602 (N_12602,N_7260,N_5831);
nand U12603 (N_12603,N_7648,N_5445);
and U12604 (N_12604,N_8442,N_6714);
and U12605 (N_12605,N_9247,N_9394);
xnor U12606 (N_12606,N_6039,N_8824);
xor U12607 (N_12607,N_9044,N_5915);
nor U12608 (N_12608,N_5365,N_6319);
or U12609 (N_12609,N_5132,N_7298);
nor U12610 (N_12610,N_5993,N_5805);
and U12611 (N_12611,N_7856,N_6838);
nor U12612 (N_12612,N_5279,N_9763);
nand U12613 (N_12613,N_9749,N_5822);
or U12614 (N_12614,N_9398,N_9860);
nand U12615 (N_12615,N_7957,N_7827);
xor U12616 (N_12616,N_5552,N_8493);
nand U12617 (N_12617,N_8120,N_8851);
or U12618 (N_12618,N_7550,N_8716);
nor U12619 (N_12619,N_8111,N_5744);
or U12620 (N_12620,N_9856,N_5041);
nor U12621 (N_12621,N_9063,N_7980);
xor U12622 (N_12622,N_5294,N_5843);
nand U12623 (N_12623,N_6572,N_6475);
nor U12624 (N_12624,N_5662,N_5447);
and U12625 (N_12625,N_9754,N_9698);
xnor U12626 (N_12626,N_9031,N_6854);
nand U12627 (N_12627,N_5446,N_7784);
nand U12628 (N_12628,N_7357,N_5007);
nand U12629 (N_12629,N_5708,N_7761);
nor U12630 (N_12630,N_9259,N_5332);
xor U12631 (N_12631,N_7331,N_6295);
nor U12632 (N_12632,N_8862,N_9995);
and U12633 (N_12633,N_9711,N_8163);
or U12634 (N_12634,N_5557,N_5326);
xnor U12635 (N_12635,N_5842,N_6353);
xnor U12636 (N_12636,N_6837,N_5755);
xnor U12637 (N_12637,N_8200,N_5950);
nor U12638 (N_12638,N_6147,N_5700);
and U12639 (N_12639,N_7814,N_9080);
and U12640 (N_12640,N_8330,N_5208);
xnor U12641 (N_12641,N_9039,N_5202);
or U12642 (N_12642,N_9541,N_6839);
xnor U12643 (N_12643,N_5171,N_5418);
nor U12644 (N_12644,N_7788,N_7352);
or U12645 (N_12645,N_8768,N_9998);
nand U12646 (N_12646,N_5391,N_6616);
and U12647 (N_12647,N_9799,N_9091);
nor U12648 (N_12648,N_6238,N_6294);
xnor U12649 (N_12649,N_7041,N_5380);
nand U12650 (N_12650,N_6061,N_6723);
nor U12651 (N_12651,N_7937,N_9181);
or U12652 (N_12652,N_5334,N_9202);
and U12653 (N_12653,N_8971,N_8955);
or U12654 (N_12654,N_5931,N_6884);
or U12655 (N_12655,N_5605,N_5958);
or U12656 (N_12656,N_8907,N_7419);
and U12657 (N_12657,N_7866,N_9217);
nor U12658 (N_12658,N_9118,N_7942);
xor U12659 (N_12659,N_7055,N_7502);
or U12660 (N_12660,N_9108,N_8682);
or U12661 (N_12661,N_6198,N_7717);
and U12662 (N_12662,N_7015,N_8169);
and U12663 (N_12663,N_5944,N_8982);
or U12664 (N_12664,N_7263,N_9820);
xor U12665 (N_12665,N_6401,N_8620);
and U12666 (N_12666,N_5243,N_7524);
nand U12667 (N_12667,N_9958,N_7089);
xor U12668 (N_12668,N_5749,N_9148);
and U12669 (N_12669,N_7983,N_5493);
or U12670 (N_12670,N_8603,N_9176);
or U12671 (N_12671,N_9117,N_8544);
and U12672 (N_12672,N_5892,N_8717);
or U12673 (N_12673,N_5484,N_5118);
or U12674 (N_12674,N_9285,N_8647);
or U12675 (N_12675,N_8912,N_5093);
xor U12676 (N_12676,N_5930,N_8678);
nor U12677 (N_12677,N_8217,N_8486);
xnor U12678 (N_12678,N_7802,N_8862);
or U12679 (N_12679,N_7621,N_9857);
xor U12680 (N_12680,N_7163,N_9582);
nand U12681 (N_12681,N_8034,N_8571);
xnor U12682 (N_12682,N_7136,N_6467);
xor U12683 (N_12683,N_9300,N_6491);
nor U12684 (N_12684,N_8913,N_9434);
or U12685 (N_12685,N_8256,N_6150);
xnor U12686 (N_12686,N_8532,N_7576);
or U12687 (N_12687,N_6015,N_6678);
and U12688 (N_12688,N_6607,N_5653);
nor U12689 (N_12689,N_6573,N_7963);
nand U12690 (N_12690,N_8633,N_8131);
or U12691 (N_12691,N_5808,N_8471);
and U12692 (N_12692,N_8185,N_9591);
nand U12693 (N_12693,N_7503,N_5337);
nand U12694 (N_12694,N_7986,N_6423);
nor U12695 (N_12695,N_8546,N_8261);
nand U12696 (N_12696,N_8273,N_7441);
and U12697 (N_12697,N_8891,N_6086);
nor U12698 (N_12698,N_7919,N_5570);
or U12699 (N_12699,N_6735,N_7550);
or U12700 (N_12700,N_6485,N_6392);
nor U12701 (N_12701,N_9482,N_5398);
nand U12702 (N_12702,N_7402,N_8974);
nor U12703 (N_12703,N_5793,N_7641);
nor U12704 (N_12704,N_8880,N_5152);
and U12705 (N_12705,N_8678,N_9477);
xor U12706 (N_12706,N_8656,N_8525);
xnor U12707 (N_12707,N_7401,N_6860);
and U12708 (N_12708,N_9022,N_8301);
nor U12709 (N_12709,N_8507,N_5864);
xor U12710 (N_12710,N_7054,N_8258);
nand U12711 (N_12711,N_6128,N_6844);
nor U12712 (N_12712,N_9325,N_8122);
nor U12713 (N_12713,N_7072,N_7831);
and U12714 (N_12714,N_6763,N_5140);
and U12715 (N_12715,N_8962,N_5921);
nor U12716 (N_12716,N_7969,N_8524);
nor U12717 (N_12717,N_9471,N_8085);
nor U12718 (N_12718,N_5226,N_7442);
or U12719 (N_12719,N_8932,N_9420);
xnor U12720 (N_12720,N_9725,N_5793);
and U12721 (N_12721,N_6321,N_9221);
and U12722 (N_12722,N_6314,N_5115);
and U12723 (N_12723,N_8533,N_7708);
xnor U12724 (N_12724,N_7900,N_5339);
or U12725 (N_12725,N_7552,N_8499);
and U12726 (N_12726,N_5339,N_6225);
nand U12727 (N_12727,N_5730,N_6593);
nor U12728 (N_12728,N_8336,N_7921);
nor U12729 (N_12729,N_9812,N_6805);
or U12730 (N_12730,N_5316,N_6672);
xor U12731 (N_12731,N_5105,N_5670);
xor U12732 (N_12732,N_7927,N_7820);
xor U12733 (N_12733,N_5959,N_7274);
or U12734 (N_12734,N_7416,N_6347);
xor U12735 (N_12735,N_8575,N_5283);
or U12736 (N_12736,N_5916,N_8222);
nand U12737 (N_12737,N_8039,N_6886);
or U12738 (N_12738,N_5481,N_6790);
nand U12739 (N_12739,N_5468,N_5521);
nor U12740 (N_12740,N_5726,N_9019);
xnor U12741 (N_12741,N_7846,N_7007);
or U12742 (N_12742,N_9836,N_6249);
or U12743 (N_12743,N_5842,N_6738);
or U12744 (N_12744,N_7025,N_9346);
nor U12745 (N_12745,N_9546,N_6225);
and U12746 (N_12746,N_8956,N_5697);
nor U12747 (N_12747,N_9921,N_9362);
nor U12748 (N_12748,N_8864,N_8733);
xnor U12749 (N_12749,N_8377,N_6644);
and U12750 (N_12750,N_6911,N_9189);
or U12751 (N_12751,N_9873,N_7025);
nand U12752 (N_12752,N_6597,N_6919);
or U12753 (N_12753,N_8279,N_5906);
or U12754 (N_12754,N_6716,N_9911);
or U12755 (N_12755,N_7244,N_7012);
xor U12756 (N_12756,N_6092,N_7402);
xor U12757 (N_12757,N_8653,N_5416);
nand U12758 (N_12758,N_9097,N_9710);
nor U12759 (N_12759,N_5538,N_7402);
or U12760 (N_12760,N_6676,N_6422);
xor U12761 (N_12761,N_9847,N_7996);
or U12762 (N_12762,N_7297,N_6504);
nand U12763 (N_12763,N_7063,N_8864);
nand U12764 (N_12764,N_7331,N_6423);
and U12765 (N_12765,N_7465,N_9803);
xnor U12766 (N_12766,N_7894,N_8527);
or U12767 (N_12767,N_7497,N_5549);
xnor U12768 (N_12768,N_9315,N_7048);
xnor U12769 (N_12769,N_9828,N_7952);
nor U12770 (N_12770,N_5668,N_6154);
xnor U12771 (N_12771,N_7686,N_7909);
nand U12772 (N_12772,N_9087,N_5081);
nand U12773 (N_12773,N_5672,N_9103);
or U12774 (N_12774,N_5128,N_9269);
nor U12775 (N_12775,N_6447,N_7102);
nand U12776 (N_12776,N_8435,N_7054);
nor U12777 (N_12777,N_6571,N_6505);
nor U12778 (N_12778,N_6148,N_9572);
nand U12779 (N_12779,N_8195,N_9614);
xnor U12780 (N_12780,N_7764,N_7174);
or U12781 (N_12781,N_7913,N_7720);
nor U12782 (N_12782,N_7713,N_6665);
and U12783 (N_12783,N_6679,N_8814);
xor U12784 (N_12784,N_9388,N_5682);
xor U12785 (N_12785,N_7293,N_7115);
xor U12786 (N_12786,N_6065,N_7487);
and U12787 (N_12787,N_8425,N_8117);
and U12788 (N_12788,N_6612,N_7163);
xnor U12789 (N_12789,N_6528,N_9137);
and U12790 (N_12790,N_6764,N_7501);
nor U12791 (N_12791,N_5671,N_6438);
nand U12792 (N_12792,N_9246,N_9367);
or U12793 (N_12793,N_8427,N_8587);
nand U12794 (N_12794,N_6582,N_9791);
and U12795 (N_12795,N_9884,N_7514);
xnor U12796 (N_12796,N_6155,N_8457);
nand U12797 (N_12797,N_8068,N_6259);
nand U12798 (N_12798,N_6413,N_8495);
or U12799 (N_12799,N_5225,N_8624);
nand U12800 (N_12800,N_7791,N_7385);
nand U12801 (N_12801,N_9358,N_7512);
xnor U12802 (N_12802,N_7631,N_6733);
xnor U12803 (N_12803,N_9537,N_8851);
nor U12804 (N_12804,N_9225,N_8865);
and U12805 (N_12805,N_5001,N_5913);
nor U12806 (N_12806,N_7795,N_8180);
nor U12807 (N_12807,N_7104,N_7739);
nand U12808 (N_12808,N_8793,N_6231);
or U12809 (N_12809,N_6824,N_5797);
xor U12810 (N_12810,N_9134,N_8062);
nor U12811 (N_12811,N_9393,N_9126);
and U12812 (N_12812,N_6826,N_7343);
nand U12813 (N_12813,N_6101,N_8811);
or U12814 (N_12814,N_9583,N_5951);
or U12815 (N_12815,N_9335,N_7601);
nor U12816 (N_12816,N_5924,N_5637);
or U12817 (N_12817,N_6037,N_7130);
or U12818 (N_12818,N_7446,N_7921);
and U12819 (N_12819,N_8516,N_6069);
nor U12820 (N_12820,N_8835,N_8148);
or U12821 (N_12821,N_9976,N_8512);
xor U12822 (N_12822,N_5860,N_9552);
xor U12823 (N_12823,N_8520,N_5766);
xor U12824 (N_12824,N_8898,N_7246);
nand U12825 (N_12825,N_9506,N_7942);
xnor U12826 (N_12826,N_6894,N_6701);
or U12827 (N_12827,N_7351,N_9113);
or U12828 (N_12828,N_7304,N_7337);
xnor U12829 (N_12829,N_7251,N_6388);
xnor U12830 (N_12830,N_9477,N_8373);
xor U12831 (N_12831,N_7095,N_7495);
nand U12832 (N_12832,N_5960,N_9322);
xor U12833 (N_12833,N_8802,N_6952);
or U12834 (N_12834,N_9455,N_6886);
or U12835 (N_12835,N_8011,N_8237);
nand U12836 (N_12836,N_7981,N_6551);
or U12837 (N_12837,N_6643,N_5023);
and U12838 (N_12838,N_7386,N_8506);
and U12839 (N_12839,N_5788,N_7647);
nand U12840 (N_12840,N_5394,N_6276);
xnor U12841 (N_12841,N_5218,N_5892);
nor U12842 (N_12842,N_7512,N_8782);
xor U12843 (N_12843,N_9080,N_6929);
nand U12844 (N_12844,N_6407,N_6291);
nand U12845 (N_12845,N_6415,N_6989);
and U12846 (N_12846,N_8072,N_7952);
nand U12847 (N_12847,N_7468,N_6489);
nor U12848 (N_12848,N_7727,N_7215);
nand U12849 (N_12849,N_9660,N_7676);
xnor U12850 (N_12850,N_9141,N_9356);
and U12851 (N_12851,N_7651,N_8300);
nor U12852 (N_12852,N_9766,N_6063);
and U12853 (N_12853,N_9026,N_7683);
nand U12854 (N_12854,N_7053,N_6271);
or U12855 (N_12855,N_6590,N_8926);
nor U12856 (N_12856,N_5218,N_5881);
nor U12857 (N_12857,N_5234,N_5739);
or U12858 (N_12858,N_7561,N_8661);
nor U12859 (N_12859,N_6496,N_8012);
nor U12860 (N_12860,N_7262,N_6756);
nand U12861 (N_12861,N_9586,N_8771);
or U12862 (N_12862,N_8599,N_7785);
xnor U12863 (N_12863,N_7961,N_8304);
and U12864 (N_12864,N_5372,N_6418);
nor U12865 (N_12865,N_8930,N_5184);
and U12866 (N_12866,N_7163,N_8339);
nor U12867 (N_12867,N_8562,N_9019);
nor U12868 (N_12868,N_7224,N_5139);
nor U12869 (N_12869,N_7478,N_7691);
xnor U12870 (N_12870,N_5538,N_9344);
nand U12871 (N_12871,N_8428,N_7953);
xor U12872 (N_12872,N_6940,N_9814);
and U12873 (N_12873,N_5571,N_9918);
or U12874 (N_12874,N_9371,N_9254);
or U12875 (N_12875,N_6860,N_5429);
nor U12876 (N_12876,N_8960,N_8661);
and U12877 (N_12877,N_7088,N_5288);
and U12878 (N_12878,N_9408,N_5438);
nand U12879 (N_12879,N_9363,N_5587);
xnor U12880 (N_12880,N_7647,N_6952);
xor U12881 (N_12881,N_7778,N_6121);
nand U12882 (N_12882,N_5212,N_8381);
and U12883 (N_12883,N_6264,N_8064);
or U12884 (N_12884,N_6573,N_9123);
and U12885 (N_12885,N_5565,N_6150);
or U12886 (N_12886,N_6260,N_7433);
nor U12887 (N_12887,N_6332,N_5999);
nand U12888 (N_12888,N_5243,N_6260);
nand U12889 (N_12889,N_7379,N_9460);
xor U12890 (N_12890,N_6070,N_5225);
xor U12891 (N_12891,N_5856,N_9251);
or U12892 (N_12892,N_5933,N_5322);
and U12893 (N_12893,N_6301,N_5114);
nor U12894 (N_12894,N_6392,N_8659);
and U12895 (N_12895,N_8723,N_6733);
and U12896 (N_12896,N_7250,N_5440);
nand U12897 (N_12897,N_5205,N_9391);
xor U12898 (N_12898,N_7632,N_9592);
xor U12899 (N_12899,N_6248,N_5981);
nand U12900 (N_12900,N_7842,N_8705);
nand U12901 (N_12901,N_6385,N_7074);
nor U12902 (N_12902,N_8299,N_9845);
xnor U12903 (N_12903,N_5090,N_9392);
or U12904 (N_12904,N_6062,N_8029);
or U12905 (N_12905,N_8267,N_7298);
nand U12906 (N_12906,N_8876,N_8589);
or U12907 (N_12907,N_8772,N_8045);
nand U12908 (N_12908,N_5789,N_9877);
xor U12909 (N_12909,N_8038,N_7450);
xnor U12910 (N_12910,N_9757,N_8965);
xnor U12911 (N_12911,N_8790,N_6692);
nor U12912 (N_12912,N_8207,N_5975);
nand U12913 (N_12913,N_5039,N_7471);
nand U12914 (N_12914,N_7153,N_6327);
and U12915 (N_12915,N_9651,N_5597);
nand U12916 (N_12916,N_6336,N_8273);
or U12917 (N_12917,N_9969,N_7304);
and U12918 (N_12918,N_6579,N_8524);
or U12919 (N_12919,N_5629,N_8447);
and U12920 (N_12920,N_6719,N_8778);
nand U12921 (N_12921,N_6512,N_7535);
or U12922 (N_12922,N_7094,N_9316);
nor U12923 (N_12923,N_9032,N_5059);
and U12924 (N_12924,N_9999,N_8877);
and U12925 (N_12925,N_7758,N_5972);
and U12926 (N_12926,N_8324,N_5796);
nand U12927 (N_12927,N_9244,N_8310);
nor U12928 (N_12928,N_8443,N_5609);
nand U12929 (N_12929,N_6375,N_9037);
xnor U12930 (N_12930,N_8088,N_5949);
and U12931 (N_12931,N_5009,N_8446);
nor U12932 (N_12932,N_9810,N_7344);
nand U12933 (N_12933,N_7648,N_7631);
or U12934 (N_12934,N_8808,N_5682);
or U12935 (N_12935,N_9011,N_7925);
and U12936 (N_12936,N_5652,N_9592);
nand U12937 (N_12937,N_6568,N_7032);
or U12938 (N_12938,N_6684,N_9212);
nand U12939 (N_12939,N_9075,N_7135);
nand U12940 (N_12940,N_8937,N_7925);
nor U12941 (N_12941,N_6706,N_7931);
and U12942 (N_12942,N_5741,N_6228);
nor U12943 (N_12943,N_5353,N_6347);
xnor U12944 (N_12944,N_6076,N_5317);
xnor U12945 (N_12945,N_9621,N_6322);
nand U12946 (N_12946,N_8696,N_6156);
xnor U12947 (N_12947,N_8003,N_8951);
nor U12948 (N_12948,N_7246,N_7085);
and U12949 (N_12949,N_6395,N_7492);
nor U12950 (N_12950,N_9845,N_6173);
nand U12951 (N_12951,N_5112,N_9167);
and U12952 (N_12952,N_6916,N_5856);
nand U12953 (N_12953,N_7010,N_6719);
and U12954 (N_12954,N_5617,N_8104);
and U12955 (N_12955,N_8000,N_7812);
and U12956 (N_12956,N_8007,N_8988);
xnor U12957 (N_12957,N_6673,N_8371);
nand U12958 (N_12958,N_5723,N_9864);
xnor U12959 (N_12959,N_6228,N_9317);
and U12960 (N_12960,N_5887,N_8917);
nor U12961 (N_12961,N_9527,N_6759);
nand U12962 (N_12962,N_7349,N_5575);
or U12963 (N_12963,N_9689,N_6826);
or U12964 (N_12964,N_5857,N_6326);
nand U12965 (N_12965,N_7939,N_8349);
nor U12966 (N_12966,N_8233,N_5707);
nand U12967 (N_12967,N_7525,N_9744);
nand U12968 (N_12968,N_5315,N_6780);
nand U12969 (N_12969,N_6817,N_6310);
xor U12970 (N_12970,N_8150,N_9696);
and U12971 (N_12971,N_6953,N_7837);
and U12972 (N_12972,N_7383,N_6381);
or U12973 (N_12973,N_5420,N_6938);
nand U12974 (N_12974,N_5584,N_8486);
nor U12975 (N_12975,N_9142,N_8736);
nand U12976 (N_12976,N_5080,N_8765);
nor U12977 (N_12977,N_5660,N_7740);
nand U12978 (N_12978,N_6523,N_9572);
xor U12979 (N_12979,N_6652,N_9535);
xor U12980 (N_12980,N_5960,N_6890);
or U12981 (N_12981,N_7679,N_9740);
xnor U12982 (N_12982,N_8164,N_8360);
or U12983 (N_12983,N_5269,N_7725);
or U12984 (N_12984,N_5018,N_9336);
nor U12985 (N_12985,N_5043,N_6035);
nor U12986 (N_12986,N_6890,N_7676);
xor U12987 (N_12987,N_7538,N_8147);
nor U12988 (N_12988,N_9522,N_6752);
xor U12989 (N_12989,N_5815,N_7538);
nand U12990 (N_12990,N_7145,N_8842);
or U12991 (N_12991,N_8679,N_9488);
and U12992 (N_12992,N_5083,N_7095);
xnor U12993 (N_12993,N_5795,N_5160);
nand U12994 (N_12994,N_6284,N_5419);
nor U12995 (N_12995,N_7885,N_9532);
nor U12996 (N_12996,N_6321,N_8108);
and U12997 (N_12997,N_5670,N_6828);
nand U12998 (N_12998,N_7331,N_9638);
nand U12999 (N_12999,N_9716,N_6372);
or U13000 (N_13000,N_7793,N_8891);
nand U13001 (N_13001,N_9810,N_5939);
xor U13002 (N_13002,N_6419,N_6088);
xnor U13003 (N_13003,N_6899,N_6676);
xnor U13004 (N_13004,N_6727,N_7379);
nand U13005 (N_13005,N_5629,N_6635);
nor U13006 (N_13006,N_9348,N_9866);
and U13007 (N_13007,N_6897,N_7136);
nand U13008 (N_13008,N_8482,N_9100);
nand U13009 (N_13009,N_7578,N_7100);
nand U13010 (N_13010,N_9931,N_8763);
xnor U13011 (N_13011,N_6206,N_7077);
nand U13012 (N_13012,N_5988,N_8346);
or U13013 (N_13013,N_9594,N_7471);
nand U13014 (N_13014,N_7334,N_9228);
nor U13015 (N_13015,N_7827,N_6977);
and U13016 (N_13016,N_6235,N_6040);
nor U13017 (N_13017,N_5513,N_9777);
xnor U13018 (N_13018,N_5653,N_5293);
or U13019 (N_13019,N_7413,N_6450);
nor U13020 (N_13020,N_6031,N_6618);
nor U13021 (N_13021,N_8600,N_9886);
nand U13022 (N_13022,N_7749,N_9651);
or U13023 (N_13023,N_7551,N_9693);
and U13024 (N_13024,N_8991,N_8117);
nor U13025 (N_13025,N_5866,N_8270);
xnor U13026 (N_13026,N_9215,N_9225);
or U13027 (N_13027,N_6857,N_7200);
xnor U13028 (N_13028,N_9714,N_6253);
xor U13029 (N_13029,N_9116,N_7457);
nor U13030 (N_13030,N_6062,N_8184);
nand U13031 (N_13031,N_5842,N_8769);
nor U13032 (N_13032,N_7787,N_6516);
or U13033 (N_13033,N_6446,N_5781);
or U13034 (N_13034,N_5756,N_6219);
xnor U13035 (N_13035,N_6091,N_6007);
or U13036 (N_13036,N_6441,N_7330);
and U13037 (N_13037,N_8707,N_5433);
and U13038 (N_13038,N_7810,N_7162);
or U13039 (N_13039,N_9744,N_8059);
xor U13040 (N_13040,N_8198,N_9046);
nand U13041 (N_13041,N_7486,N_5752);
or U13042 (N_13042,N_8775,N_7296);
xnor U13043 (N_13043,N_5476,N_5800);
nand U13044 (N_13044,N_6598,N_5175);
xnor U13045 (N_13045,N_5013,N_6706);
nor U13046 (N_13046,N_5295,N_9822);
or U13047 (N_13047,N_7548,N_9992);
nor U13048 (N_13048,N_6019,N_9149);
and U13049 (N_13049,N_6233,N_5487);
or U13050 (N_13050,N_8177,N_9475);
or U13051 (N_13051,N_5784,N_9801);
nand U13052 (N_13052,N_5953,N_8288);
and U13053 (N_13053,N_5992,N_8162);
or U13054 (N_13054,N_7449,N_5701);
xnor U13055 (N_13055,N_9076,N_5430);
xor U13056 (N_13056,N_9998,N_9481);
or U13057 (N_13057,N_6656,N_6691);
and U13058 (N_13058,N_6221,N_7405);
and U13059 (N_13059,N_7543,N_7695);
and U13060 (N_13060,N_9410,N_6887);
xor U13061 (N_13061,N_6808,N_6950);
and U13062 (N_13062,N_7948,N_9121);
nor U13063 (N_13063,N_8980,N_7684);
nand U13064 (N_13064,N_9866,N_5230);
nor U13065 (N_13065,N_5816,N_5118);
and U13066 (N_13066,N_6176,N_7407);
and U13067 (N_13067,N_8676,N_5069);
nand U13068 (N_13068,N_9943,N_7474);
nand U13069 (N_13069,N_8280,N_9115);
nand U13070 (N_13070,N_6693,N_5992);
nor U13071 (N_13071,N_8532,N_6849);
and U13072 (N_13072,N_9045,N_6791);
nand U13073 (N_13073,N_9642,N_7590);
nor U13074 (N_13074,N_7276,N_9027);
nor U13075 (N_13075,N_8545,N_6745);
xor U13076 (N_13076,N_9046,N_8804);
or U13077 (N_13077,N_8862,N_5756);
and U13078 (N_13078,N_6367,N_6608);
xor U13079 (N_13079,N_9597,N_6811);
and U13080 (N_13080,N_6628,N_5483);
and U13081 (N_13081,N_9827,N_6211);
nand U13082 (N_13082,N_5954,N_7978);
nor U13083 (N_13083,N_5906,N_9004);
nand U13084 (N_13084,N_5626,N_6726);
xor U13085 (N_13085,N_5413,N_7191);
nand U13086 (N_13086,N_7468,N_7160);
nor U13087 (N_13087,N_5820,N_9029);
nor U13088 (N_13088,N_6511,N_6647);
xnor U13089 (N_13089,N_7937,N_8863);
xnor U13090 (N_13090,N_9525,N_7266);
xnor U13091 (N_13091,N_7849,N_6847);
and U13092 (N_13092,N_7921,N_7488);
and U13093 (N_13093,N_8869,N_7148);
nor U13094 (N_13094,N_7290,N_6699);
or U13095 (N_13095,N_7490,N_8164);
and U13096 (N_13096,N_7646,N_9581);
and U13097 (N_13097,N_6091,N_8606);
xor U13098 (N_13098,N_8304,N_7440);
nand U13099 (N_13099,N_7615,N_7657);
or U13100 (N_13100,N_5015,N_6381);
nand U13101 (N_13101,N_8772,N_9730);
nor U13102 (N_13102,N_8613,N_8897);
nor U13103 (N_13103,N_9048,N_6048);
or U13104 (N_13104,N_6840,N_9816);
xnor U13105 (N_13105,N_8425,N_9453);
xor U13106 (N_13106,N_6783,N_8593);
and U13107 (N_13107,N_7743,N_8828);
nand U13108 (N_13108,N_8644,N_6573);
nand U13109 (N_13109,N_9548,N_8979);
or U13110 (N_13110,N_9267,N_7611);
and U13111 (N_13111,N_6911,N_9611);
nand U13112 (N_13112,N_7829,N_6167);
and U13113 (N_13113,N_9034,N_8115);
and U13114 (N_13114,N_7988,N_8495);
and U13115 (N_13115,N_6468,N_8185);
nand U13116 (N_13116,N_6116,N_9996);
xor U13117 (N_13117,N_7229,N_6964);
and U13118 (N_13118,N_6627,N_7967);
xnor U13119 (N_13119,N_7463,N_8883);
and U13120 (N_13120,N_8922,N_7002);
xor U13121 (N_13121,N_7566,N_7813);
nand U13122 (N_13122,N_8754,N_5990);
xor U13123 (N_13123,N_8825,N_9720);
nand U13124 (N_13124,N_5573,N_6847);
nor U13125 (N_13125,N_8134,N_7646);
and U13126 (N_13126,N_8942,N_5673);
nor U13127 (N_13127,N_7139,N_9152);
and U13128 (N_13128,N_6216,N_7299);
or U13129 (N_13129,N_8918,N_7444);
and U13130 (N_13130,N_8620,N_7908);
nand U13131 (N_13131,N_7074,N_6293);
and U13132 (N_13132,N_9271,N_8630);
or U13133 (N_13133,N_7684,N_9402);
nand U13134 (N_13134,N_7752,N_7159);
and U13135 (N_13135,N_7741,N_5498);
nand U13136 (N_13136,N_5261,N_5486);
xnor U13137 (N_13137,N_5756,N_7706);
xnor U13138 (N_13138,N_5238,N_7661);
and U13139 (N_13139,N_9011,N_7666);
and U13140 (N_13140,N_7262,N_7144);
and U13141 (N_13141,N_7578,N_8379);
or U13142 (N_13142,N_8192,N_6412);
and U13143 (N_13143,N_5411,N_5971);
nand U13144 (N_13144,N_5505,N_5226);
and U13145 (N_13145,N_7632,N_8432);
nor U13146 (N_13146,N_7374,N_9170);
nor U13147 (N_13147,N_9662,N_8788);
or U13148 (N_13148,N_5319,N_9958);
xnor U13149 (N_13149,N_9376,N_6704);
xnor U13150 (N_13150,N_7855,N_5869);
or U13151 (N_13151,N_5137,N_7253);
nor U13152 (N_13152,N_6749,N_6163);
nand U13153 (N_13153,N_5683,N_7223);
xnor U13154 (N_13154,N_6780,N_9418);
xnor U13155 (N_13155,N_6005,N_6258);
nor U13156 (N_13156,N_6999,N_6930);
nand U13157 (N_13157,N_5515,N_7198);
nand U13158 (N_13158,N_5728,N_5654);
or U13159 (N_13159,N_7363,N_9534);
or U13160 (N_13160,N_9239,N_5562);
or U13161 (N_13161,N_5898,N_9256);
and U13162 (N_13162,N_6913,N_9698);
nor U13163 (N_13163,N_7592,N_7357);
nor U13164 (N_13164,N_5498,N_7490);
and U13165 (N_13165,N_6969,N_9783);
nor U13166 (N_13166,N_5732,N_5886);
xor U13167 (N_13167,N_8105,N_5857);
or U13168 (N_13168,N_9115,N_7978);
and U13169 (N_13169,N_8313,N_6450);
and U13170 (N_13170,N_9083,N_9952);
nor U13171 (N_13171,N_9764,N_9669);
nor U13172 (N_13172,N_6886,N_7522);
xor U13173 (N_13173,N_6500,N_5005);
xor U13174 (N_13174,N_5007,N_9323);
and U13175 (N_13175,N_7339,N_5513);
nor U13176 (N_13176,N_5999,N_6977);
nor U13177 (N_13177,N_6483,N_8438);
and U13178 (N_13178,N_7003,N_6374);
nor U13179 (N_13179,N_6860,N_9051);
xnor U13180 (N_13180,N_5302,N_6949);
or U13181 (N_13181,N_9370,N_7253);
or U13182 (N_13182,N_5536,N_9086);
and U13183 (N_13183,N_9447,N_7765);
or U13184 (N_13184,N_7487,N_6472);
nor U13185 (N_13185,N_7662,N_6106);
xor U13186 (N_13186,N_6641,N_7213);
xor U13187 (N_13187,N_6937,N_6292);
nor U13188 (N_13188,N_9437,N_6346);
xor U13189 (N_13189,N_9886,N_8104);
nor U13190 (N_13190,N_8235,N_7670);
xnor U13191 (N_13191,N_8791,N_5392);
or U13192 (N_13192,N_9262,N_5145);
xor U13193 (N_13193,N_5014,N_6253);
nor U13194 (N_13194,N_9742,N_9630);
nand U13195 (N_13195,N_9580,N_6856);
or U13196 (N_13196,N_6374,N_7718);
xnor U13197 (N_13197,N_5979,N_8354);
xor U13198 (N_13198,N_7883,N_6712);
xnor U13199 (N_13199,N_8877,N_8596);
xor U13200 (N_13200,N_8511,N_6336);
nor U13201 (N_13201,N_6687,N_6009);
or U13202 (N_13202,N_8863,N_7318);
nor U13203 (N_13203,N_7341,N_9025);
and U13204 (N_13204,N_6665,N_6648);
and U13205 (N_13205,N_8890,N_6317);
and U13206 (N_13206,N_7794,N_6545);
nand U13207 (N_13207,N_6698,N_7054);
or U13208 (N_13208,N_5322,N_9784);
or U13209 (N_13209,N_7110,N_8257);
or U13210 (N_13210,N_5953,N_9256);
and U13211 (N_13211,N_5961,N_5074);
nor U13212 (N_13212,N_9479,N_7836);
xnor U13213 (N_13213,N_5449,N_7276);
nor U13214 (N_13214,N_6742,N_6826);
xnor U13215 (N_13215,N_7183,N_9899);
nor U13216 (N_13216,N_9142,N_9634);
xnor U13217 (N_13217,N_6798,N_9250);
or U13218 (N_13218,N_9237,N_5172);
and U13219 (N_13219,N_8516,N_7568);
nor U13220 (N_13220,N_5463,N_8958);
and U13221 (N_13221,N_6390,N_6310);
nor U13222 (N_13222,N_5722,N_6558);
or U13223 (N_13223,N_5542,N_9228);
xor U13224 (N_13224,N_9370,N_6002);
nor U13225 (N_13225,N_8990,N_6574);
xor U13226 (N_13226,N_8077,N_5683);
nor U13227 (N_13227,N_6461,N_5802);
nand U13228 (N_13228,N_9371,N_6838);
nor U13229 (N_13229,N_7365,N_8234);
nor U13230 (N_13230,N_7587,N_7225);
and U13231 (N_13231,N_8700,N_7348);
xnor U13232 (N_13232,N_7653,N_6792);
or U13233 (N_13233,N_7595,N_6514);
and U13234 (N_13234,N_8253,N_6545);
and U13235 (N_13235,N_9922,N_9736);
or U13236 (N_13236,N_9389,N_6945);
and U13237 (N_13237,N_9348,N_5917);
nand U13238 (N_13238,N_9163,N_9054);
nand U13239 (N_13239,N_9466,N_5571);
nand U13240 (N_13240,N_8558,N_7208);
nor U13241 (N_13241,N_9533,N_6784);
or U13242 (N_13242,N_8155,N_9149);
nand U13243 (N_13243,N_6150,N_6579);
nand U13244 (N_13244,N_7072,N_8474);
nand U13245 (N_13245,N_8203,N_8022);
nor U13246 (N_13246,N_6515,N_8167);
nand U13247 (N_13247,N_7396,N_6006);
or U13248 (N_13248,N_5836,N_7352);
nor U13249 (N_13249,N_6859,N_6962);
nand U13250 (N_13250,N_8565,N_7038);
or U13251 (N_13251,N_6418,N_9053);
nand U13252 (N_13252,N_8619,N_7196);
or U13253 (N_13253,N_7770,N_6001);
nand U13254 (N_13254,N_8650,N_5407);
nor U13255 (N_13255,N_9019,N_9191);
or U13256 (N_13256,N_9465,N_7712);
nand U13257 (N_13257,N_6671,N_8253);
and U13258 (N_13258,N_9747,N_5133);
xor U13259 (N_13259,N_5515,N_9511);
xnor U13260 (N_13260,N_7844,N_5107);
nor U13261 (N_13261,N_8194,N_9233);
xor U13262 (N_13262,N_8009,N_5977);
and U13263 (N_13263,N_6324,N_5554);
nand U13264 (N_13264,N_6772,N_8304);
nor U13265 (N_13265,N_9436,N_9365);
xnor U13266 (N_13266,N_9673,N_8283);
xnor U13267 (N_13267,N_6861,N_6248);
nand U13268 (N_13268,N_9823,N_7718);
xnor U13269 (N_13269,N_8619,N_8555);
or U13270 (N_13270,N_7991,N_5702);
and U13271 (N_13271,N_5972,N_7038);
or U13272 (N_13272,N_6965,N_6808);
and U13273 (N_13273,N_5754,N_6192);
nor U13274 (N_13274,N_8617,N_6808);
nor U13275 (N_13275,N_9769,N_8847);
xnor U13276 (N_13276,N_6416,N_5459);
xnor U13277 (N_13277,N_9163,N_5277);
or U13278 (N_13278,N_9886,N_5015);
xnor U13279 (N_13279,N_7201,N_7245);
and U13280 (N_13280,N_7757,N_5778);
or U13281 (N_13281,N_8437,N_9758);
xnor U13282 (N_13282,N_7791,N_5179);
nor U13283 (N_13283,N_7490,N_7437);
xnor U13284 (N_13284,N_8933,N_7720);
nand U13285 (N_13285,N_9248,N_8940);
and U13286 (N_13286,N_8011,N_9717);
nor U13287 (N_13287,N_5793,N_6349);
or U13288 (N_13288,N_7853,N_8545);
nand U13289 (N_13289,N_8285,N_6444);
nor U13290 (N_13290,N_9782,N_5522);
nor U13291 (N_13291,N_7372,N_5123);
xnor U13292 (N_13292,N_8263,N_7635);
and U13293 (N_13293,N_5711,N_5818);
xnor U13294 (N_13294,N_7108,N_5777);
xnor U13295 (N_13295,N_6596,N_7946);
nand U13296 (N_13296,N_8903,N_8715);
or U13297 (N_13297,N_9639,N_6322);
or U13298 (N_13298,N_6730,N_7306);
or U13299 (N_13299,N_7435,N_8857);
or U13300 (N_13300,N_9173,N_6186);
nor U13301 (N_13301,N_5138,N_9888);
xnor U13302 (N_13302,N_5462,N_5429);
and U13303 (N_13303,N_8469,N_9968);
xnor U13304 (N_13304,N_7729,N_9087);
nor U13305 (N_13305,N_9349,N_9605);
nand U13306 (N_13306,N_7015,N_6784);
nand U13307 (N_13307,N_9781,N_7944);
xor U13308 (N_13308,N_9254,N_6127);
nor U13309 (N_13309,N_9034,N_7795);
xor U13310 (N_13310,N_8861,N_5824);
or U13311 (N_13311,N_5025,N_6909);
nor U13312 (N_13312,N_8129,N_7910);
or U13313 (N_13313,N_7055,N_6627);
nand U13314 (N_13314,N_7064,N_7899);
nand U13315 (N_13315,N_6955,N_9132);
xor U13316 (N_13316,N_5908,N_6646);
nor U13317 (N_13317,N_8458,N_9381);
nand U13318 (N_13318,N_7797,N_9268);
and U13319 (N_13319,N_7484,N_5176);
xnor U13320 (N_13320,N_5132,N_9210);
nor U13321 (N_13321,N_8435,N_9539);
nor U13322 (N_13322,N_5097,N_7164);
and U13323 (N_13323,N_5229,N_8122);
and U13324 (N_13324,N_8980,N_6262);
nor U13325 (N_13325,N_7480,N_6586);
and U13326 (N_13326,N_7012,N_7006);
nor U13327 (N_13327,N_8820,N_8332);
or U13328 (N_13328,N_7559,N_5763);
nor U13329 (N_13329,N_8647,N_6759);
nor U13330 (N_13330,N_5655,N_8198);
nand U13331 (N_13331,N_6400,N_7203);
nor U13332 (N_13332,N_5507,N_7062);
nand U13333 (N_13333,N_8645,N_9427);
nor U13334 (N_13334,N_9970,N_5440);
nor U13335 (N_13335,N_6111,N_5663);
and U13336 (N_13336,N_9795,N_6271);
nor U13337 (N_13337,N_9919,N_7513);
or U13338 (N_13338,N_6726,N_7086);
xor U13339 (N_13339,N_7185,N_7275);
nand U13340 (N_13340,N_5819,N_8522);
nor U13341 (N_13341,N_9954,N_9895);
xor U13342 (N_13342,N_5964,N_5781);
xnor U13343 (N_13343,N_6509,N_9410);
nand U13344 (N_13344,N_9178,N_5770);
nand U13345 (N_13345,N_8117,N_9158);
or U13346 (N_13346,N_7370,N_7602);
or U13347 (N_13347,N_9572,N_9435);
and U13348 (N_13348,N_8736,N_8900);
nand U13349 (N_13349,N_8126,N_6666);
xor U13350 (N_13350,N_5547,N_7770);
or U13351 (N_13351,N_5297,N_9350);
nand U13352 (N_13352,N_6886,N_6666);
xnor U13353 (N_13353,N_8244,N_9203);
nand U13354 (N_13354,N_8283,N_9034);
or U13355 (N_13355,N_9403,N_6833);
nor U13356 (N_13356,N_8185,N_6571);
and U13357 (N_13357,N_7926,N_9622);
nor U13358 (N_13358,N_8136,N_5183);
xnor U13359 (N_13359,N_6510,N_9536);
nand U13360 (N_13360,N_9025,N_8866);
xnor U13361 (N_13361,N_5266,N_6749);
or U13362 (N_13362,N_6782,N_5106);
nand U13363 (N_13363,N_7755,N_6060);
nor U13364 (N_13364,N_9265,N_8019);
nand U13365 (N_13365,N_9906,N_9691);
nor U13366 (N_13366,N_6316,N_7897);
or U13367 (N_13367,N_7396,N_9981);
nor U13368 (N_13368,N_6461,N_9822);
and U13369 (N_13369,N_7471,N_5891);
xnor U13370 (N_13370,N_6101,N_9492);
and U13371 (N_13371,N_6192,N_6115);
nand U13372 (N_13372,N_8154,N_9996);
xor U13373 (N_13373,N_6200,N_7072);
and U13374 (N_13374,N_5344,N_5700);
nand U13375 (N_13375,N_6893,N_9842);
nand U13376 (N_13376,N_6794,N_7217);
or U13377 (N_13377,N_5728,N_6830);
xor U13378 (N_13378,N_9374,N_7691);
or U13379 (N_13379,N_6853,N_5877);
nor U13380 (N_13380,N_8711,N_5634);
nor U13381 (N_13381,N_5028,N_6427);
nor U13382 (N_13382,N_6537,N_5854);
and U13383 (N_13383,N_6176,N_9845);
or U13384 (N_13384,N_9779,N_8032);
or U13385 (N_13385,N_9139,N_5146);
and U13386 (N_13386,N_5110,N_5199);
nand U13387 (N_13387,N_5946,N_8564);
and U13388 (N_13388,N_6405,N_5704);
nor U13389 (N_13389,N_9093,N_7072);
and U13390 (N_13390,N_6195,N_6537);
or U13391 (N_13391,N_9903,N_6670);
xnor U13392 (N_13392,N_7778,N_5824);
xor U13393 (N_13393,N_8987,N_7768);
nor U13394 (N_13394,N_7822,N_7741);
and U13395 (N_13395,N_8048,N_8062);
and U13396 (N_13396,N_7146,N_6682);
xnor U13397 (N_13397,N_7214,N_5522);
xnor U13398 (N_13398,N_8790,N_8883);
nor U13399 (N_13399,N_7844,N_9573);
nand U13400 (N_13400,N_8161,N_6191);
and U13401 (N_13401,N_9756,N_6760);
nor U13402 (N_13402,N_5519,N_9768);
nor U13403 (N_13403,N_7016,N_7434);
and U13404 (N_13404,N_7418,N_5801);
nand U13405 (N_13405,N_8098,N_9054);
nand U13406 (N_13406,N_5111,N_5587);
nand U13407 (N_13407,N_8481,N_8069);
nand U13408 (N_13408,N_6962,N_7418);
nor U13409 (N_13409,N_6648,N_9693);
nand U13410 (N_13410,N_6206,N_5542);
nor U13411 (N_13411,N_7294,N_8635);
and U13412 (N_13412,N_9024,N_5657);
xnor U13413 (N_13413,N_6508,N_8683);
nand U13414 (N_13414,N_9188,N_8503);
xnor U13415 (N_13415,N_5964,N_7115);
and U13416 (N_13416,N_5737,N_9421);
or U13417 (N_13417,N_8704,N_8328);
nor U13418 (N_13418,N_8525,N_9187);
nor U13419 (N_13419,N_5038,N_9790);
or U13420 (N_13420,N_8744,N_7902);
and U13421 (N_13421,N_7520,N_8675);
xnor U13422 (N_13422,N_6477,N_6658);
nand U13423 (N_13423,N_6319,N_6209);
nor U13424 (N_13424,N_5799,N_6006);
nor U13425 (N_13425,N_8666,N_5117);
or U13426 (N_13426,N_9231,N_7608);
and U13427 (N_13427,N_9114,N_5629);
nand U13428 (N_13428,N_9524,N_6919);
nand U13429 (N_13429,N_7247,N_7304);
nor U13430 (N_13430,N_9173,N_7828);
and U13431 (N_13431,N_9679,N_5556);
nor U13432 (N_13432,N_9903,N_6051);
and U13433 (N_13433,N_5553,N_7254);
nand U13434 (N_13434,N_5875,N_5089);
nand U13435 (N_13435,N_5407,N_7505);
nor U13436 (N_13436,N_9150,N_8157);
xnor U13437 (N_13437,N_8445,N_5765);
nand U13438 (N_13438,N_8344,N_9897);
nor U13439 (N_13439,N_7995,N_5616);
or U13440 (N_13440,N_7618,N_8688);
or U13441 (N_13441,N_6542,N_8194);
or U13442 (N_13442,N_8653,N_6614);
and U13443 (N_13443,N_5681,N_6310);
nand U13444 (N_13444,N_9826,N_6005);
nor U13445 (N_13445,N_9235,N_8332);
xor U13446 (N_13446,N_9197,N_5781);
xor U13447 (N_13447,N_7656,N_6143);
and U13448 (N_13448,N_9483,N_9432);
xor U13449 (N_13449,N_7313,N_6815);
xnor U13450 (N_13450,N_7051,N_5988);
nor U13451 (N_13451,N_6711,N_8901);
or U13452 (N_13452,N_8020,N_9477);
nand U13453 (N_13453,N_5047,N_9265);
or U13454 (N_13454,N_5373,N_6989);
or U13455 (N_13455,N_9161,N_7388);
xnor U13456 (N_13456,N_8558,N_7251);
or U13457 (N_13457,N_5874,N_7280);
and U13458 (N_13458,N_7817,N_7864);
and U13459 (N_13459,N_6209,N_9361);
or U13460 (N_13460,N_9850,N_5231);
nor U13461 (N_13461,N_9375,N_9901);
nand U13462 (N_13462,N_7387,N_6095);
or U13463 (N_13463,N_9066,N_9903);
nand U13464 (N_13464,N_5835,N_6871);
or U13465 (N_13465,N_7958,N_6188);
and U13466 (N_13466,N_7643,N_9355);
or U13467 (N_13467,N_8039,N_7625);
xor U13468 (N_13468,N_7208,N_7593);
or U13469 (N_13469,N_7626,N_7745);
and U13470 (N_13470,N_6146,N_9878);
or U13471 (N_13471,N_6787,N_7152);
nand U13472 (N_13472,N_6393,N_6548);
xnor U13473 (N_13473,N_8516,N_5559);
and U13474 (N_13474,N_5506,N_5455);
nor U13475 (N_13475,N_8509,N_6230);
nand U13476 (N_13476,N_8217,N_5898);
and U13477 (N_13477,N_8630,N_8745);
xnor U13478 (N_13478,N_5186,N_5196);
xor U13479 (N_13479,N_6667,N_8500);
and U13480 (N_13480,N_7353,N_6142);
nor U13481 (N_13481,N_5272,N_7356);
nor U13482 (N_13482,N_5939,N_8174);
nor U13483 (N_13483,N_7729,N_9948);
nor U13484 (N_13484,N_6987,N_8214);
nor U13485 (N_13485,N_9486,N_5803);
or U13486 (N_13486,N_5949,N_5050);
nor U13487 (N_13487,N_9561,N_9643);
nand U13488 (N_13488,N_8280,N_5010);
nand U13489 (N_13489,N_7412,N_8094);
nor U13490 (N_13490,N_9953,N_8952);
and U13491 (N_13491,N_9081,N_5582);
nand U13492 (N_13492,N_7474,N_5570);
nand U13493 (N_13493,N_5288,N_8560);
nor U13494 (N_13494,N_9366,N_9932);
nor U13495 (N_13495,N_6937,N_5538);
or U13496 (N_13496,N_8313,N_9746);
nor U13497 (N_13497,N_7143,N_6547);
or U13498 (N_13498,N_6625,N_5147);
nor U13499 (N_13499,N_7722,N_8509);
and U13500 (N_13500,N_9499,N_8629);
nand U13501 (N_13501,N_5759,N_8049);
or U13502 (N_13502,N_9085,N_5786);
nand U13503 (N_13503,N_7327,N_6013);
and U13504 (N_13504,N_5098,N_6782);
or U13505 (N_13505,N_8964,N_9262);
nor U13506 (N_13506,N_6559,N_7862);
nor U13507 (N_13507,N_9581,N_9066);
and U13508 (N_13508,N_9845,N_7272);
nor U13509 (N_13509,N_5113,N_6048);
nand U13510 (N_13510,N_8866,N_6775);
nand U13511 (N_13511,N_7374,N_5031);
xor U13512 (N_13512,N_9972,N_8384);
xnor U13513 (N_13513,N_7485,N_6068);
nand U13514 (N_13514,N_6865,N_5785);
or U13515 (N_13515,N_8430,N_8455);
or U13516 (N_13516,N_9623,N_7821);
nor U13517 (N_13517,N_8470,N_9545);
and U13518 (N_13518,N_5144,N_7426);
or U13519 (N_13519,N_7104,N_8092);
or U13520 (N_13520,N_7521,N_5087);
xor U13521 (N_13521,N_6974,N_7643);
xor U13522 (N_13522,N_8967,N_5380);
and U13523 (N_13523,N_8801,N_5189);
and U13524 (N_13524,N_8286,N_9891);
nand U13525 (N_13525,N_6991,N_5086);
nand U13526 (N_13526,N_7503,N_5422);
or U13527 (N_13527,N_7798,N_5212);
xor U13528 (N_13528,N_5000,N_5645);
and U13529 (N_13529,N_9229,N_5424);
nor U13530 (N_13530,N_8423,N_9025);
and U13531 (N_13531,N_5591,N_5354);
nand U13532 (N_13532,N_5129,N_6125);
and U13533 (N_13533,N_6212,N_5820);
nor U13534 (N_13534,N_5207,N_7191);
xor U13535 (N_13535,N_8783,N_9703);
xnor U13536 (N_13536,N_6398,N_7893);
or U13537 (N_13537,N_5181,N_9882);
or U13538 (N_13538,N_9525,N_5340);
or U13539 (N_13539,N_7960,N_7090);
xor U13540 (N_13540,N_9650,N_8602);
nor U13541 (N_13541,N_6231,N_9662);
nor U13542 (N_13542,N_7984,N_9761);
nor U13543 (N_13543,N_8085,N_9165);
or U13544 (N_13544,N_5476,N_8189);
nand U13545 (N_13545,N_5139,N_6672);
and U13546 (N_13546,N_5572,N_7448);
nor U13547 (N_13547,N_8525,N_7209);
nand U13548 (N_13548,N_5753,N_9619);
nor U13549 (N_13549,N_7747,N_8702);
xor U13550 (N_13550,N_7697,N_5756);
or U13551 (N_13551,N_6360,N_5375);
nand U13552 (N_13552,N_7404,N_8890);
and U13553 (N_13553,N_9365,N_8972);
xnor U13554 (N_13554,N_7859,N_7993);
and U13555 (N_13555,N_5159,N_7884);
nor U13556 (N_13556,N_8386,N_6525);
or U13557 (N_13557,N_5498,N_5575);
and U13558 (N_13558,N_9451,N_6090);
nand U13559 (N_13559,N_8054,N_8929);
nand U13560 (N_13560,N_6669,N_7834);
nor U13561 (N_13561,N_7268,N_8267);
and U13562 (N_13562,N_9574,N_9988);
and U13563 (N_13563,N_9466,N_5849);
xnor U13564 (N_13564,N_6247,N_9310);
nor U13565 (N_13565,N_7836,N_6163);
nand U13566 (N_13566,N_9084,N_7617);
and U13567 (N_13567,N_5964,N_8144);
nand U13568 (N_13568,N_7519,N_6489);
nor U13569 (N_13569,N_6245,N_6093);
nor U13570 (N_13570,N_5605,N_7836);
xnor U13571 (N_13571,N_5642,N_5310);
xnor U13572 (N_13572,N_7876,N_9930);
nor U13573 (N_13573,N_9816,N_7723);
nand U13574 (N_13574,N_5472,N_5315);
nor U13575 (N_13575,N_6241,N_5012);
xor U13576 (N_13576,N_8470,N_9815);
nor U13577 (N_13577,N_8019,N_5170);
nor U13578 (N_13578,N_7534,N_7956);
nand U13579 (N_13579,N_8929,N_9185);
or U13580 (N_13580,N_8267,N_8701);
nor U13581 (N_13581,N_9636,N_6851);
or U13582 (N_13582,N_7032,N_7510);
xnor U13583 (N_13583,N_7570,N_5487);
xor U13584 (N_13584,N_5113,N_8870);
and U13585 (N_13585,N_6093,N_6422);
and U13586 (N_13586,N_7231,N_6898);
and U13587 (N_13587,N_6935,N_6200);
nand U13588 (N_13588,N_7776,N_7329);
xor U13589 (N_13589,N_7153,N_5787);
and U13590 (N_13590,N_7504,N_9576);
nand U13591 (N_13591,N_7922,N_5469);
or U13592 (N_13592,N_5593,N_6897);
or U13593 (N_13593,N_9906,N_9646);
nor U13594 (N_13594,N_6071,N_5370);
nand U13595 (N_13595,N_9448,N_6290);
xor U13596 (N_13596,N_9790,N_5239);
nor U13597 (N_13597,N_7236,N_7546);
and U13598 (N_13598,N_8149,N_6948);
nand U13599 (N_13599,N_9085,N_7129);
nand U13600 (N_13600,N_5084,N_5836);
or U13601 (N_13601,N_7389,N_6722);
xor U13602 (N_13602,N_9252,N_8462);
xor U13603 (N_13603,N_9075,N_5690);
or U13604 (N_13604,N_6330,N_5931);
nor U13605 (N_13605,N_7858,N_6264);
or U13606 (N_13606,N_6534,N_6995);
nor U13607 (N_13607,N_6399,N_7540);
and U13608 (N_13608,N_8407,N_9287);
xor U13609 (N_13609,N_8014,N_7124);
nand U13610 (N_13610,N_9971,N_5785);
or U13611 (N_13611,N_9448,N_7525);
nand U13612 (N_13612,N_7918,N_9225);
and U13613 (N_13613,N_7411,N_7941);
and U13614 (N_13614,N_7839,N_5174);
xnor U13615 (N_13615,N_6864,N_7434);
and U13616 (N_13616,N_8987,N_8644);
or U13617 (N_13617,N_8647,N_5869);
and U13618 (N_13618,N_6724,N_5987);
nand U13619 (N_13619,N_6070,N_8816);
nand U13620 (N_13620,N_7089,N_8579);
and U13621 (N_13621,N_6261,N_9545);
or U13622 (N_13622,N_5680,N_9945);
xnor U13623 (N_13623,N_5761,N_8497);
xor U13624 (N_13624,N_9787,N_8571);
nor U13625 (N_13625,N_7715,N_5237);
xor U13626 (N_13626,N_9646,N_5133);
xor U13627 (N_13627,N_9843,N_6580);
nand U13628 (N_13628,N_5039,N_9654);
nor U13629 (N_13629,N_7323,N_7592);
and U13630 (N_13630,N_5951,N_9923);
xor U13631 (N_13631,N_7827,N_6580);
nor U13632 (N_13632,N_7685,N_5352);
nand U13633 (N_13633,N_8611,N_7609);
nand U13634 (N_13634,N_6981,N_9888);
xor U13635 (N_13635,N_7684,N_5559);
nor U13636 (N_13636,N_8733,N_9016);
or U13637 (N_13637,N_6638,N_5277);
nor U13638 (N_13638,N_8952,N_5392);
or U13639 (N_13639,N_8953,N_7775);
xor U13640 (N_13640,N_5208,N_7460);
and U13641 (N_13641,N_5525,N_8726);
or U13642 (N_13642,N_7246,N_7129);
and U13643 (N_13643,N_9982,N_5651);
xnor U13644 (N_13644,N_9115,N_8429);
xnor U13645 (N_13645,N_9602,N_8640);
xor U13646 (N_13646,N_7666,N_9491);
xnor U13647 (N_13647,N_5684,N_9071);
xnor U13648 (N_13648,N_8080,N_5506);
or U13649 (N_13649,N_7395,N_8763);
or U13650 (N_13650,N_6842,N_5213);
nor U13651 (N_13651,N_6819,N_7618);
and U13652 (N_13652,N_8869,N_8053);
and U13653 (N_13653,N_5270,N_6425);
or U13654 (N_13654,N_6980,N_6739);
nor U13655 (N_13655,N_8013,N_7626);
xnor U13656 (N_13656,N_7708,N_5597);
nand U13657 (N_13657,N_9507,N_5993);
xnor U13658 (N_13658,N_6287,N_7107);
xnor U13659 (N_13659,N_9118,N_5573);
nor U13660 (N_13660,N_7409,N_8177);
nand U13661 (N_13661,N_6472,N_9636);
nor U13662 (N_13662,N_8919,N_6646);
and U13663 (N_13663,N_9676,N_9236);
xor U13664 (N_13664,N_8517,N_7628);
xnor U13665 (N_13665,N_8288,N_9401);
xor U13666 (N_13666,N_8163,N_9922);
nor U13667 (N_13667,N_8078,N_5356);
nand U13668 (N_13668,N_6974,N_8248);
or U13669 (N_13669,N_8671,N_5519);
or U13670 (N_13670,N_8083,N_7519);
nor U13671 (N_13671,N_6225,N_6008);
or U13672 (N_13672,N_7274,N_6884);
xor U13673 (N_13673,N_6413,N_6227);
nand U13674 (N_13674,N_5914,N_9166);
nand U13675 (N_13675,N_5542,N_9371);
nor U13676 (N_13676,N_5724,N_9963);
xnor U13677 (N_13677,N_5090,N_6811);
nor U13678 (N_13678,N_5008,N_5035);
nand U13679 (N_13679,N_8459,N_8625);
nor U13680 (N_13680,N_5847,N_6436);
nor U13681 (N_13681,N_6655,N_9884);
nand U13682 (N_13682,N_9204,N_9058);
nand U13683 (N_13683,N_5258,N_7678);
or U13684 (N_13684,N_7391,N_7757);
or U13685 (N_13685,N_7108,N_6394);
nor U13686 (N_13686,N_7354,N_5725);
and U13687 (N_13687,N_6198,N_5911);
or U13688 (N_13688,N_5778,N_5222);
and U13689 (N_13689,N_9892,N_6218);
xor U13690 (N_13690,N_6584,N_8630);
xnor U13691 (N_13691,N_9946,N_7390);
xnor U13692 (N_13692,N_5750,N_6893);
nand U13693 (N_13693,N_9994,N_5279);
and U13694 (N_13694,N_7209,N_7276);
or U13695 (N_13695,N_7438,N_5261);
nand U13696 (N_13696,N_9972,N_8580);
xnor U13697 (N_13697,N_5605,N_5946);
xnor U13698 (N_13698,N_9397,N_5592);
and U13699 (N_13699,N_7235,N_7796);
nand U13700 (N_13700,N_6067,N_6330);
and U13701 (N_13701,N_7927,N_8055);
nor U13702 (N_13702,N_5572,N_8487);
xor U13703 (N_13703,N_9756,N_6436);
nor U13704 (N_13704,N_7314,N_5890);
or U13705 (N_13705,N_8778,N_9541);
nor U13706 (N_13706,N_8442,N_6859);
or U13707 (N_13707,N_9784,N_5890);
nor U13708 (N_13708,N_9417,N_5142);
or U13709 (N_13709,N_5595,N_9140);
nand U13710 (N_13710,N_9106,N_8148);
xnor U13711 (N_13711,N_9159,N_8845);
xor U13712 (N_13712,N_9366,N_8664);
and U13713 (N_13713,N_9255,N_7556);
nor U13714 (N_13714,N_8670,N_7683);
or U13715 (N_13715,N_8207,N_7247);
nor U13716 (N_13716,N_6194,N_6110);
nand U13717 (N_13717,N_8628,N_6575);
or U13718 (N_13718,N_5974,N_6033);
nand U13719 (N_13719,N_9682,N_7331);
nand U13720 (N_13720,N_9333,N_5403);
or U13721 (N_13721,N_6389,N_9988);
nor U13722 (N_13722,N_5816,N_6391);
or U13723 (N_13723,N_5110,N_8143);
nor U13724 (N_13724,N_6870,N_9616);
or U13725 (N_13725,N_7923,N_5999);
xor U13726 (N_13726,N_8187,N_7814);
nand U13727 (N_13727,N_9666,N_6804);
or U13728 (N_13728,N_5777,N_5680);
nor U13729 (N_13729,N_7176,N_8137);
or U13730 (N_13730,N_6452,N_9934);
nor U13731 (N_13731,N_5149,N_8032);
or U13732 (N_13732,N_7768,N_9432);
or U13733 (N_13733,N_5261,N_9950);
or U13734 (N_13734,N_9295,N_8190);
and U13735 (N_13735,N_9179,N_7677);
and U13736 (N_13736,N_5534,N_5104);
xnor U13737 (N_13737,N_9012,N_5188);
xor U13738 (N_13738,N_8500,N_9624);
xnor U13739 (N_13739,N_6386,N_5191);
and U13740 (N_13740,N_5352,N_9845);
and U13741 (N_13741,N_5923,N_6065);
nand U13742 (N_13742,N_6934,N_9185);
nand U13743 (N_13743,N_9230,N_7045);
xor U13744 (N_13744,N_6989,N_8135);
or U13745 (N_13745,N_9831,N_6174);
nor U13746 (N_13746,N_9180,N_7276);
and U13747 (N_13747,N_9379,N_8927);
nor U13748 (N_13748,N_8637,N_8663);
nand U13749 (N_13749,N_5305,N_9380);
or U13750 (N_13750,N_9031,N_7651);
nor U13751 (N_13751,N_5349,N_5684);
xnor U13752 (N_13752,N_7922,N_7214);
nor U13753 (N_13753,N_6957,N_7663);
nor U13754 (N_13754,N_9332,N_8242);
nor U13755 (N_13755,N_6297,N_7457);
xnor U13756 (N_13756,N_9614,N_7172);
nor U13757 (N_13757,N_7438,N_7890);
and U13758 (N_13758,N_6526,N_7173);
nand U13759 (N_13759,N_5785,N_6545);
nand U13760 (N_13760,N_7131,N_5133);
and U13761 (N_13761,N_6760,N_5181);
or U13762 (N_13762,N_8963,N_9740);
and U13763 (N_13763,N_9912,N_6332);
xnor U13764 (N_13764,N_8829,N_5225);
nand U13765 (N_13765,N_5318,N_8893);
nor U13766 (N_13766,N_6487,N_6466);
or U13767 (N_13767,N_7083,N_8476);
and U13768 (N_13768,N_9365,N_8092);
nor U13769 (N_13769,N_8550,N_5835);
nand U13770 (N_13770,N_5681,N_5175);
and U13771 (N_13771,N_8045,N_5486);
xnor U13772 (N_13772,N_9531,N_5570);
xor U13773 (N_13773,N_9169,N_5248);
and U13774 (N_13774,N_7936,N_6027);
xor U13775 (N_13775,N_6475,N_9135);
and U13776 (N_13776,N_9110,N_6458);
xnor U13777 (N_13777,N_6897,N_5508);
nand U13778 (N_13778,N_5709,N_8517);
and U13779 (N_13779,N_8785,N_5947);
or U13780 (N_13780,N_6405,N_8458);
nand U13781 (N_13781,N_7681,N_6225);
or U13782 (N_13782,N_5630,N_5958);
nor U13783 (N_13783,N_8566,N_5083);
or U13784 (N_13784,N_8037,N_8075);
nor U13785 (N_13785,N_5015,N_7010);
and U13786 (N_13786,N_8856,N_5086);
nor U13787 (N_13787,N_8293,N_8464);
xnor U13788 (N_13788,N_5188,N_8937);
or U13789 (N_13789,N_5537,N_8620);
xnor U13790 (N_13790,N_9511,N_7171);
nand U13791 (N_13791,N_6422,N_7969);
xor U13792 (N_13792,N_5075,N_7892);
nand U13793 (N_13793,N_6367,N_8852);
xor U13794 (N_13794,N_5509,N_8959);
or U13795 (N_13795,N_9823,N_7501);
nor U13796 (N_13796,N_7310,N_7476);
nand U13797 (N_13797,N_6820,N_6526);
and U13798 (N_13798,N_5736,N_5121);
and U13799 (N_13799,N_7676,N_8261);
or U13800 (N_13800,N_8823,N_6394);
nand U13801 (N_13801,N_6272,N_7334);
and U13802 (N_13802,N_9041,N_6219);
xor U13803 (N_13803,N_9028,N_9831);
nor U13804 (N_13804,N_9390,N_9533);
or U13805 (N_13805,N_5613,N_5020);
xor U13806 (N_13806,N_9864,N_8796);
xnor U13807 (N_13807,N_5586,N_5530);
nor U13808 (N_13808,N_8416,N_7567);
nand U13809 (N_13809,N_6370,N_8656);
and U13810 (N_13810,N_5859,N_9902);
and U13811 (N_13811,N_8516,N_7430);
nor U13812 (N_13812,N_5180,N_8220);
xor U13813 (N_13813,N_7451,N_8947);
xnor U13814 (N_13814,N_5972,N_7709);
or U13815 (N_13815,N_7250,N_8639);
xor U13816 (N_13816,N_5700,N_9286);
nor U13817 (N_13817,N_5778,N_8141);
or U13818 (N_13818,N_6100,N_7982);
and U13819 (N_13819,N_9663,N_9821);
or U13820 (N_13820,N_6711,N_8458);
xnor U13821 (N_13821,N_5867,N_6170);
nor U13822 (N_13822,N_9452,N_9267);
xor U13823 (N_13823,N_6755,N_6769);
nand U13824 (N_13824,N_7468,N_9339);
and U13825 (N_13825,N_9384,N_8706);
xnor U13826 (N_13826,N_5530,N_6249);
or U13827 (N_13827,N_9696,N_9328);
nor U13828 (N_13828,N_6043,N_6653);
and U13829 (N_13829,N_7975,N_5212);
xnor U13830 (N_13830,N_5879,N_6722);
nand U13831 (N_13831,N_8194,N_7086);
or U13832 (N_13832,N_5976,N_9729);
or U13833 (N_13833,N_5036,N_9414);
or U13834 (N_13834,N_5229,N_5386);
xor U13835 (N_13835,N_7255,N_8058);
xnor U13836 (N_13836,N_5942,N_8105);
nand U13837 (N_13837,N_5116,N_8878);
nor U13838 (N_13838,N_8425,N_8026);
nor U13839 (N_13839,N_9405,N_5469);
and U13840 (N_13840,N_8687,N_7210);
and U13841 (N_13841,N_5431,N_7238);
nand U13842 (N_13842,N_9738,N_9165);
xnor U13843 (N_13843,N_5228,N_6394);
or U13844 (N_13844,N_5344,N_9348);
or U13845 (N_13845,N_8819,N_7699);
nand U13846 (N_13846,N_8676,N_8025);
nand U13847 (N_13847,N_9169,N_7544);
nand U13848 (N_13848,N_8425,N_8638);
or U13849 (N_13849,N_8359,N_6686);
nand U13850 (N_13850,N_6230,N_8410);
nor U13851 (N_13851,N_5482,N_7748);
xnor U13852 (N_13852,N_7730,N_5308);
and U13853 (N_13853,N_8633,N_8233);
nor U13854 (N_13854,N_5419,N_9532);
and U13855 (N_13855,N_9810,N_9591);
xnor U13856 (N_13856,N_6034,N_9458);
and U13857 (N_13857,N_5236,N_6221);
or U13858 (N_13858,N_5903,N_5416);
xnor U13859 (N_13859,N_5611,N_9895);
or U13860 (N_13860,N_8063,N_9268);
xor U13861 (N_13861,N_5983,N_6990);
and U13862 (N_13862,N_9234,N_9729);
nor U13863 (N_13863,N_9415,N_9896);
nor U13864 (N_13864,N_8093,N_5275);
nand U13865 (N_13865,N_9013,N_6493);
nand U13866 (N_13866,N_8187,N_9317);
or U13867 (N_13867,N_5811,N_8286);
or U13868 (N_13868,N_7690,N_8520);
nor U13869 (N_13869,N_6912,N_6146);
nor U13870 (N_13870,N_8923,N_8161);
and U13871 (N_13871,N_5995,N_7170);
nand U13872 (N_13872,N_6984,N_8930);
nand U13873 (N_13873,N_6632,N_7538);
xnor U13874 (N_13874,N_8674,N_9684);
and U13875 (N_13875,N_8801,N_5496);
nor U13876 (N_13876,N_8972,N_5811);
nor U13877 (N_13877,N_8152,N_8687);
xor U13878 (N_13878,N_7635,N_6325);
and U13879 (N_13879,N_7857,N_6735);
or U13880 (N_13880,N_8901,N_5692);
nor U13881 (N_13881,N_7222,N_5131);
nor U13882 (N_13882,N_5589,N_5220);
nand U13883 (N_13883,N_5690,N_5704);
and U13884 (N_13884,N_5125,N_6543);
nand U13885 (N_13885,N_9853,N_5254);
and U13886 (N_13886,N_7630,N_9885);
nor U13887 (N_13887,N_7253,N_9648);
and U13888 (N_13888,N_9492,N_8281);
nor U13889 (N_13889,N_8269,N_5356);
nor U13890 (N_13890,N_9130,N_9432);
nor U13891 (N_13891,N_8148,N_9512);
nand U13892 (N_13892,N_9832,N_6306);
nor U13893 (N_13893,N_9128,N_8252);
and U13894 (N_13894,N_5593,N_8936);
xor U13895 (N_13895,N_7670,N_5640);
xor U13896 (N_13896,N_5801,N_7217);
xor U13897 (N_13897,N_7423,N_9349);
or U13898 (N_13898,N_9024,N_7912);
or U13899 (N_13899,N_7692,N_6893);
xnor U13900 (N_13900,N_8243,N_8017);
nand U13901 (N_13901,N_7107,N_5463);
nor U13902 (N_13902,N_5886,N_6351);
nand U13903 (N_13903,N_6917,N_5099);
nand U13904 (N_13904,N_7016,N_9019);
nand U13905 (N_13905,N_6454,N_6562);
nor U13906 (N_13906,N_6329,N_6885);
xor U13907 (N_13907,N_6446,N_7739);
xor U13908 (N_13908,N_9599,N_7561);
or U13909 (N_13909,N_7001,N_5668);
nor U13910 (N_13910,N_7583,N_5932);
and U13911 (N_13911,N_9758,N_8266);
and U13912 (N_13912,N_7384,N_7627);
and U13913 (N_13913,N_6534,N_7990);
xnor U13914 (N_13914,N_5871,N_5047);
nor U13915 (N_13915,N_9159,N_7693);
nand U13916 (N_13916,N_8359,N_7819);
nor U13917 (N_13917,N_7384,N_5252);
or U13918 (N_13918,N_7377,N_8027);
nand U13919 (N_13919,N_9729,N_6501);
or U13920 (N_13920,N_6480,N_8715);
and U13921 (N_13921,N_7503,N_8962);
or U13922 (N_13922,N_6485,N_6765);
and U13923 (N_13923,N_6089,N_9902);
nor U13924 (N_13924,N_8923,N_8862);
or U13925 (N_13925,N_7963,N_5138);
or U13926 (N_13926,N_6549,N_7825);
nor U13927 (N_13927,N_7814,N_5381);
or U13928 (N_13928,N_7938,N_7394);
xnor U13929 (N_13929,N_8591,N_8992);
nor U13930 (N_13930,N_5313,N_6877);
and U13931 (N_13931,N_5259,N_9871);
or U13932 (N_13932,N_7201,N_7218);
and U13933 (N_13933,N_8742,N_8814);
nor U13934 (N_13934,N_8339,N_5782);
nand U13935 (N_13935,N_9785,N_6595);
nand U13936 (N_13936,N_9099,N_9690);
xor U13937 (N_13937,N_6572,N_6581);
nor U13938 (N_13938,N_9963,N_5023);
and U13939 (N_13939,N_5003,N_7013);
and U13940 (N_13940,N_5916,N_8417);
or U13941 (N_13941,N_6124,N_7724);
xnor U13942 (N_13942,N_9035,N_6040);
or U13943 (N_13943,N_7618,N_7125);
nor U13944 (N_13944,N_6193,N_6783);
xor U13945 (N_13945,N_8099,N_7950);
and U13946 (N_13946,N_9387,N_6729);
and U13947 (N_13947,N_9002,N_7272);
nor U13948 (N_13948,N_6373,N_8859);
or U13949 (N_13949,N_8993,N_5221);
nor U13950 (N_13950,N_8345,N_5919);
or U13951 (N_13951,N_7049,N_5691);
nand U13952 (N_13952,N_7210,N_6192);
nor U13953 (N_13953,N_6001,N_8520);
or U13954 (N_13954,N_8520,N_8467);
and U13955 (N_13955,N_6580,N_6502);
nand U13956 (N_13956,N_5314,N_5823);
or U13957 (N_13957,N_8060,N_7590);
and U13958 (N_13958,N_9192,N_5591);
nor U13959 (N_13959,N_9594,N_7666);
nand U13960 (N_13960,N_6218,N_6823);
or U13961 (N_13961,N_6842,N_7267);
and U13962 (N_13962,N_9239,N_7720);
or U13963 (N_13963,N_7120,N_9811);
xnor U13964 (N_13964,N_6267,N_6461);
and U13965 (N_13965,N_8719,N_7400);
or U13966 (N_13966,N_5030,N_6104);
or U13967 (N_13967,N_7275,N_8911);
or U13968 (N_13968,N_6347,N_5087);
and U13969 (N_13969,N_5906,N_8332);
nand U13970 (N_13970,N_7023,N_9460);
nand U13971 (N_13971,N_5714,N_9950);
xnor U13972 (N_13972,N_8463,N_7082);
nand U13973 (N_13973,N_5519,N_8426);
nand U13974 (N_13974,N_6969,N_6951);
and U13975 (N_13975,N_7059,N_6148);
or U13976 (N_13976,N_7078,N_5134);
xnor U13977 (N_13977,N_9191,N_8113);
and U13978 (N_13978,N_7579,N_6185);
nand U13979 (N_13979,N_9657,N_6098);
or U13980 (N_13980,N_7193,N_8177);
nor U13981 (N_13981,N_7375,N_7573);
xnor U13982 (N_13982,N_9995,N_8763);
nand U13983 (N_13983,N_6709,N_5689);
nor U13984 (N_13984,N_6101,N_7934);
nor U13985 (N_13985,N_6160,N_9977);
nand U13986 (N_13986,N_9076,N_8461);
or U13987 (N_13987,N_8492,N_6922);
or U13988 (N_13988,N_9334,N_8830);
and U13989 (N_13989,N_9657,N_8839);
nand U13990 (N_13990,N_9393,N_8908);
or U13991 (N_13991,N_9814,N_5172);
or U13992 (N_13992,N_8185,N_5187);
or U13993 (N_13993,N_6680,N_6778);
nand U13994 (N_13994,N_8832,N_5561);
and U13995 (N_13995,N_7589,N_9078);
or U13996 (N_13996,N_9733,N_6469);
xnor U13997 (N_13997,N_6380,N_9189);
xnor U13998 (N_13998,N_5304,N_7416);
xnor U13999 (N_13999,N_6734,N_5490);
nor U14000 (N_14000,N_6276,N_6148);
xor U14001 (N_14001,N_6538,N_8410);
and U14002 (N_14002,N_6136,N_8764);
nor U14003 (N_14003,N_9005,N_5943);
or U14004 (N_14004,N_7655,N_5617);
nand U14005 (N_14005,N_8142,N_8430);
nor U14006 (N_14006,N_8246,N_6884);
nor U14007 (N_14007,N_9586,N_8046);
nand U14008 (N_14008,N_7165,N_5472);
nor U14009 (N_14009,N_5468,N_5596);
and U14010 (N_14010,N_5157,N_8333);
nand U14011 (N_14011,N_6070,N_6041);
nand U14012 (N_14012,N_7044,N_5364);
xnor U14013 (N_14013,N_8079,N_6147);
nor U14014 (N_14014,N_7781,N_8326);
nand U14015 (N_14015,N_5544,N_6180);
and U14016 (N_14016,N_7988,N_8136);
and U14017 (N_14017,N_6869,N_9360);
nand U14018 (N_14018,N_5084,N_5899);
nand U14019 (N_14019,N_9322,N_6871);
and U14020 (N_14020,N_9284,N_8754);
nor U14021 (N_14021,N_7824,N_9836);
nor U14022 (N_14022,N_9866,N_6391);
nor U14023 (N_14023,N_5721,N_5669);
xnor U14024 (N_14024,N_6005,N_8027);
nand U14025 (N_14025,N_7245,N_8874);
nor U14026 (N_14026,N_6136,N_5196);
nor U14027 (N_14027,N_7969,N_5720);
or U14028 (N_14028,N_5390,N_9058);
xnor U14029 (N_14029,N_5011,N_8171);
nor U14030 (N_14030,N_7086,N_6269);
xor U14031 (N_14031,N_6015,N_7635);
nand U14032 (N_14032,N_7488,N_5069);
xnor U14033 (N_14033,N_6929,N_5869);
and U14034 (N_14034,N_7144,N_8892);
nor U14035 (N_14035,N_7722,N_6476);
nand U14036 (N_14036,N_9882,N_7927);
and U14037 (N_14037,N_7809,N_5473);
and U14038 (N_14038,N_6058,N_9736);
and U14039 (N_14039,N_9079,N_9038);
nor U14040 (N_14040,N_8740,N_9666);
or U14041 (N_14041,N_5739,N_5532);
nand U14042 (N_14042,N_7848,N_7087);
or U14043 (N_14043,N_6664,N_9004);
or U14044 (N_14044,N_6235,N_6140);
nand U14045 (N_14045,N_8746,N_9689);
or U14046 (N_14046,N_7919,N_5066);
and U14047 (N_14047,N_7132,N_6342);
nand U14048 (N_14048,N_9180,N_6229);
nand U14049 (N_14049,N_9802,N_6992);
or U14050 (N_14050,N_6755,N_8547);
and U14051 (N_14051,N_8754,N_9872);
xor U14052 (N_14052,N_7155,N_9290);
or U14053 (N_14053,N_8621,N_5600);
xor U14054 (N_14054,N_5391,N_5860);
and U14055 (N_14055,N_7476,N_7312);
nor U14056 (N_14056,N_5106,N_9116);
and U14057 (N_14057,N_8821,N_8085);
nand U14058 (N_14058,N_6250,N_7841);
nor U14059 (N_14059,N_5203,N_7510);
nor U14060 (N_14060,N_8717,N_6354);
nand U14061 (N_14061,N_8341,N_8725);
xnor U14062 (N_14062,N_9203,N_5003);
nor U14063 (N_14063,N_7658,N_9219);
and U14064 (N_14064,N_7386,N_6871);
nand U14065 (N_14065,N_8538,N_7658);
xnor U14066 (N_14066,N_8409,N_9665);
nand U14067 (N_14067,N_5607,N_9696);
nor U14068 (N_14068,N_6526,N_6886);
nand U14069 (N_14069,N_7476,N_7475);
and U14070 (N_14070,N_7424,N_8427);
xnor U14071 (N_14071,N_5277,N_9568);
nor U14072 (N_14072,N_9401,N_8085);
nand U14073 (N_14073,N_6657,N_6632);
and U14074 (N_14074,N_6276,N_7511);
nor U14075 (N_14075,N_9571,N_8844);
or U14076 (N_14076,N_9268,N_5401);
nand U14077 (N_14077,N_8034,N_9569);
and U14078 (N_14078,N_8125,N_7349);
or U14079 (N_14079,N_5686,N_9777);
or U14080 (N_14080,N_6688,N_8926);
or U14081 (N_14081,N_9967,N_7084);
xnor U14082 (N_14082,N_7759,N_6373);
nor U14083 (N_14083,N_5874,N_5940);
xnor U14084 (N_14084,N_6489,N_7586);
and U14085 (N_14085,N_9877,N_7469);
xnor U14086 (N_14086,N_7166,N_8269);
nand U14087 (N_14087,N_6714,N_5433);
nor U14088 (N_14088,N_5717,N_8047);
xnor U14089 (N_14089,N_8622,N_7328);
nor U14090 (N_14090,N_5007,N_5865);
nand U14091 (N_14091,N_6727,N_8893);
or U14092 (N_14092,N_9532,N_9495);
xor U14093 (N_14093,N_6693,N_6681);
nand U14094 (N_14094,N_8747,N_9635);
xnor U14095 (N_14095,N_9965,N_7546);
xnor U14096 (N_14096,N_9917,N_7673);
nor U14097 (N_14097,N_8265,N_5651);
or U14098 (N_14098,N_5545,N_6275);
or U14099 (N_14099,N_7609,N_8559);
and U14100 (N_14100,N_8616,N_9922);
and U14101 (N_14101,N_6922,N_6435);
or U14102 (N_14102,N_9538,N_8310);
or U14103 (N_14103,N_8023,N_6134);
xor U14104 (N_14104,N_8647,N_7404);
nor U14105 (N_14105,N_5644,N_5506);
nor U14106 (N_14106,N_9271,N_7361);
or U14107 (N_14107,N_8356,N_9719);
nand U14108 (N_14108,N_8146,N_7318);
or U14109 (N_14109,N_6378,N_9436);
or U14110 (N_14110,N_7797,N_6618);
nand U14111 (N_14111,N_7167,N_5607);
and U14112 (N_14112,N_6687,N_9101);
or U14113 (N_14113,N_6070,N_5027);
nand U14114 (N_14114,N_9613,N_5236);
xor U14115 (N_14115,N_5107,N_6916);
nand U14116 (N_14116,N_5701,N_9557);
nand U14117 (N_14117,N_9590,N_6692);
nor U14118 (N_14118,N_6542,N_9598);
and U14119 (N_14119,N_7703,N_5972);
nor U14120 (N_14120,N_5222,N_9517);
nor U14121 (N_14121,N_6775,N_6101);
and U14122 (N_14122,N_9142,N_8077);
xnor U14123 (N_14123,N_5031,N_7522);
or U14124 (N_14124,N_8969,N_7352);
and U14125 (N_14125,N_8395,N_5088);
nor U14126 (N_14126,N_7421,N_6565);
or U14127 (N_14127,N_9163,N_8063);
nor U14128 (N_14128,N_9117,N_8725);
xor U14129 (N_14129,N_9386,N_5316);
xnor U14130 (N_14130,N_9149,N_8844);
nand U14131 (N_14131,N_9930,N_7868);
nand U14132 (N_14132,N_5368,N_9168);
nand U14133 (N_14133,N_9558,N_7158);
nor U14134 (N_14134,N_9897,N_7143);
nor U14135 (N_14135,N_8368,N_5900);
or U14136 (N_14136,N_6613,N_8474);
and U14137 (N_14137,N_9578,N_8303);
xnor U14138 (N_14138,N_5200,N_6134);
xor U14139 (N_14139,N_5702,N_7199);
or U14140 (N_14140,N_5163,N_8931);
nand U14141 (N_14141,N_8082,N_8983);
xor U14142 (N_14142,N_8952,N_7174);
or U14143 (N_14143,N_9703,N_6848);
nor U14144 (N_14144,N_5732,N_5056);
and U14145 (N_14145,N_9666,N_7569);
and U14146 (N_14146,N_5786,N_9351);
and U14147 (N_14147,N_5634,N_6786);
xnor U14148 (N_14148,N_9194,N_5251);
nand U14149 (N_14149,N_6397,N_7722);
nand U14150 (N_14150,N_8688,N_6259);
nor U14151 (N_14151,N_8525,N_6435);
or U14152 (N_14152,N_8013,N_5067);
nor U14153 (N_14153,N_6178,N_9495);
xnor U14154 (N_14154,N_6239,N_8539);
xor U14155 (N_14155,N_5091,N_9646);
nand U14156 (N_14156,N_8881,N_9389);
xor U14157 (N_14157,N_6546,N_9146);
or U14158 (N_14158,N_7976,N_6584);
nand U14159 (N_14159,N_8413,N_9556);
nor U14160 (N_14160,N_8079,N_5188);
and U14161 (N_14161,N_6095,N_7857);
and U14162 (N_14162,N_7390,N_6410);
nand U14163 (N_14163,N_5056,N_6751);
xor U14164 (N_14164,N_9780,N_6782);
nand U14165 (N_14165,N_9400,N_9308);
nand U14166 (N_14166,N_5671,N_9106);
or U14167 (N_14167,N_8052,N_7328);
nand U14168 (N_14168,N_5896,N_6858);
nand U14169 (N_14169,N_8689,N_7081);
and U14170 (N_14170,N_6592,N_5701);
or U14171 (N_14171,N_6078,N_8674);
or U14172 (N_14172,N_9895,N_8195);
or U14173 (N_14173,N_9566,N_9648);
xnor U14174 (N_14174,N_8472,N_5281);
nor U14175 (N_14175,N_5396,N_6402);
or U14176 (N_14176,N_7886,N_8201);
and U14177 (N_14177,N_7531,N_5588);
or U14178 (N_14178,N_6774,N_5781);
nor U14179 (N_14179,N_9272,N_8468);
nand U14180 (N_14180,N_9279,N_8667);
xnor U14181 (N_14181,N_6849,N_8084);
xor U14182 (N_14182,N_7662,N_9204);
and U14183 (N_14183,N_6544,N_6683);
nor U14184 (N_14184,N_8896,N_7537);
nor U14185 (N_14185,N_5944,N_6178);
nor U14186 (N_14186,N_9356,N_7628);
or U14187 (N_14187,N_6622,N_8985);
and U14188 (N_14188,N_9192,N_5226);
xor U14189 (N_14189,N_6446,N_6472);
and U14190 (N_14190,N_5665,N_5392);
xor U14191 (N_14191,N_9955,N_8262);
xor U14192 (N_14192,N_9778,N_5891);
nor U14193 (N_14193,N_7736,N_5306);
and U14194 (N_14194,N_9066,N_7282);
xnor U14195 (N_14195,N_6839,N_8370);
nand U14196 (N_14196,N_5830,N_8528);
xor U14197 (N_14197,N_8715,N_6500);
nand U14198 (N_14198,N_5527,N_7614);
nor U14199 (N_14199,N_6682,N_7377);
nand U14200 (N_14200,N_5707,N_9723);
xor U14201 (N_14201,N_8596,N_6095);
nand U14202 (N_14202,N_7680,N_6656);
xnor U14203 (N_14203,N_6486,N_9381);
and U14204 (N_14204,N_8143,N_8024);
or U14205 (N_14205,N_5787,N_7766);
and U14206 (N_14206,N_9897,N_5731);
nand U14207 (N_14207,N_6105,N_6818);
nor U14208 (N_14208,N_6676,N_6504);
nand U14209 (N_14209,N_7931,N_5108);
nand U14210 (N_14210,N_8842,N_5254);
nand U14211 (N_14211,N_8613,N_7115);
nor U14212 (N_14212,N_6173,N_7683);
and U14213 (N_14213,N_5412,N_5541);
xor U14214 (N_14214,N_6694,N_5581);
nor U14215 (N_14215,N_9882,N_5320);
or U14216 (N_14216,N_7999,N_8556);
or U14217 (N_14217,N_9918,N_5629);
nand U14218 (N_14218,N_9365,N_6999);
xnor U14219 (N_14219,N_9494,N_5432);
nor U14220 (N_14220,N_6558,N_7953);
nor U14221 (N_14221,N_5246,N_6662);
and U14222 (N_14222,N_5904,N_6411);
or U14223 (N_14223,N_7496,N_8273);
xnor U14224 (N_14224,N_6384,N_8302);
or U14225 (N_14225,N_5048,N_7936);
or U14226 (N_14226,N_8747,N_5294);
nand U14227 (N_14227,N_5500,N_9367);
xor U14228 (N_14228,N_7594,N_8247);
nor U14229 (N_14229,N_9692,N_5760);
nand U14230 (N_14230,N_5497,N_7917);
and U14231 (N_14231,N_9156,N_9719);
nor U14232 (N_14232,N_6102,N_7503);
xnor U14233 (N_14233,N_8627,N_9285);
xnor U14234 (N_14234,N_8269,N_9545);
xnor U14235 (N_14235,N_5632,N_6804);
xor U14236 (N_14236,N_5582,N_6352);
nand U14237 (N_14237,N_7322,N_6840);
xnor U14238 (N_14238,N_7604,N_5482);
and U14239 (N_14239,N_9261,N_5247);
and U14240 (N_14240,N_8970,N_9768);
or U14241 (N_14241,N_8518,N_8397);
xor U14242 (N_14242,N_6489,N_6590);
xor U14243 (N_14243,N_8095,N_5477);
and U14244 (N_14244,N_9972,N_8534);
or U14245 (N_14245,N_5978,N_9060);
xor U14246 (N_14246,N_9324,N_6762);
and U14247 (N_14247,N_7063,N_8181);
nor U14248 (N_14248,N_5555,N_9401);
and U14249 (N_14249,N_6697,N_6336);
xor U14250 (N_14250,N_5183,N_7001);
nor U14251 (N_14251,N_8736,N_5769);
or U14252 (N_14252,N_7555,N_9977);
and U14253 (N_14253,N_6199,N_7525);
nand U14254 (N_14254,N_6781,N_6699);
xnor U14255 (N_14255,N_8897,N_7618);
or U14256 (N_14256,N_9552,N_8396);
xnor U14257 (N_14257,N_9604,N_8251);
xnor U14258 (N_14258,N_7503,N_8069);
or U14259 (N_14259,N_8664,N_7564);
or U14260 (N_14260,N_9544,N_9925);
nor U14261 (N_14261,N_8654,N_6386);
and U14262 (N_14262,N_8910,N_8957);
nand U14263 (N_14263,N_8585,N_9914);
and U14264 (N_14264,N_9710,N_5084);
and U14265 (N_14265,N_8453,N_9453);
nand U14266 (N_14266,N_8640,N_9107);
nor U14267 (N_14267,N_6814,N_9591);
or U14268 (N_14268,N_5032,N_6125);
or U14269 (N_14269,N_8335,N_7189);
nor U14270 (N_14270,N_6405,N_5423);
xor U14271 (N_14271,N_7434,N_8225);
nor U14272 (N_14272,N_7211,N_8665);
xnor U14273 (N_14273,N_9163,N_8158);
nand U14274 (N_14274,N_8603,N_5576);
xor U14275 (N_14275,N_7482,N_7747);
nor U14276 (N_14276,N_8577,N_8337);
xnor U14277 (N_14277,N_6249,N_9788);
xnor U14278 (N_14278,N_8637,N_8354);
nand U14279 (N_14279,N_9529,N_6305);
and U14280 (N_14280,N_6339,N_8542);
and U14281 (N_14281,N_7532,N_9810);
and U14282 (N_14282,N_9995,N_7207);
xor U14283 (N_14283,N_6868,N_6957);
nand U14284 (N_14284,N_6035,N_5293);
or U14285 (N_14285,N_5138,N_8619);
nand U14286 (N_14286,N_8054,N_7401);
nor U14287 (N_14287,N_8342,N_8846);
or U14288 (N_14288,N_7734,N_7186);
nand U14289 (N_14289,N_8940,N_6399);
or U14290 (N_14290,N_8969,N_6791);
or U14291 (N_14291,N_5637,N_5728);
xnor U14292 (N_14292,N_9611,N_9086);
or U14293 (N_14293,N_9028,N_9773);
nand U14294 (N_14294,N_9721,N_9540);
or U14295 (N_14295,N_6374,N_8573);
xnor U14296 (N_14296,N_8773,N_9112);
nor U14297 (N_14297,N_9739,N_5684);
or U14298 (N_14298,N_8094,N_9304);
or U14299 (N_14299,N_7811,N_8524);
nand U14300 (N_14300,N_5156,N_6535);
and U14301 (N_14301,N_9275,N_5443);
and U14302 (N_14302,N_5833,N_6054);
nor U14303 (N_14303,N_5195,N_7029);
xor U14304 (N_14304,N_6834,N_7221);
xor U14305 (N_14305,N_7721,N_5880);
xnor U14306 (N_14306,N_8581,N_6882);
xnor U14307 (N_14307,N_9607,N_9904);
nor U14308 (N_14308,N_8905,N_5644);
xor U14309 (N_14309,N_7548,N_5382);
xnor U14310 (N_14310,N_5380,N_9374);
or U14311 (N_14311,N_5359,N_8529);
or U14312 (N_14312,N_6275,N_8607);
or U14313 (N_14313,N_7330,N_5510);
xor U14314 (N_14314,N_5739,N_7793);
nor U14315 (N_14315,N_6839,N_8097);
nand U14316 (N_14316,N_5308,N_8251);
or U14317 (N_14317,N_5342,N_8149);
and U14318 (N_14318,N_5869,N_8364);
or U14319 (N_14319,N_5572,N_8047);
nor U14320 (N_14320,N_6622,N_5344);
nand U14321 (N_14321,N_7632,N_5065);
nor U14322 (N_14322,N_9577,N_8887);
and U14323 (N_14323,N_5068,N_7904);
xor U14324 (N_14324,N_7543,N_9564);
and U14325 (N_14325,N_6020,N_8333);
or U14326 (N_14326,N_9767,N_9331);
xor U14327 (N_14327,N_5014,N_8391);
nor U14328 (N_14328,N_9889,N_7339);
or U14329 (N_14329,N_9596,N_9170);
nand U14330 (N_14330,N_5950,N_5286);
nor U14331 (N_14331,N_6433,N_7144);
and U14332 (N_14332,N_9532,N_7364);
xnor U14333 (N_14333,N_6970,N_6638);
and U14334 (N_14334,N_9990,N_9267);
and U14335 (N_14335,N_8920,N_6475);
xor U14336 (N_14336,N_5769,N_6677);
nand U14337 (N_14337,N_7284,N_9523);
nor U14338 (N_14338,N_6144,N_7324);
or U14339 (N_14339,N_9226,N_7144);
and U14340 (N_14340,N_6793,N_8528);
nand U14341 (N_14341,N_6793,N_6584);
and U14342 (N_14342,N_7902,N_7661);
nor U14343 (N_14343,N_9447,N_9505);
and U14344 (N_14344,N_7888,N_7548);
nand U14345 (N_14345,N_8015,N_9542);
or U14346 (N_14346,N_9649,N_5037);
and U14347 (N_14347,N_5780,N_5763);
nand U14348 (N_14348,N_8802,N_9414);
xnor U14349 (N_14349,N_6162,N_5646);
nand U14350 (N_14350,N_8673,N_5320);
xor U14351 (N_14351,N_6309,N_6890);
nand U14352 (N_14352,N_7395,N_9393);
or U14353 (N_14353,N_7586,N_9493);
nand U14354 (N_14354,N_5263,N_5575);
nor U14355 (N_14355,N_9488,N_6732);
and U14356 (N_14356,N_7106,N_7786);
or U14357 (N_14357,N_8507,N_8653);
nor U14358 (N_14358,N_7188,N_7047);
or U14359 (N_14359,N_8778,N_5424);
nor U14360 (N_14360,N_8909,N_7662);
nand U14361 (N_14361,N_7345,N_5285);
nand U14362 (N_14362,N_6584,N_5836);
nand U14363 (N_14363,N_5791,N_6674);
nand U14364 (N_14364,N_6647,N_6359);
or U14365 (N_14365,N_5810,N_9275);
and U14366 (N_14366,N_7337,N_5144);
xor U14367 (N_14367,N_8732,N_6860);
nand U14368 (N_14368,N_9030,N_9796);
nor U14369 (N_14369,N_9053,N_8714);
nor U14370 (N_14370,N_9685,N_8294);
or U14371 (N_14371,N_6654,N_9107);
and U14372 (N_14372,N_6733,N_5186);
nand U14373 (N_14373,N_6560,N_9915);
xnor U14374 (N_14374,N_8588,N_5514);
or U14375 (N_14375,N_5053,N_8640);
nand U14376 (N_14376,N_8455,N_7984);
xnor U14377 (N_14377,N_9348,N_7181);
nand U14378 (N_14378,N_7583,N_9198);
or U14379 (N_14379,N_9248,N_7498);
xor U14380 (N_14380,N_7216,N_6570);
nand U14381 (N_14381,N_7800,N_8216);
nor U14382 (N_14382,N_6997,N_9954);
nand U14383 (N_14383,N_6048,N_7925);
nand U14384 (N_14384,N_9575,N_7816);
or U14385 (N_14385,N_6897,N_7489);
and U14386 (N_14386,N_7488,N_5725);
xor U14387 (N_14387,N_6034,N_6906);
or U14388 (N_14388,N_6022,N_5765);
nor U14389 (N_14389,N_5487,N_5135);
nor U14390 (N_14390,N_5496,N_6708);
xor U14391 (N_14391,N_6372,N_8448);
nor U14392 (N_14392,N_5614,N_5360);
nand U14393 (N_14393,N_6244,N_9013);
nand U14394 (N_14394,N_5553,N_5043);
xnor U14395 (N_14395,N_5190,N_9121);
and U14396 (N_14396,N_9480,N_7188);
or U14397 (N_14397,N_6885,N_5635);
nor U14398 (N_14398,N_5074,N_7681);
or U14399 (N_14399,N_5423,N_7290);
xor U14400 (N_14400,N_5420,N_9041);
and U14401 (N_14401,N_8663,N_8847);
or U14402 (N_14402,N_6999,N_8187);
nor U14403 (N_14403,N_7844,N_5448);
xnor U14404 (N_14404,N_8435,N_9799);
xnor U14405 (N_14405,N_9757,N_7097);
and U14406 (N_14406,N_8545,N_6181);
nand U14407 (N_14407,N_9369,N_8763);
xnor U14408 (N_14408,N_9763,N_7107);
nand U14409 (N_14409,N_7898,N_6813);
xnor U14410 (N_14410,N_8842,N_8491);
xnor U14411 (N_14411,N_9558,N_7234);
and U14412 (N_14412,N_7321,N_9921);
nand U14413 (N_14413,N_5763,N_8792);
nand U14414 (N_14414,N_5862,N_8571);
xnor U14415 (N_14415,N_8773,N_6298);
and U14416 (N_14416,N_9999,N_8390);
or U14417 (N_14417,N_6640,N_9654);
xor U14418 (N_14418,N_8992,N_6728);
nand U14419 (N_14419,N_6567,N_9153);
or U14420 (N_14420,N_6628,N_7032);
and U14421 (N_14421,N_7958,N_8083);
nand U14422 (N_14422,N_9881,N_7665);
xnor U14423 (N_14423,N_8139,N_8088);
or U14424 (N_14424,N_9960,N_7146);
or U14425 (N_14425,N_5455,N_9154);
xor U14426 (N_14426,N_6161,N_8814);
nand U14427 (N_14427,N_5009,N_8552);
nor U14428 (N_14428,N_5738,N_8856);
or U14429 (N_14429,N_7300,N_6760);
nand U14430 (N_14430,N_5854,N_5262);
nor U14431 (N_14431,N_5081,N_6571);
and U14432 (N_14432,N_9962,N_6773);
or U14433 (N_14433,N_6326,N_8265);
or U14434 (N_14434,N_9707,N_7282);
nor U14435 (N_14435,N_6950,N_7027);
xnor U14436 (N_14436,N_8136,N_8868);
xnor U14437 (N_14437,N_8611,N_6486);
and U14438 (N_14438,N_8171,N_9636);
and U14439 (N_14439,N_5615,N_6767);
or U14440 (N_14440,N_7696,N_8780);
nor U14441 (N_14441,N_7376,N_9392);
or U14442 (N_14442,N_5307,N_5156);
nand U14443 (N_14443,N_7997,N_5425);
and U14444 (N_14444,N_6969,N_7977);
nor U14445 (N_14445,N_5164,N_5423);
xnor U14446 (N_14446,N_9347,N_5971);
nor U14447 (N_14447,N_5166,N_6093);
xnor U14448 (N_14448,N_7435,N_6603);
nor U14449 (N_14449,N_9352,N_6892);
or U14450 (N_14450,N_9007,N_8198);
and U14451 (N_14451,N_9897,N_9049);
xor U14452 (N_14452,N_6107,N_7474);
nand U14453 (N_14453,N_9569,N_8622);
nor U14454 (N_14454,N_7793,N_9068);
xor U14455 (N_14455,N_6532,N_5060);
nand U14456 (N_14456,N_6491,N_6800);
and U14457 (N_14457,N_5246,N_9866);
nand U14458 (N_14458,N_9045,N_7336);
xor U14459 (N_14459,N_9212,N_6367);
and U14460 (N_14460,N_8135,N_5484);
and U14461 (N_14461,N_6078,N_8180);
and U14462 (N_14462,N_6250,N_6129);
nand U14463 (N_14463,N_7735,N_8287);
or U14464 (N_14464,N_6764,N_5161);
nand U14465 (N_14465,N_6061,N_9704);
nor U14466 (N_14466,N_8683,N_7529);
or U14467 (N_14467,N_7006,N_6544);
or U14468 (N_14468,N_7773,N_8147);
nand U14469 (N_14469,N_9417,N_5464);
nor U14470 (N_14470,N_8532,N_7537);
xor U14471 (N_14471,N_7443,N_9048);
xnor U14472 (N_14472,N_9410,N_6382);
nor U14473 (N_14473,N_9656,N_7701);
or U14474 (N_14474,N_5563,N_9545);
and U14475 (N_14475,N_7271,N_6575);
or U14476 (N_14476,N_5479,N_5614);
nor U14477 (N_14477,N_6610,N_7827);
xor U14478 (N_14478,N_5758,N_7815);
xnor U14479 (N_14479,N_9948,N_6624);
and U14480 (N_14480,N_5204,N_6007);
nand U14481 (N_14481,N_5161,N_6946);
xor U14482 (N_14482,N_6585,N_6102);
xor U14483 (N_14483,N_7550,N_6015);
and U14484 (N_14484,N_7485,N_8135);
nand U14485 (N_14485,N_8593,N_8927);
nor U14486 (N_14486,N_6688,N_7931);
and U14487 (N_14487,N_9947,N_9855);
or U14488 (N_14488,N_8529,N_9686);
or U14489 (N_14489,N_9613,N_5059);
nor U14490 (N_14490,N_8184,N_7338);
or U14491 (N_14491,N_9128,N_8930);
and U14492 (N_14492,N_9170,N_9348);
or U14493 (N_14493,N_5008,N_9798);
xor U14494 (N_14494,N_5204,N_9971);
or U14495 (N_14495,N_9216,N_5982);
nand U14496 (N_14496,N_5581,N_8076);
nand U14497 (N_14497,N_7245,N_8739);
and U14498 (N_14498,N_9439,N_5378);
or U14499 (N_14499,N_6252,N_6116);
xnor U14500 (N_14500,N_7536,N_7430);
xnor U14501 (N_14501,N_6327,N_8005);
and U14502 (N_14502,N_7576,N_7991);
and U14503 (N_14503,N_6429,N_9561);
nor U14504 (N_14504,N_9679,N_8931);
and U14505 (N_14505,N_6886,N_7282);
nor U14506 (N_14506,N_5893,N_8218);
nand U14507 (N_14507,N_5691,N_9836);
nand U14508 (N_14508,N_6655,N_5374);
and U14509 (N_14509,N_5261,N_7955);
and U14510 (N_14510,N_5054,N_5572);
xor U14511 (N_14511,N_8495,N_6458);
nor U14512 (N_14512,N_8104,N_7858);
nand U14513 (N_14513,N_8895,N_5723);
nor U14514 (N_14514,N_8683,N_7966);
nand U14515 (N_14515,N_6412,N_9766);
and U14516 (N_14516,N_9711,N_8566);
nor U14517 (N_14517,N_6966,N_6253);
nor U14518 (N_14518,N_5738,N_7804);
nor U14519 (N_14519,N_6983,N_6249);
nand U14520 (N_14520,N_7899,N_9392);
nor U14521 (N_14521,N_5416,N_7879);
nor U14522 (N_14522,N_8945,N_9317);
or U14523 (N_14523,N_8026,N_9431);
or U14524 (N_14524,N_8619,N_7736);
or U14525 (N_14525,N_5645,N_9418);
or U14526 (N_14526,N_7440,N_8072);
xnor U14527 (N_14527,N_9517,N_9311);
or U14528 (N_14528,N_8429,N_6407);
xnor U14529 (N_14529,N_9913,N_8554);
nor U14530 (N_14530,N_7147,N_5329);
nand U14531 (N_14531,N_6935,N_6718);
and U14532 (N_14532,N_8947,N_9090);
xor U14533 (N_14533,N_8995,N_6093);
nand U14534 (N_14534,N_5430,N_8055);
and U14535 (N_14535,N_7096,N_9017);
and U14536 (N_14536,N_6530,N_7432);
xnor U14537 (N_14537,N_7631,N_8386);
and U14538 (N_14538,N_6307,N_6144);
or U14539 (N_14539,N_8313,N_7226);
and U14540 (N_14540,N_7351,N_7990);
xnor U14541 (N_14541,N_7969,N_7918);
xor U14542 (N_14542,N_6360,N_8347);
or U14543 (N_14543,N_6899,N_6288);
and U14544 (N_14544,N_7239,N_9209);
xor U14545 (N_14545,N_8871,N_9963);
xor U14546 (N_14546,N_8285,N_7243);
or U14547 (N_14547,N_5418,N_5297);
xnor U14548 (N_14548,N_5578,N_9432);
xor U14549 (N_14549,N_5228,N_7666);
and U14550 (N_14550,N_8541,N_7848);
and U14551 (N_14551,N_8150,N_5600);
xor U14552 (N_14552,N_7372,N_5227);
and U14553 (N_14553,N_7765,N_8736);
or U14554 (N_14554,N_5609,N_6009);
xnor U14555 (N_14555,N_9311,N_6628);
xnor U14556 (N_14556,N_9305,N_8441);
and U14557 (N_14557,N_6415,N_5409);
or U14558 (N_14558,N_5732,N_9270);
xnor U14559 (N_14559,N_6561,N_8663);
or U14560 (N_14560,N_6594,N_6656);
nand U14561 (N_14561,N_8207,N_6671);
nor U14562 (N_14562,N_8255,N_8759);
nand U14563 (N_14563,N_9067,N_8740);
or U14564 (N_14564,N_8815,N_6768);
or U14565 (N_14565,N_8782,N_6418);
nor U14566 (N_14566,N_7209,N_9559);
and U14567 (N_14567,N_9114,N_5975);
and U14568 (N_14568,N_8302,N_8788);
and U14569 (N_14569,N_7804,N_8206);
and U14570 (N_14570,N_9514,N_8983);
nand U14571 (N_14571,N_7974,N_5046);
xnor U14572 (N_14572,N_7196,N_5697);
nand U14573 (N_14573,N_5334,N_5733);
nand U14574 (N_14574,N_7750,N_8304);
xor U14575 (N_14575,N_5324,N_9084);
xor U14576 (N_14576,N_7669,N_8695);
and U14577 (N_14577,N_9307,N_5925);
nand U14578 (N_14578,N_6841,N_6694);
xor U14579 (N_14579,N_6041,N_7350);
xor U14580 (N_14580,N_5291,N_5793);
nand U14581 (N_14581,N_5067,N_9602);
or U14582 (N_14582,N_6250,N_8071);
nor U14583 (N_14583,N_6406,N_5767);
xor U14584 (N_14584,N_7400,N_6595);
nor U14585 (N_14585,N_9138,N_8251);
or U14586 (N_14586,N_5112,N_5686);
and U14587 (N_14587,N_5592,N_5726);
and U14588 (N_14588,N_6998,N_7538);
nor U14589 (N_14589,N_7664,N_8978);
or U14590 (N_14590,N_9389,N_6333);
and U14591 (N_14591,N_9889,N_9093);
nand U14592 (N_14592,N_7838,N_5609);
nand U14593 (N_14593,N_6575,N_8775);
nor U14594 (N_14594,N_8399,N_7076);
nor U14595 (N_14595,N_6140,N_8573);
nand U14596 (N_14596,N_9277,N_5746);
or U14597 (N_14597,N_6541,N_5841);
nand U14598 (N_14598,N_5675,N_6810);
and U14599 (N_14599,N_6401,N_7742);
nand U14600 (N_14600,N_6291,N_7094);
nand U14601 (N_14601,N_6230,N_8614);
nand U14602 (N_14602,N_6241,N_6600);
or U14603 (N_14603,N_6529,N_7493);
nand U14604 (N_14604,N_5188,N_6294);
nor U14605 (N_14605,N_5641,N_9227);
nor U14606 (N_14606,N_7617,N_8693);
nand U14607 (N_14607,N_9920,N_6326);
nor U14608 (N_14608,N_8943,N_6203);
xor U14609 (N_14609,N_7252,N_8586);
and U14610 (N_14610,N_8640,N_6026);
or U14611 (N_14611,N_9028,N_5339);
or U14612 (N_14612,N_7396,N_5572);
and U14613 (N_14613,N_6295,N_7498);
nor U14614 (N_14614,N_8469,N_6276);
nor U14615 (N_14615,N_6157,N_7707);
nand U14616 (N_14616,N_5526,N_9635);
nor U14617 (N_14617,N_8993,N_5521);
xor U14618 (N_14618,N_7494,N_7782);
nand U14619 (N_14619,N_8642,N_6222);
nor U14620 (N_14620,N_8863,N_9271);
nand U14621 (N_14621,N_7137,N_6422);
nand U14622 (N_14622,N_5134,N_8090);
nor U14623 (N_14623,N_7458,N_5570);
or U14624 (N_14624,N_9001,N_7733);
nand U14625 (N_14625,N_5150,N_6647);
and U14626 (N_14626,N_7799,N_7868);
and U14627 (N_14627,N_9875,N_8518);
nand U14628 (N_14628,N_5472,N_7315);
and U14629 (N_14629,N_9722,N_6872);
xnor U14630 (N_14630,N_5865,N_5065);
xor U14631 (N_14631,N_9488,N_7387);
or U14632 (N_14632,N_9010,N_5949);
and U14633 (N_14633,N_5645,N_5104);
and U14634 (N_14634,N_7974,N_5214);
or U14635 (N_14635,N_9729,N_9740);
nand U14636 (N_14636,N_8808,N_9390);
or U14637 (N_14637,N_7030,N_7553);
nand U14638 (N_14638,N_6678,N_6417);
nor U14639 (N_14639,N_9289,N_8771);
nor U14640 (N_14640,N_9849,N_6586);
xor U14641 (N_14641,N_9991,N_5219);
and U14642 (N_14642,N_5552,N_7782);
or U14643 (N_14643,N_9324,N_9686);
xnor U14644 (N_14644,N_9830,N_9834);
or U14645 (N_14645,N_9922,N_6331);
xor U14646 (N_14646,N_9900,N_8637);
xor U14647 (N_14647,N_6681,N_9202);
xor U14648 (N_14648,N_6759,N_6126);
and U14649 (N_14649,N_7300,N_9133);
or U14650 (N_14650,N_6178,N_8416);
nor U14651 (N_14651,N_5446,N_6218);
and U14652 (N_14652,N_8748,N_5825);
and U14653 (N_14653,N_9148,N_8109);
or U14654 (N_14654,N_7717,N_7512);
nor U14655 (N_14655,N_5274,N_6806);
or U14656 (N_14656,N_5723,N_6476);
nor U14657 (N_14657,N_8184,N_6245);
nand U14658 (N_14658,N_7741,N_8135);
nor U14659 (N_14659,N_7430,N_9388);
xnor U14660 (N_14660,N_5694,N_5676);
xor U14661 (N_14661,N_9528,N_6788);
and U14662 (N_14662,N_6975,N_5924);
or U14663 (N_14663,N_5940,N_7376);
xor U14664 (N_14664,N_7469,N_6401);
xnor U14665 (N_14665,N_7733,N_7204);
xnor U14666 (N_14666,N_7537,N_8945);
or U14667 (N_14667,N_9029,N_6245);
and U14668 (N_14668,N_6574,N_5343);
nand U14669 (N_14669,N_8850,N_8626);
xor U14670 (N_14670,N_7505,N_9972);
and U14671 (N_14671,N_8955,N_9027);
nor U14672 (N_14672,N_5530,N_9966);
or U14673 (N_14673,N_7122,N_9719);
or U14674 (N_14674,N_7920,N_9952);
or U14675 (N_14675,N_7325,N_6281);
nand U14676 (N_14676,N_6295,N_6524);
and U14677 (N_14677,N_6189,N_7026);
or U14678 (N_14678,N_5397,N_6058);
xor U14679 (N_14679,N_7221,N_8434);
nand U14680 (N_14680,N_6149,N_5803);
or U14681 (N_14681,N_7584,N_5266);
nand U14682 (N_14682,N_6529,N_6660);
and U14683 (N_14683,N_5261,N_5184);
and U14684 (N_14684,N_6752,N_7705);
or U14685 (N_14685,N_6428,N_7396);
nand U14686 (N_14686,N_5092,N_5450);
or U14687 (N_14687,N_7340,N_6943);
nor U14688 (N_14688,N_8789,N_9875);
nor U14689 (N_14689,N_7765,N_5295);
xnor U14690 (N_14690,N_8238,N_6502);
or U14691 (N_14691,N_7359,N_9987);
nand U14692 (N_14692,N_8583,N_7710);
nand U14693 (N_14693,N_9299,N_5708);
and U14694 (N_14694,N_6745,N_7231);
or U14695 (N_14695,N_9263,N_5239);
and U14696 (N_14696,N_5129,N_5652);
nor U14697 (N_14697,N_9263,N_8213);
and U14698 (N_14698,N_5558,N_8190);
nor U14699 (N_14699,N_5008,N_8784);
nor U14700 (N_14700,N_9890,N_7035);
nor U14701 (N_14701,N_6686,N_7563);
or U14702 (N_14702,N_7025,N_6940);
nor U14703 (N_14703,N_8058,N_9373);
and U14704 (N_14704,N_8097,N_7613);
nand U14705 (N_14705,N_5045,N_8305);
nand U14706 (N_14706,N_9584,N_7191);
xnor U14707 (N_14707,N_8042,N_8505);
xor U14708 (N_14708,N_5577,N_7084);
or U14709 (N_14709,N_7106,N_8907);
xor U14710 (N_14710,N_7818,N_8675);
nor U14711 (N_14711,N_5793,N_5267);
nand U14712 (N_14712,N_9688,N_5842);
and U14713 (N_14713,N_7661,N_9079);
and U14714 (N_14714,N_9770,N_5076);
or U14715 (N_14715,N_8776,N_6934);
or U14716 (N_14716,N_8391,N_6435);
and U14717 (N_14717,N_9665,N_6988);
nor U14718 (N_14718,N_5951,N_7463);
xor U14719 (N_14719,N_7151,N_5786);
and U14720 (N_14720,N_8197,N_8632);
and U14721 (N_14721,N_9111,N_5331);
nor U14722 (N_14722,N_7606,N_8853);
or U14723 (N_14723,N_9589,N_5184);
and U14724 (N_14724,N_6794,N_7740);
nor U14725 (N_14725,N_6306,N_5290);
nor U14726 (N_14726,N_5758,N_6979);
nor U14727 (N_14727,N_7416,N_6111);
nor U14728 (N_14728,N_8302,N_8391);
nand U14729 (N_14729,N_9828,N_8918);
xnor U14730 (N_14730,N_9775,N_7939);
and U14731 (N_14731,N_7761,N_7371);
nor U14732 (N_14732,N_5275,N_7764);
nand U14733 (N_14733,N_9335,N_6187);
and U14734 (N_14734,N_9545,N_6033);
or U14735 (N_14735,N_7155,N_8674);
and U14736 (N_14736,N_8933,N_8832);
or U14737 (N_14737,N_8454,N_6524);
and U14738 (N_14738,N_8814,N_7848);
xor U14739 (N_14739,N_9443,N_7962);
and U14740 (N_14740,N_9861,N_9004);
nand U14741 (N_14741,N_5390,N_7347);
or U14742 (N_14742,N_7064,N_6201);
or U14743 (N_14743,N_9533,N_6266);
nand U14744 (N_14744,N_9503,N_5228);
nand U14745 (N_14745,N_5459,N_7865);
xnor U14746 (N_14746,N_7185,N_7846);
or U14747 (N_14747,N_7973,N_6309);
and U14748 (N_14748,N_5238,N_6176);
nor U14749 (N_14749,N_8510,N_6135);
or U14750 (N_14750,N_6312,N_9426);
or U14751 (N_14751,N_6160,N_7941);
nor U14752 (N_14752,N_6508,N_9290);
xor U14753 (N_14753,N_8683,N_7124);
nand U14754 (N_14754,N_7623,N_9302);
and U14755 (N_14755,N_7006,N_9032);
nor U14756 (N_14756,N_9832,N_9868);
and U14757 (N_14757,N_7074,N_7735);
and U14758 (N_14758,N_9268,N_9789);
nor U14759 (N_14759,N_6414,N_6030);
nor U14760 (N_14760,N_8834,N_6945);
and U14761 (N_14761,N_9692,N_9089);
or U14762 (N_14762,N_7839,N_7924);
xor U14763 (N_14763,N_7818,N_7603);
nand U14764 (N_14764,N_9737,N_6388);
xnor U14765 (N_14765,N_6629,N_5738);
nor U14766 (N_14766,N_7301,N_8176);
or U14767 (N_14767,N_9075,N_6009);
and U14768 (N_14768,N_9839,N_7934);
nand U14769 (N_14769,N_6431,N_7736);
or U14770 (N_14770,N_7904,N_6484);
xnor U14771 (N_14771,N_9224,N_5314);
nand U14772 (N_14772,N_7832,N_6894);
or U14773 (N_14773,N_7258,N_5151);
and U14774 (N_14774,N_7031,N_6778);
nor U14775 (N_14775,N_8557,N_8341);
or U14776 (N_14776,N_8122,N_7616);
nand U14777 (N_14777,N_8054,N_9782);
nor U14778 (N_14778,N_8572,N_6409);
nand U14779 (N_14779,N_7922,N_6136);
nor U14780 (N_14780,N_8295,N_9304);
xnor U14781 (N_14781,N_7252,N_6701);
nand U14782 (N_14782,N_6440,N_8244);
and U14783 (N_14783,N_5980,N_5515);
nand U14784 (N_14784,N_8339,N_5107);
xor U14785 (N_14785,N_8937,N_7164);
nand U14786 (N_14786,N_8996,N_5527);
or U14787 (N_14787,N_8455,N_9559);
nor U14788 (N_14788,N_8589,N_5087);
xnor U14789 (N_14789,N_8913,N_7868);
xor U14790 (N_14790,N_5540,N_5066);
xor U14791 (N_14791,N_5783,N_7577);
and U14792 (N_14792,N_5262,N_9743);
xor U14793 (N_14793,N_7125,N_6285);
nor U14794 (N_14794,N_7380,N_8456);
nand U14795 (N_14795,N_5926,N_6705);
nor U14796 (N_14796,N_6563,N_8938);
xor U14797 (N_14797,N_8954,N_9945);
xor U14798 (N_14798,N_9243,N_6864);
nor U14799 (N_14799,N_7857,N_9996);
or U14800 (N_14800,N_7764,N_6867);
and U14801 (N_14801,N_5807,N_9189);
or U14802 (N_14802,N_9649,N_6668);
nand U14803 (N_14803,N_8772,N_6532);
or U14804 (N_14804,N_6620,N_6495);
xnor U14805 (N_14805,N_6949,N_9384);
nand U14806 (N_14806,N_5371,N_5872);
xor U14807 (N_14807,N_9924,N_5790);
xor U14808 (N_14808,N_8385,N_5483);
and U14809 (N_14809,N_8932,N_7182);
nor U14810 (N_14810,N_8719,N_8640);
xnor U14811 (N_14811,N_9370,N_6517);
or U14812 (N_14812,N_9958,N_8762);
and U14813 (N_14813,N_7429,N_6372);
nor U14814 (N_14814,N_6265,N_7931);
nand U14815 (N_14815,N_7212,N_6917);
or U14816 (N_14816,N_9130,N_9161);
nand U14817 (N_14817,N_5541,N_5007);
or U14818 (N_14818,N_7557,N_8124);
nand U14819 (N_14819,N_6262,N_7627);
and U14820 (N_14820,N_8537,N_8554);
xor U14821 (N_14821,N_5616,N_9776);
nor U14822 (N_14822,N_7787,N_7960);
or U14823 (N_14823,N_9725,N_8738);
or U14824 (N_14824,N_8775,N_5258);
xor U14825 (N_14825,N_6740,N_6310);
and U14826 (N_14826,N_9838,N_8325);
nand U14827 (N_14827,N_6702,N_9324);
xor U14828 (N_14828,N_5857,N_7576);
and U14829 (N_14829,N_7329,N_6071);
nor U14830 (N_14830,N_6632,N_5648);
nand U14831 (N_14831,N_9256,N_9455);
or U14832 (N_14832,N_5627,N_9843);
and U14833 (N_14833,N_7296,N_7512);
nand U14834 (N_14834,N_5902,N_8104);
xnor U14835 (N_14835,N_6302,N_6023);
and U14836 (N_14836,N_6326,N_9171);
and U14837 (N_14837,N_5247,N_8720);
or U14838 (N_14838,N_6567,N_5112);
nand U14839 (N_14839,N_6126,N_5625);
and U14840 (N_14840,N_9433,N_9598);
xor U14841 (N_14841,N_9085,N_7659);
or U14842 (N_14842,N_6484,N_8223);
xor U14843 (N_14843,N_6955,N_6214);
nor U14844 (N_14844,N_5078,N_7906);
or U14845 (N_14845,N_6661,N_8706);
xnor U14846 (N_14846,N_8211,N_5525);
or U14847 (N_14847,N_6570,N_8811);
nand U14848 (N_14848,N_5596,N_9535);
nand U14849 (N_14849,N_6429,N_5023);
nor U14850 (N_14850,N_7494,N_9314);
or U14851 (N_14851,N_6231,N_8321);
and U14852 (N_14852,N_5411,N_8383);
or U14853 (N_14853,N_5890,N_6986);
xor U14854 (N_14854,N_6733,N_6925);
xnor U14855 (N_14855,N_7502,N_8623);
xnor U14856 (N_14856,N_8155,N_8300);
nor U14857 (N_14857,N_8750,N_7492);
nor U14858 (N_14858,N_6237,N_7731);
nand U14859 (N_14859,N_7676,N_7486);
xnor U14860 (N_14860,N_5265,N_6618);
or U14861 (N_14861,N_6305,N_9096);
nor U14862 (N_14862,N_7117,N_7423);
xor U14863 (N_14863,N_8266,N_8966);
or U14864 (N_14864,N_8444,N_6516);
or U14865 (N_14865,N_5534,N_8973);
and U14866 (N_14866,N_8196,N_5052);
and U14867 (N_14867,N_5411,N_5338);
or U14868 (N_14868,N_6363,N_7354);
xnor U14869 (N_14869,N_5931,N_5673);
nor U14870 (N_14870,N_9871,N_9540);
or U14871 (N_14871,N_6812,N_9358);
nor U14872 (N_14872,N_6984,N_8991);
xnor U14873 (N_14873,N_9417,N_8653);
xnor U14874 (N_14874,N_9752,N_5099);
or U14875 (N_14875,N_5988,N_8366);
or U14876 (N_14876,N_7742,N_8879);
and U14877 (N_14877,N_6047,N_5864);
nand U14878 (N_14878,N_7014,N_6634);
nor U14879 (N_14879,N_8642,N_5820);
or U14880 (N_14880,N_8823,N_9427);
xor U14881 (N_14881,N_8338,N_9213);
xnor U14882 (N_14882,N_8960,N_9306);
and U14883 (N_14883,N_9092,N_7559);
nor U14884 (N_14884,N_6477,N_8401);
and U14885 (N_14885,N_9385,N_7982);
nand U14886 (N_14886,N_5221,N_5789);
xor U14887 (N_14887,N_9852,N_8336);
and U14888 (N_14888,N_8904,N_5056);
and U14889 (N_14889,N_7274,N_5285);
nor U14890 (N_14890,N_7068,N_7465);
nor U14891 (N_14891,N_5329,N_8410);
and U14892 (N_14892,N_9745,N_7111);
xor U14893 (N_14893,N_8224,N_8242);
nor U14894 (N_14894,N_9334,N_6032);
xnor U14895 (N_14895,N_6711,N_5907);
nor U14896 (N_14896,N_8355,N_8027);
and U14897 (N_14897,N_7162,N_9245);
nand U14898 (N_14898,N_9521,N_5640);
or U14899 (N_14899,N_9525,N_9428);
xor U14900 (N_14900,N_5156,N_5966);
nand U14901 (N_14901,N_9417,N_8428);
nand U14902 (N_14902,N_8134,N_7902);
nor U14903 (N_14903,N_7419,N_8722);
nand U14904 (N_14904,N_7731,N_5117);
xnor U14905 (N_14905,N_9442,N_9878);
and U14906 (N_14906,N_7139,N_7458);
and U14907 (N_14907,N_6466,N_6426);
nor U14908 (N_14908,N_7682,N_5340);
xor U14909 (N_14909,N_5103,N_6301);
and U14910 (N_14910,N_9140,N_9220);
and U14911 (N_14911,N_7469,N_6479);
nor U14912 (N_14912,N_9500,N_9667);
or U14913 (N_14913,N_9130,N_6757);
xor U14914 (N_14914,N_8625,N_8804);
and U14915 (N_14915,N_5514,N_8498);
xor U14916 (N_14916,N_6353,N_9694);
nand U14917 (N_14917,N_9582,N_9282);
nor U14918 (N_14918,N_7006,N_5914);
and U14919 (N_14919,N_7747,N_8559);
or U14920 (N_14920,N_6446,N_8929);
nor U14921 (N_14921,N_9779,N_7429);
nand U14922 (N_14922,N_8849,N_8670);
nand U14923 (N_14923,N_8409,N_6339);
or U14924 (N_14924,N_5551,N_8388);
nor U14925 (N_14925,N_7624,N_7838);
or U14926 (N_14926,N_7576,N_9672);
nor U14927 (N_14927,N_5200,N_6857);
nand U14928 (N_14928,N_5167,N_6435);
nand U14929 (N_14929,N_8216,N_8403);
nand U14930 (N_14930,N_9784,N_9643);
nor U14931 (N_14931,N_8673,N_6643);
or U14932 (N_14932,N_7505,N_5951);
and U14933 (N_14933,N_7561,N_8989);
and U14934 (N_14934,N_5303,N_5007);
or U14935 (N_14935,N_6611,N_9288);
and U14936 (N_14936,N_8768,N_5868);
or U14937 (N_14937,N_6030,N_6241);
nor U14938 (N_14938,N_5451,N_9844);
nor U14939 (N_14939,N_7364,N_8745);
xor U14940 (N_14940,N_9256,N_7587);
nor U14941 (N_14941,N_5399,N_9606);
or U14942 (N_14942,N_6813,N_6379);
or U14943 (N_14943,N_6176,N_9447);
or U14944 (N_14944,N_7450,N_6677);
or U14945 (N_14945,N_8180,N_9136);
and U14946 (N_14946,N_7737,N_9261);
or U14947 (N_14947,N_5417,N_5581);
nor U14948 (N_14948,N_6628,N_9002);
and U14949 (N_14949,N_9158,N_9573);
xnor U14950 (N_14950,N_8701,N_7746);
or U14951 (N_14951,N_6895,N_5595);
or U14952 (N_14952,N_5549,N_8806);
or U14953 (N_14953,N_9412,N_6526);
nor U14954 (N_14954,N_6007,N_8043);
and U14955 (N_14955,N_7009,N_5607);
nor U14956 (N_14956,N_5970,N_6334);
and U14957 (N_14957,N_8465,N_8291);
and U14958 (N_14958,N_8499,N_7492);
nor U14959 (N_14959,N_8134,N_7453);
and U14960 (N_14960,N_9097,N_9013);
nor U14961 (N_14961,N_7082,N_6361);
nor U14962 (N_14962,N_6702,N_6274);
nand U14963 (N_14963,N_8243,N_9575);
nand U14964 (N_14964,N_7601,N_9100);
nand U14965 (N_14965,N_9747,N_5166);
xnor U14966 (N_14966,N_7433,N_6417);
xnor U14967 (N_14967,N_7803,N_7068);
xnor U14968 (N_14968,N_5663,N_9137);
nand U14969 (N_14969,N_9981,N_9417);
or U14970 (N_14970,N_7887,N_8003);
or U14971 (N_14971,N_6487,N_9608);
nor U14972 (N_14972,N_8428,N_7864);
and U14973 (N_14973,N_6835,N_7209);
or U14974 (N_14974,N_7914,N_9899);
or U14975 (N_14975,N_7770,N_9702);
xor U14976 (N_14976,N_6769,N_6142);
nor U14977 (N_14977,N_7003,N_5494);
or U14978 (N_14978,N_6639,N_6537);
nor U14979 (N_14979,N_8898,N_7322);
nor U14980 (N_14980,N_7787,N_8444);
xnor U14981 (N_14981,N_5364,N_9582);
xnor U14982 (N_14982,N_7799,N_8346);
and U14983 (N_14983,N_9453,N_9353);
nor U14984 (N_14984,N_5283,N_6126);
xnor U14985 (N_14985,N_5599,N_6613);
and U14986 (N_14986,N_7651,N_8079);
xor U14987 (N_14987,N_9518,N_6194);
or U14988 (N_14988,N_8812,N_8033);
or U14989 (N_14989,N_7419,N_5469);
and U14990 (N_14990,N_8663,N_9547);
nand U14991 (N_14991,N_6307,N_6640);
or U14992 (N_14992,N_8179,N_5297);
nand U14993 (N_14993,N_8590,N_6866);
nand U14994 (N_14994,N_6699,N_9849);
or U14995 (N_14995,N_7872,N_9071);
or U14996 (N_14996,N_5901,N_7324);
or U14997 (N_14997,N_8820,N_7353);
nor U14998 (N_14998,N_6361,N_5257);
and U14999 (N_14999,N_9051,N_7104);
nor UO_0 (O_0,N_13913,N_14931);
xor UO_1 (O_1,N_10814,N_13678);
and UO_2 (O_2,N_10732,N_10036);
nor UO_3 (O_3,N_12629,N_10920);
nand UO_4 (O_4,N_14276,N_14257);
nand UO_5 (O_5,N_13623,N_11337);
or UO_6 (O_6,N_14070,N_10476);
and UO_7 (O_7,N_10287,N_12017);
xnor UO_8 (O_8,N_12053,N_11668);
and UO_9 (O_9,N_12148,N_14682);
xnor UO_10 (O_10,N_10808,N_12465);
nor UO_11 (O_11,N_12990,N_14845);
xor UO_12 (O_12,N_11299,N_14964);
nand UO_13 (O_13,N_11913,N_14130);
xor UO_14 (O_14,N_12807,N_14537);
xor UO_15 (O_15,N_10396,N_14983);
and UO_16 (O_16,N_10751,N_14227);
nand UO_17 (O_17,N_14837,N_14427);
or UO_18 (O_18,N_10576,N_10000);
and UO_19 (O_19,N_13332,N_14401);
nand UO_20 (O_20,N_10674,N_12342);
or UO_21 (O_21,N_11980,N_10900);
xnor UO_22 (O_22,N_12490,N_14881);
and UO_23 (O_23,N_12652,N_12212);
nor UO_24 (O_24,N_11765,N_14029);
nor UO_25 (O_25,N_13590,N_13447);
nor UO_26 (O_26,N_10663,N_11308);
and UO_27 (O_27,N_13306,N_13656);
nor UO_28 (O_28,N_10182,N_12753);
or UO_29 (O_29,N_11602,N_13734);
nor UO_30 (O_30,N_14763,N_14455);
xnor UO_31 (O_31,N_13503,N_14065);
and UO_32 (O_32,N_14638,N_14811);
and UO_33 (O_33,N_13709,N_12472);
nand UO_34 (O_34,N_12969,N_13414);
and UO_35 (O_35,N_11554,N_13452);
nand UO_36 (O_36,N_12256,N_10088);
nor UO_37 (O_37,N_14096,N_13801);
and UO_38 (O_38,N_10274,N_12929);
nor UO_39 (O_39,N_12254,N_12089);
and UO_40 (O_40,N_11423,N_11859);
xor UO_41 (O_41,N_11739,N_14431);
nor UO_42 (O_42,N_10778,N_13796);
nand UO_43 (O_43,N_14386,N_12247);
nor UO_44 (O_44,N_12500,N_11475);
or UO_45 (O_45,N_13339,N_11039);
nand UO_46 (O_46,N_13952,N_13568);
or UO_47 (O_47,N_11797,N_12427);
nor UO_48 (O_48,N_10312,N_12888);
nand UO_49 (O_49,N_13640,N_12641);
nand UO_50 (O_50,N_11855,N_13108);
or UO_51 (O_51,N_11688,N_12917);
and UO_52 (O_52,N_10589,N_13934);
xor UO_53 (O_53,N_14511,N_14879);
xor UO_54 (O_54,N_14712,N_11922);
xnor UO_55 (O_55,N_12746,N_13340);
xor UO_56 (O_56,N_13591,N_10745);
nand UO_57 (O_57,N_10143,N_13750);
xnor UO_58 (O_58,N_13685,N_13384);
xor UO_59 (O_59,N_13944,N_11832);
nand UO_60 (O_60,N_11249,N_11182);
nand UO_61 (O_61,N_12931,N_11111);
and UO_62 (O_62,N_10275,N_13786);
and UO_63 (O_63,N_13860,N_10819);
nand UO_64 (O_64,N_13410,N_14397);
or UO_65 (O_65,N_14760,N_13136);
xor UO_66 (O_66,N_11824,N_12161);
xor UO_67 (O_67,N_11338,N_13105);
nand UO_68 (O_68,N_12671,N_11802);
nand UO_69 (O_69,N_13090,N_13784);
xor UO_70 (O_70,N_13900,N_10615);
nand UO_71 (O_71,N_14373,N_10480);
or UO_72 (O_72,N_12369,N_12850);
nand UO_73 (O_73,N_10262,N_10716);
xor UO_74 (O_74,N_12589,N_14339);
nor UO_75 (O_75,N_10942,N_11643);
or UO_76 (O_76,N_13998,N_12559);
nor UO_77 (O_77,N_14060,N_13547);
nor UO_78 (O_78,N_14578,N_10191);
nand UO_79 (O_79,N_14774,N_14010);
xor UO_80 (O_80,N_12496,N_11636);
or UO_81 (O_81,N_12631,N_13157);
and UO_82 (O_82,N_13299,N_13641);
nand UO_83 (O_83,N_12595,N_12441);
or UO_84 (O_84,N_12993,N_10153);
or UO_85 (O_85,N_12285,N_14362);
nand UO_86 (O_86,N_13084,N_12003);
or UO_87 (O_87,N_13872,N_14254);
nand UO_88 (O_88,N_13807,N_12337);
nand UO_89 (O_89,N_13488,N_13033);
or UO_90 (O_90,N_10201,N_12123);
nand UO_91 (O_91,N_10181,N_14176);
xor UO_92 (O_92,N_12389,N_11473);
or UO_93 (O_93,N_13195,N_13395);
or UO_94 (O_94,N_10828,N_11310);
or UO_95 (O_95,N_11831,N_12109);
nand UO_96 (O_96,N_13767,N_14572);
nor UO_97 (O_97,N_13513,N_14945);
and UO_98 (O_98,N_10498,N_10352);
nand UO_99 (O_99,N_13617,N_13983);
xor UO_100 (O_100,N_11053,N_10199);
xnor UO_101 (O_101,N_14909,N_11549);
xor UO_102 (O_102,N_13230,N_13476);
and UO_103 (O_103,N_14253,N_11270);
and UO_104 (O_104,N_12101,N_14219);
xor UO_105 (O_105,N_14528,N_11428);
nor UO_106 (O_106,N_13828,N_11984);
nor UO_107 (O_107,N_10838,N_14777);
nor UO_108 (O_108,N_14803,N_14988);
and UO_109 (O_109,N_13560,N_12902);
nor UO_110 (O_110,N_11751,N_14531);
and UO_111 (O_111,N_14884,N_11864);
nand UO_112 (O_112,N_10404,N_12755);
xor UO_113 (O_113,N_14678,N_12223);
or UO_114 (O_114,N_10180,N_10975);
nand UO_115 (O_115,N_11497,N_14066);
and UO_116 (O_116,N_14943,N_13017);
nor UO_117 (O_117,N_14753,N_14894);
nand UO_118 (O_118,N_12258,N_11481);
nand UO_119 (O_119,N_12548,N_14178);
or UO_120 (O_120,N_11564,N_11525);
nor UO_121 (O_121,N_11761,N_14140);
nand UO_122 (O_122,N_12105,N_13267);
nor UO_123 (O_123,N_12230,N_12196);
or UO_124 (O_124,N_11145,N_11102);
xnor UO_125 (O_125,N_11694,N_11231);
or UO_126 (O_126,N_13619,N_13464);
nand UO_127 (O_127,N_13958,N_12047);
nor UO_128 (O_128,N_12396,N_14004);
nor UO_129 (O_129,N_12848,N_10956);
nand UO_130 (O_130,N_14888,N_11457);
and UO_131 (O_131,N_12371,N_14598);
nor UO_132 (O_132,N_13394,N_14392);
nand UO_133 (O_133,N_13917,N_13927);
xnor UO_134 (O_134,N_10534,N_11384);
nand UO_135 (O_135,N_10881,N_14039);
nor UO_136 (O_136,N_10815,N_10358);
and UO_137 (O_137,N_10512,N_14037);
and UO_138 (O_138,N_12795,N_12423);
nor UO_139 (O_139,N_10760,N_10782);
xnor UO_140 (O_140,N_14105,N_10200);
nand UO_141 (O_141,N_12562,N_13542);
and UO_142 (O_142,N_10679,N_12949);
and UO_143 (O_143,N_11031,N_11301);
nor UO_144 (O_144,N_11520,N_13960);
and UO_145 (O_145,N_13215,N_14053);
nand UO_146 (O_146,N_10629,N_12493);
nand UO_147 (O_147,N_13126,N_12645);
and UO_148 (O_148,N_12892,N_10423);
nor UO_149 (O_149,N_14525,N_10853);
xnor UO_150 (O_150,N_13080,N_12853);
xor UO_151 (O_151,N_10223,N_14833);
nor UO_152 (O_152,N_13803,N_10151);
nand UO_153 (O_153,N_13889,N_13779);
nor UO_154 (O_154,N_12772,N_14300);
nor UO_155 (O_155,N_12740,N_10090);
nor UO_156 (O_156,N_12665,N_14443);
xor UO_157 (O_157,N_10177,N_11376);
and UO_158 (O_158,N_13581,N_10770);
xor UO_159 (O_159,N_13248,N_12222);
nand UO_160 (O_160,N_10327,N_13101);
nor UO_161 (O_161,N_12666,N_13558);
nor UO_162 (O_162,N_12514,N_13642);
or UO_163 (O_163,N_14027,N_13325);
and UO_164 (O_164,N_10192,N_12452);
nor UO_165 (O_165,N_10696,N_13873);
nand UO_166 (O_166,N_13615,N_11028);
or UO_167 (O_167,N_12617,N_13219);
nor UO_168 (O_168,N_12082,N_14900);
or UO_169 (O_169,N_10039,N_14034);
xor UO_170 (O_170,N_12055,N_11247);
xnor UO_171 (O_171,N_14666,N_13774);
nand UO_172 (O_172,N_13695,N_11996);
nor UO_173 (O_173,N_11854,N_11025);
xor UO_174 (O_174,N_11395,N_13100);
nor UO_175 (O_175,N_14069,N_10718);
xor UO_176 (O_176,N_11970,N_13578);
xor UO_177 (O_177,N_10162,N_13139);
nand UO_178 (O_178,N_13841,N_11902);
nand UO_179 (O_179,N_14372,N_11628);
xor UO_180 (O_180,N_11402,N_11411);
or UO_181 (O_181,N_12482,N_11330);
or UO_182 (O_182,N_12074,N_11657);
and UO_183 (O_183,N_14938,N_12612);
xor UO_184 (O_184,N_10218,N_14051);
nand UO_185 (O_185,N_12728,N_10744);
nand UO_186 (O_186,N_12533,N_12937);
xor UO_187 (O_187,N_12150,N_13565);
nand UO_188 (O_188,N_13022,N_10329);
and UO_189 (O_189,N_14168,N_14293);
and UO_190 (O_190,N_13652,N_10284);
nor UO_191 (O_191,N_14395,N_12213);
nor UO_192 (O_192,N_12777,N_12171);
and UO_193 (O_193,N_11105,N_10582);
and UO_194 (O_194,N_12682,N_10767);
nor UO_195 (O_195,N_11256,N_12635);
xor UO_196 (O_196,N_10935,N_10306);
and UO_197 (O_197,N_13111,N_14658);
xor UO_198 (O_198,N_10373,N_14814);
xnor UO_199 (O_199,N_13583,N_14901);
and UO_200 (O_200,N_12163,N_14167);
and UO_201 (O_201,N_10707,N_12973);
or UO_202 (O_202,N_13275,N_13448);
and UO_203 (O_203,N_14442,N_13599);
xnor UO_204 (O_204,N_10713,N_11511);
xnor UO_205 (O_205,N_11393,N_11945);
nand UO_206 (O_206,N_14655,N_11676);
nor UO_207 (O_207,N_14458,N_14017);
nand UO_208 (O_208,N_13835,N_11168);
nand UO_209 (O_209,N_11509,N_14152);
or UO_210 (O_210,N_10443,N_10933);
nor UO_211 (O_211,N_14137,N_11581);
and UO_212 (O_212,N_13320,N_13506);
nand UO_213 (O_213,N_12729,N_10810);
and UO_214 (O_214,N_10469,N_10461);
nor UO_215 (O_215,N_13659,N_11314);
and UO_216 (O_216,N_12063,N_14277);
nand UO_217 (O_217,N_11313,N_14011);
and UO_218 (O_218,N_12873,N_12450);
and UO_219 (O_219,N_14118,N_12042);
nor UO_220 (O_220,N_14143,N_11507);
or UO_221 (O_221,N_12275,N_11071);
nand UO_222 (O_222,N_14716,N_14805);
nand UO_223 (O_223,N_12556,N_11758);
and UO_224 (O_224,N_14692,N_10585);
nor UO_225 (O_225,N_10765,N_10890);
or UO_226 (O_226,N_10290,N_13785);
nor UO_227 (O_227,N_13886,N_14074);
xnor UO_228 (O_228,N_11164,N_10502);
nand UO_229 (O_229,N_13305,N_11563);
nand UO_230 (O_230,N_13456,N_11504);
xnor UO_231 (O_231,N_13871,N_14503);
nand UO_232 (O_232,N_11038,N_13301);
or UO_233 (O_233,N_11926,N_14788);
and UO_234 (O_234,N_12032,N_14998);
xor UO_235 (O_235,N_10166,N_10539);
or UO_236 (O_236,N_14327,N_13517);
and UO_237 (O_237,N_14388,N_10069);
or UO_238 (O_238,N_13415,N_12779);
or UO_239 (O_239,N_13224,N_10103);
and UO_240 (O_240,N_13666,N_10425);
and UO_241 (O_241,N_12207,N_13711);
nor UO_242 (O_242,N_11325,N_11479);
nand UO_243 (O_243,N_14807,N_10195);
nand UO_244 (O_244,N_12741,N_14083);
and UO_245 (O_245,N_11538,N_14106);
xnor UO_246 (O_246,N_14061,N_13021);
or UO_247 (O_247,N_12430,N_14331);
nand UO_248 (O_248,N_12355,N_12374);
nand UO_249 (O_249,N_11024,N_14723);
and UO_250 (O_250,N_13367,N_14131);
nand UO_251 (O_251,N_14918,N_11919);
and UO_252 (O_252,N_12153,N_10472);
xor UO_253 (O_253,N_12431,N_12698);
xnor UO_254 (O_254,N_13397,N_13259);
and UO_255 (O_255,N_11262,N_10785);
or UO_256 (O_256,N_14098,N_14342);
nor UO_257 (O_257,N_11850,N_11904);
or UO_258 (O_258,N_14101,N_14247);
nor UO_259 (O_259,N_13526,N_14145);
nor UO_260 (O_260,N_11652,N_12471);
nor UO_261 (O_261,N_13516,N_11813);
and UO_262 (O_262,N_10059,N_11326);
xor UO_263 (O_263,N_11655,N_14432);
or UO_264 (O_264,N_12236,N_12013);
or UO_265 (O_265,N_12844,N_11702);
xor UO_266 (O_266,N_12051,N_13840);
xnor UO_267 (O_267,N_11344,N_14942);
nor UO_268 (O_268,N_11928,N_13811);
nand UO_269 (O_269,N_13481,N_11429);
nand UO_270 (O_270,N_10105,N_14564);
nor UO_271 (O_271,N_10918,N_14206);
xnor UO_272 (O_272,N_10726,N_10431);
or UO_273 (O_273,N_12766,N_10735);
nand UO_274 (O_274,N_11414,N_10865);
or UO_275 (O_275,N_12154,N_12476);
and UO_276 (O_276,N_13266,N_14163);
xnor UO_277 (O_277,N_14025,N_10981);
and UO_278 (O_278,N_14225,N_11772);
nor UO_279 (O_279,N_11448,N_10660);
or UO_280 (O_280,N_10030,N_10394);
or UO_281 (O_281,N_13610,N_12276);
xnor UO_282 (O_282,N_13477,N_13016);
xor UO_283 (O_283,N_10145,N_11513);
or UO_284 (O_284,N_12404,N_11756);
and UO_285 (O_285,N_13005,N_13915);
xor UO_286 (O_286,N_13881,N_13999);
and UO_287 (O_287,N_11020,N_13713);
and UO_288 (O_288,N_13975,N_11838);
nor UO_289 (O_289,N_11352,N_12749);
xor UO_290 (O_290,N_10254,N_14369);
nand UO_291 (O_291,N_11673,N_14050);
nor UO_292 (O_292,N_12650,N_12913);
nor UO_293 (O_293,N_14809,N_13928);
nand UO_294 (O_294,N_13588,N_13650);
xor UO_295 (O_295,N_10349,N_12605);
nor UO_296 (O_296,N_13967,N_14992);
nand UO_297 (O_297,N_11472,N_13984);
xnor UO_298 (O_298,N_14660,N_12478);
xor UO_299 (O_299,N_12859,N_11350);
xnor UO_300 (O_300,N_10973,N_13552);
nand UO_301 (O_301,N_11542,N_14530);
nand UO_302 (O_302,N_14195,N_10376);
or UO_303 (O_303,N_10296,N_11154);
nand UO_304 (O_304,N_10687,N_12056);
or UO_305 (O_305,N_12819,N_11196);
xor UO_306 (O_306,N_14209,N_11742);
nand UO_307 (O_307,N_10673,N_12667);
and UO_308 (O_308,N_10340,N_12068);
xnor UO_309 (O_309,N_13616,N_11016);
nand UO_310 (O_310,N_11749,N_11903);
or UO_311 (O_311,N_10821,N_14473);
nor UO_312 (O_312,N_13777,N_10100);
or UO_313 (O_313,N_14343,N_10113);
and UO_314 (O_314,N_10164,N_10882);
or UO_315 (O_315,N_12370,N_11822);
and UO_316 (O_316,N_14450,N_10783);
nor UO_317 (O_317,N_11620,N_11740);
and UO_318 (O_318,N_10816,N_12965);
nor UO_319 (O_319,N_13327,N_10407);
xor UO_320 (O_320,N_12540,N_13269);
xnor UO_321 (O_321,N_13728,N_14370);
nor UO_322 (O_322,N_12985,N_14380);
xor UO_323 (O_323,N_13164,N_12709);
nor UO_324 (O_324,N_10840,N_10096);
nand UO_325 (O_325,N_10347,N_10831);
and UO_326 (O_326,N_10864,N_10174);
nor UO_327 (O_327,N_11773,N_14711);
or UO_328 (O_328,N_10773,N_14645);
and UO_329 (O_329,N_13632,N_10027);
xnor UO_330 (O_330,N_11239,N_13374);
nor UO_331 (O_331,N_12599,N_11748);
nor UO_332 (O_332,N_10946,N_13968);
or UO_333 (O_333,N_14498,N_10302);
nor UO_334 (O_334,N_11887,N_10388);
xnor UO_335 (O_335,N_13400,N_12662);
or UO_336 (O_336,N_10965,N_12241);
and UO_337 (O_337,N_14434,N_13523);
xnor UO_338 (O_338,N_12194,N_10074);
nand UO_339 (O_339,N_12865,N_14196);
xor UO_340 (O_340,N_14231,N_12498);
and UO_341 (O_341,N_11604,N_10487);
and UO_342 (O_342,N_14835,N_11345);
xnor UO_343 (O_343,N_12994,N_12321);
xnor UO_344 (O_344,N_10859,N_11993);
or UO_345 (O_345,N_14566,N_10658);
and UO_346 (O_346,N_10695,N_12198);
nor UO_347 (O_347,N_13323,N_14595);
and UO_348 (O_348,N_10325,N_10102);
nand UO_349 (O_349,N_12925,N_13858);
or UO_350 (O_350,N_13726,N_10610);
nor UO_351 (O_351,N_13330,N_14844);
and UO_352 (O_352,N_11381,N_12976);
and UO_353 (O_353,N_14007,N_11356);
xnor UO_354 (O_354,N_11536,N_13392);
nor UO_355 (O_355,N_11439,N_12552);
nor UO_356 (O_356,N_14796,N_11910);
nand UO_357 (O_357,N_13502,N_13334);
and UO_358 (O_358,N_14399,N_12255);
xnor UO_359 (O_359,N_13361,N_14691);
xor UO_360 (O_360,N_13183,N_13722);
nand UO_361 (O_361,N_10951,N_12934);
nand UO_362 (O_362,N_12299,N_13196);
nor UO_363 (O_363,N_13031,N_10441);
nand UO_364 (O_364,N_13708,N_11340);
and UO_365 (O_365,N_13187,N_13972);
or UO_366 (O_366,N_11149,N_10276);
xnor UO_367 (O_367,N_12348,N_12084);
or UO_368 (O_368,N_12422,N_10852);
xnor UO_369 (O_369,N_11323,N_12601);
and UO_370 (O_370,N_11933,N_14628);
and UO_371 (O_371,N_11543,N_11784);
nor UO_372 (O_372,N_11498,N_14023);
and UO_373 (O_373,N_10639,N_10072);
nand UO_374 (O_374,N_11449,N_12884);
nand UO_375 (O_375,N_13935,N_12845);
and UO_376 (O_376,N_11659,N_11043);
or UO_377 (O_377,N_13351,N_11026);
and UO_378 (O_378,N_12200,N_12497);
nor UO_379 (O_379,N_13814,N_11807);
or UO_380 (O_380,N_12083,N_13413);
nand UO_381 (O_381,N_14393,N_10006);
and UO_382 (O_382,N_12336,N_13707);
or UO_383 (O_383,N_12095,N_11261);
and UO_384 (O_384,N_13119,N_10304);
nand UO_385 (O_385,N_14776,N_14138);
xnor UO_386 (O_386,N_10125,N_13142);
nor UO_387 (O_387,N_13497,N_11721);
and UO_388 (O_388,N_11021,N_10089);
and UO_389 (O_389,N_11377,N_11221);
xnor UO_390 (O_390,N_14926,N_10281);
and UO_391 (O_391,N_12111,N_14786);
nor UO_392 (O_392,N_12693,N_12188);
and UO_393 (O_393,N_10099,N_12346);
xnor UO_394 (O_394,N_14221,N_11422);
nor UO_395 (O_395,N_13754,N_14794);
and UO_396 (O_396,N_14089,N_14937);
and UO_397 (O_397,N_12229,N_13049);
and UO_398 (O_398,N_10621,N_11432);
and UO_399 (O_399,N_10507,N_13058);
or UO_400 (O_400,N_11521,N_11117);
nor UO_401 (O_401,N_10501,N_11845);
and UO_402 (O_402,N_14030,N_12376);
nand UO_403 (O_403,N_14516,N_13721);
xnor UO_404 (O_404,N_12757,N_14217);
nand UO_405 (O_405,N_13628,N_14663);
and UO_406 (O_406,N_10455,N_12201);
nor UO_407 (O_407,N_11701,N_13226);
and UO_408 (O_408,N_11973,N_11767);
nor UO_409 (O_409,N_11397,N_11911);
nor UO_410 (O_410,N_10738,N_14895);
xor UO_411 (O_411,N_12778,N_11906);
xor UO_412 (O_412,N_14771,N_11011);
nor UO_413 (O_413,N_14127,N_14991);
nand UO_414 (O_414,N_14383,N_14368);
xor UO_415 (O_415,N_10070,N_11526);
xnor UO_416 (O_416,N_13315,N_11883);
xnor UO_417 (O_417,N_13598,N_12918);
nand UO_418 (O_418,N_11569,N_10987);
nand UO_419 (O_419,N_10129,N_11420);
nand UO_420 (O_420,N_11198,N_14644);
and UO_421 (O_421,N_12209,N_13647);
or UO_422 (O_422,N_12311,N_13776);
nand UO_423 (O_423,N_12900,N_10228);
xnor UO_424 (O_424,N_10283,N_12048);
and UO_425 (O_425,N_12218,N_14191);
and UO_426 (O_426,N_14204,N_10781);
nor UO_427 (O_427,N_11500,N_13437);
xnor UO_428 (O_428,N_14085,N_13895);
nand UO_429 (O_429,N_10688,N_12542);
nand UO_430 (O_430,N_14291,N_14951);
xnor UO_431 (O_431,N_13156,N_14181);
and UO_432 (O_432,N_12412,N_11212);
or UO_433 (O_433,N_11339,N_11800);
and UO_434 (O_434,N_13646,N_13696);
and UO_435 (O_435,N_11760,N_12278);
nand UO_436 (O_436,N_10463,N_12767);
and UO_437 (O_437,N_14561,N_10969);
nand UO_438 (O_438,N_11425,N_13863);
nor UO_439 (O_439,N_11090,N_11588);
xor UO_440 (O_440,N_10769,N_13203);
or UO_441 (O_441,N_10733,N_13252);
nand UO_442 (O_442,N_13788,N_10126);
or UO_443 (O_443,N_12491,N_14724);
xnor UO_444 (O_444,N_11645,N_10652);
or UO_445 (O_445,N_13633,N_10389);
or UO_446 (O_446,N_10637,N_13760);
or UO_447 (O_447,N_10953,N_14235);
nor UO_448 (O_448,N_12265,N_14569);
and UO_449 (O_449,N_14797,N_13727);
nand UO_450 (O_450,N_14579,N_13044);
or UO_451 (O_451,N_10702,N_14026);
and UO_452 (O_452,N_11770,N_11811);
nand UO_453 (O_453,N_10884,N_13894);
and UO_454 (O_454,N_12103,N_12119);
nor UO_455 (O_455,N_10874,N_10470);
xnor UO_456 (O_456,N_12245,N_13775);
and UO_457 (O_457,N_10545,N_11994);
and UO_458 (O_458,N_13307,N_10677);
xor UO_459 (O_459,N_12801,N_14205);
nor UO_460 (O_460,N_12350,N_14749);
xnor UO_461 (O_461,N_12453,N_10233);
and UO_462 (O_462,N_13579,N_10260);
or UO_463 (O_463,N_10414,N_11036);
xnor UO_464 (O_464,N_12618,N_11950);
nor UO_465 (O_465,N_10635,N_12602);
nor UO_466 (O_466,N_14878,N_13385);
nand UO_467 (O_467,N_13372,N_14433);
nor UO_468 (O_468,N_13071,N_12899);
or UO_469 (O_469,N_11958,N_14553);
and UO_470 (O_470,N_10742,N_12227);
nand UO_471 (O_471,N_13989,N_10966);
nor UO_472 (O_472,N_13849,N_11259);
xor UO_473 (O_473,N_13924,N_10988);
xnor UO_474 (O_474,N_14258,N_12978);
and UO_475 (O_475,N_14479,N_12185);
and UO_476 (O_476,N_10598,N_12027);
nor UO_477 (O_477,N_12489,N_14501);
xor UO_478 (O_478,N_13208,N_14412);
and UO_479 (O_479,N_14850,N_10906);
nor UO_480 (O_480,N_14430,N_13660);
or UO_481 (O_481,N_14604,N_11759);
nor UO_482 (O_482,N_13377,N_11754);
nand UO_483 (O_483,N_12249,N_13303);
or UO_484 (O_484,N_11332,N_14904);
xnor UO_485 (O_485,N_12228,N_10035);
nand UO_486 (O_486,N_11237,N_11115);
or UO_487 (O_487,N_13450,N_14962);
and UO_488 (O_488,N_10997,N_13862);
or UO_489 (O_489,N_12232,N_10509);
xnor UO_490 (O_490,N_13605,N_14325);
or UO_491 (O_491,N_14993,N_14255);
nor UO_492 (O_492,N_13997,N_11921);
and UO_493 (O_493,N_14082,N_11430);
or UO_494 (O_494,N_10259,N_14863);
nand UO_495 (O_495,N_10448,N_14475);
or UO_496 (O_496,N_12705,N_14585);
xor UO_497 (O_497,N_11715,N_12817);
or UO_498 (O_498,N_13236,N_14187);
or UO_499 (O_499,N_12785,N_13684);
and UO_500 (O_500,N_11131,N_12781);
nor UO_501 (O_501,N_11210,N_14701);
and UO_502 (O_502,N_14675,N_10456);
nand UO_503 (O_503,N_11979,N_13519);
nand UO_504 (O_504,N_12016,N_12686);
xor UO_505 (O_505,N_12463,N_10593);
nor UO_506 (O_506,N_13318,N_12761);
or UO_507 (O_507,N_11576,N_13172);
xnor UO_508 (O_508,N_10157,N_10780);
nor UO_509 (O_509,N_14199,N_10646);
or UO_510 (O_510,N_14256,N_11216);
and UO_511 (O_511,N_13087,N_13427);
nand UO_512 (O_512,N_12521,N_13461);
nand UO_513 (O_513,N_13042,N_13585);
nand UO_514 (O_514,N_10493,N_13431);
and UO_515 (O_515,N_12938,N_10542);
xnor UO_516 (O_516,N_14629,N_11317);
xnor UO_517 (O_517,N_13015,N_10665);
and UO_518 (O_518,N_14478,N_10812);
nor UO_519 (O_519,N_12710,N_13887);
xor UO_520 (O_520,N_14982,N_13050);
nand UO_521 (O_521,N_13027,N_12166);
nor UO_522 (O_522,N_13942,N_12950);
and UO_523 (O_523,N_13573,N_10623);
nor UO_524 (O_524,N_11551,N_13757);
nor UO_525 (O_525,N_13748,N_14366);
nand UO_526 (O_526,N_14560,N_11743);
nor UO_527 (O_527,N_13355,N_11665);
nand UO_528 (O_528,N_14073,N_12141);
nand UO_529 (O_529,N_10360,N_10893);
or UO_530 (O_530,N_12157,N_14999);
or UO_531 (O_531,N_12732,N_13322);
nor UO_532 (O_532,N_13296,N_12972);
and UO_533 (O_533,N_11027,N_14289);
nor UO_534 (O_534,N_12863,N_12292);
xnor UO_535 (O_535,N_12683,N_14336);
nor UO_536 (O_536,N_14332,N_12952);
nand UO_537 (O_537,N_13380,N_12847);
nand UO_538 (O_538,N_10402,N_13936);
or UO_539 (O_539,N_12368,N_12060);
nor UO_540 (O_540,N_10588,N_10060);
and UO_541 (O_541,N_14363,N_14446);
nor UO_542 (O_542,N_11019,N_11433);
nor UO_543 (O_543,N_10194,N_12948);
xor UO_544 (O_544,N_11985,N_13036);
and UO_545 (O_545,N_13563,N_14155);
nand UO_546 (O_546,N_13393,N_11794);
xnor UO_547 (O_547,N_14018,N_11172);
or UO_548 (O_548,N_13109,N_14139);
and UO_549 (O_549,N_10761,N_11777);
xnor UO_550 (O_550,N_14480,N_11017);
xor UO_551 (O_551,N_10627,N_10514);
or UO_552 (O_552,N_14402,N_12638);
and UO_553 (O_553,N_14936,N_10938);
xnor UO_554 (O_554,N_13486,N_14650);
or UO_555 (O_555,N_14154,N_14281);
xor UO_556 (O_556,N_13882,N_10154);
nand UO_557 (O_557,N_10451,N_10056);
and UO_558 (O_558,N_11867,N_10179);
and UO_559 (O_559,N_14486,N_13081);
xnor UO_560 (O_560,N_14398,N_13770);
nand UO_561 (O_561,N_11671,N_14463);
or UO_562 (O_562,N_13797,N_12910);
and UO_563 (O_563,N_11342,N_10520);
or UO_564 (O_564,N_13761,N_11218);
and UO_565 (O_565,N_12359,N_13765);
or UO_566 (O_566,N_13831,N_14815);
nand UO_567 (O_567,N_11983,N_12751);
xnor UO_568 (O_568,N_11963,N_10432);
or UO_569 (O_569,N_10731,N_13753);
nor UO_570 (O_570,N_13712,N_14057);
xor UO_571 (O_571,N_12685,N_10672);
and UO_572 (O_572,N_14059,N_12069);
xnor UO_573 (O_573,N_14587,N_11897);
xor UO_574 (O_574,N_10319,N_10709);
and UO_575 (O_575,N_13832,N_14526);
xnor UO_576 (O_576,N_13494,N_14129);
nand UO_577 (O_577,N_13870,N_14957);
and UO_578 (O_578,N_14738,N_12524);
and UO_579 (O_579,N_13546,N_13045);
and UO_580 (O_580,N_13867,N_10772);
or UO_581 (O_581,N_13527,N_12663);
nand UO_582 (O_582,N_10790,N_14622);
and UO_583 (O_583,N_11534,N_10604);
nand UO_584 (O_584,N_11865,N_11382);
and UO_585 (O_585,N_10631,N_11837);
nand UO_586 (O_586,N_12739,N_11437);
nor UO_587 (O_587,N_11503,N_11992);
xnor UO_588 (O_588,N_13823,N_12031);
xnor UO_589 (O_589,N_11491,N_12543);
xnor UO_590 (O_590,N_14976,N_10899);
xor UO_591 (O_591,N_13213,N_13978);
xor UO_592 (O_592,N_12676,N_10570);
and UO_593 (O_593,N_12409,N_14947);
xnor UO_594 (O_594,N_10205,N_14005);
or UO_595 (O_595,N_11987,N_12014);
or UO_596 (O_596,N_10650,N_10108);
and UO_597 (O_597,N_11771,N_10107);
and UO_598 (O_598,N_11846,N_10564);
nor UO_599 (O_599,N_10230,N_12386);
nand UO_600 (O_600,N_14429,N_11092);
nor UO_601 (O_601,N_12217,N_10904);
and UO_602 (O_602,N_11757,N_10298);
xor UO_603 (O_603,N_11692,N_11076);
and UO_604 (O_604,N_10042,N_12515);
nor UO_605 (O_605,N_14899,N_10186);
nor UO_606 (O_606,N_12352,N_14409);
and UO_607 (O_607,N_11646,N_11675);
and UO_608 (O_608,N_14320,N_13041);
xnor UO_609 (O_609,N_12561,N_14707);
and UO_610 (O_610,N_14464,N_11078);
and UO_611 (O_611,N_12623,N_12246);
or UO_612 (O_612,N_13537,N_11143);
nor UO_613 (O_613,N_14064,N_10255);
xor UO_614 (O_614,N_10937,N_11574);
xnor UO_615 (O_615,N_12724,N_10568);
xnor UO_616 (O_616,N_11699,N_14893);
and UO_617 (O_617,N_13890,N_12410);
nor UO_618 (O_618,N_14471,N_14457);
xnor UO_619 (O_619,N_13676,N_13223);
nor UO_620 (O_620,N_12928,N_13509);
xnor UO_621 (O_621,N_13679,N_14111);
xor UO_622 (O_622,N_11949,N_13996);
xnor UO_623 (O_623,N_13602,N_10123);
nand UO_624 (O_624,N_14621,N_14268);
nand UO_625 (O_625,N_14353,N_10983);
or UO_626 (O_626,N_13498,N_14941);
xor UO_627 (O_627,N_14672,N_13724);
nand UO_628 (O_628,N_11208,N_12681);
xnor UO_629 (O_629,N_11009,N_12216);
xor UO_630 (O_630,N_11515,N_12018);
xnor UO_631 (O_631,N_12481,N_10062);
or UO_632 (O_632,N_12791,N_11065);
and UO_633 (O_633,N_14832,N_13151);
nand UO_634 (O_634,N_13480,N_10711);
and UO_635 (O_635,N_12916,N_11140);
xor UO_636 (O_636,N_14646,N_11427);
and UO_637 (O_637,N_10348,N_11637);
nand UO_638 (O_638,N_11683,N_14185);
nand UO_639 (O_639,N_13859,N_14077);
and UO_640 (O_640,N_10040,N_13216);
and UO_641 (O_641,N_11264,N_13557);
and UO_642 (O_642,N_11708,N_12523);
nor UO_643 (O_643,N_14539,N_10714);
and UO_644 (O_644,N_13815,N_14174);
nor UO_645 (O_645,N_11209,N_14159);
nand UO_646 (O_646,N_13120,N_13561);
nor UO_647 (O_647,N_10410,N_12567);
or UO_648 (O_648,N_11141,N_14403);
xor UO_649 (O_649,N_11181,N_14274);
xor UO_650 (O_650,N_11860,N_11627);
nor UO_651 (O_651,N_14698,N_10548);
or UO_652 (O_652,N_12165,N_13950);
or UO_653 (O_653,N_10076,N_12881);
nand UO_654 (O_654,N_10144,N_13116);
or UO_655 (O_655,N_13010,N_13356);
or UO_656 (O_656,N_13816,N_12309);
or UO_657 (O_657,N_14472,N_10892);
nand UO_658 (O_658,N_12722,N_11736);
or UO_659 (O_659,N_14804,N_13199);
nand UO_660 (O_660,N_14170,N_14656);
nand UO_661 (O_661,N_12597,N_10251);
xor UO_662 (O_662,N_12799,N_14272);
or UO_663 (O_663,N_13364,N_13655);
xnor UO_664 (O_664,N_14673,N_10655);
xor UO_665 (O_665,N_14136,N_12982);
nor UO_666 (O_666,N_14889,N_14169);
or UO_667 (O_667,N_14853,N_13148);
nor UO_668 (O_668,N_13663,N_14377);
and UO_669 (O_669,N_14615,N_11953);
xnor UO_670 (O_670,N_12189,N_13851);
nand UO_671 (O_671,N_14492,N_10929);
and UO_672 (O_672,N_14375,N_11306);
nand UO_673 (O_673,N_12981,N_11829);
xnor UO_674 (O_674,N_13034,N_11070);
nor UO_675 (O_675,N_12464,N_13255);
or UO_676 (O_676,N_11403,N_14908);
nand UO_677 (O_677,N_14445,N_14509);
nand UO_678 (O_678,N_11056,N_10691);
nand UO_679 (O_679,N_10943,N_10947);
and UO_680 (O_680,N_14667,N_10178);
nor UO_681 (O_681,N_12224,N_13282);
or UO_682 (O_682,N_11886,N_11785);
or UO_683 (O_683,N_11677,N_10095);
or UO_684 (O_684,N_11912,N_12270);
or UO_685 (O_685,N_10285,N_11798);
nor UO_686 (O_686,N_10131,N_12563);
nand UO_687 (O_687,N_12029,N_11871);
nor UO_688 (O_688,N_10341,N_10384);
xnor UO_689 (O_689,N_10333,N_13543);
xnor UO_690 (O_690,N_14456,N_12252);
or UO_691 (O_691,N_10395,N_12588);
and UO_692 (O_692,N_12445,N_14687);
nand UO_693 (O_693,N_13121,N_10560);
nor UO_694 (O_694,N_13792,N_13706);
nor UO_695 (O_695,N_10478,N_14997);
nand UO_696 (O_696,N_14282,N_12233);
and UO_697 (O_697,N_12137,N_12145);
xor UO_698 (O_698,N_12759,N_11649);
or UO_699 (O_699,N_13802,N_13990);
nand UO_700 (O_700,N_13294,N_10620);
nand UO_701 (O_701,N_12687,N_10662);
nor UO_702 (O_702,N_11790,N_10948);
and UO_703 (O_703,N_12039,N_12187);
and UO_704 (O_704,N_13499,N_12673);
xnor UO_705 (O_705,N_14086,N_13645);
nor UO_706 (O_706,N_12357,N_14875);
or UO_707 (O_707,N_11002,N_13342);
nor UO_708 (O_708,N_13154,N_12387);
xor UO_709 (O_709,N_11492,N_12182);
nor UO_710 (O_710,N_10720,N_14474);
nand UO_711 (O_711,N_14189,N_11579);
nand UO_712 (O_712,N_14499,N_12933);
and UO_713 (O_713,N_12360,N_12958);
nor UO_714 (O_714,N_13988,N_11848);
nor UO_715 (O_715,N_13359,N_14260);
xnor UO_716 (O_716,N_14848,N_12438);
xnor UO_717 (O_717,N_11585,N_10823);
nor UO_718 (O_718,N_11891,N_14347);
xor UO_719 (O_719,N_14680,N_14319);
nand UO_720 (O_720,N_10875,N_10422);
nand UO_721 (O_721,N_11192,N_10656);
and UO_722 (O_722,N_11392,N_13620);
or UO_723 (O_723,N_12298,N_10010);
nand UO_724 (O_724,N_11804,N_11874);
or UO_725 (O_725,N_13308,N_11328);
nand UO_726 (O_726,N_11013,N_12146);
and UO_727 (O_727,N_12090,N_11480);
nor UO_728 (O_728,N_12874,N_13280);
xor UO_729 (O_729,N_13751,N_13495);
and UO_730 (O_730,N_11696,N_10492);
xnor UO_731 (O_731,N_13107,N_12259);
or UO_732 (O_732,N_14785,N_13210);
and UO_733 (O_733,N_14194,N_10499);
xor UO_734 (O_734,N_12956,N_10558);
nor UO_735 (O_735,N_11296,N_10038);
xnor UO_736 (O_736,N_10483,N_13930);
xnor UO_737 (O_737,N_14827,N_10566);
or UO_738 (O_738,N_11488,N_12804);
or UO_739 (O_739,N_14640,N_13540);
xnor UO_740 (O_740,N_10149,N_11647);
nor UO_741 (O_741,N_14183,N_11291);
xor UO_742 (O_742,N_12707,N_11799);
and UO_743 (O_743,N_11123,N_14690);
or UO_744 (O_744,N_10992,N_14969);
nand UO_745 (O_745,N_12486,N_10979);
or UO_746 (O_746,N_14824,N_13250);
or UO_747 (O_747,N_11081,N_13262);
xor UO_748 (O_748,N_11939,N_14965);
xor UO_749 (O_749,N_10541,N_11200);
xor UO_750 (O_750,N_13411,N_11440);
xor UO_751 (O_751,N_12239,N_10699);
nor UO_752 (O_752,N_12637,N_11531);
nand UO_753 (O_753,N_11617,N_13324);
or UO_754 (O_754,N_12058,N_14583);
and UO_755 (O_755,N_12551,N_14766);
and UO_756 (O_756,N_11762,N_11745);
xnor UO_757 (O_757,N_12405,N_10681);
or UO_758 (O_758,N_12536,N_11570);
and UO_759 (O_759,N_12932,N_14406);
nand UO_760 (O_760,N_14165,N_12211);
xnor UO_761 (O_761,N_13854,N_11819);
nor UO_762 (O_762,N_11246,N_14576);
nand UO_763 (O_763,N_10366,N_13904);
xnor UO_764 (O_764,N_11286,N_13812);
nor UO_765 (O_765,N_11827,N_14177);
or UO_766 (O_766,N_10268,N_11889);
nor UO_767 (O_767,N_10097,N_13261);
nand UO_768 (O_768,N_13455,N_14203);
and UO_769 (O_769,N_12625,N_12923);
and UO_770 (O_770,N_11890,N_14795);
nor UO_771 (O_771,N_14197,N_12820);
nor UO_772 (O_772,N_14076,N_13194);
xor UO_773 (O_773,N_12114,N_14784);
and UO_774 (O_774,N_12843,N_12281);
and UO_775 (O_775,N_13980,N_12886);
nor UO_776 (O_776,N_11137,N_10221);
nor UO_777 (O_777,N_13238,N_13662);
xor UO_778 (O_778,N_12962,N_10028);
or UO_779 (O_779,N_14540,N_11577);
or UO_780 (O_780,N_11379,N_11691);
and UO_781 (O_781,N_14313,N_11358);
xnor UO_782 (O_782,N_11737,N_12926);
or UO_783 (O_783,N_11923,N_11290);
xnor UO_784 (O_784,N_13769,N_11641);
nand UO_785 (O_785,N_13956,N_14928);
nor UO_786 (O_786,N_13501,N_12272);
or UO_787 (O_787,N_10762,N_10955);
or UO_788 (O_788,N_14153,N_11611);
nor UO_789 (O_789,N_14791,N_13099);
or UO_790 (O_790,N_10116,N_11522);
xnor UO_791 (O_791,N_13404,N_12893);
xor UO_792 (O_792,N_14624,N_12720);
nor UO_793 (O_793,N_10872,N_13205);
and UO_794 (O_794,N_11315,N_12429);
nor UO_795 (O_795,N_11805,N_11580);
and UO_796 (O_796,N_14755,N_13191);
xor UO_797 (O_797,N_14437,N_14953);
nand UO_798 (O_798,N_12578,N_13175);
and UO_799 (O_799,N_12718,N_12323);
nor UO_800 (O_800,N_13809,N_10618);
and UO_801 (O_801,N_12977,N_13673);
nor UO_802 (O_802,N_13220,N_11490);
nand UO_803 (O_803,N_11700,N_11241);
nand UO_804 (O_804,N_14634,N_14686);
nand UO_805 (O_805,N_11251,N_11986);
nor UO_806 (O_806,N_11997,N_12684);
nand UO_807 (O_807,N_11957,N_13435);
and UO_808 (O_808,N_11001,N_14593);
nand UO_809 (O_809,N_11385,N_11976);
and UO_810 (O_810,N_10087,N_10657);
and UO_811 (O_811,N_14337,N_10474);
or UO_812 (O_812,N_10556,N_11112);
and UO_813 (O_813,N_10106,N_12444);
nand UO_814 (O_814,N_10424,N_10613);
nor UO_815 (O_815,N_11505,N_10270);
xnor UO_816 (O_816,N_12240,N_10009);
or UO_817 (O_817,N_11260,N_10150);
nand UO_818 (O_818,N_12038,N_10537);
xnor UO_819 (O_819,N_11174,N_12046);
and UO_820 (O_820,N_12439,N_11788);
or UO_821 (O_821,N_11621,N_10996);
nor UO_822 (O_822,N_12026,N_11801);
and UO_823 (O_823,N_12077,N_10141);
nor UO_824 (O_824,N_10550,N_13667);
and UO_825 (O_825,N_11362,N_13626);
or UO_826 (O_826,N_14705,N_13295);
nor UO_827 (O_827,N_13193,N_12499);
and UO_828 (O_828,N_12573,N_11327);
or UO_829 (O_829,N_10741,N_11732);
or UO_830 (O_830,N_14514,N_12351);
nor UO_831 (O_831,N_13885,N_13864);
nand UO_832 (O_832,N_10447,N_12901);
or UO_833 (O_833,N_10845,N_13672);
xnor UO_834 (O_834,N_11808,N_10382);
nand UO_835 (O_835,N_14597,N_14146);
nand UO_836 (O_836,N_14567,N_11725);
or UO_837 (O_837,N_10429,N_11755);
nand UO_838 (O_838,N_14745,N_14902);
xor UO_839 (O_839,N_10147,N_12723);
and UO_840 (O_840,N_11018,N_11774);
nand UO_841 (O_841,N_11276,N_10266);
nor UO_842 (O_842,N_11840,N_13491);
xor UO_843 (O_843,N_11465,N_12773);
xor UO_844 (O_844,N_10363,N_10743);
or UO_845 (O_845,N_11127,N_14328);
xnor UO_846 (O_846,N_10051,N_12126);
nand UO_847 (O_847,N_13861,N_10571);
nand UO_848 (O_848,N_10481,N_11610);
xor UO_849 (O_849,N_14215,N_13593);
xor UO_850 (O_850,N_10213,N_14448);
and UO_851 (O_851,N_12266,N_12574);
xor UO_852 (O_852,N_13970,N_13603);
xnor UO_853 (O_853,N_12457,N_11723);
xor UO_854 (O_854,N_13576,N_13402);
and UO_855 (O_855,N_10734,N_13171);
nor UO_856 (O_856,N_11046,N_12987);
nand UO_857 (O_857,N_14404,N_13948);
and UO_858 (O_858,N_10649,N_14513);
xnor UO_859 (O_859,N_12475,N_13925);
nand UO_860 (O_860,N_14813,N_14156);
nand UO_861 (O_861,N_14022,N_11894);
or UO_862 (O_862,N_12854,N_12384);
and UO_863 (O_863,N_12697,N_14647);
and UO_864 (O_864,N_12798,N_12647);
nor UO_865 (O_865,N_13845,N_11292);
and UO_866 (O_866,N_12535,N_11455);
nand UO_867 (O_867,N_14424,N_10413);
and UO_868 (O_868,N_13493,N_10342);
xor UO_869 (O_869,N_13287,N_14271);
xnor UO_870 (O_870,N_12094,N_11791);
nand UO_871 (O_871,N_12144,N_13733);
nor UO_872 (O_872,N_11936,N_14789);
or UO_873 (O_873,N_13054,N_11418);
nor UO_874 (O_874,N_10112,N_14324);
and UO_875 (O_875,N_13333,N_14657);
or UO_876 (O_876,N_10320,N_14157);
xnor UO_877 (O_877,N_10393,N_10642);
xor UO_878 (O_878,N_10496,N_14559);
xor UO_879 (O_879,N_10265,N_11978);
and UO_880 (O_880,N_13371,N_14823);
or UO_881 (O_881,N_10703,N_10957);
nand UO_882 (O_882,N_11364,N_14104);
nor UO_883 (O_883,N_14590,N_12313);
or UO_884 (O_884,N_10314,N_14378);
nor UO_885 (O_885,N_10023,N_10804);
and UO_886 (O_886,N_11951,N_11459);
xnor UO_887 (O_887,N_10883,N_12530);
nand UO_888 (O_888,N_14974,N_10888);
nor UO_889 (O_889,N_11116,N_12818);
and UO_890 (O_890,N_11178,N_11280);
nor UO_891 (O_891,N_10161,N_10210);
and UO_892 (O_892,N_13130,N_10120);
nand UO_893 (O_893,N_10345,N_11062);
or UO_894 (O_894,N_12823,N_12808);
nand UO_895 (O_895,N_10168,N_12586);
xor UO_896 (O_896,N_11245,N_13310);
and UO_897 (O_897,N_13515,N_13791);
nand UO_898 (O_898,N_11079,N_12403);
and UO_899 (O_899,N_14266,N_13009);
or UO_900 (O_900,N_13490,N_11682);
and UO_901 (O_901,N_12484,N_13412);
nor UO_902 (O_902,N_13454,N_10533);
nand UO_903 (O_903,N_10110,N_12519);
xor UO_904 (O_904,N_10119,N_13284);
xnor UO_905 (O_905,N_10500,N_13441);
nand UO_906 (O_906,N_10752,N_12315);
nand UO_907 (O_907,N_13365,N_13434);
nor UO_908 (O_908,N_11825,N_13534);
nor UO_909 (O_909,N_10641,N_13624);
xnor UO_910 (O_910,N_12541,N_13152);
or UO_911 (O_911,N_12343,N_13436);
nor UO_912 (O_912,N_11630,N_11562);
nand UO_913 (O_913,N_12702,N_13114);
xor UO_914 (O_914,N_11060,N_10561);
nor UO_915 (O_915,N_12507,N_11224);
xnor UO_916 (O_916,N_11353,N_10235);
and UO_917 (O_917,N_13048,N_12951);
nand UO_918 (O_918,N_11190,N_13460);
or UO_919 (O_919,N_10338,N_13458);
nand UO_920 (O_920,N_10288,N_13634);
nor UO_921 (O_921,N_10405,N_10412);
nand UO_922 (O_922,N_10915,N_12167);
or UO_923 (O_923,N_10197,N_13606);
nand UO_924 (O_924,N_13097,N_13020);
nand UO_925 (O_925,N_11969,N_14417);
xor UO_926 (O_926,N_11240,N_11369);
or UO_927 (O_927,N_12112,N_13103);
and UO_928 (O_928,N_11205,N_10239);
and UO_929 (O_929,N_10928,N_11304);
nand UO_930 (O_930,N_13995,N_14834);
and UO_931 (O_931,N_10829,N_13549);
nor UO_932 (O_932,N_12480,N_11284);
and UO_933 (O_933,N_11532,N_13745);
and UO_934 (O_934,N_11499,N_13766);
nand UO_935 (O_935,N_14846,N_14550);
nand UO_936 (O_936,N_12365,N_14435);
xnor UO_937 (O_937,N_14790,N_10894);
nor UO_938 (O_938,N_10442,N_13680);
xnor UO_939 (O_939,N_10190,N_11565);
and UO_940 (O_940,N_12565,N_11868);
or UO_941 (O_941,N_12004,N_11999);
xor UO_942 (O_942,N_10428,N_11421);
nor UO_943 (O_943,N_11875,N_13469);
and UO_944 (O_944,N_14508,N_12920);
or UO_945 (O_945,N_11217,N_12242);
and UO_946 (O_946,N_11098,N_13161);
xnor UO_947 (O_947,N_12885,N_12072);
and UO_948 (O_948,N_12159,N_11955);
xnor UO_949 (O_949,N_10369,N_10315);
nor UO_950 (O_950,N_11666,N_14410);
nand UO_951 (O_951,N_13833,N_10256);
xor UO_952 (O_952,N_14986,N_12708);
nand UO_953 (O_953,N_12529,N_12656);
nor UO_954 (O_954,N_11768,N_10581);
nor UO_955 (O_955,N_11780,N_14751);
nand UO_956 (O_956,N_11460,N_12362);
nand UO_957 (O_957,N_14264,N_11977);
and UO_958 (O_958,N_14800,N_14842);
nor UO_959 (O_959,N_12192,N_12830);
xor UO_960 (O_960,N_12943,N_11287);
xor UO_961 (O_961,N_14841,N_12415);
or UO_962 (O_962,N_11592,N_13004);
or UO_963 (O_963,N_14665,N_13459);
nor UO_964 (O_964,N_12468,N_13290);
or UO_965 (O_965,N_11228,N_12367);
and UO_966 (O_966,N_13865,N_12640);
and UO_967 (O_967,N_11724,N_11177);
or UO_968 (O_968,N_12379,N_12043);
xnor UO_969 (O_969,N_12915,N_14110);
and UO_970 (O_970,N_13820,N_14269);
xor UO_971 (O_971,N_11341,N_14488);
and UO_972 (O_972,N_13752,N_13600);
nand UO_973 (O_973,N_12846,N_12226);
nor UO_974 (O_974,N_10704,N_10844);
nand UO_975 (O_975,N_10538,N_11512);
or UO_976 (O_976,N_11003,N_12467);
nor UO_977 (O_977,N_10227,N_14979);
nand UO_978 (O_978,N_10416,N_10729);
nor UO_979 (O_979,N_12372,N_12733);
nand UO_980 (O_980,N_10843,N_14267);
and UO_981 (O_981,N_13341,N_14662);
and UO_982 (O_982,N_11489,N_14972);
nor UO_983 (O_983,N_14323,N_13635);
nor UO_984 (O_984,N_10249,N_13638);
nand UO_985 (O_985,N_13227,N_10127);
or UO_986 (O_986,N_14013,N_12399);
nand UO_987 (O_987,N_11964,N_14575);
xnor UO_988 (O_988,N_14226,N_13740);
nor UO_989 (O_989,N_14669,N_12711);
xnor UO_990 (O_990,N_12195,N_14415);
or UO_991 (O_991,N_11300,N_12328);
and UO_992 (O_992,N_10659,N_12590);
or UO_993 (O_993,N_11728,N_10519);
or UO_994 (O_994,N_10453,N_13032);
xnor UO_995 (O_995,N_11661,N_14808);
and UO_996 (O_996,N_11471,N_12366);
or UO_997 (O_997,N_13061,N_10616);
nand UO_998 (O_998,N_14133,N_14596);
nor UO_999 (O_999,N_12670,N_14147);
nor UO_1000 (O_1000,N_10667,N_11389);
and UO_1001 (O_1001,N_12485,N_10640);
nand UO_1002 (O_1002,N_10377,N_11000);
xor UO_1003 (O_1003,N_10913,N_10886);
xnor UO_1004 (O_1004,N_12619,N_11124);
and UO_1005 (O_1005,N_10877,N_14107);
or UO_1006 (O_1006,N_14944,N_12880);
or UO_1007 (O_1007,N_11468,N_14636);
and UO_1008 (O_1008,N_10494,N_12325);
nand UO_1009 (O_1009,N_10878,N_11707);
or UO_1010 (O_1010,N_10516,N_13987);
nand UO_1011 (O_1011,N_14541,N_12456);
xor UO_1012 (O_1012,N_14460,N_10016);
xnor UO_1013 (O_1013,N_14496,N_10569);
nor UO_1014 (O_1014,N_11857,N_10375);
nand UO_1015 (O_1015,N_14115,N_12414);
nand UO_1016 (O_1016,N_12110,N_11753);
xnor UO_1017 (O_1017,N_14088,N_14439);
xnor UO_1018 (O_1018,N_10037,N_14536);
nand UO_1019 (O_1019,N_10385,N_14820);
or UO_1020 (O_1020,N_10459,N_11608);
nand UO_1021 (O_1021,N_12946,N_10737);
nand UO_1022 (O_1022,N_13073,N_12878);
nor UO_1023 (O_1023,N_11099,N_14112);
xnor UO_1024 (O_1024,N_14006,N_14954);
and UO_1025 (O_1025,N_10322,N_14538);
xor UO_1026 (O_1026,N_13716,N_11373);
or UO_1027 (O_1027,N_11042,N_11626);
and UO_1028 (O_1028,N_10004,N_13068);
and UO_1029 (O_1029,N_11918,N_11467);
and UO_1030 (O_1030,N_13062,N_13123);
or UO_1031 (O_1031,N_12797,N_14505);
xnor UO_1032 (O_1032,N_13955,N_11399);
and UO_1033 (O_1033,N_10603,N_13992);
nand UO_1034 (O_1034,N_13291,N_13329);
or UO_1035 (O_1035,N_11689,N_14603);
xnor UO_1036 (O_1036,N_12234,N_14494);
xnor UO_1037 (O_1037,N_12296,N_11972);
nand UO_1038 (O_1038,N_13144,N_13577);
nor UO_1039 (O_1039,N_12015,N_14887);
nand UO_1040 (O_1040,N_13582,N_11321);
and UO_1041 (O_1041,N_12989,N_12826);
nand UO_1042 (O_1042,N_12436,N_10547);
and UO_1043 (O_1043,N_13188,N_13170);
xor UO_1044 (O_1044,N_11049,N_11252);
and UO_1045 (O_1045,N_12282,N_10977);
or UO_1046 (O_1046,N_12314,N_14828);
and UO_1047 (O_1047,N_14912,N_12528);
and UO_1048 (O_1048,N_12054,N_11101);
or UO_1049 (O_1049,N_10939,N_12426);
and UO_1050 (O_1050,N_12780,N_10307);
xor UO_1051 (O_1051,N_13601,N_13921);
or UO_1052 (O_1052,N_13609,N_13842);
nor UO_1053 (O_1053,N_14461,N_11834);
xor UO_1054 (O_1054,N_13878,N_10562);
nand UO_1055 (O_1055,N_13768,N_11166);
nor UO_1056 (O_1056,N_12139,N_14764);
xnor UO_1057 (O_1057,N_14768,N_10014);
and UO_1058 (O_1058,N_11914,N_11662);
xnor UO_1059 (O_1059,N_14333,N_14003);
or UO_1060 (O_1060,N_11316,N_13957);
xnor UO_1061 (O_1061,N_10856,N_12000);
or UO_1062 (O_1062,N_13463,N_12118);
or UO_1063 (O_1063,N_11900,N_13846);
nand UO_1064 (O_1064,N_14960,N_13649);
nor UO_1065 (O_1065,N_13720,N_11151);
nand UO_1066 (O_1066,N_13790,N_13025);
or UO_1067 (O_1067,N_13702,N_10986);
xnor UO_1068 (O_1068,N_12087,N_12059);
and UO_1069 (O_1069,N_10356,N_13511);
nand UO_1070 (O_1070,N_12609,N_12219);
nor UO_1071 (O_1071,N_10049,N_13098);
nor UO_1072 (O_1072,N_14913,N_12836);
and UO_1073 (O_1073,N_12443,N_14002);
nor UO_1074 (O_1074,N_13625,N_12462);
and UO_1075 (O_1075,N_11184,N_11211);
or UO_1076 (O_1076,N_13403,N_14001);
and UO_1077 (O_1077,N_13949,N_13289);
or UO_1078 (O_1078,N_13370,N_14151);
and UO_1079 (O_1079,N_10080,N_12857);
or UO_1080 (O_1080,N_10170,N_10850);
xnor UO_1081 (O_1081,N_11640,N_12649);
and UO_1082 (O_1082,N_12834,N_11663);
and UO_1083 (O_1083,N_14917,N_14874);
and UO_1084 (O_1084,N_13190,N_13639);
and UO_1085 (O_1085,N_10188,N_12754);
xor UO_1086 (O_1086,N_11173,N_11089);
nor UO_1087 (O_1087,N_11876,N_10830);
or UO_1088 (O_1088,N_10048,N_11121);
nand UO_1089 (O_1089,N_12544,N_12790);
and UO_1090 (O_1090,N_10390,N_10482);
xnor UO_1091 (O_1091,N_11147,N_13409);
xnor UO_1092 (O_1092,N_14482,N_12303);
and UO_1093 (O_1093,N_14522,N_10497);
xor UO_1094 (O_1094,N_14933,N_11372);
and UO_1095 (O_1095,N_10117,N_13420);
and UO_1096 (O_1096,N_13177,N_13462);
xnor UO_1097 (O_1097,N_10580,N_11594);
xnor UO_1098 (O_1098,N_11368,N_10891);
and UO_1099 (O_1099,N_13953,N_12382);
xnor UO_1100 (O_1100,N_11082,N_11651);
xnor UO_1101 (O_1101,N_12919,N_11153);
and UO_1102 (O_1102,N_10071,N_11722);
nor UO_1103 (O_1103,N_13969,N_12181);
nor UO_1104 (O_1104,N_13799,N_12206);
xnor UO_1105 (O_1105,N_12147,N_10220);
and UO_1106 (O_1106,N_10066,N_11022);
xnor UO_1107 (O_1107,N_11658,N_11040);
or UO_1108 (O_1108,N_10300,N_14009);
xnor UO_1109 (O_1109,N_13550,N_14321);
and UO_1110 (O_1110,N_11254,N_14818);
nand UO_1111 (O_1111,N_14306,N_10651);
xor UO_1112 (O_1112,N_11954,N_14854);
xnor UO_1113 (O_1113,N_14829,N_13440);
or UO_1114 (O_1114,N_10795,N_10002);
nand UO_1115 (O_1115,N_12940,N_11690);
xor UO_1116 (O_1116,N_14102,N_10044);
nor UO_1117 (O_1117,N_11597,N_10295);
or UO_1118 (O_1118,N_11578,N_12655);
nand UO_1119 (O_1119,N_12510,N_10139);
or UO_1120 (O_1120,N_11250,N_13533);
nor UO_1121 (O_1121,N_11442,N_10206);
and UO_1122 (O_1122,N_10867,N_14602);
xor UO_1123 (O_1123,N_10668,N_12816);
or UO_1124 (O_1124,N_13764,N_13040);
nand UO_1125 (O_1125,N_14847,N_14523);
and UO_1126 (O_1126,N_11387,N_13694);
xor UO_1127 (O_1127,N_14092,N_12138);
nand UO_1128 (O_1128,N_10506,N_10898);
nor UO_1129 (O_1129,N_13222,N_11464);
xor UO_1130 (O_1130,N_13719,N_11213);
or UO_1131 (O_1131,N_13939,N_13349);
nand UO_1132 (O_1132,N_13074,N_14775);
or UO_1133 (O_1133,N_11917,N_13051);
xor UO_1134 (O_1134,N_10033,N_13974);
xor UO_1135 (O_1135,N_14714,N_11975);
nand UO_1136 (O_1136,N_14040,N_14588);
nor UO_1137 (O_1137,N_10863,N_13847);
nand UO_1138 (O_1138,N_11319,N_11843);
or UO_1139 (O_1139,N_13553,N_12974);
xnor UO_1140 (O_1140,N_13256,N_13067);
and UO_1141 (O_1141,N_12549,N_12717);
or UO_1142 (O_1142,N_14632,N_13681);
nand UO_1143 (O_1143,N_10670,N_10999);
nand UO_1144 (O_1144,N_10064,N_10132);
or UO_1145 (O_1145,N_12294,N_14238);
or UO_1146 (O_1146,N_10303,N_13937);
and UO_1147 (O_1147,N_11279,N_10786);
nor UO_1148 (O_1148,N_11631,N_11058);
nor UO_1149 (O_1149,N_11833,N_10555);
nor UO_1150 (O_1150,N_11967,N_12262);
xor UO_1151 (O_1151,N_11590,N_14731);
and UO_1152 (O_1152,N_11114,N_10601);
and UO_1153 (O_1153,N_12964,N_14364);
xnor UO_1154 (O_1154,N_12726,N_10401);
and UO_1155 (O_1155,N_12364,N_10690);
and UO_1156 (O_1156,N_11396,N_13023);
nand UO_1157 (O_1157,N_14920,N_14551);
and UO_1158 (O_1158,N_12596,N_11125);
nand UO_1159 (O_1159,N_13855,N_11962);
xnor UO_1160 (O_1160,N_10204,N_10403);
nor UO_1161 (O_1161,N_10994,N_12210);
or UO_1162 (O_1162,N_11066,N_12648);
or UO_1163 (O_1163,N_12253,N_14664);
or UO_1164 (O_1164,N_10435,N_11553);
and UO_1165 (O_1165,N_12164,N_12257);
nor UO_1166 (O_1166,N_12546,N_12413);
xnor UO_1167 (O_1167,N_13853,N_12175);
and UO_1168 (O_1168,N_12293,N_12839);
or UO_1169 (O_1169,N_13035,N_12713);
and UO_1170 (O_1170,N_10022,N_10792);
nor UO_1171 (O_1171,N_11729,N_10896);
and UO_1172 (O_1172,N_11678,N_12307);
and UO_1173 (O_1173,N_11010,N_13478);
nand UO_1174 (O_1174,N_12388,N_10293);
nand UO_1175 (O_1175,N_12289,N_14243);
and UO_1176 (O_1176,N_10930,N_12872);
nor UO_1177 (O_1177,N_12743,N_12286);
xor UO_1178 (O_1178,N_14357,N_10291);
nor UO_1179 (O_1179,N_14273,N_10636);
nand UO_1180 (O_1180,N_13852,N_12851);
or UO_1181 (O_1181,N_11776,N_11552);
or UO_1182 (O_1182,N_12566,N_11982);
or UO_1183 (O_1183,N_10527,N_11469);
nand UO_1184 (O_1184,N_11295,N_11720);
xor UO_1185 (O_1185,N_14346,N_13424);
nand UO_1186 (O_1186,N_14056,N_12025);
nand UO_1187 (O_1187,N_12380,N_10803);
nand UO_1188 (O_1188,N_14208,N_11718);
nor UO_1189 (O_1189,N_13407,N_10475);
nor UO_1190 (O_1190,N_10600,N_13512);
xor UO_1191 (O_1191,N_14668,N_13982);
nand UO_1192 (O_1192,N_10774,N_13086);
or UO_1193 (O_1193,N_14198,N_10269);
nor UO_1194 (O_1194,N_13055,N_10895);
and UO_1195 (O_1195,N_10854,N_12052);
and UO_1196 (O_1196,N_10202,N_13134);
or UO_1197 (O_1197,N_13566,N_13169);
nand UO_1198 (O_1198,N_11156,N_13743);
and UO_1199 (O_1199,N_10418,N_12924);
and UO_1200 (O_1200,N_14661,N_14616);
or UO_1201 (O_1201,N_14886,N_14141);
and UO_1202 (O_1202,N_14554,N_10277);
xnor UO_1203 (O_1203,N_10626,N_12279);
and UO_1204 (O_1204,N_13787,N_13039);
nand UO_1205 (O_1205,N_10836,N_13965);
xnor UO_1206 (O_1206,N_10224,N_12483);
or UO_1207 (O_1207,N_12134,N_12912);
nand UO_1208 (O_1208,N_14563,N_13869);
and UO_1209 (O_1209,N_14817,N_13910);
nor UO_1210 (O_1210,N_11596,N_14172);
or UO_1211 (O_1211,N_11139,N_13309);
nand UO_1212 (O_1212,N_11410,N_14611);
xnor UO_1213 (O_1213,N_11187,N_10515);
nand UO_1214 (O_1214,N_12783,N_13271);
nor UO_1215 (O_1215,N_11204,N_14641);
or UO_1216 (O_1216,N_12764,N_13442);
and UO_1217 (O_1217,N_11841,N_13946);
or UO_1218 (O_1218,N_11680,N_14618);
or UO_1219 (O_1219,N_12809,N_14422);
nor UO_1220 (O_1220,N_11556,N_14890);
and UO_1221 (O_1221,N_10985,N_10971);
or UO_1222 (O_1222,N_14985,N_11568);
and UO_1223 (O_1223,N_12010,N_11095);
nor UO_1224 (O_1224,N_10927,N_12244);
nand UO_1225 (O_1225,N_12106,N_13795);
or UO_1226 (O_1226,N_13531,N_14233);
nand UO_1227 (O_1227,N_11119,N_11451);
or UO_1228 (O_1228,N_10351,N_10379);
and UO_1229 (O_1229,N_13263,N_12538);
or UO_1230 (O_1230,N_14444,N_14171);
xor UO_1231 (O_1231,N_13981,N_10297);
and UO_1232 (O_1232,N_14067,N_11072);
nand UO_1233 (O_1233,N_14391,N_13254);
or UO_1234 (O_1234,N_14758,N_14591);
xnor UO_1235 (O_1235,N_11584,N_12659);
or UO_1236 (O_1236,N_11817,N_13231);
and UO_1237 (O_1237,N_10225,N_10171);
xnor UO_1238 (O_1238,N_11365,N_14201);
and UO_1239 (O_1239,N_14524,N_11803);
nor UO_1240 (O_1240,N_10330,N_14290);
nand UO_1241 (O_1241,N_14868,N_11087);
nand UO_1242 (O_1242,N_11880,N_11188);
xnor UO_1243 (O_1243,N_12719,N_10421);
or UO_1244 (O_1244,N_14120,N_12067);
nand UO_1245 (O_1245,N_13143,N_11598);
nor UO_1246 (O_1246,N_14084,N_13741);
or UO_1247 (O_1247,N_11322,N_14748);
nand UO_1248 (O_1248,N_10807,N_12966);
and UO_1249 (O_1249,N_12604,N_13755);
or UO_1250 (O_1250,N_10380,N_11226);
nand UO_1251 (O_1251,N_10806,N_10788);
and UO_1252 (O_1252,N_11175,N_13379);
nor UO_1253 (O_1253,N_10193,N_10318);
nor UO_1254 (O_1254,N_14605,N_10628);
nor UO_1255 (O_1255,N_14589,N_14179);
or UO_1256 (O_1256,N_14989,N_12075);
nand UO_1257 (O_1257,N_12221,N_10909);
and UO_1258 (O_1258,N_10954,N_12550);
xnor UO_1259 (O_1259,N_12033,N_14055);
nor UO_1260 (O_1260,N_14099,N_11255);
or UO_1261 (O_1261,N_14856,N_13559);
or UO_1262 (O_1262,N_13518,N_11555);
or UO_1263 (O_1263,N_10599,N_14873);
and UO_1264 (O_1264,N_10398,N_10919);
nand UO_1265 (O_1265,N_11863,N_11648);
nand UO_1266 (O_1266,N_12341,N_10305);
or UO_1267 (O_1267,N_13938,N_10754);
xnor UO_1268 (O_1268,N_13562,N_14700);
and UO_1269 (O_1269,N_13382,N_10209);
or UO_1270 (O_1270,N_10532,N_10286);
xor UO_1271 (O_1271,N_11766,N_14477);
xnor UO_1272 (O_1272,N_10339,N_11360);
xnor UO_1273 (O_1273,N_13538,N_14695);
xnor UO_1274 (O_1274,N_12575,N_11586);
and UO_1275 (O_1275,N_13485,N_10183);
xnor UO_1276 (O_1276,N_12725,N_14135);
xor UO_1277 (O_1277,N_13539,N_11077);
and UO_1278 (O_1278,N_11591,N_14911);
nor UO_1279 (O_1279,N_11929,N_11514);
or UO_1280 (O_1280,N_11877,N_14288);
or UO_1281 (O_1281,N_14996,N_12998);
xnor UO_1282 (O_1282,N_10011,N_13133);
or UO_1283 (O_1283,N_12613,N_11068);
xor UO_1284 (O_1284,N_10094,N_13047);
nor UO_1285 (O_1285,N_10211,N_14283);
nor UO_1286 (O_1286,N_14126,N_14396);
nand UO_1287 (O_1287,N_12080,N_10557);
and UO_1288 (O_1288,N_11191,N_11282);
nand UO_1289 (O_1289,N_13131,N_11519);
xor UO_1290 (O_1290,N_11947,N_10536);
xnor UO_1291 (O_1291,N_10647,N_11494);
or UO_1292 (O_1292,N_12517,N_13417);
nand UO_1293 (O_1293,N_14175,N_12297);
nor UO_1294 (O_1294,N_10587,N_11035);
xnor UO_1295 (O_1295,N_13686,N_13235);
xor UO_1296 (O_1296,N_11815,N_14994);
xor UO_1297 (O_1297,N_12947,N_13954);
nand UO_1298 (O_1298,N_11267,N_11667);
and UO_1299 (O_1299,N_14298,N_13118);
and UO_1300 (O_1300,N_10530,N_10926);
and UO_1301 (O_1301,N_13019,N_13386);
or UO_1302 (O_1302,N_11920,N_14041);
and UO_1303 (O_1303,N_14218,N_12858);
nand UO_1304 (O_1304,N_13185,N_10583);
xor UO_1305 (O_1305,N_14295,N_10169);
or UO_1306 (O_1306,N_11100,N_14610);
nor UO_1307 (O_1307,N_10749,N_12449);
or UO_1308 (O_1308,N_13731,N_11478);
xor UO_1309 (O_1309,N_14248,N_14558);
nand UO_1310 (O_1310,N_11885,N_14689);
and UO_1311 (O_1311,N_14880,N_11573);
nor UO_1312 (O_1312,N_12391,N_10438);
or UO_1313 (O_1313,N_12628,N_11075);
or UO_1314 (O_1314,N_12770,N_11717);
and UO_1315 (O_1315,N_14967,N_13076);
xor UO_1316 (O_1316,N_13158,N_11435);
nor UO_1317 (O_1317,N_10832,N_12040);
and UO_1318 (O_1318,N_11697,N_12011);
nand UO_1319 (O_1319,N_13496,N_11938);
nand UO_1320 (O_1320,N_11441,N_13908);
or UO_1321 (O_1321,N_10510,N_10746);
and UO_1322 (O_1322,N_10156,N_13060);
xor UO_1323 (O_1323,N_14555,N_13258);
xnor UO_1324 (O_1324,N_10146,N_12395);
nand UO_1325 (O_1325,N_11961,N_13094);
nor UO_1326 (O_1326,N_14643,N_13244);
xnor UO_1327 (O_1327,N_10486,N_14801);
nand UO_1328 (O_1328,N_13574,N_13614);
xnor UO_1329 (O_1329,N_11548,N_14862);
nand UO_1330 (O_1330,N_13470,N_10155);
nor UO_1331 (O_1331,N_11935,N_11858);
and UO_1332 (O_1332,N_13736,N_10847);
nand UO_1333 (O_1333,N_12995,N_13141);
nor UO_1334 (O_1334,N_10058,N_12107);
or UO_1335 (O_1335,N_14188,N_11558);
or UO_1336 (O_1336,N_13059,N_12975);
nand UO_1337 (O_1337,N_14821,N_13246);
or UO_1338 (O_1338,N_12996,N_11735);
nand UO_1339 (O_1339,N_14356,N_11704);
and UO_1340 (O_1340,N_14308,N_10354);
nor UO_1341 (O_1341,N_10406,N_14491);
and UO_1342 (O_1342,N_10995,N_10092);
xnor UO_1343 (O_1343,N_14354,N_14617);
and UO_1344 (O_1344,N_11281,N_12841);
nor UO_1345 (O_1345,N_11165,N_14932);
xor UO_1346 (O_1346,N_10471,N_13167);
xor UO_1347 (O_1347,N_14286,N_14568);
and UO_1348 (O_1348,N_11674,N_10420);
or UO_1349 (O_1349,N_12564,N_13780);
or UO_1350 (O_1350,N_10489,N_14311);
nor UO_1351 (O_1351,N_10855,N_13689);
or UO_1352 (O_1352,N_12890,N_13817);
and UO_1353 (O_1353,N_12832,N_10324);
nor UO_1354 (O_1354,N_12448,N_14612);
and UO_1355 (O_1355,N_14428,N_12534);
and UO_1356 (O_1356,N_12911,N_14038);
nor UO_1357 (O_1357,N_12131,N_12378);
and UO_1358 (O_1358,N_11882,N_10911);
or UO_1359 (O_1359,N_13268,N_14977);
nand UO_1360 (O_1360,N_10245,N_13693);
or UO_1361 (O_1361,N_13698,N_11644);
and UO_1362 (O_1362,N_13510,N_14754);
nand UO_1363 (O_1363,N_14822,N_11530);
nor UO_1364 (O_1364,N_11363,N_13066);
or UO_1365 (O_1365,N_12458,N_14091);
and UO_1366 (O_1366,N_10584,N_14742);
and UO_1367 (O_1367,N_14510,N_14799);
xnor UO_1368 (O_1368,N_14021,N_10759);
or UO_1369 (O_1369,N_12155,N_14389);
nand UO_1370 (O_1370,N_10708,N_11444);
or UO_1371 (O_1371,N_11916,N_13827);
and UO_1372 (O_1372,N_10248,N_10579);
and UO_1373 (O_1373,N_10907,N_13742);
nor UO_1374 (O_1374,N_11351,N_11404);
nor UO_1375 (O_1375,N_14016,N_12140);
and UO_1376 (O_1376,N_12358,N_12021);
nor UO_1377 (O_1377,N_10540,N_12331);
and UO_1378 (O_1378,N_12805,N_13749);
nor UO_1379 (O_1379,N_13398,N_13146);
nand UO_1380 (O_1380,N_13423,N_13532);
nand UO_1381 (O_1381,N_12273,N_14718);
or UO_1382 (O_1382,N_14772,N_14935);
nor UO_1383 (O_1383,N_11816,N_13251);
and UO_1384 (O_1384,N_10370,N_12009);
and UO_1385 (O_1385,N_10721,N_14674);
nand UO_1386 (O_1386,N_13228,N_10316);
or UO_1387 (O_1387,N_13328,N_13467);
xor UO_1388 (O_1388,N_10238,N_14344);
nand UO_1389 (O_1389,N_12170,N_13918);
nor UO_1390 (O_1390,N_12028,N_11288);
nand UO_1391 (O_1391,N_11271,N_13536);
nor UO_1392 (O_1392,N_14239,N_11483);
or UO_1393 (O_1393,N_13848,N_13947);
xnor UO_1394 (O_1394,N_10609,N_14653);
nor UO_1395 (O_1395,N_11091,N_11229);
nor UO_1396 (O_1396,N_13856,N_10974);
or UO_1397 (O_1397,N_10273,N_12511);
xor UO_1398 (O_1398,N_11320,N_13675);
nand UO_1399 (O_1399,N_10876,N_13608);
nor UO_1400 (O_1400,N_10091,N_10196);
nand UO_1401 (O_1401,N_11851,N_13011);
nor UO_1402 (O_1402,N_12704,N_13013);
xor UO_1403 (O_1403,N_10368,N_14770);
xor UO_1404 (O_1404,N_13489,N_13064);
xor UO_1405 (O_1405,N_13201,N_14855);
nor UO_1406 (O_1406,N_10350,N_11714);
nand UO_1407 (O_1407,N_10114,N_11810);
or UO_1408 (O_1408,N_12251,N_12158);
or UO_1409 (O_1409,N_12883,N_10837);
xnor UO_1410 (O_1410,N_12871,N_14542);
xnor UO_1411 (O_1411,N_12942,N_11567);
and UO_1412 (O_1412,N_14094,N_14164);
nor UO_1413 (O_1413,N_14279,N_11069);
or UO_1414 (O_1414,N_11730,N_14517);
nand UO_1415 (O_1415,N_12992,N_13418);
xnor UO_1416 (O_1416,N_11155,N_12581);
or UO_1417 (O_1417,N_10901,N_13703);
or UO_1418 (O_1418,N_12945,N_13979);
nand UO_1419 (O_1419,N_10596,N_10391);
or UO_1420 (O_1420,N_13457,N_11593);
xnor UO_1421 (O_1421,N_11625,N_10294);
nor UO_1422 (O_1422,N_10109,N_10756);
or UO_1423 (O_1423,N_11051,N_12860);
nand UO_1424 (O_1424,N_10694,N_11856);
and UO_1425 (O_1425,N_14704,N_11820);
or UO_1426 (O_1426,N_13416,N_12160);
or UO_1427 (O_1427,N_12793,N_14739);
or UO_1428 (O_1428,N_14441,N_14440);
and UO_1429 (O_1429,N_10173,N_10573);
xor UO_1430 (O_1430,N_12231,N_14261);
and UO_1431 (O_1431,N_14278,N_13257);
nand UO_1432 (O_1432,N_11366,N_12831);
nor UO_1433 (O_1433,N_14980,N_13483);
or UO_1434 (O_1434,N_10378,N_14214);
xor UO_1435 (O_1435,N_11719,N_14423);
nor UO_1436 (O_1436,N_14125,N_12970);
nor UO_1437 (O_1437,N_14360,N_12288);
nor UO_1438 (O_1438,N_13747,N_14028);
and UO_1439 (O_1439,N_10897,N_13357);
nand UO_1440 (O_1440,N_12908,N_11083);
or UO_1441 (O_1441,N_14161,N_14114);
or UO_1442 (O_1442,N_13668,N_14684);
nand UO_1443 (O_1443,N_14338,N_10622);
nor UO_1444 (O_1444,N_12081,N_13444);
or UO_1445 (O_1445,N_13162,N_13399);
or UO_1446 (O_1446,N_13991,N_13313);
xnor UO_1447 (O_1447,N_10710,N_14259);
xnor UO_1448 (O_1448,N_11779,N_14546);
or UO_1449 (O_1449,N_13880,N_12580);
or UO_1450 (O_1450,N_11495,N_13571);
or UO_1451 (O_1451,N_11946,N_11624);
xnor UO_1452 (O_1452,N_14470,N_10964);
nand UO_1453 (O_1453,N_14232,N_14210);
xor UO_1454 (O_1454,N_11135,N_14916);
and UO_1455 (O_1455,N_13919,N_14759);
nor UO_1456 (O_1456,N_10666,N_12758);
and UO_1457 (O_1457,N_11419,N_11446);
xor UO_1458 (O_1458,N_14309,N_13249);
and UO_1459 (O_1459,N_14497,N_11289);
or UO_1460 (O_1460,N_13352,N_12600);
nor UO_1461 (O_1461,N_12474,N_14905);
xor UO_1462 (O_1462,N_14462,N_11041);
xnor UO_1463 (O_1463,N_11359,N_13279);
nand UO_1464 (O_1464,N_12076,N_11741);
nor UO_1465 (O_1465,N_10237,N_13321);
or UO_1466 (O_1466,N_12537,N_11158);
xnor UO_1467 (O_1467,N_11844,N_10552);
xor UO_1468 (O_1468,N_13376,N_11786);
or UO_1469 (O_1469,N_10079,N_13125);
nor UO_1470 (O_1470,N_12469,N_11795);
nor UO_1471 (O_1471,N_10063,N_14637);
or UO_1472 (O_1472,N_14959,N_11274);
xnor UO_1473 (O_1473,N_13643,N_12921);
or UO_1474 (O_1474,N_14355,N_11518);
or UO_1475 (O_1475,N_14121,N_14651);
or UO_1476 (O_1476,N_12585,N_12284);
nor UO_1477 (O_1477,N_13426,N_14426);
xnor UO_1478 (O_1478,N_12593,N_11710);
xor UO_1479 (O_1479,N_13482,N_13671);
xor UO_1480 (O_1480,N_14186,N_14606);
or UO_1481 (O_1481,N_14693,N_14405);
nor UO_1482 (O_1482,N_13525,N_13419);
and UO_1483 (O_1483,N_11493,N_10554);
nand UO_1484 (O_1484,N_10905,N_14549);
nor UO_1485 (O_1485,N_13117,N_14556);
or UO_1486 (O_1486,N_10522,N_12269);
and UO_1487 (O_1487,N_13008,N_13825);
and UO_1488 (O_1488,N_13408,N_11266);
nand UO_1489 (O_1489,N_12385,N_13052);
nand UO_1490 (O_1490,N_10381,N_10458);
nand UO_1491 (O_1491,N_14507,N_12020);
nand UO_1492 (O_1492,N_13670,N_14476);
and UO_1493 (O_1493,N_13916,N_10535);
nand UO_1494 (O_1494,N_14382,N_12505);
nand UO_1495 (O_1495,N_11575,N_11023);
nand UO_1496 (O_1496,N_11527,N_13951);
nand UO_1497 (O_1497,N_11206,N_13368);
nor UO_1498 (O_1498,N_14123,N_12700);
nand UO_1499 (O_1499,N_11203,N_10970);
xor UO_1500 (O_1500,N_14955,N_14930);
and UO_1501 (O_1501,N_13973,N_12283);
xor UO_1502 (O_1502,N_12738,N_12419);
nor UO_1503 (O_1503,N_12802,N_10334);
or UO_1504 (O_1504,N_14914,N_13725);
nand UO_1505 (O_1505,N_14978,N_14614);
and UO_1506 (O_1506,N_12787,N_13528);
xor UO_1507 (O_1507,N_14242,N_11711);
xor UO_1508 (O_1508,N_12174,N_14387);
or UO_1509 (O_1509,N_13621,N_11940);
and UO_1510 (O_1510,N_11642,N_10607);
nand UO_1511 (O_1511,N_12762,N_14361);
nor UO_1512 (O_1512,N_10755,N_14453);
nand UO_1513 (O_1513,N_10768,N_11302);
xnor UO_1514 (O_1514,N_11601,N_14708);
nand UO_1515 (O_1515,N_11653,N_13866);
and UO_1516 (O_1516,N_12136,N_10057);
xnor UO_1517 (O_1517,N_11731,N_10104);
nor UO_1518 (O_1518,N_11899,N_12261);
xor UO_1519 (O_1519,N_11305,N_11222);
and UO_1520 (O_1520,N_14314,N_12582);
or UO_1521 (O_1521,N_11108,N_11048);
xnor UO_1522 (O_1522,N_11293,N_12088);
nand UO_1523 (O_1523,N_13336,N_13691);
nor UO_1524 (O_1524,N_12983,N_13772);
or UO_1525 (O_1525,N_14158,N_10007);
nor UO_1526 (O_1526,N_13406,N_11193);
nor UO_1527 (O_1527,N_13278,N_10617);
and UO_1528 (O_1528,N_11669,N_11307);
nor UO_1529 (O_1529,N_14079,N_14987);
or UO_1530 (O_1530,N_11612,N_14045);
or UO_1531 (O_1531,N_11059,N_10870);
and UO_1532 (O_1532,N_11879,N_12312);
xnor UO_1533 (O_1533,N_13206,N_14465);
and UO_1534 (O_1534,N_12318,N_11547);
nor UO_1535 (O_1535,N_10163,N_12121);
xnor UO_1536 (O_1536,N_12280,N_11160);
and UO_1537 (O_1537,N_10264,N_10779);
xnor UO_1538 (O_1538,N_10465,N_14166);
and UO_1539 (O_1539,N_10775,N_14548);
xnor UO_1540 (O_1540,N_12437,N_12113);
xnor UO_1541 (O_1541,N_14743,N_10910);
nor UO_1542 (O_1542,N_11214,N_11605);
nand UO_1543 (O_1543,N_12714,N_14782);
and UO_1544 (O_1544,N_13630,N_13178);
nand UO_1545 (O_1545,N_10940,N_13783);
or UO_1546 (O_1546,N_10705,N_12736);
and UO_1547 (O_1547,N_10184,N_14535);
xnor UO_1548 (O_1548,N_12861,N_14036);
nand UO_1549 (O_1549,N_14527,N_14044);
nand UO_1550 (O_1550,N_10241,N_10602);
and UO_1551 (O_1551,N_14341,N_13683);
nand UO_1552 (O_1552,N_13926,N_12577);
nor UO_1553 (O_1553,N_11884,N_10932);
or UO_1554 (O_1554,N_10521,N_13106);
and UO_1555 (O_1555,N_11937,N_12488);
nand UO_1556 (O_1556,N_13363,N_11600);
nor UO_1557 (O_1557,N_13985,N_11836);
nor UO_1558 (O_1558,N_12744,N_14236);
nand UO_1559 (O_1559,N_12789,N_14049);
xnor UO_1560 (O_1560,N_14849,N_13302);
and UO_1561 (O_1561,N_11324,N_12291);
and UO_1562 (O_1562,N_11346,N_13388);
or UO_1563 (O_1563,N_13818,N_13879);
or UO_1564 (O_1564,N_14103,N_10263);
and UO_1565 (O_1565,N_12607,N_14345);
and UO_1566 (O_1566,N_13153,N_14310);
nor UO_1567 (O_1567,N_11233,N_14802);
and UO_1568 (O_1568,N_12381,N_14318);
xor UO_1569 (O_1569,N_10046,N_13443);
or UO_1570 (O_1570,N_14594,N_13758);
xor UO_1571 (O_1571,N_14113,N_13700);
nand UO_1572 (O_1572,N_12434,N_10700);
or UO_1573 (O_1573,N_12398,N_10077);
or UO_1574 (O_1574,N_13166,N_11716);
and UO_1575 (O_1575,N_12906,N_14806);
nor UO_1576 (O_1576,N_13430,N_14825);
nand UO_1577 (O_1577,N_10252,N_10093);
nand UO_1578 (O_1578,N_13564,N_10430);
or UO_1579 (O_1579,N_10809,N_14515);
or UO_1580 (O_1580,N_11783,N_12814);
nand UO_1581 (O_1581,N_11995,N_14599);
nand UO_1582 (O_1582,N_11603,N_11781);
nor UO_1583 (O_1583,N_12756,N_11450);
and UO_1584 (O_1584,N_11050,N_14365);
and UO_1585 (O_1585,N_11956,N_11583);
xor UO_1586 (O_1586,N_12421,N_14836);
xnor UO_1587 (O_1587,N_10243,N_13389);
and UO_1588 (O_1588,N_12721,N_13548);
nor UO_1589 (O_1589,N_13551,N_12361);
or UO_1590 (O_1590,N_13326,N_10437);
or UO_1591 (O_1591,N_13507,N_14425);
nand UO_1592 (O_1592,N_12967,N_14237);
xnor UO_1593 (O_1593,N_12875,N_10078);
nand UO_1594 (O_1594,N_13304,N_14609);
and UO_1595 (O_1595,N_13115,N_10525);
nor UO_1596 (O_1596,N_12961,N_14414);
and UO_1597 (O_1597,N_14830,N_13701);
or UO_1598 (O_1598,N_13580,N_12308);
or UO_1599 (O_1599,N_10034,N_10575);
or UO_1600 (O_1600,N_13892,N_12828);
or UO_1601 (O_1601,N_11073,N_10591);
nand UO_1602 (O_1602,N_11615,N_10914);
or UO_1603 (O_1603,N_11609,N_11118);
nor UO_1604 (O_1604,N_12674,N_12024);
and UO_1605 (O_1605,N_12420,N_10355);
or UO_1606 (O_1606,N_11052,N_10015);
nand UO_1607 (O_1607,N_10902,N_10246);
or UO_1608 (O_1608,N_14294,N_12335);
xor UO_1609 (O_1609,N_10549,N_13281);
nor UO_1610 (O_1610,N_10343,N_10466);
nor UO_1611 (O_1611,N_12006,N_12295);
xor UO_1612 (O_1612,N_12326,N_14840);
or UO_1613 (O_1613,N_10614,N_10053);
nor UO_1614 (O_1614,N_10282,N_13810);
xnor UO_1615 (O_1615,N_12503,N_12290);
nor UO_1616 (O_1616,N_11183,N_13723);
nor UO_1617 (O_1617,N_14750,N_12428);
nand UO_1618 (O_1618,N_11809,N_14490);
nor UO_1619 (O_1619,N_10941,N_11199);
nand UO_1620 (O_1620,N_10712,N_14019);
nor UO_1621 (O_1621,N_14626,N_11971);
xnor UO_1622 (O_1622,N_12324,N_11242);
nor UO_1623 (O_1623,N_11454,N_12688);
nand UO_1624 (O_1624,N_12277,N_10267);
nor UO_1625 (O_1625,N_12782,N_12513);
nor UO_1626 (O_1626,N_10137,N_14838);
xnor UO_1627 (O_1627,N_11303,N_13362);
nor UO_1628 (O_1628,N_11839,N_11849);
nor UO_1629 (O_1629,N_12699,N_11438);
xor UO_1630 (O_1630,N_12771,N_12416);
xnor UO_1631 (O_1631,N_10925,N_12383);
nand UO_1632 (O_1632,N_11508,N_12442);
and UO_1633 (O_1633,N_14518,N_11207);
nor UO_1634 (O_1634,N_13920,N_10817);
nor UO_1635 (O_1635,N_13128,N_14767);
nand UO_1636 (O_1636,N_11599,N_13335);
and UO_1637 (O_1637,N_10698,N_10724);
xor UO_1638 (O_1638,N_12338,N_11272);
xor UO_1639 (O_1639,N_14359,N_13140);
nor UO_1640 (O_1640,N_11243,N_13179);
xnor UO_1641 (O_1641,N_13253,N_10485);
nor UO_1642 (O_1642,N_10991,N_10408);
and UO_1643 (O_1643,N_14620,N_11107);
nand UO_1644 (O_1644,N_14861,N_10446);
nand UO_1645 (O_1645,N_13468,N_13690);
nor UO_1646 (O_1646,N_12672,N_12852);
xnor UO_1647 (O_1647,N_10822,N_11309);
or UO_1648 (O_1648,N_11273,N_14949);
nor UO_1649 (O_1649,N_11664,N_10212);
xor UO_1650 (O_1650,N_11485,N_13834);
nor UO_1651 (O_1651,N_11484,N_12401);
xor UO_1652 (O_1652,N_14608,N_13465);
xor UO_1653 (O_1653,N_14970,N_12560);
nand UO_1654 (O_1654,N_14934,N_10777);
xor UO_1655 (O_1655,N_13283,N_12520);
nor UO_1656 (O_1656,N_13718,N_10490);
nand UO_1657 (O_1657,N_13520,N_13217);
and UO_1658 (O_1658,N_12678,N_11792);
and UO_1659 (O_1659,N_14975,N_14042);
xnor UO_1660 (O_1660,N_14780,N_14317);
or UO_1661 (O_1661,N_14374,N_10445);
xor UO_1662 (O_1662,N_10242,N_12895);
nand UO_1663 (O_1663,N_11763,N_12078);
nand UO_1664 (O_1664,N_14939,N_11782);
xnor UO_1665 (O_1665,N_10950,N_13669);
nand UO_1666 (O_1666,N_10771,N_13445);
nor UO_1667 (O_1667,N_12620,N_12310);
or UO_1668 (O_1668,N_10849,N_14184);
nor UO_1669 (O_1669,N_11870,N_10887);
nand UO_1670 (O_1670,N_11367,N_12454);
or UO_1671 (O_1671,N_10758,N_10869);
or UO_1672 (O_1672,N_11619,N_12569);
xnor UO_1673 (O_1673,N_10862,N_10565);
nand UO_1674 (O_1674,N_12984,N_13293);
or UO_1675 (O_1675,N_12742,N_13637);
and UO_1676 (O_1676,N_12091,N_12152);
or UO_1677 (O_1677,N_13466,N_12402);
or UO_1678 (O_1678,N_12330,N_11974);
and UO_1679 (O_1679,N_12679,N_11927);
or UO_1680 (O_1680,N_14570,N_12130);
or UO_1681 (O_1681,N_13432,N_13821);
nor UO_1682 (O_1682,N_14683,N_12214);
nor UO_1683 (O_1683,N_14798,N_11405);
nand UO_1684 (O_1684,N_11161,N_11004);
and UO_1685 (O_1685,N_11727,N_10326);
or UO_1686 (O_1686,N_11634,N_14927);
nor UO_1687 (O_1687,N_12689,N_11104);
or UO_1688 (O_1688,N_13492,N_10577);
nand UO_1689 (O_1689,N_10873,N_10383);
nor UO_1690 (O_1690,N_12568,N_14946);
and UO_1691 (O_1691,N_11150,N_14090);
nand UO_1692 (O_1692,N_14483,N_12632);
nor UO_1693 (O_1693,N_11965,N_11616);
nor UO_1694 (O_1694,N_14348,N_14779);
and UO_1695 (O_1695,N_14349,N_11901);
and UO_1696 (O_1696,N_11501,N_13383);
nor UO_1697 (O_1697,N_13096,N_11516);
nand UO_1698 (O_1698,N_13976,N_13535);
nor UO_1699 (O_1699,N_10680,N_14866);
xor UO_1700 (O_1700,N_10337,N_11400);
nand UO_1701 (O_1701,N_13212,N_13651);
nand UO_1702 (O_1702,N_13449,N_14922);
nand UO_1703 (O_1703,N_11086,N_14633);
nand UO_1704 (O_1704,N_13627,N_13288);
or UO_1705 (O_1705,N_14925,N_13664);
nand UO_1706 (O_1706,N_14757,N_10392);
and UO_1707 (O_1707,N_14843,N_11374);
or UO_1708 (O_1708,N_10372,N_11796);
and UO_1709 (O_1709,N_12501,N_12098);
nand UO_1710 (O_1710,N_12451,N_12999);
or UO_1711 (O_1711,N_14316,N_10972);
xor UO_1712 (O_1712,N_10085,N_14600);
and UO_1713 (O_1713,N_12748,N_12473);
xnor UO_1714 (O_1714,N_11826,N_12997);
nand UO_1715 (O_1715,N_11343,N_12690);
xnor UO_1716 (O_1716,N_10086,N_14162);
nor UO_1717 (O_1717,N_10921,N_13053);
xor UO_1718 (O_1718,N_11219,N_10130);
xor UO_1719 (O_1719,N_12306,N_13595);
nor UO_1720 (O_1720,N_13104,N_13521);
xor UO_1721 (O_1721,N_11169,N_14134);
nor UO_1722 (O_1722,N_13276,N_10730);
or UO_1723 (O_1723,N_11110,N_11544);
or UO_1724 (O_1724,N_13314,N_12425);
or UO_1725 (O_1725,N_11639,N_13083);
nor UO_1726 (O_1726,N_13186,N_10984);
and UO_1727 (O_1727,N_13145,N_14400);
or UO_1728 (O_1728,N_12968,N_14619);
xnor UO_1729 (O_1729,N_11932,N_14787);
xnor UO_1730 (O_1730,N_10311,N_11227);
or UO_1731 (O_1731,N_13159,N_14627);
nand UO_1732 (O_1732,N_12769,N_14148);
xnor UO_1733 (O_1733,N_12339,N_10719);
or UO_1734 (O_1734,N_10633,N_11088);
xnor UO_1735 (O_1735,N_14240,N_11537);
nor UO_1736 (O_1736,N_14419,N_14963);
or UO_1737 (O_1737,N_12571,N_13241);
and UO_1738 (O_1738,N_13001,N_13242);
or UO_1739 (O_1739,N_12156,N_13192);
nor UO_1740 (O_1740,N_13923,N_12545);
or UO_1741 (O_1741,N_10728,N_11991);
nor UO_1742 (O_1742,N_14921,N_10572);
xor UO_1743 (O_1743,N_13350,N_11853);
and UO_1744 (O_1744,N_13665,N_14411);
or UO_1745 (O_1745,N_10528,N_14407);
and UO_1746 (O_1746,N_10444,N_14299);
and UO_1747 (O_1747,N_13857,N_12927);
and UO_1748 (O_1748,N_10118,N_14910);
nor UO_1749 (O_1749,N_14447,N_13837);
xor UO_1750 (O_1750,N_12125,N_13260);
and UO_1751 (O_1751,N_14812,N_14046);
or UO_1752 (O_1752,N_13401,N_14697);
or UO_1753 (O_1753,N_11063,N_11746);
or UO_1754 (O_1754,N_11189,N_13688);
nor UO_1755 (O_1755,N_12768,N_12394);
nand UO_1756 (O_1756,N_13245,N_12642);
nand UO_1757 (O_1757,N_11443,N_14213);
nor UO_1758 (O_1758,N_14839,N_12838);
or UO_1759 (O_1759,N_14816,N_10152);
nand UO_1760 (O_1760,N_10644,N_13135);
or UO_1761 (O_1761,N_11633,N_12694);
nand UO_1762 (O_1762,N_12870,N_11888);
xnor UO_1763 (O_1763,N_11180,N_10805);
or UO_1764 (O_1764,N_12102,N_10426);
nand UO_1765 (O_1765,N_10468,N_11878);
and UO_1766 (O_1766,N_13661,N_13029);
and UO_1767 (O_1767,N_11431,N_14584);
or UO_1768 (O_1768,N_13607,N_13358);
or UO_1769 (O_1769,N_14031,N_11152);
xor UO_1770 (O_1770,N_10976,N_12887);
and UO_1771 (O_1771,N_13069,N_12019);
nor UO_1772 (O_1772,N_10003,N_12248);
and UO_1773 (O_1773,N_14047,N_14736);
xor UO_1774 (O_1774,N_10590,N_14851);
or UO_1775 (O_1775,N_11487,N_13247);
nand UO_1776 (O_1776,N_12208,N_11197);
xnor UO_1777 (O_1777,N_10397,N_14532);
xnor UO_1778 (O_1778,N_10982,N_11029);
or UO_1779 (O_1779,N_11263,N_11847);
xor UO_1780 (O_1780,N_14100,N_12587);
or UO_1781 (O_1781,N_13072,N_10653);
and UO_1782 (O_1782,N_14109,N_12532);
and UO_1783 (O_1783,N_12260,N_11862);
xor UO_1784 (O_1784,N_13541,N_11136);
and UO_1785 (O_1785,N_12572,N_13594);
and UO_1786 (O_1786,N_10387,N_12737);
xnor UO_1787 (O_1787,N_10798,N_14263);
and UO_1788 (O_1788,N_13782,N_10959);
nand UO_1789 (O_1789,N_11453,N_11371);
and UO_1790 (O_1790,N_13572,N_14190);
or UO_1791 (O_1791,N_13347,N_12173);
or UO_1792 (O_1792,N_11398,N_12598);
nand UO_1793 (O_1793,N_14670,N_14906);
xnor UO_1794 (O_1794,N_10134,N_12905);
xor UO_1795 (O_1795,N_14696,N_12712);
xor UO_1796 (O_1796,N_10748,N_14180);
xor UO_1797 (O_1797,N_14284,N_10050);
and UO_1798 (O_1798,N_14211,N_11378);
nor UO_1799 (O_1799,N_14981,N_11613);
nand UO_1800 (O_1800,N_10018,N_13353);
or UO_1801 (O_1801,N_11257,N_10608);
xnor UO_1802 (O_1802,N_12494,N_12877);
nand UO_1803 (O_1803,N_12008,N_10111);
or UO_1804 (O_1804,N_12815,N_14725);
nor UO_1805 (O_1805,N_10081,N_12070);
and UO_1806 (O_1806,N_10960,N_12238);
or UO_1807 (O_1807,N_14574,N_12356);
or UO_1808 (O_1808,N_14728,N_12855);
nand UO_1809 (O_1809,N_10834,N_10128);
nor UO_1810 (O_1810,N_14489,N_14860);
nor UO_1811 (O_1811,N_14312,N_12810);
nand UO_1812 (O_1812,N_10648,N_14676);
or UO_1813 (O_1813,N_10203,N_11539);
nand UO_1814 (O_1814,N_12243,N_10839);
xnor UO_1815 (O_1815,N_11122,N_10924);
or UO_1816 (O_1816,N_11687,N_10664);
xnor UO_1817 (O_1817,N_11931,N_13173);
nand UO_1818 (O_1818,N_11744,N_10949);
nand UO_1819 (O_1819,N_14063,N_12487);
and UO_1820 (O_1820,N_11818,N_10142);
and UO_1821 (O_1821,N_11012,N_10952);
nand UO_1822 (O_1822,N_12730,N_13070);
nand UO_1823 (O_1823,N_13687,N_14858);
or UO_1824 (O_1824,N_12104,N_10917);
and UO_1825 (O_1825,N_10851,N_13674);
or UO_1826 (O_1826,N_11194,N_12007);
and UO_1827 (O_1827,N_11698,N_13555);
nand UO_1828 (O_1828,N_12300,N_11146);
nand UO_1829 (O_1829,N_14071,N_14035);
and UO_1830 (O_1830,N_10717,N_13028);
nand UO_1831 (O_1831,N_13000,N_10504);
nand UO_1832 (O_1832,N_14966,N_11988);
nor UO_1833 (O_1833,N_10176,N_11806);
nor UO_1834 (O_1834,N_13762,N_12504);
nor UO_1835 (O_1835,N_13433,N_12614);
nor UO_1836 (O_1836,N_13089,N_10747);
nor UO_1837 (O_1837,N_14573,N_14438);
or UO_1838 (O_1838,N_11202,N_14950);
nor UO_1839 (O_1839,N_14119,N_13421);
nand UO_1840 (O_1840,N_12050,N_11007);
and UO_1841 (O_1841,N_12073,N_11960);
nand UO_1842 (O_1842,N_11852,N_10323);
nor UO_1843 (O_1843,N_11566,N_13658);
nor UO_1844 (O_1844,N_11528,N_12735);
or UO_1845 (O_1845,N_11842,N_13273);
or UO_1846 (O_1846,N_11895,N_12477);
xnor UO_1847 (O_1847,N_10961,N_13850);
xor UO_1848 (O_1848,N_11775,N_13063);
or UO_1849 (O_1849,N_10794,N_12001);
nand UO_1850 (O_1850,N_11336,N_10253);
nor UO_1851 (O_1851,N_10784,N_14702);
nand UO_1852 (O_1852,N_14350,N_14054);
nand UO_1853 (O_1853,N_12045,N_11738);
and UO_1854 (O_1854,N_11294,N_11517);
nand UO_1855 (O_1855,N_13095,N_10578);
nor UO_1856 (O_1856,N_10292,N_12406);
xnor UO_1857 (O_1857,N_12116,N_10543);
or UO_1858 (O_1858,N_13773,N_12349);
nand UO_1859 (O_1859,N_12302,N_10136);
or UO_1860 (O_1860,N_11277,N_10313);
xnor UO_1861 (O_1861,N_13149,N_14519);
nand UO_1862 (O_1862,N_12812,N_13018);
xor UO_1863 (O_1863,N_11998,N_14495);
nand UO_1864 (O_1864,N_13198,N_12179);
xnor UO_1865 (O_1865,N_11560,N_13065);
xor UO_1866 (O_1866,N_11278,N_13911);
and UO_1867 (O_1867,N_12071,N_10317);
and UO_1868 (O_1868,N_14292,N_14781);
xnor UO_1869 (O_1869,N_14735,N_14487);
xor UO_1870 (O_1870,N_14715,N_14826);
or UO_1871 (O_1871,N_12177,N_13763);
xnor UO_1872 (O_1872,N_10722,N_13348);
xnor UO_1873 (O_1873,N_10793,N_11235);
or UO_1874 (O_1874,N_13345,N_10012);
or UO_1875 (O_1875,N_14990,N_10133);
nor UO_1876 (O_1876,N_14351,N_11390);
and UO_1877 (O_1877,N_14859,N_12100);
xnor UO_1878 (O_1878,N_12654,N_10820);
nand UO_1879 (O_1879,N_13586,N_11185);
or UO_1880 (O_1880,N_12264,N_14117);
and UO_1881 (O_1881,N_12914,N_12955);
or UO_1882 (O_1882,N_12960,N_12639);
or UO_1883 (O_1883,N_10857,N_14072);
nand UO_1884 (O_1884,N_12347,N_12591);
xnor UO_1885 (O_1885,N_14506,N_10301);
nand UO_1886 (O_1886,N_12124,N_13057);
xnor UO_1887 (O_1887,N_14940,N_12646);
xnor UO_1888 (O_1888,N_12745,N_10367);
xor UO_1889 (O_1889,N_10400,N_14948);
xor UO_1890 (O_1890,N_14307,N_11258);
xnor UO_1891 (O_1891,N_13529,N_12133);
nor UO_1892 (O_1892,N_12301,N_11113);
or UO_1893 (O_1893,N_14330,N_12304);
or UO_1894 (O_1894,N_12856,N_14746);
nor UO_1895 (O_1895,N_11614,N_13160);
nor UO_1896 (O_1896,N_12539,N_12199);
and UO_1897 (O_1897,N_13127,N_14710);
or UO_1898 (O_1898,N_10045,N_12909);
and UO_1899 (O_1899,N_14648,N_12190);
nor UO_1900 (O_1900,N_10563,N_12186);
nor UO_1901 (O_1901,N_12516,N_12747);
nand UO_1902 (O_1902,N_14852,N_13091);
xor UO_1903 (O_1903,N_12030,N_14334);
and UO_1904 (O_1904,N_14012,N_12065);
nand UO_1905 (O_1905,N_11881,N_12630);
and UO_1906 (O_1906,N_14793,N_10047);
nor UO_1907 (O_1907,N_12579,N_12954);
and UO_1908 (O_1908,N_13422,N_14652);
nand UO_1909 (O_1909,N_13959,N_10135);
or UO_1910 (O_1910,N_10240,N_11054);
xor UO_1911 (O_1911,N_13082,N_13906);
or UO_1912 (O_1912,N_10544,N_14384);
xor UO_1913 (O_1913,N_12035,N_12658);
and UO_1914 (O_1914,N_12172,N_14659);
nand UO_1915 (O_1915,N_12005,N_11130);
nor UO_1916 (O_1916,N_11535,N_11006);
or UO_1917 (O_1917,N_13704,N_13077);
xor UO_1918 (O_1918,N_12099,N_13204);
and UO_1919 (O_1919,N_14582,N_11989);
nor UO_1920 (O_1920,N_13221,N_11734);
and UO_1921 (O_1921,N_14592,N_13207);
nor UO_1922 (O_1922,N_14773,N_11787);
and UO_1923 (O_1923,N_14631,N_14625);
nand UO_1924 (O_1924,N_12867,N_10989);
nor UO_1925 (O_1925,N_10310,N_14581);
and UO_1926 (O_1926,N_12959,N_10835);
nand UO_1927 (O_1927,N_13554,N_12907);
nor UO_1928 (O_1928,N_10518,N_12727);
or UO_1929 (O_1929,N_10124,N_12044);
nand UO_1930 (O_1930,N_12526,N_10024);
and UO_1931 (O_1931,N_14871,N_12461);
and UO_1932 (O_1932,N_12235,N_13163);
nand UO_1933 (O_1933,N_10685,N_14467);
nor UO_1934 (O_1934,N_12446,N_12151);
or UO_1935 (O_1935,N_12800,N_11348);
or UO_1936 (O_1936,N_11789,N_14193);
or UO_1937 (O_1937,N_14870,N_12622);
or UO_1938 (O_1938,N_13798,N_12041);
nor UO_1939 (O_1939,N_12433,N_10800);
and UO_1940 (O_1940,N_10701,N_12803);
nand UO_1941 (O_1941,N_12143,N_10084);
xnor UO_1942 (O_1942,N_11436,N_12466);
or UO_1943 (O_1943,N_13137,N_11269);
xor UO_1944 (O_1944,N_14502,N_14729);
nand UO_1945 (O_1945,N_11408,N_14635);
nor UO_1946 (O_1946,N_12837,N_10175);
or UO_1947 (O_1947,N_10824,N_11253);
xor UO_1948 (O_1948,N_14681,N_10594);
or UO_1949 (O_1949,N_12129,N_11386);
or UO_1950 (O_1950,N_12864,N_14709);
and UO_1951 (O_1951,N_10148,N_11571);
nand UO_1952 (O_1952,N_13884,N_14192);
nor UO_1953 (O_1953,N_13429,N_12576);
nor UO_1954 (O_1954,N_12354,N_14058);
and UO_1955 (O_1955,N_11045,N_13896);
nor UO_1956 (O_1956,N_11828,N_12127);
nor UO_1957 (O_1957,N_13002,N_13165);
or UO_1958 (O_1958,N_11908,N_14730);
or UO_1959 (O_1959,N_13806,N_10439);
or UO_1960 (O_1960,N_12896,N_11275);
xnor UO_1961 (O_1961,N_11162,N_14737);
xor UO_1962 (O_1962,N_11703,N_11093);
xnor UO_1963 (O_1963,N_10846,N_10858);
xnor UO_1964 (O_1964,N_13618,N_10503);
nand UO_1965 (O_1965,N_12034,N_14481);
or UO_1966 (O_1966,N_14654,N_11171);
and UO_1967 (O_1967,N_14207,N_12287);
nand UO_1968 (O_1968,N_11814,N_11893);
or UO_1969 (O_1969,N_14394,N_10922);
nor UO_1970 (O_1970,N_14452,N_12340);
nor UO_1971 (O_1971,N_14335,N_13405);
nand UO_1972 (O_1972,N_12849,N_14732);
nand UO_1973 (O_1973,N_13931,N_10833);
nand UO_1974 (O_1974,N_13286,N_12930);
and UO_1975 (O_1975,N_10517,N_13829);
or UO_1976 (O_1976,N_13830,N_13264);
or UO_1977 (O_1977,N_11589,N_13504);
nor UO_1978 (O_1978,N_12250,N_14896);
nor UO_1979 (O_1979,N_11297,N_10811);
or UO_1980 (O_1980,N_14305,N_12827);
nor UO_1981 (O_1981,N_12651,N_13239);
xnor UO_1982 (O_1982,N_10244,N_12408);
or UO_1983 (O_1983,N_11477,N_13006);
xor UO_1984 (O_1984,N_10799,N_11179);
nor UO_1985 (O_1985,N_14097,N_13274);
or UO_1986 (O_1986,N_14897,N_10796);
xor UO_1987 (O_1987,N_12603,N_14128);
nand UO_1988 (O_1988,N_13229,N_14275);
xnor UO_1989 (O_1989,N_12935,N_11034);
nor UO_1990 (O_1990,N_13147,N_13901);
xor UO_1991 (O_1991,N_12036,N_13391);
nand UO_1992 (O_1992,N_14883,N_12621);
xnor UO_1993 (O_1993,N_13907,N_13813);
and UO_1994 (O_1994,N_11394,N_14876);
and UO_1995 (O_1995,N_13710,N_12202);
or UO_1996 (O_1996,N_13138,N_10068);
xor UO_1997 (O_1997,N_14095,N_12022);
nor UO_1998 (O_1998,N_11861,N_12963);
nor UO_1999 (O_1999,N_12677,N_14033);
endmodule