module basic_500_3000_500_15_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_332,In_197);
or U1 (N_1,In_135,In_394);
nand U2 (N_2,In_447,In_130);
and U3 (N_3,In_419,In_439);
nor U4 (N_4,In_106,In_281);
or U5 (N_5,In_466,In_349);
nor U6 (N_6,In_15,In_102);
nand U7 (N_7,In_23,In_198);
or U8 (N_8,In_423,In_443);
nand U9 (N_9,In_188,In_495);
or U10 (N_10,In_313,In_55);
nor U11 (N_11,In_403,In_206);
nand U12 (N_12,In_73,In_211);
nor U13 (N_13,In_382,In_243);
nand U14 (N_14,In_355,In_136);
nand U15 (N_15,In_484,In_167);
or U16 (N_16,In_263,In_255);
nor U17 (N_17,In_497,In_336);
nor U18 (N_18,In_462,In_290);
and U19 (N_19,In_125,In_318);
and U20 (N_20,In_45,In_414);
nor U21 (N_21,In_486,In_7);
and U22 (N_22,In_182,In_129);
and U23 (N_23,In_294,In_433);
or U24 (N_24,In_343,In_253);
or U25 (N_25,In_276,In_489);
nand U26 (N_26,In_221,In_444);
or U27 (N_27,In_446,In_227);
and U28 (N_28,In_464,In_63);
and U29 (N_29,In_87,In_226);
nand U30 (N_30,In_105,In_233);
or U31 (N_31,In_375,In_64);
and U32 (N_32,In_53,In_5);
or U33 (N_33,In_454,In_360);
or U34 (N_34,In_448,In_393);
nor U35 (N_35,In_289,In_149);
and U36 (N_36,In_97,In_66);
nand U37 (N_37,In_426,In_244);
or U38 (N_38,In_417,In_398);
nand U39 (N_39,In_117,In_401);
nand U40 (N_40,In_316,In_99);
nand U41 (N_41,In_101,In_264);
nor U42 (N_42,In_202,In_96);
nand U43 (N_43,In_242,In_492);
and U44 (N_44,In_100,In_111);
nor U45 (N_45,In_402,In_212);
and U46 (N_46,In_72,In_374);
nand U47 (N_47,In_71,In_147);
or U48 (N_48,In_388,In_164);
and U49 (N_49,In_474,In_119);
and U50 (N_50,In_452,In_341);
nand U51 (N_51,In_321,In_168);
or U52 (N_52,In_75,In_59);
nand U53 (N_53,In_399,In_249);
and U54 (N_54,In_293,In_335);
and U55 (N_55,In_68,In_225);
nor U56 (N_56,In_104,In_410);
nand U57 (N_57,In_421,In_425);
nand U58 (N_58,In_21,In_109);
nand U59 (N_59,In_488,In_257);
and U60 (N_60,In_9,In_422);
nand U61 (N_61,In_37,In_69);
or U62 (N_62,In_113,In_438);
or U63 (N_63,In_451,In_493);
xor U64 (N_64,In_62,In_481);
or U65 (N_65,In_77,In_286);
nand U66 (N_66,In_376,In_259);
or U67 (N_67,In_265,In_78);
or U68 (N_68,In_480,In_114);
nor U69 (N_69,In_17,In_261);
or U70 (N_70,In_159,In_371);
nor U71 (N_71,In_51,In_381);
nor U72 (N_72,In_163,In_347);
nand U73 (N_73,In_224,In_496);
or U74 (N_74,In_103,In_469);
and U75 (N_75,In_232,In_40);
and U76 (N_76,In_258,In_431);
nand U77 (N_77,In_120,In_282);
nor U78 (N_78,In_20,In_247);
nand U79 (N_79,In_358,In_161);
nor U80 (N_80,In_12,In_76);
nand U81 (N_81,In_95,In_187);
nor U82 (N_82,In_445,In_123);
nand U83 (N_83,In_373,In_179);
nand U84 (N_84,In_222,In_329);
nor U85 (N_85,In_334,In_262);
or U86 (N_86,In_86,In_141);
or U87 (N_87,In_256,In_396);
nor U88 (N_88,In_353,In_291);
and U89 (N_89,In_169,In_352);
nor U90 (N_90,In_178,In_116);
nor U91 (N_91,In_406,In_390);
nor U92 (N_92,In_298,In_144);
nor U93 (N_93,In_94,In_412);
and U94 (N_94,In_380,In_366);
nand U95 (N_95,In_81,In_440);
and U96 (N_96,In_326,In_342);
nand U97 (N_97,In_277,In_465);
and U98 (N_98,In_460,In_369);
nor U99 (N_99,In_171,In_311);
and U100 (N_100,In_42,In_296);
or U101 (N_101,In_333,In_67);
or U102 (N_102,In_453,In_237);
nor U103 (N_103,In_301,In_83);
and U104 (N_104,In_207,In_199);
and U105 (N_105,In_485,In_145);
nor U106 (N_106,In_209,In_300);
nand U107 (N_107,In_153,In_194);
or U108 (N_108,In_476,In_272);
and U109 (N_109,In_200,In_218);
nor U110 (N_110,In_6,In_35);
nor U111 (N_111,In_165,In_387);
and U112 (N_112,In_467,In_112);
or U113 (N_113,In_190,In_11);
and U114 (N_114,In_471,In_328);
and U115 (N_115,In_459,In_345);
xor U116 (N_116,In_362,In_499);
nor U117 (N_117,In_30,In_475);
or U118 (N_118,In_133,In_404);
or U119 (N_119,In_18,In_208);
nor U120 (N_120,In_395,In_43);
and U121 (N_121,In_49,In_266);
or U122 (N_122,In_430,In_148);
nor U123 (N_123,In_191,In_82);
or U124 (N_124,In_304,In_154);
and U125 (N_125,In_93,In_463);
nand U126 (N_126,In_241,In_47);
and U127 (N_127,In_240,In_160);
or U128 (N_128,In_46,In_456);
nor U129 (N_129,In_434,In_418);
or U130 (N_130,In_437,In_274);
nand U131 (N_131,In_391,In_379);
nand U132 (N_132,In_204,In_140);
or U133 (N_133,In_91,In_107);
nand U134 (N_134,In_323,In_340);
and U135 (N_135,In_288,In_359);
nand U136 (N_136,In_70,In_48);
and U137 (N_137,In_121,In_108);
nand U138 (N_138,In_386,In_56);
nand U139 (N_139,In_442,In_384);
nor U140 (N_140,In_213,In_473);
and U141 (N_141,In_248,In_432);
or U142 (N_142,In_468,In_477);
and U143 (N_143,In_24,In_201);
or U144 (N_144,In_483,In_142);
xor U145 (N_145,In_220,In_184);
nand U146 (N_146,In_383,In_348);
or U147 (N_147,In_429,In_65);
nand U148 (N_148,In_405,In_315);
or U149 (N_149,In_155,In_354);
nand U150 (N_150,In_268,In_230);
or U151 (N_151,In_312,In_181);
and U152 (N_152,In_314,In_238);
or U153 (N_153,In_41,In_90);
nor U154 (N_154,In_88,In_118);
or U155 (N_155,In_357,In_267);
nor U156 (N_156,In_458,In_368);
or U157 (N_157,In_4,In_28);
and U158 (N_158,In_435,In_472);
nor U159 (N_159,In_32,In_193);
and U160 (N_160,In_205,In_292);
and U161 (N_161,In_372,In_303);
and U162 (N_162,In_494,In_305);
and U163 (N_163,In_151,In_415);
or U164 (N_164,In_370,In_210);
and U165 (N_165,In_498,In_400);
or U166 (N_166,In_344,In_52);
nor U167 (N_167,In_175,In_223);
and U168 (N_168,In_339,In_307);
nand U169 (N_169,In_356,In_351);
nand U170 (N_170,In_306,In_14);
nor U171 (N_171,In_367,In_13);
or U172 (N_172,In_350,In_16);
or U173 (N_173,In_162,In_215);
and U174 (N_174,In_457,In_0);
and U175 (N_175,In_441,In_424);
or U176 (N_176,In_31,In_166);
nor U177 (N_177,In_57,In_278);
or U178 (N_178,In_299,In_309);
nor U179 (N_179,In_363,In_150);
and U180 (N_180,In_110,In_411);
and U181 (N_181,In_10,In_269);
nor U182 (N_182,In_127,In_58);
or U183 (N_183,In_25,In_216);
or U184 (N_184,In_479,In_377);
nand U185 (N_185,In_38,In_490);
or U186 (N_186,In_491,In_280);
and U187 (N_187,In_214,In_128);
nor U188 (N_188,In_361,In_337);
nand U189 (N_189,In_33,In_324);
nand U190 (N_190,In_170,In_39);
nor U191 (N_191,In_196,In_34);
nand U192 (N_192,In_392,In_29);
nor U193 (N_193,In_177,In_285);
or U194 (N_194,In_420,In_60);
and U195 (N_195,In_450,In_310);
or U196 (N_196,In_260,In_449);
or U197 (N_197,In_79,In_320);
or U198 (N_198,In_364,In_436);
nor U199 (N_199,In_176,In_461);
nand U200 (N_200,N_85,In_22);
and U201 (N_201,N_65,In_252);
or U202 (N_202,In_19,N_114);
nand U203 (N_203,In_134,N_53);
nand U204 (N_204,N_88,In_254);
or U205 (N_205,In_283,In_158);
nand U206 (N_206,N_72,N_48);
nor U207 (N_207,N_70,N_138);
or U208 (N_208,N_142,N_59);
nand U209 (N_209,In_287,In_346);
nand U210 (N_210,In_251,N_165);
xnor U211 (N_211,In_327,N_144);
nand U212 (N_212,N_29,N_185);
nor U213 (N_213,N_160,N_135);
nor U214 (N_214,In_186,N_179);
or U215 (N_215,N_153,N_116);
nand U216 (N_216,N_1,In_229);
or U217 (N_217,In_54,In_409);
nand U218 (N_218,N_7,N_36);
nand U219 (N_219,In_131,In_397);
and U220 (N_220,N_118,N_181);
nor U221 (N_221,N_171,N_63);
or U222 (N_222,N_75,In_156);
or U223 (N_223,N_126,N_146);
nand U224 (N_224,N_134,N_25);
nand U225 (N_225,N_52,N_6);
nand U226 (N_226,In_234,N_77);
and U227 (N_227,N_189,In_389);
nor U228 (N_228,N_166,N_109);
or U229 (N_229,In_407,N_95);
nand U230 (N_230,N_168,In_239);
nand U231 (N_231,N_129,In_44);
and U232 (N_232,N_123,N_12);
or U233 (N_233,In_317,N_92);
nand U234 (N_234,N_190,N_67);
or U235 (N_235,N_32,N_84);
or U236 (N_236,N_55,N_151);
or U237 (N_237,In_478,In_115);
xor U238 (N_238,In_192,N_128);
nand U239 (N_239,N_73,N_45);
and U240 (N_240,N_4,In_3);
nand U241 (N_241,N_58,N_161);
nand U242 (N_242,N_30,In_143);
and U243 (N_243,N_16,In_246);
or U244 (N_244,N_89,In_1);
nand U245 (N_245,N_5,N_40);
or U246 (N_246,In_330,In_183);
or U247 (N_247,N_9,In_180);
or U248 (N_248,N_164,N_94);
and U249 (N_249,N_149,N_19);
nand U250 (N_250,N_197,N_132);
or U251 (N_251,N_103,N_112);
nor U252 (N_252,In_219,N_157);
nand U253 (N_253,N_91,N_80);
and U254 (N_254,In_195,N_131);
or U255 (N_255,N_97,In_416);
nand U256 (N_256,N_120,N_17);
or U257 (N_257,N_76,N_83);
and U258 (N_258,N_121,In_139);
nand U259 (N_259,N_56,N_162);
nand U260 (N_260,In_231,N_198);
or U261 (N_261,In_487,N_35);
nor U262 (N_262,In_27,N_98);
and U263 (N_263,N_154,In_245);
or U264 (N_264,In_235,N_108);
nor U265 (N_265,N_196,In_284);
or U266 (N_266,In_61,N_159);
and U267 (N_267,In_8,N_148);
nand U268 (N_268,N_145,N_199);
nand U269 (N_269,N_195,In_74);
or U270 (N_270,In_295,N_133);
nand U271 (N_271,In_378,N_51);
nor U272 (N_272,N_106,N_158);
or U273 (N_273,N_170,N_10);
nand U274 (N_274,N_42,N_104);
or U275 (N_275,In_385,In_122);
nor U276 (N_276,In_172,N_127);
nand U277 (N_277,N_175,N_79);
or U278 (N_278,In_455,N_100);
and U279 (N_279,N_41,N_172);
nor U280 (N_280,N_2,N_44);
or U281 (N_281,In_482,N_82);
nand U282 (N_282,N_62,N_46);
and U283 (N_283,In_308,N_74);
nor U284 (N_284,N_174,In_126);
and U285 (N_285,N_81,N_22);
nand U286 (N_286,N_143,N_191);
or U287 (N_287,In_470,N_3);
nor U288 (N_288,In_325,In_185);
and U289 (N_289,In_273,In_174);
nor U290 (N_290,N_130,N_28);
and U291 (N_291,N_173,N_13);
and U292 (N_292,In_279,N_34);
or U293 (N_293,N_194,N_136);
and U294 (N_294,In_297,N_90);
or U295 (N_295,N_139,In_275);
nor U296 (N_296,N_93,N_0);
or U297 (N_297,In_236,N_21);
nor U298 (N_298,N_61,N_122);
nand U299 (N_299,N_8,N_37);
nand U300 (N_300,In_157,N_50);
xor U301 (N_301,N_107,N_105);
nor U302 (N_302,In_124,N_193);
nor U303 (N_303,N_57,In_132);
nor U304 (N_304,N_113,In_408);
or U305 (N_305,In_85,N_167);
and U306 (N_306,N_54,N_169);
and U307 (N_307,N_176,In_26);
nor U308 (N_308,In_146,N_125);
nor U309 (N_309,N_119,In_365);
or U310 (N_310,N_69,N_124);
or U311 (N_311,N_47,N_26);
nor U312 (N_312,N_99,N_60);
and U313 (N_313,In_92,In_138);
and U314 (N_314,N_184,N_102);
nand U315 (N_315,N_15,In_250);
or U316 (N_316,In_270,N_20);
and U317 (N_317,N_68,N_111);
and U318 (N_318,N_180,In_80);
nand U319 (N_319,In_98,N_43);
nor U320 (N_320,N_86,In_84);
or U321 (N_321,In_331,N_96);
and U322 (N_322,N_31,In_322);
nand U323 (N_323,N_39,In_228);
nor U324 (N_324,N_110,N_152);
or U325 (N_325,N_192,In_217);
nand U326 (N_326,In_271,N_117);
nand U327 (N_327,In_319,N_156);
and U328 (N_328,N_64,N_101);
and U329 (N_329,In_427,In_413);
nor U330 (N_330,In_302,In_189);
nand U331 (N_331,In_173,N_163);
xnor U332 (N_332,N_14,N_49);
or U333 (N_333,N_155,N_78);
and U334 (N_334,In_203,N_137);
nand U335 (N_335,N_38,In_137);
nor U336 (N_336,N_182,N_187);
nand U337 (N_337,N_115,N_140);
or U338 (N_338,In_36,N_188);
or U339 (N_339,In_89,N_27);
or U340 (N_340,N_147,In_338);
nand U341 (N_341,N_178,N_33);
nor U342 (N_342,N_23,N_87);
nand U343 (N_343,In_428,N_66);
or U344 (N_344,In_2,N_71);
nand U345 (N_345,In_50,N_183);
nor U346 (N_346,In_152,N_18);
nand U347 (N_347,N_186,N_24);
xnor U348 (N_348,N_141,N_150);
and U349 (N_349,N_177,N_11);
nand U350 (N_350,N_12,N_177);
nand U351 (N_351,In_322,In_234);
nor U352 (N_352,In_84,N_19);
nor U353 (N_353,In_413,In_137);
nand U354 (N_354,N_129,In_245);
and U355 (N_355,N_8,In_416);
or U356 (N_356,N_32,N_164);
nand U357 (N_357,N_92,N_5);
and U358 (N_358,N_58,N_167);
or U359 (N_359,In_44,N_6);
nor U360 (N_360,In_157,In_98);
nor U361 (N_361,N_151,In_8);
and U362 (N_362,In_322,In_378);
or U363 (N_363,In_455,N_175);
nor U364 (N_364,N_196,N_91);
and U365 (N_365,N_89,N_168);
and U366 (N_366,In_180,In_74);
nor U367 (N_367,N_65,N_190);
nand U368 (N_368,N_98,N_31);
or U369 (N_369,In_235,N_151);
nor U370 (N_370,N_116,N_50);
nand U371 (N_371,In_44,In_80);
and U372 (N_372,N_114,In_413);
and U373 (N_373,N_112,N_56);
nand U374 (N_374,N_197,N_140);
or U375 (N_375,N_160,N_90);
nor U376 (N_376,N_142,N_114);
and U377 (N_377,N_60,N_50);
nand U378 (N_378,N_193,N_75);
nor U379 (N_379,In_254,N_4);
nor U380 (N_380,N_111,N_66);
nor U381 (N_381,N_74,N_14);
nand U382 (N_382,In_455,In_235);
nand U383 (N_383,N_192,N_94);
or U384 (N_384,N_65,N_81);
nand U385 (N_385,N_37,In_427);
xnor U386 (N_386,N_1,N_32);
nand U387 (N_387,In_273,In_228);
nor U388 (N_388,N_20,N_120);
nor U389 (N_389,In_139,N_95);
or U390 (N_390,N_73,N_180);
nand U391 (N_391,In_409,In_185);
or U392 (N_392,N_176,N_181);
nor U393 (N_393,N_60,In_385);
or U394 (N_394,N_126,In_428);
nor U395 (N_395,N_30,N_120);
and U396 (N_396,In_124,N_20);
or U397 (N_397,N_41,N_139);
nor U398 (N_398,N_191,N_145);
or U399 (N_399,In_61,In_180);
and U400 (N_400,N_374,N_215);
nand U401 (N_401,N_366,N_247);
nand U402 (N_402,N_240,N_267);
and U403 (N_403,N_370,N_228);
nand U404 (N_404,N_233,N_386);
or U405 (N_405,N_363,N_308);
or U406 (N_406,N_229,N_316);
nor U407 (N_407,N_383,N_312);
xnor U408 (N_408,N_270,N_382);
nor U409 (N_409,N_379,N_209);
nand U410 (N_410,N_389,N_290);
nand U411 (N_411,N_277,N_265);
nand U412 (N_412,N_221,N_348);
or U413 (N_413,N_291,N_395);
or U414 (N_414,N_361,N_331);
nand U415 (N_415,N_202,N_318);
nand U416 (N_416,N_253,N_293);
and U417 (N_417,N_230,N_214);
or U418 (N_418,N_213,N_394);
nor U419 (N_419,N_268,N_239);
nand U420 (N_420,N_231,N_281);
nor U421 (N_421,N_325,N_345);
nand U422 (N_422,N_241,N_332);
nor U423 (N_423,N_393,N_340);
and U424 (N_424,N_355,N_380);
nand U425 (N_425,N_310,N_372);
and U426 (N_426,N_269,N_203);
nand U427 (N_427,N_341,N_257);
nand U428 (N_428,N_222,N_200);
nand U429 (N_429,N_208,N_384);
nand U430 (N_430,N_349,N_245);
nand U431 (N_431,N_242,N_304);
nand U432 (N_432,N_365,N_398);
or U433 (N_433,N_210,N_359);
and U434 (N_434,N_299,N_309);
nand U435 (N_435,N_252,N_217);
nand U436 (N_436,N_360,N_313);
nor U437 (N_437,N_298,N_212);
nor U438 (N_438,N_323,N_235);
nand U439 (N_439,N_258,N_224);
or U440 (N_440,N_385,N_282);
nor U441 (N_441,N_305,N_362);
and U442 (N_442,N_338,N_296);
and U443 (N_443,N_333,N_324);
or U444 (N_444,N_292,N_356);
and U445 (N_445,N_289,N_330);
nand U446 (N_446,N_220,N_250);
nor U447 (N_447,N_278,N_314);
nand U448 (N_448,N_205,N_223);
or U449 (N_449,N_399,N_378);
nor U450 (N_450,N_300,N_227);
xor U451 (N_451,N_396,N_339);
or U452 (N_452,N_315,N_284);
and U453 (N_453,N_322,N_280);
nand U454 (N_454,N_216,N_263);
nand U455 (N_455,N_327,N_354);
nand U456 (N_456,N_367,N_294);
or U457 (N_457,N_364,N_259);
nor U458 (N_458,N_352,N_271);
nor U459 (N_459,N_273,N_243);
and U460 (N_460,N_343,N_285);
nor U461 (N_461,N_204,N_306);
nand U462 (N_462,N_369,N_201);
xnor U463 (N_463,N_387,N_336);
or U464 (N_464,N_353,N_328);
nor U465 (N_465,N_207,N_254);
nor U466 (N_466,N_334,N_218);
nand U467 (N_467,N_237,N_264);
nand U468 (N_468,N_274,N_329);
or U469 (N_469,N_236,N_342);
nor U470 (N_470,N_392,N_260);
nor U471 (N_471,N_219,N_373);
nor U472 (N_472,N_286,N_307);
nor U473 (N_473,N_319,N_301);
and U474 (N_474,N_283,N_251);
or U475 (N_475,N_261,N_266);
nor U476 (N_476,N_232,N_248);
nand U477 (N_477,N_344,N_377);
nand U478 (N_478,N_287,N_226);
nor U479 (N_479,N_255,N_238);
nor U480 (N_480,N_371,N_311);
nand U481 (N_481,N_297,N_279);
nor U482 (N_482,N_276,N_256);
and U483 (N_483,N_244,N_295);
nand U484 (N_484,N_390,N_346);
nor U485 (N_485,N_375,N_376);
nor U486 (N_486,N_326,N_368);
or U487 (N_487,N_302,N_351);
nor U488 (N_488,N_317,N_275);
nor U489 (N_489,N_272,N_288);
nand U490 (N_490,N_225,N_321);
nand U491 (N_491,N_303,N_350);
or U492 (N_492,N_206,N_337);
nor U493 (N_493,N_211,N_391);
nand U494 (N_494,N_335,N_347);
nor U495 (N_495,N_262,N_234);
and U496 (N_496,N_357,N_388);
or U497 (N_497,N_381,N_320);
nand U498 (N_498,N_358,N_397);
and U499 (N_499,N_246,N_249);
or U500 (N_500,N_394,N_226);
nand U501 (N_501,N_256,N_265);
nand U502 (N_502,N_236,N_248);
nor U503 (N_503,N_309,N_358);
and U504 (N_504,N_222,N_305);
nor U505 (N_505,N_244,N_207);
nand U506 (N_506,N_303,N_290);
and U507 (N_507,N_349,N_221);
and U508 (N_508,N_348,N_212);
nand U509 (N_509,N_393,N_253);
nor U510 (N_510,N_216,N_376);
nand U511 (N_511,N_392,N_253);
and U512 (N_512,N_275,N_319);
nor U513 (N_513,N_363,N_248);
or U514 (N_514,N_278,N_312);
or U515 (N_515,N_206,N_324);
and U516 (N_516,N_257,N_275);
and U517 (N_517,N_355,N_265);
and U518 (N_518,N_344,N_353);
or U519 (N_519,N_200,N_226);
nand U520 (N_520,N_280,N_333);
nor U521 (N_521,N_378,N_204);
or U522 (N_522,N_343,N_379);
nand U523 (N_523,N_362,N_342);
nor U524 (N_524,N_228,N_232);
nand U525 (N_525,N_391,N_217);
and U526 (N_526,N_364,N_277);
nor U527 (N_527,N_327,N_225);
and U528 (N_528,N_382,N_348);
or U529 (N_529,N_291,N_230);
nor U530 (N_530,N_330,N_234);
and U531 (N_531,N_329,N_315);
or U532 (N_532,N_272,N_205);
and U533 (N_533,N_246,N_363);
and U534 (N_534,N_256,N_285);
nor U535 (N_535,N_269,N_354);
or U536 (N_536,N_203,N_274);
nor U537 (N_537,N_251,N_200);
nor U538 (N_538,N_323,N_321);
or U539 (N_539,N_328,N_373);
nor U540 (N_540,N_300,N_361);
nand U541 (N_541,N_262,N_220);
and U542 (N_542,N_398,N_372);
and U543 (N_543,N_325,N_253);
nand U544 (N_544,N_378,N_265);
or U545 (N_545,N_355,N_244);
and U546 (N_546,N_329,N_398);
nand U547 (N_547,N_397,N_249);
or U548 (N_548,N_219,N_286);
or U549 (N_549,N_279,N_250);
or U550 (N_550,N_359,N_228);
and U551 (N_551,N_351,N_342);
nor U552 (N_552,N_327,N_214);
and U553 (N_553,N_255,N_371);
nor U554 (N_554,N_285,N_293);
nor U555 (N_555,N_304,N_206);
nand U556 (N_556,N_327,N_341);
and U557 (N_557,N_227,N_333);
or U558 (N_558,N_360,N_300);
and U559 (N_559,N_266,N_299);
nor U560 (N_560,N_234,N_200);
nand U561 (N_561,N_375,N_342);
nor U562 (N_562,N_367,N_316);
and U563 (N_563,N_299,N_350);
nor U564 (N_564,N_313,N_222);
and U565 (N_565,N_285,N_284);
or U566 (N_566,N_216,N_357);
nand U567 (N_567,N_360,N_386);
nor U568 (N_568,N_201,N_254);
and U569 (N_569,N_294,N_334);
or U570 (N_570,N_314,N_321);
nand U571 (N_571,N_287,N_332);
nand U572 (N_572,N_362,N_368);
and U573 (N_573,N_301,N_210);
nand U574 (N_574,N_367,N_392);
or U575 (N_575,N_297,N_264);
nor U576 (N_576,N_213,N_305);
nor U577 (N_577,N_238,N_383);
nand U578 (N_578,N_337,N_284);
and U579 (N_579,N_338,N_382);
or U580 (N_580,N_205,N_243);
nand U581 (N_581,N_303,N_358);
nand U582 (N_582,N_232,N_237);
nand U583 (N_583,N_201,N_284);
nand U584 (N_584,N_251,N_214);
or U585 (N_585,N_221,N_227);
xor U586 (N_586,N_210,N_221);
and U587 (N_587,N_265,N_328);
nor U588 (N_588,N_340,N_286);
nor U589 (N_589,N_241,N_292);
and U590 (N_590,N_282,N_212);
and U591 (N_591,N_389,N_272);
and U592 (N_592,N_379,N_204);
or U593 (N_593,N_322,N_387);
nand U594 (N_594,N_344,N_294);
or U595 (N_595,N_371,N_329);
and U596 (N_596,N_396,N_398);
and U597 (N_597,N_332,N_229);
and U598 (N_598,N_241,N_317);
or U599 (N_599,N_319,N_270);
or U600 (N_600,N_554,N_400);
or U601 (N_601,N_530,N_503);
nand U602 (N_602,N_517,N_402);
nor U603 (N_603,N_483,N_599);
or U604 (N_604,N_509,N_588);
nor U605 (N_605,N_424,N_591);
nor U606 (N_606,N_597,N_521);
and U607 (N_607,N_555,N_584);
nor U608 (N_608,N_566,N_516);
or U609 (N_609,N_482,N_570);
nand U610 (N_610,N_439,N_539);
nand U611 (N_611,N_568,N_518);
or U612 (N_612,N_438,N_550);
nor U613 (N_613,N_575,N_500);
and U614 (N_614,N_479,N_593);
nor U615 (N_615,N_468,N_458);
and U616 (N_616,N_450,N_556);
nor U617 (N_617,N_589,N_508);
and U618 (N_618,N_443,N_525);
or U619 (N_619,N_466,N_401);
nand U620 (N_620,N_552,N_463);
or U621 (N_621,N_428,N_426);
nor U622 (N_622,N_414,N_563);
nand U623 (N_623,N_523,N_418);
nor U624 (N_624,N_553,N_551);
or U625 (N_625,N_411,N_471);
nand U626 (N_626,N_557,N_486);
or U627 (N_627,N_491,N_538);
nor U628 (N_628,N_582,N_461);
nor U629 (N_629,N_453,N_452);
or U630 (N_630,N_487,N_449);
nand U631 (N_631,N_595,N_583);
or U632 (N_632,N_533,N_545);
or U633 (N_633,N_574,N_501);
and U634 (N_634,N_544,N_534);
or U635 (N_635,N_577,N_592);
and U636 (N_636,N_416,N_474);
or U637 (N_637,N_447,N_524);
or U638 (N_638,N_565,N_511);
nand U639 (N_639,N_576,N_484);
nor U640 (N_640,N_560,N_526);
nor U641 (N_641,N_430,N_493);
or U642 (N_642,N_531,N_462);
xor U643 (N_643,N_548,N_497);
nand U644 (N_644,N_489,N_448);
nand U645 (N_645,N_422,N_569);
nor U646 (N_646,N_454,N_480);
and U647 (N_647,N_413,N_561);
nor U648 (N_648,N_433,N_481);
nand U649 (N_649,N_455,N_415);
nor U650 (N_650,N_547,N_507);
nor U651 (N_651,N_512,N_571);
nand U652 (N_652,N_535,N_440);
and U653 (N_653,N_578,N_549);
or U654 (N_654,N_485,N_496);
nor U655 (N_655,N_543,N_436);
or U656 (N_656,N_540,N_541);
nand U657 (N_657,N_510,N_409);
nor U658 (N_658,N_514,N_594);
or U659 (N_659,N_457,N_558);
nor U660 (N_660,N_598,N_567);
or U661 (N_661,N_527,N_506);
nand U662 (N_662,N_442,N_513);
or U663 (N_663,N_412,N_590);
and U664 (N_664,N_580,N_498);
or U665 (N_665,N_403,N_532);
nor U666 (N_666,N_579,N_407);
and U667 (N_667,N_420,N_417);
nor U668 (N_668,N_460,N_476);
nor U669 (N_669,N_446,N_528);
nand U670 (N_670,N_419,N_515);
nand U671 (N_671,N_475,N_562);
and U672 (N_672,N_410,N_519);
nor U673 (N_673,N_444,N_441);
and U674 (N_674,N_472,N_451);
nor U675 (N_675,N_477,N_505);
and U676 (N_676,N_459,N_502);
and U677 (N_677,N_542,N_469);
nand U678 (N_678,N_536,N_470);
nor U679 (N_679,N_573,N_437);
and U680 (N_680,N_596,N_456);
nand U681 (N_681,N_435,N_408);
and U682 (N_682,N_564,N_490);
and U683 (N_683,N_445,N_429);
and U684 (N_684,N_587,N_405);
nor U685 (N_685,N_529,N_478);
nor U686 (N_686,N_520,N_432);
nand U687 (N_687,N_546,N_434);
and U688 (N_688,N_406,N_499);
or U689 (N_689,N_495,N_473);
and U690 (N_690,N_504,N_464);
nand U691 (N_691,N_421,N_425);
and U692 (N_692,N_586,N_467);
nor U693 (N_693,N_537,N_465);
or U694 (N_694,N_494,N_404);
nand U695 (N_695,N_581,N_423);
nor U696 (N_696,N_559,N_427);
nor U697 (N_697,N_572,N_492);
nand U698 (N_698,N_431,N_488);
and U699 (N_699,N_585,N_522);
or U700 (N_700,N_485,N_483);
nand U701 (N_701,N_557,N_474);
nor U702 (N_702,N_487,N_471);
or U703 (N_703,N_435,N_559);
and U704 (N_704,N_409,N_516);
nor U705 (N_705,N_519,N_440);
nor U706 (N_706,N_499,N_561);
and U707 (N_707,N_494,N_471);
nand U708 (N_708,N_475,N_434);
and U709 (N_709,N_439,N_533);
nand U710 (N_710,N_490,N_505);
and U711 (N_711,N_537,N_596);
nor U712 (N_712,N_548,N_550);
and U713 (N_713,N_411,N_564);
or U714 (N_714,N_490,N_556);
nor U715 (N_715,N_430,N_593);
or U716 (N_716,N_424,N_442);
or U717 (N_717,N_464,N_443);
nand U718 (N_718,N_482,N_496);
nand U719 (N_719,N_562,N_494);
nor U720 (N_720,N_507,N_599);
nand U721 (N_721,N_465,N_478);
nor U722 (N_722,N_536,N_505);
nand U723 (N_723,N_415,N_542);
or U724 (N_724,N_407,N_503);
and U725 (N_725,N_478,N_410);
and U726 (N_726,N_461,N_408);
nand U727 (N_727,N_528,N_539);
nor U728 (N_728,N_418,N_479);
and U729 (N_729,N_598,N_594);
and U730 (N_730,N_449,N_403);
nor U731 (N_731,N_527,N_583);
or U732 (N_732,N_578,N_572);
nor U733 (N_733,N_412,N_456);
nor U734 (N_734,N_551,N_447);
nand U735 (N_735,N_559,N_500);
or U736 (N_736,N_462,N_459);
and U737 (N_737,N_476,N_440);
or U738 (N_738,N_575,N_477);
nor U739 (N_739,N_407,N_596);
nand U740 (N_740,N_537,N_529);
nand U741 (N_741,N_485,N_428);
nand U742 (N_742,N_416,N_427);
nor U743 (N_743,N_596,N_415);
nor U744 (N_744,N_580,N_522);
and U745 (N_745,N_522,N_553);
and U746 (N_746,N_592,N_572);
and U747 (N_747,N_504,N_446);
xnor U748 (N_748,N_510,N_436);
or U749 (N_749,N_585,N_537);
and U750 (N_750,N_482,N_565);
nor U751 (N_751,N_523,N_410);
nand U752 (N_752,N_509,N_458);
or U753 (N_753,N_489,N_521);
or U754 (N_754,N_554,N_478);
nand U755 (N_755,N_418,N_540);
nor U756 (N_756,N_489,N_403);
and U757 (N_757,N_423,N_431);
nor U758 (N_758,N_535,N_515);
and U759 (N_759,N_573,N_568);
nor U760 (N_760,N_530,N_577);
nor U761 (N_761,N_484,N_518);
or U762 (N_762,N_547,N_541);
nand U763 (N_763,N_553,N_427);
or U764 (N_764,N_593,N_444);
and U765 (N_765,N_535,N_405);
or U766 (N_766,N_471,N_406);
nor U767 (N_767,N_553,N_406);
and U768 (N_768,N_535,N_517);
or U769 (N_769,N_599,N_575);
nor U770 (N_770,N_487,N_470);
or U771 (N_771,N_584,N_498);
or U772 (N_772,N_552,N_521);
nand U773 (N_773,N_457,N_577);
nor U774 (N_774,N_403,N_408);
and U775 (N_775,N_400,N_471);
nand U776 (N_776,N_544,N_553);
nand U777 (N_777,N_597,N_594);
or U778 (N_778,N_413,N_522);
nand U779 (N_779,N_511,N_475);
or U780 (N_780,N_513,N_521);
or U781 (N_781,N_451,N_522);
nor U782 (N_782,N_439,N_586);
and U783 (N_783,N_531,N_496);
or U784 (N_784,N_443,N_569);
or U785 (N_785,N_574,N_505);
nor U786 (N_786,N_406,N_493);
and U787 (N_787,N_537,N_579);
xor U788 (N_788,N_455,N_432);
or U789 (N_789,N_553,N_410);
or U790 (N_790,N_413,N_487);
nand U791 (N_791,N_519,N_514);
nor U792 (N_792,N_538,N_550);
and U793 (N_793,N_525,N_528);
nor U794 (N_794,N_442,N_485);
and U795 (N_795,N_442,N_478);
nor U796 (N_796,N_441,N_439);
and U797 (N_797,N_448,N_505);
or U798 (N_798,N_546,N_549);
or U799 (N_799,N_492,N_441);
nor U800 (N_800,N_608,N_771);
nand U801 (N_801,N_690,N_756);
and U802 (N_802,N_793,N_719);
and U803 (N_803,N_634,N_665);
nand U804 (N_804,N_692,N_680);
and U805 (N_805,N_654,N_648);
nor U806 (N_806,N_704,N_782);
and U807 (N_807,N_770,N_701);
nor U808 (N_808,N_600,N_739);
nand U809 (N_809,N_722,N_682);
or U810 (N_810,N_645,N_610);
nand U811 (N_811,N_711,N_699);
nor U812 (N_812,N_751,N_688);
and U813 (N_813,N_742,N_700);
and U814 (N_814,N_694,N_785);
or U815 (N_815,N_725,N_633);
and U816 (N_816,N_732,N_681);
or U817 (N_817,N_664,N_728);
nand U818 (N_818,N_629,N_741);
nand U819 (N_819,N_609,N_638);
or U820 (N_820,N_754,N_765);
and U821 (N_821,N_768,N_602);
and U822 (N_822,N_729,N_651);
nor U823 (N_823,N_677,N_621);
or U824 (N_824,N_753,N_639);
nor U825 (N_825,N_641,N_749);
nor U826 (N_826,N_781,N_685);
nand U827 (N_827,N_662,N_646);
and U828 (N_828,N_750,N_684);
or U829 (N_829,N_792,N_713);
nor U830 (N_830,N_702,N_775);
nand U831 (N_831,N_767,N_642);
nor U832 (N_832,N_637,N_720);
or U833 (N_833,N_693,N_604);
and U834 (N_834,N_655,N_743);
or U835 (N_835,N_780,N_687);
nor U836 (N_836,N_628,N_661);
xor U837 (N_837,N_656,N_675);
nor U838 (N_838,N_716,N_607);
nand U839 (N_839,N_683,N_616);
and U840 (N_840,N_735,N_709);
nor U841 (N_841,N_674,N_737);
nand U842 (N_842,N_738,N_710);
or U843 (N_843,N_601,N_772);
or U844 (N_844,N_606,N_733);
and U845 (N_845,N_786,N_620);
nor U846 (N_846,N_669,N_740);
and U847 (N_847,N_672,N_673);
or U848 (N_848,N_640,N_766);
xnor U849 (N_849,N_717,N_652);
and U850 (N_850,N_676,N_774);
nor U851 (N_851,N_653,N_763);
or U852 (N_852,N_623,N_707);
nand U853 (N_853,N_776,N_791);
and U854 (N_854,N_698,N_691);
nor U855 (N_855,N_708,N_773);
or U856 (N_856,N_764,N_614);
nor U857 (N_857,N_647,N_745);
and U858 (N_858,N_796,N_611);
nor U859 (N_859,N_667,N_736);
or U860 (N_860,N_794,N_626);
or U861 (N_861,N_613,N_649);
or U862 (N_862,N_744,N_618);
nand U863 (N_863,N_630,N_678);
and U864 (N_864,N_779,N_718);
and U865 (N_865,N_797,N_712);
nand U866 (N_866,N_715,N_723);
nor U867 (N_867,N_727,N_714);
nor U868 (N_868,N_705,N_657);
and U869 (N_869,N_612,N_721);
and U870 (N_870,N_635,N_658);
nand U871 (N_871,N_636,N_758);
nor U872 (N_872,N_783,N_650);
or U873 (N_873,N_617,N_679);
and U874 (N_874,N_644,N_752);
or U875 (N_875,N_760,N_747);
nor U876 (N_876,N_746,N_790);
and U877 (N_877,N_670,N_799);
nand U878 (N_878,N_731,N_668);
nand U879 (N_879,N_784,N_666);
nor U880 (N_880,N_777,N_659);
and U881 (N_881,N_631,N_761);
nand U882 (N_882,N_706,N_757);
nand U883 (N_883,N_632,N_622);
nor U884 (N_884,N_748,N_625);
nand U885 (N_885,N_795,N_759);
nand U886 (N_886,N_695,N_769);
nor U887 (N_887,N_788,N_686);
nand U888 (N_888,N_762,N_671);
and U889 (N_889,N_778,N_726);
nand U890 (N_890,N_627,N_605);
or U891 (N_891,N_734,N_624);
and U892 (N_892,N_663,N_703);
or U893 (N_893,N_660,N_789);
or U894 (N_894,N_787,N_697);
nor U895 (N_895,N_615,N_619);
and U896 (N_896,N_724,N_755);
nand U897 (N_897,N_603,N_730);
and U898 (N_898,N_696,N_643);
and U899 (N_899,N_798,N_689);
nand U900 (N_900,N_673,N_728);
nor U901 (N_901,N_733,N_771);
and U902 (N_902,N_707,N_647);
nand U903 (N_903,N_705,N_714);
nand U904 (N_904,N_646,N_703);
nor U905 (N_905,N_779,N_748);
nand U906 (N_906,N_762,N_781);
or U907 (N_907,N_754,N_730);
or U908 (N_908,N_729,N_751);
or U909 (N_909,N_687,N_645);
and U910 (N_910,N_656,N_633);
nand U911 (N_911,N_779,N_612);
nor U912 (N_912,N_619,N_684);
nor U913 (N_913,N_627,N_739);
and U914 (N_914,N_654,N_777);
and U915 (N_915,N_726,N_786);
nor U916 (N_916,N_784,N_785);
nand U917 (N_917,N_756,N_674);
and U918 (N_918,N_745,N_650);
or U919 (N_919,N_699,N_697);
nand U920 (N_920,N_781,N_663);
nand U921 (N_921,N_690,N_694);
or U922 (N_922,N_782,N_707);
or U923 (N_923,N_723,N_612);
or U924 (N_924,N_676,N_637);
or U925 (N_925,N_692,N_634);
or U926 (N_926,N_720,N_755);
nor U927 (N_927,N_680,N_605);
and U928 (N_928,N_649,N_603);
nand U929 (N_929,N_720,N_764);
nor U930 (N_930,N_782,N_660);
and U931 (N_931,N_765,N_726);
nor U932 (N_932,N_607,N_788);
nor U933 (N_933,N_661,N_745);
or U934 (N_934,N_721,N_739);
or U935 (N_935,N_754,N_716);
or U936 (N_936,N_770,N_631);
or U937 (N_937,N_702,N_757);
or U938 (N_938,N_619,N_623);
and U939 (N_939,N_717,N_625);
or U940 (N_940,N_612,N_710);
or U941 (N_941,N_646,N_620);
or U942 (N_942,N_744,N_679);
nor U943 (N_943,N_638,N_628);
or U944 (N_944,N_635,N_641);
nand U945 (N_945,N_792,N_709);
nor U946 (N_946,N_654,N_655);
or U947 (N_947,N_660,N_702);
or U948 (N_948,N_683,N_720);
and U949 (N_949,N_604,N_700);
nor U950 (N_950,N_640,N_609);
nand U951 (N_951,N_718,N_618);
or U952 (N_952,N_623,N_780);
nor U953 (N_953,N_709,N_650);
or U954 (N_954,N_720,N_714);
and U955 (N_955,N_773,N_646);
and U956 (N_956,N_781,N_758);
nand U957 (N_957,N_667,N_640);
nand U958 (N_958,N_631,N_765);
and U959 (N_959,N_630,N_695);
and U960 (N_960,N_628,N_602);
nor U961 (N_961,N_704,N_736);
nor U962 (N_962,N_773,N_784);
nand U963 (N_963,N_756,N_703);
and U964 (N_964,N_782,N_729);
and U965 (N_965,N_796,N_709);
nand U966 (N_966,N_680,N_728);
nand U967 (N_967,N_629,N_726);
and U968 (N_968,N_788,N_694);
nor U969 (N_969,N_648,N_795);
nand U970 (N_970,N_705,N_770);
nor U971 (N_971,N_716,N_786);
and U972 (N_972,N_724,N_727);
xor U973 (N_973,N_675,N_764);
and U974 (N_974,N_786,N_634);
or U975 (N_975,N_787,N_713);
and U976 (N_976,N_793,N_628);
nor U977 (N_977,N_755,N_768);
xnor U978 (N_978,N_653,N_730);
or U979 (N_979,N_719,N_614);
and U980 (N_980,N_668,N_786);
or U981 (N_981,N_797,N_783);
and U982 (N_982,N_779,N_603);
or U983 (N_983,N_735,N_696);
nand U984 (N_984,N_702,N_680);
and U985 (N_985,N_777,N_727);
nor U986 (N_986,N_780,N_709);
or U987 (N_987,N_772,N_733);
nor U988 (N_988,N_630,N_774);
nand U989 (N_989,N_702,N_726);
nor U990 (N_990,N_601,N_645);
and U991 (N_991,N_723,N_663);
nor U992 (N_992,N_687,N_663);
xor U993 (N_993,N_639,N_729);
and U994 (N_994,N_690,N_765);
nor U995 (N_995,N_647,N_770);
nand U996 (N_996,N_653,N_626);
nor U997 (N_997,N_699,N_611);
or U998 (N_998,N_630,N_745);
nor U999 (N_999,N_671,N_711);
and U1000 (N_1000,N_886,N_890);
nor U1001 (N_1001,N_896,N_961);
and U1002 (N_1002,N_989,N_857);
nor U1003 (N_1003,N_999,N_913);
nand U1004 (N_1004,N_940,N_816);
and U1005 (N_1005,N_992,N_967);
and U1006 (N_1006,N_912,N_942);
nand U1007 (N_1007,N_956,N_848);
or U1008 (N_1008,N_963,N_981);
and U1009 (N_1009,N_906,N_858);
and U1010 (N_1010,N_859,N_914);
nor U1011 (N_1011,N_900,N_899);
nor U1012 (N_1012,N_991,N_819);
nand U1013 (N_1013,N_960,N_926);
nand U1014 (N_1014,N_964,N_864);
and U1015 (N_1015,N_946,N_995);
nor U1016 (N_1016,N_852,N_983);
nor U1017 (N_1017,N_953,N_868);
nor U1018 (N_1018,N_888,N_826);
nand U1019 (N_1019,N_892,N_823);
or U1020 (N_1020,N_903,N_834);
nand U1021 (N_1021,N_941,N_936);
and U1022 (N_1022,N_811,N_951);
or U1023 (N_1023,N_959,N_802);
nor U1024 (N_1024,N_915,N_856);
nand U1025 (N_1025,N_968,N_844);
nand U1026 (N_1026,N_817,N_980);
nor U1027 (N_1027,N_815,N_882);
nand U1028 (N_1028,N_846,N_840);
and U1029 (N_1029,N_904,N_814);
nand U1030 (N_1030,N_966,N_939);
nand U1031 (N_1031,N_931,N_962);
or U1032 (N_1032,N_894,N_803);
nand U1033 (N_1033,N_937,N_997);
and U1034 (N_1034,N_982,N_893);
nor U1035 (N_1035,N_849,N_873);
or U1036 (N_1036,N_998,N_821);
nor U1037 (N_1037,N_979,N_854);
nand U1038 (N_1038,N_809,N_812);
and U1039 (N_1039,N_925,N_869);
or U1040 (N_1040,N_944,N_820);
nor U1041 (N_1041,N_993,N_870);
nand U1042 (N_1042,N_808,N_924);
and U1043 (N_1043,N_883,N_898);
nand U1044 (N_1044,N_813,N_822);
or U1045 (N_1045,N_974,N_985);
nor U1046 (N_1046,N_838,N_928);
or U1047 (N_1047,N_806,N_850);
nand U1048 (N_1048,N_837,N_972);
nand U1049 (N_1049,N_911,N_860);
nand U1050 (N_1050,N_818,N_996);
nor U1051 (N_1051,N_880,N_832);
and U1052 (N_1052,N_975,N_845);
nor U1053 (N_1053,N_824,N_950);
nor U1054 (N_1054,N_976,N_862);
nor U1055 (N_1055,N_807,N_987);
or U1056 (N_1056,N_943,N_895);
nand U1057 (N_1057,N_842,N_805);
or U1058 (N_1058,N_843,N_923);
and U1059 (N_1059,N_917,N_905);
and U1060 (N_1060,N_839,N_947);
nor U1061 (N_1061,N_969,N_831);
nor U1062 (N_1062,N_855,N_938);
and U1063 (N_1063,N_994,N_910);
nand U1064 (N_1064,N_800,N_986);
and U1065 (N_1065,N_828,N_970);
nor U1066 (N_1066,N_830,N_861);
nand U1067 (N_1067,N_804,N_934);
or U1068 (N_1068,N_881,N_930);
nand U1069 (N_1069,N_867,N_909);
or U1070 (N_1070,N_884,N_954);
or U1071 (N_1071,N_948,N_908);
and U1072 (N_1072,N_847,N_851);
or U1073 (N_1073,N_889,N_874);
and U1074 (N_1074,N_835,N_865);
nor U1075 (N_1075,N_825,N_878);
or U1076 (N_1076,N_901,N_907);
and U1077 (N_1077,N_891,N_916);
nor U1078 (N_1078,N_902,N_984);
nor U1079 (N_1079,N_920,N_927);
nand U1080 (N_1080,N_918,N_952);
nor U1081 (N_1081,N_876,N_922);
and U1082 (N_1082,N_990,N_875);
nor U1083 (N_1083,N_841,N_949);
nand U1084 (N_1084,N_836,N_866);
nand U1085 (N_1085,N_810,N_871);
xor U1086 (N_1086,N_973,N_879);
nor U1087 (N_1087,N_945,N_957);
and U1088 (N_1088,N_897,N_958);
or U1089 (N_1089,N_971,N_829);
nor U1090 (N_1090,N_877,N_977);
nor U1091 (N_1091,N_932,N_887);
nor U1092 (N_1092,N_919,N_935);
nand U1093 (N_1093,N_827,N_872);
and U1094 (N_1094,N_978,N_921);
xnor U1095 (N_1095,N_988,N_965);
nand U1096 (N_1096,N_933,N_833);
nand U1097 (N_1097,N_929,N_885);
or U1098 (N_1098,N_863,N_955);
or U1099 (N_1099,N_801,N_853);
nand U1100 (N_1100,N_800,N_804);
and U1101 (N_1101,N_999,N_919);
and U1102 (N_1102,N_984,N_831);
or U1103 (N_1103,N_880,N_953);
nor U1104 (N_1104,N_815,N_982);
nor U1105 (N_1105,N_873,N_872);
or U1106 (N_1106,N_833,N_818);
or U1107 (N_1107,N_871,N_949);
nor U1108 (N_1108,N_875,N_869);
and U1109 (N_1109,N_875,N_824);
or U1110 (N_1110,N_958,N_942);
and U1111 (N_1111,N_888,N_962);
nor U1112 (N_1112,N_833,N_875);
or U1113 (N_1113,N_845,N_833);
and U1114 (N_1114,N_868,N_846);
nor U1115 (N_1115,N_990,N_912);
nor U1116 (N_1116,N_965,N_879);
nand U1117 (N_1117,N_947,N_835);
nand U1118 (N_1118,N_806,N_882);
nor U1119 (N_1119,N_870,N_996);
and U1120 (N_1120,N_956,N_829);
nor U1121 (N_1121,N_939,N_835);
and U1122 (N_1122,N_981,N_912);
or U1123 (N_1123,N_957,N_914);
nand U1124 (N_1124,N_973,N_951);
and U1125 (N_1125,N_880,N_819);
and U1126 (N_1126,N_871,N_862);
or U1127 (N_1127,N_834,N_999);
nor U1128 (N_1128,N_832,N_934);
or U1129 (N_1129,N_850,N_886);
and U1130 (N_1130,N_957,N_862);
nor U1131 (N_1131,N_978,N_971);
and U1132 (N_1132,N_828,N_929);
nor U1133 (N_1133,N_936,N_888);
nand U1134 (N_1134,N_843,N_976);
or U1135 (N_1135,N_986,N_863);
nand U1136 (N_1136,N_990,N_937);
and U1137 (N_1137,N_862,N_972);
or U1138 (N_1138,N_993,N_887);
nand U1139 (N_1139,N_966,N_885);
nand U1140 (N_1140,N_843,N_835);
nand U1141 (N_1141,N_971,N_821);
and U1142 (N_1142,N_958,N_844);
nor U1143 (N_1143,N_827,N_856);
nor U1144 (N_1144,N_891,N_840);
nor U1145 (N_1145,N_978,N_956);
or U1146 (N_1146,N_916,N_881);
nand U1147 (N_1147,N_980,N_896);
nand U1148 (N_1148,N_968,N_874);
or U1149 (N_1149,N_832,N_814);
or U1150 (N_1150,N_916,N_852);
nand U1151 (N_1151,N_943,N_814);
nor U1152 (N_1152,N_930,N_827);
nand U1153 (N_1153,N_811,N_855);
nor U1154 (N_1154,N_935,N_844);
and U1155 (N_1155,N_810,N_998);
nand U1156 (N_1156,N_900,N_970);
nor U1157 (N_1157,N_990,N_843);
and U1158 (N_1158,N_928,N_980);
xor U1159 (N_1159,N_944,N_927);
or U1160 (N_1160,N_898,N_945);
nand U1161 (N_1161,N_881,N_863);
nor U1162 (N_1162,N_814,N_865);
nor U1163 (N_1163,N_918,N_849);
and U1164 (N_1164,N_875,N_837);
and U1165 (N_1165,N_914,N_959);
nor U1166 (N_1166,N_860,N_902);
and U1167 (N_1167,N_879,N_877);
or U1168 (N_1168,N_858,N_842);
nor U1169 (N_1169,N_828,N_825);
nor U1170 (N_1170,N_916,N_978);
nor U1171 (N_1171,N_913,N_953);
nor U1172 (N_1172,N_938,N_805);
nand U1173 (N_1173,N_895,N_853);
nor U1174 (N_1174,N_803,N_996);
or U1175 (N_1175,N_961,N_849);
and U1176 (N_1176,N_976,N_951);
nor U1177 (N_1177,N_902,N_955);
nor U1178 (N_1178,N_906,N_984);
or U1179 (N_1179,N_985,N_821);
nand U1180 (N_1180,N_935,N_873);
and U1181 (N_1181,N_999,N_863);
or U1182 (N_1182,N_912,N_989);
and U1183 (N_1183,N_958,N_957);
nor U1184 (N_1184,N_995,N_953);
nor U1185 (N_1185,N_931,N_910);
and U1186 (N_1186,N_924,N_869);
nor U1187 (N_1187,N_805,N_833);
nand U1188 (N_1188,N_849,N_937);
nand U1189 (N_1189,N_845,N_909);
or U1190 (N_1190,N_997,N_862);
nor U1191 (N_1191,N_897,N_927);
or U1192 (N_1192,N_994,N_842);
or U1193 (N_1193,N_979,N_894);
nor U1194 (N_1194,N_943,N_834);
and U1195 (N_1195,N_934,N_917);
and U1196 (N_1196,N_967,N_995);
nand U1197 (N_1197,N_908,N_832);
and U1198 (N_1198,N_941,N_981);
or U1199 (N_1199,N_870,N_920);
nor U1200 (N_1200,N_1161,N_1019);
and U1201 (N_1201,N_1159,N_1026);
nor U1202 (N_1202,N_1078,N_1086);
and U1203 (N_1203,N_1122,N_1193);
and U1204 (N_1204,N_1123,N_1119);
and U1205 (N_1205,N_1035,N_1110);
nor U1206 (N_1206,N_1134,N_1047);
nand U1207 (N_1207,N_1091,N_1165);
nand U1208 (N_1208,N_1156,N_1188);
and U1209 (N_1209,N_1011,N_1151);
nand U1210 (N_1210,N_1039,N_1009);
and U1211 (N_1211,N_1109,N_1059);
and U1212 (N_1212,N_1032,N_1192);
nand U1213 (N_1213,N_1031,N_1195);
and U1214 (N_1214,N_1147,N_1094);
nor U1215 (N_1215,N_1008,N_1021);
nor U1216 (N_1216,N_1145,N_1184);
and U1217 (N_1217,N_1093,N_1092);
nand U1218 (N_1218,N_1173,N_1155);
nor U1219 (N_1219,N_1014,N_1000);
nand U1220 (N_1220,N_1117,N_1022);
or U1221 (N_1221,N_1044,N_1172);
and U1222 (N_1222,N_1133,N_1171);
nor U1223 (N_1223,N_1075,N_1007);
and U1224 (N_1224,N_1001,N_1163);
or U1225 (N_1225,N_1115,N_1095);
or U1226 (N_1226,N_1062,N_1182);
nand U1227 (N_1227,N_1004,N_1118);
and U1228 (N_1228,N_1038,N_1183);
nand U1229 (N_1229,N_1049,N_1170);
nor U1230 (N_1230,N_1116,N_1037);
and U1231 (N_1231,N_1025,N_1131);
or U1232 (N_1232,N_1056,N_1186);
xor U1233 (N_1233,N_1088,N_1154);
or U1234 (N_1234,N_1098,N_1187);
nor U1235 (N_1235,N_1160,N_1104);
and U1236 (N_1236,N_1157,N_1130);
and U1237 (N_1237,N_1111,N_1042);
nand U1238 (N_1238,N_1189,N_1143);
or U1239 (N_1239,N_1112,N_1089);
nand U1240 (N_1240,N_1051,N_1064);
nand U1241 (N_1241,N_1177,N_1146);
and U1242 (N_1242,N_1176,N_1190);
and U1243 (N_1243,N_1029,N_1139);
and U1244 (N_1244,N_1140,N_1027);
and U1245 (N_1245,N_1196,N_1061);
nand U1246 (N_1246,N_1033,N_1071);
nor U1247 (N_1247,N_1072,N_1180);
nand U1248 (N_1248,N_1137,N_1012);
or U1249 (N_1249,N_1144,N_1028);
and U1250 (N_1250,N_1066,N_1178);
nor U1251 (N_1251,N_1197,N_1158);
nand U1252 (N_1252,N_1079,N_1181);
nor U1253 (N_1253,N_1106,N_1010);
or U1254 (N_1254,N_1135,N_1076);
nor U1255 (N_1255,N_1053,N_1030);
and U1256 (N_1256,N_1002,N_1141);
or U1257 (N_1257,N_1199,N_1073);
or U1258 (N_1258,N_1142,N_1103);
nand U1259 (N_1259,N_1082,N_1149);
nor U1260 (N_1260,N_1048,N_1191);
or U1261 (N_1261,N_1058,N_1136);
nand U1262 (N_1262,N_1174,N_1099);
nand U1263 (N_1263,N_1138,N_1126);
and U1264 (N_1264,N_1108,N_1179);
nand U1265 (N_1265,N_1120,N_1070);
nand U1266 (N_1266,N_1100,N_1175);
or U1267 (N_1267,N_1166,N_1150);
nand U1268 (N_1268,N_1081,N_1065);
or U1269 (N_1269,N_1164,N_1050);
nor U1270 (N_1270,N_1045,N_1097);
nor U1271 (N_1271,N_1152,N_1013);
and U1272 (N_1272,N_1069,N_1107);
and U1273 (N_1273,N_1080,N_1023);
or U1274 (N_1274,N_1167,N_1169);
nor U1275 (N_1275,N_1043,N_1084);
nand U1276 (N_1276,N_1067,N_1168);
or U1277 (N_1277,N_1068,N_1162);
nand U1278 (N_1278,N_1024,N_1128);
and U1279 (N_1279,N_1090,N_1132);
and U1280 (N_1280,N_1198,N_1114);
and U1281 (N_1281,N_1036,N_1148);
or U1282 (N_1282,N_1034,N_1185);
or U1283 (N_1283,N_1153,N_1060);
nand U1284 (N_1284,N_1055,N_1105);
or U1285 (N_1285,N_1096,N_1006);
nor U1286 (N_1286,N_1015,N_1057);
nor U1287 (N_1287,N_1003,N_1054);
nand U1288 (N_1288,N_1020,N_1040);
nor U1289 (N_1289,N_1016,N_1125);
nor U1290 (N_1290,N_1085,N_1077);
nand U1291 (N_1291,N_1083,N_1129);
nand U1292 (N_1292,N_1005,N_1121);
nor U1293 (N_1293,N_1102,N_1101);
nor U1294 (N_1294,N_1052,N_1127);
or U1295 (N_1295,N_1087,N_1017);
nand U1296 (N_1296,N_1018,N_1041);
or U1297 (N_1297,N_1124,N_1113);
nor U1298 (N_1298,N_1046,N_1063);
or U1299 (N_1299,N_1074,N_1194);
nand U1300 (N_1300,N_1140,N_1111);
and U1301 (N_1301,N_1151,N_1091);
or U1302 (N_1302,N_1062,N_1037);
or U1303 (N_1303,N_1047,N_1089);
or U1304 (N_1304,N_1159,N_1029);
and U1305 (N_1305,N_1102,N_1100);
or U1306 (N_1306,N_1094,N_1189);
and U1307 (N_1307,N_1092,N_1053);
nand U1308 (N_1308,N_1143,N_1119);
nand U1309 (N_1309,N_1082,N_1001);
xnor U1310 (N_1310,N_1020,N_1138);
nand U1311 (N_1311,N_1109,N_1060);
and U1312 (N_1312,N_1054,N_1112);
nor U1313 (N_1313,N_1154,N_1092);
and U1314 (N_1314,N_1127,N_1093);
nand U1315 (N_1315,N_1095,N_1069);
nand U1316 (N_1316,N_1022,N_1089);
nand U1317 (N_1317,N_1191,N_1032);
nor U1318 (N_1318,N_1051,N_1033);
nor U1319 (N_1319,N_1112,N_1080);
nor U1320 (N_1320,N_1119,N_1155);
and U1321 (N_1321,N_1004,N_1157);
xor U1322 (N_1322,N_1120,N_1023);
nor U1323 (N_1323,N_1073,N_1197);
nor U1324 (N_1324,N_1037,N_1170);
nand U1325 (N_1325,N_1188,N_1187);
and U1326 (N_1326,N_1093,N_1002);
or U1327 (N_1327,N_1192,N_1130);
nand U1328 (N_1328,N_1044,N_1054);
or U1329 (N_1329,N_1124,N_1147);
and U1330 (N_1330,N_1198,N_1135);
nor U1331 (N_1331,N_1031,N_1111);
and U1332 (N_1332,N_1169,N_1066);
nand U1333 (N_1333,N_1176,N_1125);
and U1334 (N_1334,N_1193,N_1002);
nand U1335 (N_1335,N_1191,N_1137);
or U1336 (N_1336,N_1175,N_1099);
or U1337 (N_1337,N_1140,N_1168);
and U1338 (N_1338,N_1109,N_1015);
nand U1339 (N_1339,N_1033,N_1178);
and U1340 (N_1340,N_1067,N_1106);
and U1341 (N_1341,N_1072,N_1192);
and U1342 (N_1342,N_1148,N_1033);
nand U1343 (N_1343,N_1151,N_1071);
nor U1344 (N_1344,N_1150,N_1033);
or U1345 (N_1345,N_1064,N_1080);
or U1346 (N_1346,N_1071,N_1144);
or U1347 (N_1347,N_1143,N_1193);
nor U1348 (N_1348,N_1075,N_1146);
or U1349 (N_1349,N_1152,N_1000);
and U1350 (N_1350,N_1055,N_1182);
nor U1351 (N_1351,N_1189,N_1089);
nor U1352 (N_1352,N_1005,N_1034);
and U1353 (N_1353,N_1054,N_1056);
nand U1354 (N_1354,N_1191,N_1076);
nor U1355 (N_1355,N_1110,N_1055);
nand U1356 (N_1356,N_1157,N_1125);
and U1357 (N_1357,N_1058,N_1075);
nand U1358 (N_1358,N_1033,N_1137);
nor U1359 (N_1359,N_1144,N_1130);
and U1360 (N_1360,N_1066,N_1064);
or U1361 (N_1361,N_1156,N_1193);
nand U1362 (N_1362,N_1150,N_1081);
and U1363 (N_1363,N_1048,N_1056);
nor U1364 (N_1364,N_1063,N_1194);
nor U1365 (N_1365,N_1139,N_1049);
and U1366 (N_1366,N_1008,N_1110);
and U1367 (N_1367,N_1156,N_1150);
nand U1368 (N_1368,N_1078,N_1002);
or U1369 (N_1369,N_1136,N_1195);
nor U1370 (N_1370,N_1094,N_1127);
nor U1371 (N_1371,N_1069,N_1102);
and U1372 (N_1372,N_1189,N_1137);
nor U1373 (N_1373,N_1090,N_1072);
nor U1374 (N_1374,N_1084,N_1160);
nor U1375 (N_1375,N_1147,N_1177);
or U1376 (N_1376,N_1048,N_1081);
nand U1377 (N_1377,N_1028,N_1027);
nor U1378 (N_1378,N_1050,N_1027);
nand U1379 (N_1379,N_1132,N_1110);
nand U1380 (N_1380,N_1035,N_1127);
or U1381 (N_1381,N_1089,N_1033);
nand U1382 (N_1382,N_1143,N_1135);
nand U1383 (N_1383,N_1166,N_1167);
nor U1384 (N_1384,N_1096,N_1079);
nand U1385 (N_1385,N_1009,N_1073);
or U1386 (N_1386,N_1077,N_1038);
and U1387 (N_1387,N_1102,N_1155);
nand U1388 (N_1388,N_1121,N_1003);
nor U1389 (N_1389,N_1064,N_1147);
or U1390 (N_1390,N_1013,N_1199);
and U1391 (N_1391,N_1165,N_1124);
nor U1392 (N_1392,N_1195,N_1085);
or U1393 (N_1393,N_1077,N_1010);
nor U1394 (N_1394,N_1122,N_1060);
xor U1395 (N_1395,N_1013,N_1028);
or U1396 (N_1396,N_1034,N_1114);
nor U1397 (N_1397,N_1064,N_1087);
and U1398 (N_1398,N_1051,N_1024);
or U1399 (N_1399,N_1097,N_1191);
nor U1400 (N_1400,N_1348,N_1248);
nor U1401 (N_1401,N_1218,N_1328);
or U1402 (N_1402,N_1246,N_1376);
nand U1403 (N_1403,N_1399,N_1202);
or U1404 (N_1404,N_1339,N_1265);
and U1405 (N_1405,N_1310,N_1277);
nor U1406 (N_1406,N_1278,N_1252);
or U1407 (N_1407,N_1304,N_1393);
nor U1408 (N_1408,N_1261,N_1333);
or U1409 (N_1409,N_1314,N_1327);
nor U1410 (N_1410,N_1309,N_1317);
and U1411 (N_1411,N_1302,N_1268);
nor U1412 (N_1412,N_1282,N_1274);
xor U1413 (N_1413,N_1290,N_1242);
nand U1414 (N_1414,N_1208,N_1292);
nor U1415 (N_1415,N_1276,N_1330);
nand U1416 (N_1416,N_1212,N_1335);
or U1417 (N_1417,N_1345,N_1236);
and U1418 (N_1418,N_1269,N_1307);
and U1419 (N_1419,N_1211,N_1293);
and U1420 (N_1420,N_1286,N_1321);
nand U1421 (N_1421,N_1390,N_1240);
or U1422 (N_1422,N_1209,N_1262);
or U1423 (N_1423,N_1326,N_1256);
nand U1424 (N_1424,N_1312,N_1254);
nand U1425 (N_1425,N_1331,N_1241);
or U1426 (N_1426,N_1350,N_1264);
nand U1427 (N_1427,N_1382,N_1398);
nand U1428 (N_1428,N_1200,N_1377);
and U1429 (N_1429,N_1353,N_1358);
nor U1430 (N_1430,N_1371,N_1344);
and U1431 (N_1431,N_1210,N_1340);
and U1432 (N_1432,N_1396,N_1365);
or U1433 (N_1433,N_1315,N_1392);
nor U1434 (N_1434,N_1324,N_1383);
nor U1435 (N_1435,N_1283,N_1354);
nor U1436 (N_1436,N_1338,N_1225);
nor U1437 (N_1437,N_1366,N_1291);
or U1438 (N_1438,N_1267,N_1323);
or U1439 (N_1439,N_1311,N_1359);
nor U1440 (N_1440,N_1332,N_1351);
or U1441 (N_1441,N_1303,N_1250);
nor U1442 (N_1442,N_1280,N_1271);
nand U1443 (N_1443,N_1281,N_1375);
and U1444 (N_1444,N_1285,N_1362);
nor U1445 (N_1445,N_1299,N_1381);
or U1446 (N_1446,N_1205,N_1319);
and U1447 (N_1447,N_1329,N_1336);
nand U1448 (N_1448,N_1203,N_1227);
or U1449 (N_1449,N_1325,N_1334);
nor U1450 (N_1450,N_1217,N_1222);
or U1451 (N_1451,N_1387,N_1201);
nand U1452 (N_1452,N_1235,N_1226);
nand U1453 (N_1453,N_1395,N_1287);
nand U1454 (N_1454,N_1361,N_1229);
and U1455 (N_1455,N_1284,N_1249);
and U1456 (N_1456,N_1369,N_1368);
and U1457 (N_1457,N_1305,N_1373);
and U1458 (N_1458,N_1379,N_1394);
or U1459 (N_1459,N_1320,N_1337);
nand U1460 (N_1460,N_1363,N_1237);
and U1461 (N_1461,N_1367,N_1273);
or U1462 (N_1462,N_1389,N_1385);
and U1463 (N_1463,N_1215,N_1322);
nor U1464 (N_1464,N_1380,N_1206);
nor U1465 (N_1465,N_1253,N_1220);
and U1466 (N_1466,N_1388,N_1306);
nor U1467 (N_1467,N_1247,N_1232);
and U1468 (N_1468,N_1272,N_1295);
and U1469 (N_1469,N_1296,N_1297);
nand U1470 (N_1470,N_1370,N_1355);
nand U1471 (N_1471,N_1260,N_1341);
nand U1472 (N_1472,N_1239,N_1228);
or U1473 (N_1473,N_1391,N_1275);
or U1474 (N_1474,N_1374,N_1386);
and U1475 (N_1475,N_1216,N_1233);
and U1476 (N_1476,N_1397,N_1289);
and U1477 (N_1477,N_1251,N_1263);
nand U1478 (N_1478,N_1372,N_1349);
nand U1479 (N_1479,N_1357,N_1238);
or U1480 (N_1480,N_1313,N_1213);
or U1481 (N_1481,N_1270,N_1207);
or U1482 (N_1482,N_1257,N_1258);
nand U1483 (N_1483,N_1316,N_1360);
or U1484 (N_1484,N_1346,N_1378);
and U1485 (N_1485,N_1234,N_1243);
or U1486 (N_1486,N_1223,N_1300);
nor U1487 (N_1487,N_1279,N_1342);
nor U1488 (N_1488,N_1288,N_1230);
or U1489 (N_1489,N_1221,N_1219);
or U1490 (N_1490,N_1259,N_1266);
or U1491 (N_1491,N_1244,N_1255);
nor U1492 (N_1492,N_1224,N_1347);
and U1493 (N_1493,N_1356,N_1318);
nor U1494 (N_1494,N_1301,N_1384);
and U1495 (N_1495,N_1298,N_1294);
nor U1496 (N_1496,N_1352,N_1214);
nor U1497 (N_1497,N_1245,N_1231);
nor U1498 (N_1498,N_1343,N_1308);
and U1499 (N_1499,N_1364,N_1204);
nor U1500 (N_1500,N_1329,N_1373);
nor U1501 (N_1501,N_1364,N_1347);
nand U1502 (N_1502,N_1202,N_1286);
or U1503 (N_1503,N_1278,N_1366);
nor U1504 (N_1504,N_1272,N_1296);
or U1505 (N_1505,N_1345,N_1217);
or U1506 (N_1506,N_1380,N_1240);
nor U1507 (N_1507,N_1304,N_1368);
nor U1508 (N_1508,N_1241,N_1228);
nand U1509 (N_1509,N_1351,N_1358);
nor U1510 (N_1510,N_1306,N_1349);
nor U1511 (N_1511,N_1384,N_1351);
nor U1512 (N_1512,N_1397,N_1376);
or U1513 (N_1513,N_1267,N_1255);
or U1514 (N_1514,N_1245,N_1285);
and U1515 (N_1515,N_1358,N_1290);
and U1516 (N_1516,N_1208,N_1302);
and U1517 (N_1517,N_1396,N_1210);
and U1518 (N_1518,N_1344,N_1364);
and U1519 (N_1519,N_1293,N_1273);
or U1520 (N_1520,N_1380,N_1207);
or U1521 (N_1521,N_1228,N_1314);
xor U1522 (N_1522,N_1314,N_1334);
nand U1523 (N_1523,N_1303,N_1300);
or U1524 (N_1524,N_1273,N_1398);
or U1525 (N_1525,N_1215,N_1297);
and U1526 (N_1526,N_1383,N_1395);
and U1527 (N_1527,N_1272,N_1208);
or U1528 (N_1528,N_1307,N_1297);
or U1529 (N_1529,N_1311,N_1223);
and U1530 (N_1530,N_1292,N_1239);
nor U1531 (N_1531,N_1239,N_1225);
nor U1532 (N_1532,N_1282,N_1306);
and U1533 (N_1533,N_1225,N_1348);
nand U1534 (N_1534,N_1372,N_1235);
or U1535 (N_1535,N_1204,N_1394);
nor U1536 (N_1536,N_1212,N_1322);
and U1537 (N_1537,N_1229,N_1291);
or U1538 (N_1538,N_1392,N_1353);
and U1539 (N_1539,N_1378,N_1334);
nand U1540 (N_1540,N_1254,N_1250);
and U1541 (N_1541,N_1288,N_1355);
nor U1542 (N_1542,N_1210,N_1380);
nand U1543 (N_1543,N_1235,N_1263);
nand U1544 (N_1544,N_1210,N_1200);
nand U1545 (N_1545,N_1318,N_1377);
nor U1546 (N_1546,N_1355,N_1258);
nor U1547 (N_1547,N_1393,N_1379);
nor U1548 (N_1548,N_1223,N_1335);
nor U1549 (N_1549,N_1267,N_1235);
and U1550 (N_1550,N_1348,N_1304);
or U1551 (N_1551,N_1226,N_1246);
nor U1552 (N_1552,N_1386,N_1399);
or U1553 (N_1553,N_1398,N_1340);
or U1554 (N_1554,N_1294,N_1297);
nor U1555 (N_1555,N_1392,N_1247);
nor U1556 (N_1556,N_1250,N_1398);
nand U1557 (N_1557,N_1204,N_1342);
or U1558 (N_1558,N_1221,N_1381);
or U1559 (N_1559,N_1228,N_1326);
xor U1560 (N_1560,N_1252,N_1361);
and U1561 (N_1561,N_1369,N_1288);
nand U1562 (N_1562,N_1282,N_1204);
nor U1563 (N_1563,N_1250,N_1200);
xnor U1564 (N_1564,N_1399,N_1368);
nand U1565 (N_1565,N_1253,N_1340);
nor U1566 (N_1566,N_1230,N_1332);
and U1567 (N_1567,N_1393,N_1293);
or U1568 (N_1568,N_1310,N_1289);
and U1569 (N_1569,N_1360,N_1321);
or U1570 (N_1570,N_1318,N_1229);
and U1571 (N_1571,N_1350,N_1289);
nand U1572 (N_1572,N_1358,N_1256);
and U1573 (N_1573,N_1204,N_1283);
and U1574 (N_1574,N_1224,N_1250);
nand U1575 (N_1575,N_1291,N_1394);
and U1576 (N_1576,N_1226,N_1339);
nor U1577 (N_1577,N_1316,N_1231);
nor U1578 (N_1578,N_1300,N_1292);
nand U1579 (N_1579,N_1292,N_1303);
or U1580 (N_1580,N_1390,N_1362);
nor U1581 (N_1581,N_1220,N_1233);
nor U1582 (N_1582,N_1381,N_1320);
nand U1583 (N_1583,N_1249,N_1285);
nand U1584 (N_1584,N_1310,N_1205);
nand U1585 (N_1585,N_1258,N_1267);
or U1586 (N_1586,N_1320,N_1282);
and U1587 (N_1587,N_1390,N_1397);
or U1588 (N_1588,N_1269,N_1289);
nand U1589 (N_1589,N_1217,N_1215);
and U1590 (N_1590,N_1258,N_1329);
and U1591 (N_1591,N_1216,N_1296);
nor U1592 (N_1592,N_1231,N_1325);
nor U1593 (N_1593,N_1314,N_1342);
nand U1594 (N_1594,N_1292,N_1347);
nand U1595 (N_1595,N_1227,N_1366);
or U1596 (N_1596,N_1293,N_1220);
or U1597 (N_1597,N_1392,N_1241);
nand U1598 (N_1598,N_1333,N_1285);
nand U1599 (N_1599,N_1207,N_1334);
and U1600 (N_1600,N_1569,N_1553);
and U1601 (N_1601,N_1487,N_1456);
and U1602 (N_1602,N_1431,N_1516);
and U1603 (N_1603,N_1450,N_1568);
nor U1604 (N_1604,N_1508,N_1503);
or U1605 (N_1605,N_1537,N_1510);
nand U1606 (N_1606,N_1547,N_1417);
and U1607 (N_1607,N_1590,N_1478);
nand U1608 (N_1608,N_1593,N_1464);
nor U1609 (N_1609,N_1545,N_1551);
nand U1610 (N_1610,N_1484,N_1595);
nand U1611 (N_1611,N_1408,N_1495);
nor U1612 (N_1612,N_1423,N_1578);
and U1613 (N_1613,N_1474,N_1564);
or U1614 (N_1614,N_1556,N_1505);
nor U1615 (N_1615,N_1559,N_1514);
xor U1616 (N_1616,N_1570,N_1411);
and U1617 (N_1617,N_1511,N_1438);
nor U1618 (N_1618,N_1531,N_1504);
nand U1619 (N_1619,N_1506,N_1546);
and U1620 (N_1620,N_1498,N_1482);
nand U1621 (N_1621,N_1414,N_1419);
and U1622 (N_1622,N_1557,N_1558);
and U1623 (N_1623,N_1433,N_1522);
or U1624 (N_1624,N_1497,N_1410);
nand U1625 (N_1625,N_1589,N_1437);
and U1626 (N_1626,N_1402,N_1457);
or U1627 (N_1627,N_1562,N_1481);
nor U1628 (N_1628,N_1581,N_1526);
or U1629 (N_1629,N_1421,N_1413);
and U1630 (N_1630,N_1565,N_1502);
nor U1631 (N_1631,N_1420,N_1528);
and U1632 (N_1632,N_1462,N_1523);
nand U1633 (N_1633,N_1405,N_1567);
nor U1634 (N_1634,N_1428,N_1499);
nand U1635 (N_1635,N_1486,N_1576);
nand U1636 (N_1636,N_1401,N_1451);
nand U1637 (N_1637,N_1573,N_1594);
nand U1638 (N_1638,N_1415,N_1473);
and U1639 (N_1639,N_1465,N_1521);
or U1640 (N_1640,N_1403,N_1580);
or U1641 (N_1641,N_1540,N_1472);
nor U1642 (N_1642,N_1449,N_1582);
xor U1643 (N_1643,N_1579,N_1538);
nand U1644 (N_1644,N_1517,N_1574);
and U1645 (N_1645,N_1445,N_1548);
and U1646 (N_1646,N_1552,N_1544);
and U1647 (N_1647,N_1571,N_1572);
nand U1648 (N_1648,N_1598,N_1424);
or U1649 (N_1649,N_1448,N_1429);
or U1650 (N_1650,N_1549,N_1461);
nor U1651 (N_1651,N_1454,N_1446);
and U1652 (N_1652,N_1587,N_1555);
nor U1653 (N_1653,N_1409,N_1422);
nand U1654 (N_1654,N_1535,N_1542);
nor U1655 (N_1655,N_1539,N_1533);
nand U1656 (N_1656,N_1443,N_1494);
or U1657 (N_1657,N_1507,N_1501);
and U1658 (N_1658,N_1527,N_1566);
and U1659 (N_1659,N_1467,N_1460);
or U1660 (N_1660,N_1475,N_1599);
nor U1661 (N_1661,N_1541,N_1550);
or U1662 (N_1662,N_1468,N_1561);
nor U1663 (N_1663,N_1407,N_1585);
and U1664 (N_1664,N_1416,N_1434);
nand U1665 (N_1665,N_1532,N_1418);
and U1666 (N_1666,N_1404,N_1534);
nand U1667 (N_1667,N_1515,N_1469);
or U1668 (N_1668,N_1512,N_1441);
nand U1669 (N_1669,N_1432,N_1436);
nor U1670 (N_1670,N_1476,N_1463);
or U1671 (N_1671,N_1584,N_1586);
or U1672 (N_1672,N_1525,N_1524);
and U1673 (N_1673,N_1492,N_1440);
nand U1674 (N_1674,N_1477,N_1560);
xor U1675 (N_1675,N_1543,N_1493);
nand U1676 (N_1676,N_1442,N_1453);
nor U1677 (N_1677,N_1513,N_1496);
and U1678 (N_1678,N_1488,N_1577);
nor U1679 (N_1679,N_1518,N_1466);
nor U1680 (N_1680,N_1489,N_1447);
or U1681 (N_1681,N_1400,N_1455);
nand U1682 (N_1682,N_1596,N_1563);
or U1683 (N_1683,N_1435,N_1591);
or U1684 (N_1684,N_1597,N_1529);
nor U1685 (N_1685,N_1412,N_1480);
xor U1686 (N_1686,N_1536,N_1575);
or U1687 (N_1687,N_1471,N_1426);
nor U1688 (N_1688,N_1509,N_1490);
nand U1689 (N_1689,N_1483,N_1470);
or U1690 (N_1690,N_1588,N_1439);
and U1691 (N_1691,N_1425,N_1519);
or U1692 (N_1692,N_1583,N_1459);
or U1693 (N_1693,N_1530,N_1554);
nand U1694 (N_1694,N_1430,N_1479);
or U1695 (N_1695,N_1427,N_1406);
nand U1696 (N_1696,N_1491,N_1520);
nor U1697 (N_1697,N_1500,N_1452);
nor U1698 (N_1698,N_1592,N_1458);
or U1699 (N_1699,N_1485,N_1444);
or U1700 (N_1700,N_1530,N_1499);
nor U1701 (N_1701,N_1457,N_1533);
or U1702 (N_1702,N_1551,N_1520);
nand U1703 (N_1703,N_1597,N_1426);
nand U1704 (N_1704,N_1476,N_1450);
nand U1705 (N_1705,N_1594,N_1565);
nand U1706 (N_1706,N_1410,N_1594);
nor U1707 (N_1707,N_1521,N_1496);
nor U1708 (N_1708,N_1432,N_1588);
nand U1709 (N_1709,N_1564,N_1532);
nand U1710 (N_1710,N_1544,N_1465);
or U1711 (N_1711,N_1551,N_1524);
or U1712 (N_1712,N_1400,N_1492);
and U1713 (N_1713,N_1594,N_1578);
and U1714 (N_1714,N_1453,N_1494);
or U1715 (N_1715,N_1445,N_1402);
nor U1716 (N_1716,N_1494,N_1495);
or U1717 (N_1717,N_1491,N_1526);
nor U1718 (N_1718,N_1406,N_1547);
nand U1719 (N_1719,N_1526,N_1593);
and U1720 (N_1720,N_1468,N_1593);
nor U1721 (N_1721,N_1512,N_1429);
nand U1722 (N_1722,N_1482,N_1591);
or U1723 (N_1723,N_1432,N_1548);
and U1724 (N_1724,N_1547,N_1403);
nor U1725 (N_1725,N_1571,N_1436);
nand U1726 (N_1726,N_1548,N_1500);
nor U1727 (N_1727,N_1482,N_1414);
nor U1728 (N_1728,N_1446,N_1476);
or U1729 (N_1729,N_1403,N_1538);
nor U1730 (N_1730,N_1542,N_1536);
nor U1731 (N_1731,N_1546,N_1417);
nand U1732 (N_1732,N_1459,N_1590);
nand U1733 (N_1733,N_1545,N_1492);
or U1734 (N_1734,N_1549,N_1435);
nor U1735 (N_1735,N_1528,N_1515);
nand U1736 (N_1736,N_1590,N_1406);
nand U1737 (N_1737,N_1577,N_1472);
nor U1738 (N_1738,N_1510,N_1405);
nor U1739 (N_1739,N_1444,N_1435);
or U1740 (N_1740,N_1597,N_1515);
nor U1741 (N_1741,N_1588,N_1410);
and U1742 (N_1742,N_1553,N_1415);
nand U1743 (N_1743,N_1559,N_1433);
and U1744 (N_1744,N_1438,N_1574);
nand U1745 (N_1745,N_1518,N_1585);
nand U1746 (N_1746,N_1447,N_1480);
nand U1747 (N_1747,N_1424,N_1400);
nand U1748 (N_1748,N_1496,N_1569);
or U1749 (N_1749,N_1483,N_1422);
and U1750 (N_1750,N_1523,N_1528);
nor U1751 (N_1751,N_1462,N_1598);
nor U1752 (N_1752,N_1554,N_1479);
and U1753 (N_1753,N_1562,N_1537);
nand U1754 (N_1754,N_1576,N_1457);
and U1755 (N_1755,N_1501,N_1427);
nand U1756 (N_1756,N_1438,N_1513);
nand U1757 (N_1757,N_1546,N_1541);
and U1758 (N_1758,N_1444,N_1510);
nand U1759 (N_1759,N_1525,N_1436);
and U1760 (N_1760,N_1583,N_1412);
or U1761 (N_1761,N_1565,N_1592);
or U1762 (N_1762,N_1428,N_1418);
or U1763 (N_1763,N_1420,N_1544);
nand U1764 (N_1764,N_1435,N_1556);
and U1765 (N_1765,N_1446,N_1542);
and U1766 (N_1766,N_1441,N_1456);
nor U1767 (N_1767,N_1518,N_1537);
and U1768 (N_1768,N_1580,N_1466);
xor U1769 (N_1769,N_1412,N_1545);
nor U1770 (N_1770,N_1516,N_1459);
or U1771 (N_1771,N_1530,N_1545);
nand U1772 (N_1772,N_1529,N_1402);
xor U1773 (N_1773,N_1511,N_1471);
nand U1774 (N_1774,N_1405,N_1528);
nand U1775 (N_1775,N_1569,N_1495);
or U1776 (N_1776,N_1568,N_1546);
and U1777 (N_1777,N_1454,N_1403);
and U1778 (N_1778,N_1506,N_1410);
nor U1779 (N_1779,N_1462,N_1433);
nand U1780 (N_1780,N_1539,N_1400);
and U1781 (N_1781,N_1569,N_1521);
nand U1782 (N_1782,N_1594,N_1424);
nor U1783 (N_1783,N_1425,N_1458);
nand U1784 (N_1784,N_1403,N_1423);
and U1785 (N_1785,N_1418,N_1459);
or U1786 (N_1786,N_1529,N_1467);
and U1787 (N_1787,N_1492,N_1578);
nand U1788 (N_1788,N_1593,N_1503);
nor U1789 (N_1789,N_1515,N_1539);
nor U1790 (N_1790,N_1568,N_1497);
or U1791 (N_1791,N_1599,N_1519);
or U1792 (N_1792,N_1507,N_1451);
nor U1793 (N_1793,N_1557,N_1465);
nand U1794 (N_1794,N_1460,N_1492);
or U1795 (N_1795,N_1536,N_1446);
nor U1796 (N_1796,N_1528,N_1423);
and U1797 (N_1797,N_1487,N_1523);
nor U1798 (N_1798,N_1571,N_1546);
and U1799 (N_1799,N_1490,N_1587);
nor U1800 (N_1800,N_1714,N_1746);
or U1801 (N_1801,N_1645,N_1620);
nand U1802 (N_1802,N_1650,N_1696);
or U1803 (N_1803,N_1667,N_1658);
nand U1804 (N_1804,N_1784,N_1671);
nor U1805 (N_1805,N_1765,N_1711);
and U1806 (N_1806,N_1649,N_1723);
and U1807 (N_1807,N_1771,N_1797);
nor U1808 (N_1808,N_1615,N_1624);
or U1809 (N_1809,N_1605,N_1754);
or U1810 (N_1810,N_1672,N_1724);
or U1811 (N_1811,N_1769,N_1703);
and U1812 (N_1812,N_1721,N_1648);
and U1813 (N_1813,N_1708,N_1761);
nor U1814 (N_1814,N_1735,N_1747);
and U1815 (N_1815,N_1734,N_1799);
nand U1816 (N_1816,N_1767,N_1783);
or U1817 (N_1817,N_1713,N_1674);
nor U1818 (N_1818,N_1792,N_1760);
nand U1819 (N_1819,N_1640,N_1638);
or U1820 (N_1820,N_1749,N_1676);
nand U1821 (N_1821,N_1633,N_1603);
or U1822 (N_1822,N_1618,N_1675);
and U1823 (N_1823,N_1610,N_1704);
nor U1824 (N_1824,N_1741,N_1685);
nand U1825 (N_1825,N_1611,N_1694);
nor U1826 (N_1826,N_1722,N_1635);
nor U1827 (N_1827,N_1758,N_1634);
nor U1828 (N_1828,N_1623,N_1643);
or U1829 (N_1829,N_1636,N_1774);
nor U1830 (N_1830,N_1701,N_1727);
nor U1831 (N_1831,N_1600,N_1653);
nor U1832 (N_1832,N_1778,N_1743);
and U1833 (N_1833,N_1693,N_1656);
and U1834 (N_1834,N_1730,N_1790);
or U1835 (N_1835,N_1719,N_1604);
nor U1836 (N_1836,N_1728,N_1773);
nor U1837 (N_1837,N_1751,N_1788);
nand U1838 (N_1838,N_1742,N_1732);
and U1839 (N_1839,N_1786,N_1678);
nand U1840 (N_1840,N_1630,N_1764);
or U1841 (N_1841,N_1698,N_1716);
nand U1842 (N_1842,N_1775,N_1745);
nor U1843 (N_1843,N_1744,N_1686);
or U1844 (N_1844,N_1625,N_1641);
or U1845 (N_1845,N_1700,N_1683);
and U1846 (N_1846,N_1613,N_1660);
and U1847 (N_1847,N_1748,N_1669);
and U1848 (N_1848,N_1717,N_1617);
nor U1849 (N_1849,N_1687,N_1776);
nor U1850 (N_1850,N_1677,N_1791);
and U1851 (N_1851,N_1628,N_1632);
and U1852 (N_1852,N_1740,N_1795);
nand U1853 (N_1853,N_1720,N_1782);
or U1854 (N_1854,N_1762,N_1659);
nand U1855 (N_1855,N_1607,N_1709);
nor U1856 (N_1856,N_1681,N_1781);
and U1857 (N_1857,N_1794,N_1750);
or U1858 (N_1858,N_1770,N_1601);
nand U1859 (N_1859,N_1699,N_1766);
and U1860 (N_1860,N_1668,N_1705);
nand U1861 (N_1861,N_1602,N_1697);
and U1862 (N_1862,N_1639,N_1657);
nor U1863 (N_1863,N_1768,N_1666);
and U1864 (N_1864,N_1779,N_1780);
and U1865 (N_1865,N_1759,N_1757);
nor U1866 (N_1866,N_1637,N_1796);
nand U1867 (N_1867,N_1789,N_1665);
or U1868 (N_1868,N_1715,N_1739);
or U1869 (N_1869,N_1661,N_1712);
nor U1870 (N_1870,N_1707,N_1619);
and U1871 (N_1871,N_1752,N_1654);
nand U1872 (N_1872,N_1798,N_1662);
nand U1873 (N_1873,N_1793,N_1725);
and U1874 (N_1874,N_1647,N_1690);
or U1875 (N_1875,N_1627,N_1753);
and U1876 (N_1876,N_1729,N_1689);
nand U1877 (N_1877,N_1691,N_1692);
and U1878 (N_1878,N_1738,N_1644);
or U1879 (N_1879,N_1622,N_1688);
nand U1880 (N_1880,N_1663,N_1655);
nand U1881 (N_1881,N_1680,N_1737);
nand U1882 (N_1882,N_1626,N_1642);
nor U1883 (N_1883,N_1621,N_1670);
nor U1884 (N_1884,N_1756,N_1777);
nor U1885 (N_1885,N_1706,N_1616);
or U1886 (N_1886,N_1646,N_1726);
or U1887 (N_1887,N_1787,N_1629);
or U1888 (N_1888,N_1718,N_1652);
nand U1889 (N_1889,N_1682,N_1684);
nand U1890 (N_1890,N_1695,N_1710);
or U1891 (N_1891,N_1763,N_1631);
nor U1892 (N_1892,N_1731,N_1736);
nand U1893 (N_1893,N_1679,N_1673);
nor U1894 (N_1894,N_1606,N_1651);
nand U1895 (N_1895,N_1755,N_1612);
nor U1896 (N_1896,N_1785,N_1614);
nor U1897 (N_1897,N_1733,N_1702);
nor U1898 (N_1898,N_1608,N_1772);
xnor U1899 (N_1899,N_1609,N_1664);
nor U1900 (N_1900,N_1604,N_1697);
nor U1901 (N_1901,N_1612,N_1648);
nand U1902 (N_1902,N_1688,N_1709);
nand U1903 (N_1903,N_1653,N_1645);
or U1904 (N_1904,N_1636,N_1603);
or U1905 (N_1905,N_1717,N_1653);
and U1906 (N_1906,N_1714,N_1729);
nor U1907 (N_1907,N_1620,N_1763);
nand U1908 (N_1908,N_1776,N_1775);
and U1909 (N_1909,N_1790,N_1713);
or U1910 (N_1910,N_1760,N_1712);
nand U1911 (N_1911,N_1651,N_1713);
nand U1912 (N_1912,N_1746,N_1739);
and U1913 (N_1913,N_1798,N_1736);
or U1914 (N_1914,N_1763,N_1779);
or U1915 (N_1915,N_1670,N_1740);
or U1916 (N_1916,N_1633,N_1793);
or U1917 (N_1917,N_1651,N_1755);
nand U1918 (N_1918,N_1679,N_1736);
nand U1919 (N_1919,N_1677,N_1624);
nand U1920 (N_1920,N_1730,N_1661);
or U1921 (N_1921,N_1625,N_1792);
or U1922 (N_1922,N_1688,N_1658);
and U1923 (N_1923,N_1715,N_1733);
nand U1924 (N_1924,N_1695,N_1697);
nor U1925 (N_1925,N_1628,N_1732);
nor U1926 (N_1926,N_1703,N_1659);
nand U1927 (N_1927,N_1655,N_1660);
nand U1928 (N_1928,N_1620,N_1742);
and U1929 (N_1929,N_1713,N_1668);
or U1930 (N_1930,N_1678,N_1703);
and U1931 (N_1931,N_1648,N_1758);
nand U1932 (N_1932,N_1634,N_1707);
or U1933 (N_1933,N_1660,N_1682);
nor U1934 (N_1934,N_1767,N_1695);
nor U1935 (N_1935,N_1645,N_1628);
nor U1936 (N_1936,N_1684,N_1696);
nor U1937 (N_1937,N_1785,N_1610);
or U1938 (N_1938,N_1728,N_1721);
or U1939 (N_1939,N_1688,N_1760);
and U1940 (N_1940,N_1687,N_1706);
nor U1941 (N_1941,N_1614,N_1777);
and U1942 (N_1942,N_1685,N_1670);
or U1943 (N_1943,N_1771,N_1757);
nand U1944 (N_1944,N_1782,N_1766);
and U1945 (N_1945,N_1731,N_1775);
or U1946 (N_1946,N_1759,N_1698);
and U1947 (N_1947,N_1792,N_1713);
xor U1948 (N_1948,N_1755,N_1745);
or U1949 (N_1949,N_1629,N_1784);
nor U1950 (N_1950,N_1795,N_1615);
nand U1951 (N_1951,N_1768,N_1620);
nor U1952 (N_1952,N_1605,N_1663);
and U1953 (N_1953,N_1623,N_1788);
nor U1954 (N_1954,N_1712,N_1633);
or U1955 (N_1955,N_1777,N_1695);
and U1956 (N_1956,N_1606,N_1740);
or U1957 (N_1957,N_1631,N_1651);
and U1958 (N_1958,N_1772,N_1605);
and U1959 (N_1959,N_1726,N_1740);
nand U1960 (N_1960,N_1782,N_1729);
xor U1961 (N_1961,N_1634,N_1638);
nand U1962 (N_1962,N_1780,N_1774);
nor U1963 (N_1963,N_1780,N_1651);
nor U1964 (N_1964,N_1630,N_1799);
nand U1965 (N_1965,N_1743,N_1782);
nor U1966 (N_1966,N_1717,N_1619);
nand U1967 (N_1967,N_1787,N_1775);
and U1968 (N_1968,N_1622,N_1620);
nand U1969 (N_1969,N_1695,N_1791);
nor U1970 (N_1970,N_1725,N_1787);
or U1971 (N_1971,N_1763,N_1604);
xor U1972 (N_1972,N_1742,N_1771);
and U1973 (N_1973,N_1675,N_1623);
or U1974 (N_1974,N_1700,N_1606);
nor U1975 (N_1975,N_1614,N_1644);
nor U1976 (N_1976,N_1759,N_1673);
nand U1977 (N_1977,N_1744,N_1761);
nand U1978 (N_1978,N_1741,N_1669);
and U1979 (N_1979,N_1711,N_1759);
nand U1980 (N_1980,N_1721,N_1688);
nor U1981 (N_1981,N_1766,N_1700);
and U1982 (N_1982,N_1778,N_1621);
or U1983 (N_1983,N_1628,N_1706);
nand U1984 (N_1984,N_1780,N_1636);
or U1985 (N_1985,N_1707,N_1748);
and U1986 (N_1986,N_1692,N_1667);
and U1987 (N_1987,N_1724,N_1794);
or U1988 (N_1988,N_1661,N_1695);
or U1989 (N_1989,N_1765,N_1683);
nor U1990 (N_1990,N_1786,N_1704);
nand U1991 (N_1991,N_1685,N_1649);
or U1992 (N_1992,N_1756,N_1674);
nor U1993 (N_1993,N_1791,N_1652);
nor U1994 (N_1994,N_1700,N_1655);
or U1995 (N_1995,N_1680,N_1609);
or U1996 (N_1996,N_1605,N_1609);
and U1997 (N_1997,N_1676,N_1696);
and U1998 (N_1998,N_1736,N_1726);
nand U1999 (N_1999,N_1621,N_1673);
nand U2000 (N_2000,N_1846,N_1949);
nor U2001 (N_2001,N_1838,N_1959);
and U2002 (N_2002,N_1890,N_1939);
and U2003 (N_2003,N_1800,N_1879);
nand U2004 (N_2004,N_1969,N_1851);
or U2005 (N_2005,N_1983,N_1968);
nand U2006 (N_2006,N_1875,N_1935);
or U2007 (N_2007,N_1813,N_1901);
nor U2008 (N_2008,N_1945,N_1926);
nor U2009 (N_2009,N_1853,N_1805);
nor U2010 (N_2010,N_1874,N_1927);
or U2011 (N_2011,N_1859,N_1924);
nand U2012 (N_2012,N_1881,N_1946);
nand U2013 (N_2013,N_1810,N_1819);
nand U2014 (N_2014,N_1942,N_1826);
and U2015 (N_2015,N_1914,N_1920);
nor U2016 (N_2016,N_1913,N_1937);
and U2017 (N_2017,N_1982,N_1812);
and U2018 (N_2018,N_1957,N_1991);
or U2019 (N_2019,N_1828,N_1801);
and U2020 (N_2020,N_1947,N_1895);
or U2021 (N_2021,N_1887,N_1970);
and U2022 (N_2022,N_1900,N_1839);
and U2023 (N_2023,N_1941,N_1965);
nand U2024 (N_2024,N_1882,N_1817);
and U2025 (N_2025,N_1876,N_1902);
nand U2026 (N_2026,N_1896,N_1886);
nor U2027 (N_2027,N_1940,N_1993);
nor U2028 (N_2028,N_1972,N_1842);
or U2029 (N_2029,N_1840,N_1827);
nor U2030 (N_2030,N_1986,N_1824);
xnor U2031 (N_2031,N_1866,N_1845);
and U2032 (N_2032,N_1919,N_1952);
or U2033 (N_2033,N_1889,N_1815);
and U2034 (N_2034,N_1932,N_1960);
nor U2035 (N_2035,N_1884,N_1974);
nor U2036 (N_2036,N_1861,N_1962);
or U2037 (N_2037,N_1871,N_1858);
nand U2038 (N_2038,N_1831,N_1903);
nor U2039 (N_2039,N_1976,N_1943);
and U2040 (N_2040,N_1823,N_1880);
or U2041 (N_2041,N_1835,N_1860);
or U2042 (N_2042,N_1916,N_1888);
nand U2043 (N_2043,N_1917,N_1883);
or U2044 (N_2044,N_1911,N_1843);
and U2045 (N_2045,N_1865,N_1996);
and U2046 (N_2046,N_1904,N_1837);
nand U2047 (N_2047,N_1862,N_1873);
nor U2048 (N_2048,N_1921,N_1966);
nand U2049 (N_2049,N_1809,N_1822);
and U2050 (N_2050,N_1808,N_1953);
and U2051 (N_2051,N_1869,N_1816);
nand U2052 (N_2052,N_1997,N_1973);
nor U2053 (N_2053,N_1908,N_1967);
or U2054 (N_2054,N_1802,N_1971);
nor U2055 (N_2055,N_1832,N_1867);
or U2056 (N_2056,N_1847,N_1998);
and U2057 (N_2057,N_1877,N_1820);
nand U2058 (N_2058,N_1849,N_1915);
or U2059 (N_2059,N_1897,N_1933);
xor U2060 (N_2060,N_1961,N_1855);
and U2061 (N_2061,N_1885,N_1893);
or U2062 (N_2062,N_1841,N_1850);
nor U2063 (N_2063,N_1990,N_1891);
and U2064 (N_2064,N_1954,N_1868);
nand U2065 (N_2065,N_1950,N_1811);
nand U2066 (N_2066,N_1892,N_1995);
nor U2067 (N_2067,N_1825,N_1930);
and U2068 (N_2068,N_1856,N_1907);
nor U2069 (N_2069,N_1989,N_1964);
nand U2070 (N_2070,N_1872,N_1948);
or U2071 (N_2071,N_1818,N_1999);
nand U2072 (N_2072,N_1980,N_1898);
or U2073 (N_2073,N_1936,N_1803);
nand U2074 (N_2074,N_1981,N_1956);
nand U2075 (N_2075,N_1977,N_1906);
or U2076 (N_2076,N_1804,N_1821);
xnor U2077 (N_2077,N_1984,N_1878);
and U2078 (N_2078,N_1929,N_1864);
and U2079 (N_2079,N_1994,N_1848);
and U2080 (N_2080,N_1992,N_1979);
or U2081 (N_2081,N_1830,N_1833);
nor U2082 (N_2082,N_1923,N_1863);
xor U2083 (N_2083,N_1988,N_1834);
xor U2084 (N_2084,N_1938,N_1925);
nand U2085 (N_2085,N_1814,N_1909);
and U2086 (N_2086,N_1870,N_1905);
or U2087 (N_2087,N_1934,N_1958);
nor U2088 (N_2088,N_1806,N_1829);
and U2089 (N_2089,N_1852,N_1854);
nor U2090 (N_2090,N_1899,N_1836);
or U2091 (N_2091,N_1944,N_1978);
or U2092 (N_2092,N_1955,N_1987);
or U2093 (N_2093,N_1807,N_1912);
nor U2094 (N_2094,N_1951,N_1928);
and U2095 (N_2095,N_1931,N_1910);
nand U2096 (N_2096,N_1857,N_1844);
nor U2097 (N_2097,N_1918,N_1894);
nor U2098 (N_2098,N_1922,N_1975);
or U2099 (N_2099,N_1985,N_1963);
and U2100 (N_2100,N_1944,N_1915);
or U2101 (N_2101,N_1961,N_1946);
or U2102 (N_2102,N_1808,N_1933);
and U2103 (N_2103,N_1808,N_1960);
nand U2104 (N_2104,N_1880,N_1973);
nand U2105 (N_2105,N_1836,N_1915);
nand U2106 (N_2106,N_1839,N_1815);
nand U2107 (N_2107,N_1896,N_1842);
and U2108 (N_2108,N_1969,N_1868);
or U2109 (N_2109,N_1993,N_1947);
and U2110 (N_2110,N_1935,N_1898);
or U2111 (N_2111,N_1972,N_1846);
nor U2112 (N_2112,N_1802,N_1937);
and U2113 (N_2113,N_1930,N_1855);
nor U2114 (N_2114,N_1883,N_1946);
or U2115 (N_2115,N_1951,N_1930);
or U2116 (N_2116,N_1956,N_1941);
or U2117 (N_2117,N_1819,N_1804);
nor U2118 (N_2118,N_1848,N_1983);
nor U2119 (N_2119,N_1843,N_1992);
and U2120 (N_2120,N_1852,N_1806);
and U2121 (N_2121,N_1989,N_1816);
nor U2122 (N_2122,N_1809,N_1882);
nor U2123 (N_2123,N_1922,N_1851);
nand U2124 (N_2124,N_1971,N_1898);
xor U2125 (N_2125,N_1916,N_1875);
nor U2126 (N_2126,N_1946,N_1868);
or U2127 (N_2127,N_1889,N_1860);
nand U2128 (N_2128,N_1851,N_1829);
and U2129 (N_2129,N_1833,N_1820);
nand U2130 (N_2130,N_1852,N_1977);
nor U2131 (N_2131,N_1952,N_1999);
nor U2132 (N_2132,N_1924,N_1805);
nor U2133 (N_2133,N_1843,N_1887);
nor U2134 (N_2134,N_1870,N_1837);
nor U2135 (N_2135,N_1834,N_1931);
nand U2136 (N_2136,N_1904,N_1955);
or U2137 (N_2137,N_1878,N_1926);
nand U2138 (N_2138,N_1897,N_1944);
nor U2139 (N_2139,N_1930,N_1979);
and U2140 (N_2140,N_1880,N_1833);
and U2141 (N_2141,N_1863,N_1876);
nor U2142 (N_2142,N_1820,N_1945);
or U2143 (N_2143,N_1938,N_1954);
and U2144 (N_2144,N_1966,N_1898);
nand U2145 (N_2145,N_1910,N_1832);
nand U2146 (N_2146,N_1806,N_1932);
nand U2147 (N_2147,N_1801,N_1988);
or U2148 (N_2148,N_1990,N_1975);
and U2149 (N_2149,N_1914,N_1995);
nand U2150 (N_2150,N_1805,N_1836);
and U2151 (N_2151,N_1840,N_1992);
nand U2152 (N_2152,N_1912,N_1946);
or U2153 (N_2153,N_1852,N_1954);
and U2154 (N_2154,N_1844,N_1813);
and U2155 (N_2155,N_1904,N_1839);
nand U2156 (N_2156,N_1819,N_1850);
or U2157 (N_2157,N_1845,N_1803);
nor U2158 (N_2158,N_1976,N_1893);
and U2159 (N_2159,N_1945,N_1856);
nand U2160 (N_2160,N_1866,N_1990);
nand U2161 (N_2161,N_1869,N_1955);
nor U2162 (N_2162,N_1802,N_1836);
and U2163 (N_2163,N_1860,N_1844);
or U2164 (N_2164,N_1978,N_1851);
nand U2165 (N_2165,N_1803,N_1960);
nor U2166 (N_2166,N_1938,N_1803);
nor U2167 (N_2167,N_1866,N_1824);
nand U2168 (N_2168,N_1914,N_1884);
or U2169 (N_2169,N_1910,N_1920);
nor U2170 (N_2170,N_1806,N_1862);
and U2171 (N_2171,N_1875,N_1850);
nor U2172 (N_2172,N_1945,N_1938);
or U2173 (N_2173,N_1956,N_1944);
and U2174 (N_2174,N_1991,N_1946);
and U2175 (N_2175,N_1863,N_1973);
nor U2176 (N_2176,N_1948,N_1927);
nand U2177 (N_2177,N_1931,N_1912);
nand U2178 (N_2178,N_1823,N_1804);
nor U2179 (N_2179,N_1887,N_1883);
nand U2180 (N_2180,N_1949,N_1863);
and U2181 (N_2181,N_1881,N_1952);
nand U2182 (N_2182,N_1800,N_1849);
nor U2183 (N_2183,N_1801,N_1885);
and U2184 (N_2184,N_1924,N_1837);
nand U2185 (N_2185,N_1830,N_1832);
nand U2186 (N_2186,N_1875,N_1982);
and U2187 (N_2187,N_1956,N_1846);
nand U2188 (N_2188,N_1931,N_1884);
nand U2189 (N_2189,N_1927,N_1837);
nor U2190 (N_2190,N_1950,N_1978);
nor U2191 (N_2191,N_1984,N_1813);
or U2192 (N_2192,N_1862,N_1909);
or U2193 (N_2193,N_1968,N_1835);
nand U2194 (N_2194,N_1800,N_1838);
nand U2195 (N_2195,N_1836,N_1959);
or U2196 (N_2196,N_1835,N_1867);
nor U2197 (N_2197,N_1892,N_1916);
xor U2198 (N_2198,N_1966,N_1872);
xnor U2199 (N_2199,N_1845,N_1887);
and U2200 (N_2200,N_2063,N_2170);
and U2201 (N_2201,N_2091,N_2160);
nor U2202 (N_2202,N_2052,N_2132);
or U2203 (N_2203,N_2039,N_2106);
or U2204 (N_2204,N_2119,N_2121);
and U2205 (N_2205,N_2064,N_2152);
nand U2206 (N_2206,N_2089,N_2023);
or U2207 (N_2207,N_2027,N_2000);
and U2208 (N_2208,N_2129,N_2149);
xor U2209 (N_2209,N_2017,N_2105);
or U2210 (N_2210,N_2024,N_2042);
nand U2211 (N_2211,N_2186,N_2071);
or U2212 (N_2212,N_2179,N_2151);
nor U2213 (N_2213,N_2146,N_2067);
nor U2214 (N_2214,N_2101,N_2093);
nand U2215 (N_2215,N_2150,N_2158);
and U2216 (N_2216,N_2002,N_2060);
or U2217 (N_2217,N_2109,N_2174);
and U2218 (N_2218,N_2161,N_2081);
and U2219 (N_2219,N_2140,N_2133);
nand U2220 (N_2220,N_2034,N_2153);
or U2221 (N_2221,N_2198,N_2036);
nand U2222 (N_2222,N_2007,N_2187);
nor U2223 (N_2223,N_2041,N_2053);
or U2224 (N_2224,N_2073,N_2092);
nor U2225 (N_2225,N_2022,N_2137);
nand U2226 (N_2226,N_2005,N_2190);
nand U2227 (N_2227,N_2199,N_2100);
or U2228 (N_2228,N_2154,N_2131);
nand U2229 (N_2229,N_2026,N_2175);
nor U2230 (N_2230,N_2029,N_2094);
nand U2231 (N_2231,N_2085,N_2114);
nor U2232 (N_2232,N_2192,N_2176);
or U2233 (N_2233,N_2118,N_2057);
nand U2234 (N_2234,N_2122,N_2080);
nor U2235 (N_2235,N_2163,N_2172);
or U2236 (N_2236,N_2130,N_2010);
nand U2237 (N_2237,N_2145,N_2079);
nor U2238 (N_2238,N_2072,N_2123);
or U2239 (N_2239,N_2183,N_2135);
nor U2240 (N_2240,N_2098,N_2021);
nor U2241 (N_2241,N_2068,N_2189);
and U2242 (N_2242,N_2178,N_2008);
and U2243 (N_2243,N_2086,N_2103);
xnor U2244 (N_2244,N_2075,N_2082);
or U2245 (N_2245,N_2194,N_2004);
and U2246 (N_2246,N_2025,N_2043);
nand U2247 (N_2247,N_2185,N_2003);
and U2248 (N_2248,N_2049,N_2127);
or U2249 (N_2249,N_2076,N_2001);
and U2250 (N_2250,N_2097,N_2142);
or U2251 (N_2251,N_2035,N_2045);
nand U2252 (N_2252,N_2125,N_2083);
and U2253 (N_2253,N_2197,N_2088);
nand U2254 (N_2254,N_2048,N_2028);
nor U2255 (N_2255,N_2102,N_2013);
nand U2256 (N_2256,N_2104,N_2037);
xor U2257 (N_2257,N_2099,N_2196);
and U2258 (N_2258,N_2031,N_2018);
nor U2259 (N_2259,N_2164,N_2087);
nor U2260 (N_2260,N_2156,N_2056);
nor U2261 (N_2261,N_2096,N_2011);
or U2262 (N_2262,N_2120,N_2032);
or U2263 (N_2263,N_2012,N_2117);
nand U2264 (N_2264,N_2074,N_2165);
nor U2265 (N_2265,N_2110,N_2126);
nand U2266 (N_2266,N_2143,N_2157);
or U2267 (N_2267,N_2040,N_2180);
or U2268 (N_2268,N_2033,N_2065);
and U2269 (N_2269,N_2016,N_2193);
nor U2270 (N_2270,N_2019,N_2182);
and U2271 (N_2271,N_2167,N_2195);
and U2272 (N_2272,N_2020,N_2090);
or U2273 (N_2273,N_2046,N_2141);
nor U2274 (N_2274,N_2173,N_2191);
nand U2275 (N_2275,N_2134,N_2038);
and U2276 (N_2276,N_2015,N_2077);
and U2277 (N_2277,N_2171,N_2116);
or U2278 (N_2278,N_2061,N_2069);
nand U2279 (N_2279,N_2138,N_2047);
or U2280 (N_2280,N_2166,N_2006);
and U2281 (N_2281,N_2155,N_2112);
nor U2282 (N_2282,N_2177,N_2009);
or U2283 (N_2283,N_2169,N_2062);
nor U2284 (N_2284,N_2078,N_2128);
or U2285 (N_2285,N_2014,N_2066);
or U2286 (N_2286,N_2111,N_2054);
nand U2287 (N_2287,N_2159,N_2070);
nand U2288 (N_2288,N_2115,N_2188);
and U2289 (N_2289,N_2148,N_2136);
nor U2290 (N_2290,N_2181,N_2058);
or U2291 (N_2291,N_2107,N_2044);
or U2292 (N_2292,N_2147,N_2084);
nor U2293 (N_2293,N_2162,N_2030);
or U2294 (N_2294,N_2055,N_2168);
and U2295 (N_2295,N_2139,N_2095);
xor U2296 (N_2296,N_2059,N_2124);
nor U2297 (N_2297,N_2051,N_2113);
nor U2298 (N_2298,N_2184,N_2108);
or U2299 (N_2299,N_2144,N_2050);
nor U2300 (N_2300,N_2137,N_2072);
nand U2301 (N_2301,N_2135,N_2010);
or U2302 (N_2302,N_2087,N_2152);
or U2303 (N_2303,N_2102,N_2185);
nand U2304 (N_2304,N_2181,N_2095);
nor U2305 (N_2305,N_2022,N_2183);
and U2306 (N_2306,N_2183,N_2078);
nand U2307 (N_2307,N_2008,N_2144);
and U2308 (N_2308,N_2023,N_2012);
and U2309 (N_2309,N_2025,N_2141);
nand U2310 (N_2310,N_2164,N_2096);
nor U2311 (N_2311,N_2111,N_2165);
and U2312 (N_2312,N_2138,N_2103);
nor U2313 (N_2313,N_2063,N_2113);
nor U2314 (N_2314,N_2129,N_2114);
nor U2315 (N_2315,N_2044,N_2077);
nor U2316 (N_2316,N_2063,N_2184);
or U2317 (N_2317,N_2151,N_2073);
nand U2318 (N_2318,N_2119,N_2192);
nand U2319 (N_2319,N_2074,N_2005);
nand U2320 (N_2320,N_2104,N_2070);
nor U2321 (N_2321,N_2178,N_2091);
nand U2322 (N_2322,N_2060,N_2138);
and U2323 (N_2323,N_2132,N_2063);
and U2324 (N_2324,N_2125,N_2055);
or U2325 (N_2325,N_2101,N_2117);
or U2326 (N_2326,N_2182,N_2197);
or U2327 (N_2327,N_2116,N_2035);
nor U2328 (N_2328,N_2165,N_2039);
and U2329 (N_2329,N_2049,N_2067);
and U2330 (N_2330,N_2162,N_2137);
nand U2331 (N_2331,N_2045,N_2130);
nor U2332 (N_2332,N_2003,N_2161);
and U2333 (N_2333,N_2008,N_2161);
nor U2334 (N_2334,N_2046,N_2109);
nand U2335 (N_2335,N_2124,N_2092);
or U2336 (N_2336,N_2074,N_2046);
and U2337 (N_2337,N_2095,N_2112);
nor U2338 (N_2338,N_2006,N_2029);
nor U2339 (N_2339,N_2048,N_2020);
nand U2340 (N_2340,N_2074,N_2144);
nor U2341 (N_2341,N_2171,N_2075);
nand U2342 (N_2342,N_2173,N_2098);
nand U2343 (N_2343,N_2198,N_2055);
and U2344 (N_2344,N_2075,N_2021);
nand U2345 (N_2345,N_2045,N_2164);
and U2346 (N_2346,N_2060,N_2174);
and U2347 (N_2347,N_2028,N_2053);
or U2348 (N_2348,N_2051,N_2127);
nor U2349 (N_2349,N_2032,N_2126);
nand U2350 (N_2350,N_2056,N_2071);
nor U2351 (N_2351,N_2074,N_2038);
nor U2352 (N_2352,N_2151,N_2077);
nand U2353 (N_2353,N_2000,N_2109);
and U2354 (N_2354,N_2045,N_2030);
nand U2355 (N_2355,N_2106,N_2045);
nand U2356 (N_2356,N_2048,N_2014);
or U2357 (N_2357,N_2162,N_2117);
and U2358 (N_2358,N_2071,N_2085);
and U2359 (N_2359,N_2142,N_2108);
nand U2360 (N_2360,N_2175,N_2044);
nor U2361 (N_2361,N_2000,N_2046);
or U2362 (N_2362,N_2106,N_2161);
nand U2363 (N_2363,N_2153,N_2185);
nor U2364 (N_2364,N_2083,N_2148);
nor U2365 (N_2365,N_2049,N_2019);
or U2366 (N_2366,N_2113,N_2058);
xor U2367 (N_2367,N_2072,N_2075);
and U2368 (N_2368,N_2030,N_2037);
nand U2369 (N_2369,N_2131,N_2084);
or U2370 (N_2370,N_2125,N_2124);
xnor U2371 (N_2371,N_2072,N_2136);
nor U2372 (N_2372,N_2141,N_2148);
nand U2373 (N_2373,N_2126,N_2101);
or U2374 (N_2374,N_2088,N_2180);
or U2375 (N_2375,N_2125,N_2062);
or U2376 (N_2376,N_2043,N_2058);
nand U2377 (N_2377,N_2119,N_2118);
and U2378 (N_2378,N_2182,N_2183);
nor U2379 (N_2379,N_2051,N_2086);
nor U2380 (N_2380,N_2058,N_2068);
nand U2381 (N_2381,N_2143,N_2049);
and U2382 (N_2382,N_2091,N_2000);
nand U2383 (N_2383,N_2168,N_2035);
and U2384 (N_2384,N_2140,N_2001);
nand U2385 (N_2385,N_2105,N_2076);
and U2386 (N_2386,N_2122,N_2102);
and U2387 (N_2387,N_2110,N_2116);
or U2388 (N_2388,N_2143,N_2067);
and U2389 (N_2389,N_2196,N_2169);
nor U2390 (N_2390,N_2040,N_2092);
nand U2391 (N_2391,N_2171,N_2193);
nand U2392 (N_2392,N_2017,N_2129);
nand U2393 (N_2393,N_2057,N_2170);
and U2394 (N_2394,N_2144,N_2119);
nor U2395 (N_2395,N_2036,N_2147);
nor U2396 (N_2396,N_2100,N_2003);
nor U2397 (N_2397,N_2121,N_2092);
or U2398 (N_2398,N_2052,N_2046);
nor U2399 (N_2399,N_2075,N_2106);
and U2400 (N_2400,N_2254,N_2276);
nand U2401 (N_2401,N_2331,N_2241);
and U2402 (N_2402,N_2346,N_2257);
nor U2403 (N_2403,N_2217,N_2306);
and U2404 (N_2404,N_2291,N_2215);
and U2405 (N_2405,N_2232,N_2314);
and U2406 (N_2406,N_2295,N_2228);
nor U2407 (N_2407,N_2329,N_2239);
and U2408 (N_2408,N_2310,N_2327);
and U2409 (N_2409,N_2333,N_2352);
or U2410 (N_2410,N_2202,N_2261);
nand U2411 (N_2411,N_2277,N_2376);
nand U2412 (N_2412,N_2201,N_2390);
or U2413 (N_2413,N_2203,N_2209);
or U2414 (N_2414,N_2235,N_2282);
and U2415 (N_2415,N_2392,N_2339);
or U2416 (N_2416,N_2321,N_2384);
nand U2417 (N_2417,N_2238,N_2284);
and U2418 (N_2418,N_2388,N_2233);
or U2419 (N_2419,N_2389,N_2328);
nand U2420 (N_2420,N_2391,N_2326);
and U2421 (N_2421,N_2371,N_2305);
nor U2422 (N_2422,N_2317,N_2367);
or U2423 (N_2423,N_2380,N_2296);
nand U2424 (N_2424,N_2385,N_2332);
and U2425 (N_2425,N_2207,N_2256);
nor U2426 (N_2426,N_2301,N_2292);
nand U2427 (N_2427,N_2298,N_2344);
and U2428 (N_2428,N_2365,N_2323);
and U2429 (N_2429,N_2262,N_2288);
nor U2430 (N_2430,N_2330,N_2347);
and U2431 (N_2431,N_2294,N_2253);
and U2432 (N_2432,N_2274,N_2275);
nor U2433 (N_2433,N_2297,N_2267);
nor U2434 (N_2434,N_2299,N_2303);
nor U2435 (N_2435,N_2393,N_2386);
and U2436 (N_2436,N_2210,N_2236);
or U2437 (N_2437,N_2377,N_2312);
and U2438 (N_2438,N_2363,N_2338);
and U2439 (N_2439,N_2378,N_2366);
and U2440 (N_2440,N_2381,N_2372);
nand U2441 (N_2441,N_2316,N_2287);
or U2442 (N_2442,N_2362,N_2319);
nor U2443 (N_2443,N_2258,N_2357);
or U2444 (N_2444,N_2399,N_2247);
or U2445 (N_2445,N_2204,N_2350);
and U2446 (N_2446,N_2243,N_2374);
xor U2447 (N_2447,N_2320,N_2250);
or U2448 (N_2448,N_2227,N_2221);
nor U2449 (N_2449,N_2396,N_2370);
and U2450 (N_2450,N_2272,N_2349);
nor U2451 (N_2451,N_2355,N_2208);
nor U2452 (N_2452,N_2345,N_2226);
nor U2453 (N_2453,N_2279,N_2356);
nor U2454 (N_2454,N_2206,N_2283);
nor U2455 (N_2455,N_2231,N_2251);
or U2456 (N_2456,N_2341,N_2200);
nand U2457 (N_2457,N_2337,N_2219);
nand U2458 (N_2458,N_2373,N_2269);
nor U2459 (N_2459,N_2340,N_2216);
nand U2460 (N_2460,N_2265,N_2273);
or U2461 (N_2461,N_2334,N_2260);
or U2462 (N_2462,N_2259,N_2214);
or U2463 (N_2463,N_2281,N_2307);
nor U2464 (N_2464,N_2335,N_2240);
and U2465 (N_2465,N_2230,N_2395);
nor U2466 (N_2466,N_2218,N_2234);
and U2467 (N_2467,N_2354,N_2224);
or U2468 (N_2468,N_2394,N_2325);
nor U2469 (N_2469,N_2220,N_2278);
and U2470 (N_2470,N_2249,N_2322);
nand U2471 (N_2471,N_2271,N_2364);
nor U2472 (N_2472,N_2369,N_2311);
or U2473 (N_2473,N_2222,N_2290);
nand U2474 (N_2474,N_2293,N_2289);
xnor U2475 (N_2475,N_2324,N_2398);
and U2476 (N_2476,N_2382,N_2211);
and U2477 (N_2477,N_2318,N_2212);
nor U2478 (N_2478,N_2263,N_2383);
nand U2479 (N_2479,N_2351,N_2387);
and U2480 (N_2480,N_2308,N_2264);
or U2481 (N_2481,N_2309,N_2343);
nor U2482 (N_2482,N_2246,N_2286);
or U2483 (N_2483,N_2313,N_2223);
or U2484 (N_2484,N_2358,N_2353);
or U2485 (N_2485,N_2348,N_2242);
or U2486 (N_2486,N_2245,N_2205);
and U2487 (N_2487,N_2336,N_2280);
nor U2488 (N_2488,N_2375,N_2368);
nor U2489 (N_2489,N_2266,N_2225);
and U2490 (N_2490,N_2361,N_2229);
or U2491 (N_2491,N_2213,N_2268);
and U2492 (N_2492,N_2315,N_2397);
or U2493 (N_2493,N_2244,N_2359);
nor U2494 (N_2494,N_2304,N_2300);
or U2495 (N_2495,N_2360,N_2248);
and U2496 (N_2496,N_2379,N_2285);
nand U2497 (N_2497,N_2270,N_2252);
and U2498 (N_2498,N_2255,N_2302);
and U2499 (N_2499,N_2342,N_2237);
and U2500 (N_2500,N_2351,N_2223);
nor U2501 (N_2501,N_2312,N_2254);
or U2502 (N_2502,N_2225,N_2228);
and U2503 (N_2503,N_2232,N_2302);
and U2504 (N_2504,N_2370,N_2288);
and U2505 (N_2505,N_2322,N_2243);
nor U2506 (N_2506,N_2294,N_2374);
and U2507 (N_2507,N_2358,N_2222);
xnor U2508 (N_2508,N_2332,N_2362);
and U2509 (N_2509,N_2363,N_2216);
or U2510 (N_2510,N_2238,N_2272);
nor U2511 (N_2511,N_2207,N_2322);
or U2512 (N_2512,N_2295,N_2296);
and U2513 (N_2513,N_2219,N_2363);
nor U2514 (N_2514,N_2341,N_2334);
xor U2515 (N_2515,N_2285,N_2366);
nor U2516 (N_2516,N_2207,N_2335);
and U2517 (N_2517,N_2306,N_2283);
or U2518 (N_2518,N_2312,N_2215);
nand U2519 (N_2519,N_2220,N_2290);
or U2520 (N_2520,N_2348,N_2394);
nand U2521 (N_2521,N_2389,N_2360);
and U2522 (N_2522,N_2336,N_2327);
nand U2523 (N_2523,N_2312,N_2399);
or U2524 (N_2524,N_2239,N_2319);
nor U2525 (N_2525,N_2297,N_2360);
nor U2526 (N_2526,N_2287,N_2240);
nor U2527 (N_2527,N_2341,N_2298);
nor U2528 (N_2528,N_2297,N_2212);
or U2529 (N_2529,N_2269,N_2256);
nand U2530 (N_2530,N_2328,N_2215);
or U2531 (N_2531,N_2368,N_2322);
nor U2532 (N_2532,N_2259,N_2319);
and U2533 (N_2533,N_2339,N_2272);
or U2534 (N_2534,N_2266,N_2324);
and U2535 (N_2535,N_2300,N_2298);
or U2536 (N_2536,N_2236,N_2348);
and U2537 (N_2537,N_2217,N_2281);
nor U2538 (N_2538,N_2352,N_2348);
nor U2539 (N_2539,N_2206,N_2316);
and U2540 (N_2540,N_2228,N_2366);
nand U2541 (N_2541,N_2383,N_2362);
nor U2542 (N_2542,N_2232,N_2265);
and U2543 (N_2543,N_2375,N_2392);
and U2544 (N_2544,N_2244,N_2352);
nand U2545 (N_2545,N_2379,N_2392);
nand U2546 (N_2546,N_2212,N_2222);
nor U2547 (N_2547,N_2320,N_2358);
nand U2548 (N_2548,N_2338,N_2395);
nor U2549 (N_2549,N_2314,N_2339);
or U2550 (N_2550,N_2203,N_2241);
nand U2551 (N_2551,N_2203,N_2237);
and U2552 (N_2552,N_2304,N_2220);
and U2553 (N_2553,N_2369,N_2363);
nand U2554 (N_2554,N_2203,N_2234);
nand U2555 (N_2555,N_2363,N_2204);
or U2556 (N_2556,N_2222,N_2258);
nor U2557 (N_2557,N_2370,N_2399);
or U2558 (N_2558,N_2331,N_2204);
and U2559 (N_2559,N_2364,N_2245);
and U2560 (N_2560,N_2254,N_2365);
nand U2561 (N_2561,N_2348,N_2388);
and U2562 (N_2562,N_2336,N_2210);
and U2563 (N_2563,N_2272,N_2228);
and U2564 (N_2564,N_2314,N_2294);
and U2565 (N_2565,N_2227,N_2281);
and U2566 (N_2566,N_2392,N_2374);
nand U2567 (N_2567,N_2387,N_2261);
nor U2568 (N_2568,N_2386,N_2329);
and U2569 (N_2569,N_2323,N_2271);
or U2570 (N_2570,N_2285,N_2331);
and U2571 (N_2571,N_2372,N_2379);
and U2572 (N_2572,N_2234,N_2266);
nor U2573 (N_2573,N_2311,N_2338);
nor U2574 (N_2574,N_2214,N_2394);
nor U2575 (N_2575,N_2269,N_2282);
nand U2576 (N_2576,N_2398,N_2351);
or U2577 (N_2577,N_2334,N_2398);
nor U2578 (N_2578,N_2286,N_2239);
nand U2579 (N_2579,N_2362,N_2295);
nand U2580 (N_2580,N_2242,N_2306);
or U2581 (N_2581,N_2358,N_2327);
nor U2582 (N_2582,N_2210,N_2348);
or U2583 (N_2583,N_2254,N_2210);
and U2584 (N_2584,N_2233,N_2380);
or U2585 (N_2585,N_2220,N_2235);
and U2586 (N_2586,N_2201,N_2292);
nand U2587 (N_2587,N_2387,N_2333);
nor U2588 (N_2588,N_2358,N_2373);
or U2589 (N_2589,N_2395,N_2318);
nor U2590 (N_2590,N_2306,N_2218);
or U2591 (N_2591,N_2353,N_2251);
nand U2592 (N_2592,N_2359,N_2302);
or U2593 (N_2593,N_2218,N_2373);
or U2594 (N_2594,N_2215,N_2202);
nor U2595 (N_2595,N_2211,N_2222);
nand U2596 (N_2596,N_2383,N_2388);
and U2597 (N_2597,N_2232,N_2210);
or U2598 (N_2598,N_2367,N_2250);
nor U2599 (N_2599,N_2377,N_2300);
nor U2600 (N_2600,N_2437,N_2575);
and U2601 (N_2601,N_2582,N_2448);
or U2602 (N_2602,N_2506,N_2441);
or U2603 (N_2603,N_2539,N_2503);
nand U2604 (N_2604,N_2570,N_2598);
nor U2605 (N_2605,N_2561,N_2492);
nand U2606 (N_2606,N_2595,N_2404);
nand U2607 (N_2607,N_2566,N_2593);
nand U2608 (N_2608,N_2471,N_2428);
and U2609 (N_2609,N_2421,N_2535);
and U2610 (N_2610,N_2417,N_2543);
nor U2611 (N_2611,N_2475,N_2466);
nand U2612 (N_2612,N_2559,N_2552);
or U2613 (N_2613,N_2479,N_2555);
and U2614 (N_2614,N_2451,N_2487);
nor U2615 (N_2615,N_2414,N_2517);
nand U2616 (N_2616,N_2569,N_2418);
or U2617 (N_2617,N_2488,N_2528);
nand U2618 (N_2618,N_2591,N_2402);
nor U2619 (N_2619,N_2450,N_2502);
nand U2620 (N_2620,N_2573,N_2519);
or U2621 (N_2621,N_2473,N_2459);
nor U2622 (N_2622,N_2435,N_2438);
or U2623 (N_2623,N_2453,N_2556);
and U2624 (N_2624,N_2589,N_2571);
nor U2625 (N_2625,N_2516,N_2518);
nor U2626 (N_2626,N_2526,N_2544);
nand U2627 (N_2627,N_2538,N_2482);
nor U2628 (N_2628,N_2554,N_2520);
or U2629 (N_2629,N_2588,N_2585);
or U2630 (N_2630,N_2486,N_2449);
nor U2631 (N_2631,N_2424,N_2496);
nand U2632 (N_2632,N_2413,N_2501);
and U2633 (N_2633,N_2423,N_2574);
and U2634 (N_2634,N_2549,N_2599);
nand U2635 (N_2635,N_2587,N_2467);
or U2636 (N_2636,N_2403,N_2465);
nand U2637 (N_2637,N_2509,N_2490);
or U2638 (N_2638,N_2444,N_2411);
or U2639 (N_2639,N_2527,N_2532);
nand U2640 (N_2640,N_2523,N_2495);
nand U2641 (N_2641,N_2463,N_2551);
and U2642 (N_2642,N_2430,N_2415);
nor U2643 (N_2643,N_2489,N_2483);
nand U2644 (N_2644,N_2447,N_2581);
or U2645 (N_2645,N_2420,N_2474);
or U2646 (N_2646,N_2458,N_2578);
and U2647 (N_2647,N_2443,N_2577);
nand U2648 (N_2648,N_2480,N_2550);
and U2649 (N_2649,N_2565,N_2542);
and U2650 (N_2650,N_2477,N_2434);
or U2651 (N_2651,N_2553,N_2514);
and U2652 (N_2652,N_2425,N_2405);
nor U2653 (N_2653,N_2469,N_2512);
or U2654 (N_2654,N_2497,N_2472);
nand U2655 (N_2655,N_2536,N_2427);
and U2656 (N_2656,N_2433,N_2500);
and U2657 (N_2657,N_2562,N_2505);
nor U2658 (N_2658,N_2476,N_2521);
nor U2659 (N_2659,N_2454,N_2510);
or U2660 (N_2660,N_2478,N_2568);
nand U2661 (N_2661,N_2560,N_2586);
nand U2662 (N_2662,N_2592,N_2557);
xnor U2663 (N_2663,N_2432,N_2440);
and U2664 (N_2664,N_2460,N_2445);
or U2665 (N_2665,N_2422,N_2546);
nor U2666 (N_2666,N_2407,N_2409);
nor U2667 (N_2667,N_2590,N_2485);
nand U2668 (N_2668,N_2563,N_2533);
or U2669 (N_2669,N_2456,N_2484);
and U2670 (N_2670,N_2442,N_2494);
nor U2671 (N_2671,N_2596,N_2547);
nor U2672 (N_2672,N_2515,N_2498);
or U2673 (N_2673,N_2491,N_2499);
and U2674 (N_2674,N_2541,N_2493);
and U2675 (N_2675,N_2545,N_2530);
nand U2676 (N_2676,N_2400,N_2576);
nand U2677 (N_2677,N_2548,N_2529);
and U2678 (N_2678,N_2426,N_2419);
and U2679 (N_2679,N_2412,N_2406);
nand U2680 (N_2680,N_2558,N_2584);
nor U2681 (N_2681,N_2522,N_2508);
nand U2682 (N_2682,N_2567,N_2583);
or U2683 (N_2683,N_2534,N_2564);
nand U2684 (N_2684,N_2468,N_2408);
nor U2685 (N_2685,N_2461,N_2525);
nor U2686 (N_2686,N_2531,N_2416);
nand U2687 (N_2687,N_2540,N_2572);
or U2688 (N_2688,N_2511,N_2462);
nor U2689 (N_2689,N_2580,N_2431);
nor U2690 (N_2690,N_2470,N_2457);
nor U2691 (N_2691,N_2597,N_2439);
nand U2692 (N_2692,N_2481,N_2537);
nand U2693 (N_2693,N_2452,N_2594);
and U2694 (N_2694,N_2464,N_2429);
or U2695 (N_2695,N_2513,N_2436);
nand U2696 (N_2696,N_2401,N_2507);
nand U2697 (N_2697,N_2455,N_2410);
and U2698 (N_2698,N_2446,N_2504);
nand U2699 (N_2699,N_2579,N_2524);
nand U2700 (N_2700,N_2410,N_2539);
or U2701 (N_2701,N_2583,N_2566);
xnor U2702 (N_2702,N_2500,N_2546);
nor U2703 (N_2703,N_2414,N_2502);
and U2704 (N_2704,N_2417,N_2581);
and U2705 (N_2705,N_2510,N_2435);
nor U2706 (N_2706,N_2585,N_2519);
nor U2707 (N_2707,N_2434,N_2511);
or U2708 (N_2708,N_2540,N_2403);
or U2709 (N_2709,N_2533,N_2427);
and U2710 (N_2710,N_2506,N_2478);
and U2711 (N_2711,N_2555,N_2543);
nand U2712 (N_2712,N_2558,N_2518);
and U2713 (N_2713,N_2443,N_2583);
and U2714 (N_2714,N_2570,N_2514);
nor U2715 (N_2715,N_2577,N_2432);
nor U2716 (N_2716,N_2494,N_2438);
nor U2717 (N_2717,N_2454,N_2418);
and U2718 (N_2718,N_2409,N_2469);
nand U2719 (N_2719,N_2574,N_2547);
or U2720 (N_2720,N_2416,N_2401);
nand U2721 (N_2721,N_2531,N_2451);
nor U2722 (N_2722,N_2418,N_2534);
nor U2723 (N_2723,N_2518,N_2507);
or U2724 (N_2724,N_2514,N_2419);
or U2725 (N_2725,N_2549,N_2501);
and U2726 (N_2726,N_2498,N_2570);
nor U2727 (N_2727,N_2466,N_2495);
and U2728 (N_2728,N_2552,N_2437);
or U2729 (N_2729,N_2448,N_2470);
and U2730 (N_2730,N_2433,N_2459);
nor U2731 (N_2731,N_2553,N_2533);
nand U2732 (N_2732,N_2470,N_2437);
nand U2733 (N_2733,N_2541,N_2560);
nor U2734 (N_2734,N_2461,N_2526);
and U2735 (N_2735,N_2489,N_2475);
xor U2736 (N_2736,N_2435,N_2460);
nand U2737 (N_2737,N_2413,N_2519);
nand U2738 (N_2738,N_2479,N_2490);
or U2739 (N_2739,N_2538,N_2498);
nor U2740 (N_2740,N_2464,N_2456);
nor U2741 (N_2741,N_2523,N_2546);
or U2742 (N_2742,N_2539,N_2552);
and U2743 (N_2743,N_2467,N_2569);
nor U2744 (N_2744,N_2421,N_2485);
and U2745 (N_2745,N_2565,N_2560);
nand U2746 (N_2746,N_2424,N_2494);
or U2747 (N_2747,N_2434,N_2407);
nand U2748 (N_2748,N_2557,N_2503);
or U2749 (N_2749,N_2481,N_2413);
or U2750 (N_2750,N_2512,N_2572);
nor U2751 (N_2751,N_2431,N_2525);
nor U2752 (N_2752,N_2520,N_2530);
nand U2753 (N_2753,N_2406,N_2447);
nand U2754 (N_2754,N_2508,N_2513);
and U2755 (N_2755,N_2562,N_2544);
and U2756 (N_2756,N_2437,N_2443);
or U2757 (N_2757,N_2408,N_2545);
nand U2758 (N_2758,N_2554,N_2410);
or U2759 (N_2759,N_2445,N_2420);
nor U2760 (N_2760,N_2582,N_2431);
nor U2761 (N_2761,N_2512,N_2574);
or U2762 (N_2762,N_2498,N_2552);
and U2763 (N_2763,N_2570,N_2559);
nand U2764 (N_2764,N_2459,N_2479);
or U2765 (N_2765,N_2564,N_2421);
nand U2766 (N_2766,N_2443,N_2595);
nor U2767 (N_2767,N_2586,N_2444);
or U2768 (N_2768,N_2400,N_2559);
nand U2769 (N_2769,N_2594,N_2537);
and U2770 (N_2770,N_2584,N_2559);
nand U2771 (N_2771,N_2416,N_2480);
or U2772 (N_2772,N_2587,N_2511);
nor U2773 (N_2773,N_2524,N_2462);
nor U2774 (N_2774,N_2472,N_2552);
and U2775 (N_2775,N_2566,N_2576);
nor U2776 (N_2776,N_2459,N_2595);
or U2777 (N_2777,N_2509,N_2469);
nand U2778 (N_2778,N_2445,N_2432);
nor U2779 (N_2779,N_2414,N_2576);
nor U2780 (N_2780,N_2418,N_2570);
nand U2781 (N_2781,N_2549,N_2499);
and U2782 (N_2782,N_2597,N_2525);
and U2783 (N_2783,N_2549,N_2547);
or U2784 (N_2784,N_2457,N_2574);
and U2785 (N_2785,N_2504,N_2461);
or U2786 (N_2786,N_2513,N_2591);
and U2787 (N_2787,N_2436,N_2518);
and U2788 (N_2788,N_2550,N_2563);
or U2789 (N_2789,N_2451,N_2426);
or U2790 (N_2790,N_2563,N_2572);
nand U2791 (N_2791,N_2518,N_2483);
nand U2792 (N_2792,N_2446,N_2518);
or U2793 (N_2793,N_2542,N_2443);
nand U2794 (N_2794,N_2463,N_2426);
nand U2795 (N_2795,N_2514,N_2569);
nor U2796 (N_2796,N_2547,N_2458);
or U2797 (N_2797,N_2401,N_2522);
and U2798 (N_2798,N_2433,N_2525);
or U2799 (N_2799,N_2459,N_2550);
or U2800 (N_2800,N_2680,N_2618);
nand U2801 (N_2801,N_2741,N_2636);
nor U2802 (N_2802,N_2734,N_2639);
xor U2803 (N_2803,N_2656,N_2771);
nor U2804 (N_2804,N_2774,N_2731);
and U2805 (N_2805,N_2772,N_2723);
and U2806 (N_2806,N_2782,N_2726);
or U2807 (N_2807,N_2705,N_2742);
nand U2808 (N_2808,N_2706,N_2709);
nand U2809 (N_2809,N_2681,N_2783);
and U2810 (N_2810,N_2688,N_2780);
nor U2811 (N_2811,N_2630,N_2662);
and U2812 (N_2812,N_2673,N_2665);
or U2813 (N_2813,N_2602,N_2622);
and U2814 (N_2814,N_2744,N_2659);
or U2815 (N_2815,N_2703,N_2762);
and U2816 (N_2816,N_2693,N_2773);
or U2817 (N_2817,N_2788,N_2716);
nor U2818 (N_2818,N_2607,N_2747);
nand U2819 (N_2819,N_2635,N_2672);
or U2820 (N_2820,N_2616,N_2613);
nor U2821 (N_2821,N_2603,N_2696);
and U2822 (N_2822,N_2612,N_2689);
nor U2823 (N_2823,N_2694,N_2752);
nor U2824 (N_2824,N_2751,N_2700);
nand U2825 (N_2825,N_2713,N_2712);
nor U2826 (N_2826,N_2768,N_2617);
nand U2827 (N_2827,N_2701,N_2759);
nand U2828 (N_2828,N_2798,N_2642);
or U2829 (N_2829,N_2609,N_2683);
nand U2830 (N_2830,N_2736,N_2675);
and U2831 (N_2831,N_2753,N_2769);
nand U2832 (N_2832,N_2770,N_2757);
nor U2833 (N_2833,N_2644,N_2685);
or U2834 (N_2834,N_2754,N_2760);
or U2835 (N_2835,N_2614,N_2715);
and U2836 (N_2836,N_2725,N_2748);
and U2837 (N_2837,N_2678,N_2641);
nand U2838 (N_2838,N_2746,N_2648);
and U2839 (N_2839,N_2649,N_2724);
or U2840 (N_2840,N_2745,N_2714);
and U2841 (N_2841,N_2632,N_2755);
nor U2842 (N_2842,N_2796,N_2797);
nand U2843 (N_2843,N_2676,N_2727);
or U2844 (N_2844,N_2652,N_2721);
and U2845 (N_2845,N_2638,N_2664);
nand U2846 (N_2846,N_2695,N_2634);
nand U2847 (N_2847,N_2601,N_2739);
nor U2848 (N_2848,N_2625,N_2795);
nand U2849 (N_2849,N_2657,N_2767);
nor U2850 (N_2850,N_2738,N_2799);
and U2851 (N_2851,N_2667,N_2729);
and U2852 (N_2852,N_2720,N_2779);
and U2853 (N_2853,N_2655,N_2776);
and U2854 (N_2854,N_2697,N_2777);
nand U2855 (N_2855,N_2620,N_2606);
and U2856 (N_2856,N_2784,N_2750);
or U2857 (N_2857,N_2710,N_2669);
nor U2858 (N_2858,N_2698,N_2766);
nand U2859 (N_2859,N_2605,N_2666);
nand U2860 (N_2860,N_2735,N_2728);
xor U2861 (N_2861,N_2781,N_2787);
or U2862 (N_2862,N_2791,N_2692);
or U2863 (N_2863,N_2686,N_2786);
nand U2864 (N_2864,N_2711,N_2790);
nor U2865 (N_2865,N_2624,N_2637);
nand U2866 (N_2866,N_2627,N_2682);
nand U2867 (N_2867,N_2761,N_2619);
nand U2868 (N_2868,N_2704,N_2650);
and U2869 (N_2869,N_2764,N_2792);
and U2870 (N_2870,N_2654,N_2775);
nand U2871 (N_2871,N_2611,N_2633);
or U2872 (N_2872,N_2621,N_2604);
or U2873 (N_2873,N_2658,N_2737);
nor U2874 (N_2874,N_2749,N_2743);
and U2875 (N_2875,N_2793,N_2629);
nor U2876 (N_2876,N_2719,N_2785);
nand U2877 (N_2877,N_2702,N_2668);
nand U2878 (N_2878,N_2679,N_2718);
nor U2879 (N_2879,N_2756,N_2643);
nor U2880 (N_2880,N_2626,N_2647);
nand U2881 (N_2881,N_2687,N_2730);
and U2882 (N_2882,N_2663,N_2653);
nand U2883 (N_2883,N_2758,N_2684);
nor U2884 (N_2884,N_2740,N_2651);
or U2885 (N_2885,N_2660,N_2646);
nand U2886 (N_2886,N_2623,N_2699);
nand U2887 (N_2887,N_2628,N_2661);
nor U2888 (N_2888,N_2690,N_2671);
nand U2889 (N_2889,N_2732,N_2640);
nor U2890 (N_2890,N_2765,N_2707);
nor U2891 (N_2891,N_2645,N_2691);
nor U2892 (N_2892,N_2670,N_2789);
and U2893 (N_2893,N_2708,N_2615);
and U2894 (N_2894,N_2794,N_2674);
and U2895 (N_2895,N_2631,N_2763);
or U2896 (N_2896,N_2722,N_2610);
nor U2897 (N_2897,N_2600,N_2608);
nor U2898 (N_2898,N_2733,N_2677);
or U2899 (N_2899,N_2778,N_2717);
nor U2900 (N_2900,N_2632,N_2601);
and U2901 (N_2901,N_2790,N_2752);
nand U2902 (N_2902,N_2636,N_2789);
nor U2903 (N_2903,N_2771,N_2631);
nor U2904 (N_2904,N_2796,N_2637);
nor U2905 (N_2905,N_2781,N_2732);
nor U2906 (N_2906,N_2607,N_2639);
or U2907 (N_2907,N_2627,N_2674);
and U2908 (N_2908,N_2604,N_2646);
and U2909 (N_2909,N_2773,N_2695);
or U2910 (N_2910,N_2670,N_2759);
nand U2911 (N_2911,N_2749,N_2612);
and U2912 (N_2912,N_2724,N_2689);
and U2913 (N_2913,N_2692,N_2765);
nand U2914 (N_2914,N_2638,N_2697);
and U2915 (N_2915,N_2665,N_2609);
nand U2916 (N_2916,N_2639,N_2686);
or U2917 (N_2917,N_2786,N_2767);
nor U2918 (N_2918,N_2634,N_2698);
nor U2919 (N_2919,N_2648,N_2671);
nand U2920 (N_2920,N_2611,N_2648);
and U2921 (N_2921,N_2748,N_2741);
or U2922 (N_2922,N_2722,N_2729);
and U2923 (N_2923,N_2786,N_2783);
nor U2924 (N_2924,N_2700,N_2693);
and U2925 (N_2925,N_2675,N_2789);
or U2926 (N_2926,N_2726,N_2686);
and U2927 (N_2927,N_2784,N_2677);
nor U2928 (N_2928,N_2668,N_2754);
nor U2929 (N_2929,N_2763,N_2641);
nand U2930 (N_2930,N_2798,N_2711);
nor U2931 (N_2931,N_2734,N_2702);
or U2932 (N_2932,N_2747,N_2774);
and U2933 (N_2933,N_2797,N_2656);
nor U2934 (N_2934,N_2622,N_2690);
or U2935 (N_2935,N_2663,N_2717);
nor U2936 (N_2936,N_2672,N_2666);
nor U2937 (N_2937,N_2734,N_2601);
and U2938 (N_2938,N_2600,N_2621);
nand U2939 (N_2939,N_2660,N_2656);
or U2940 (N_2940,N_2702,N_2721);
xnor U2941 (N_2941,N_2752,N_2606);
nand U2942 (N_2942,N_2733,N_2676);
nand U2943 (N_2943,N_2792,N_2737);
or U2944 (N_2944,N_2780,N_2713);
and U2945 (N_2945,N_2763,N_2745);
and U2946 (N_2946,N_2679,N_2729);
and U2947 (N_2947,N_2692,N_2628);
or U2948 (N_2948,N_2777,N_2711);
or U2949 (N_2949,N_2626,N_2747);
or U2950 (N_2950,N_2676,N_2784);
nor U2951 (N_2951,N_2701,N_2601);
or U2952 (N_2952,N_2647,N_2693);
and U2953 (N_2953,N_2702,N_2762);
or U2954 (N_2954,N_2682,N_2677);
and U2955 (N_2955,N_2608,N_2674);
nor U2956 (N_2956,N_2761,N_2679);
and U2957 (N_2957,N_2798,N_2694);
xnor U2958 (N_2958,N_2792,N_2682);
and U2959 (N_2959,N_2708,N_2664);
nand U2960 (N_2960,N_2716,N_2636);
and U2961 (N_2961,N_2735,N_2727);
nor U2962 (N_2962,N_2617,N_2722);
nor U2963 (N_2963,N_2681,N_2788);
and U2964 (N_2964,N_2673,N_2656);
nand U2965 (N_2965,N_2631,N_2776);
nor U2966 (N_2966,N_2748,N_2735);
nand U2967 (N_2967,N_2708,N_2606);
nor U2968 (N_2968,N_2787,N_2635);
and U2969 (N_2969,N_2696,N_2656);
nor U2970 (N_2970,N_2687,N_2710);
nand U2971 (N_2971,N_2646,N_2720);
and U2972 (N_2972,N_2757,N_2662);
or U2973 (N_2973,N_2770,N_2675);
nor U2974 (N_2974,N_2764,N_2619);
and U2975 (N_2975,N_2701,N_2669);
nand U2976 (N_2976,N_2623,N_2784);
nand U2977 (N_2977,N_2603,N_2682);
nor U2978 (N_2978,N_2772,N_2680);
nor U2979 (N_2979,N_2617,N_2737);
nand U2980 (N_2980,N_2646,N_2618);
nand U2981 (N_2981,N_2711,N_2782);
or U2982 (N_2982,N_2712,N_2777);
nor U2983 (N_2983,N_2775,N_2736);
nand U2984 (N_2984,N_2784,N_2647);
and U2985 (N_2985,N_2778,N_2650);
or U2986 (N_2986,N_2747,N_2627);
and U2987 (N_2987,N_2689,N_2653);
or U2988 (N_2988,N_2698,N_2744);
nor U2989 (N_2989,N_2760,N_2763);
or U2990 (N_2990,N_2763,N_2623);
or U2991 (N_2991,N_2791,N_2735);
and U2992 (N_2992,N_2736,N_2755);
or U2993 (N_2993,N_2612,N_2787);
or U2994 (N_2994,N_2670,N_2749);
and U2995 (N_2995,N_2688,N_2756);
nand U2996 (N_2996,N_2638,N_2609);
and U2997 (N_2997,N_2776,N_2755);
and U2998 (N_2998,N_2675,N_2793);
or U2999 (N_2999,N_2773,N_2642);
and UO_0 (O_0,N_2950,N_2823);
or UO_1 (O_1,N_2843,N_2824);
nor UO_2 (O_2,N_2967,N_2826);
nand UO_3 (O_3,N_2845,N_2833);
or UO_4 (O_4,N_2949,N_2985);
nor UO_5 (O_5,N_2954,N_2996);
nor UO_6 (O_6,N_2803,N_2986);
or UO_7 (O_7,N_2841,N_2957);
nor UO_8 (O_8,N_2953,N_2972);
nor UO_9 (O_9,N_2887,N_2875);
or UO_10 (O_10,N_2800,N_2931);
nand UO_11 (O_11,N_2825,N_2910);
nor UO_12 (O_12,N_2956,N_2854);
nor UO_13 (O_13,N_2959,N_2849);
nor UO_14 (O_14,N_2810,N_2816);
or UO_15 (O_15,N_2888,N_2905);
nor UO_16 (O_16,N_2869,N_2817);
and UO_17 (O_17,N_2873,N_2928);
nand UO_18 (O_18,N_2966,N_2984);
and UO_19 (O_19,N_2885,N_2999);
nand UO_20 (O_20,N_2813,N_2870);
nor UO_21 (O_21,N_2815,N_2915);
nand UO_22 (O_22,N_2937,N_2947);
and UO_23 (O_23,N_2912,N_2983);
or UO_24 (O_24,N_2866,N_2840);
or UO_25 (O_25,N_2934,N_2863);
nor UO_26 (O_26,N_2926,N_2965);
or UO_27 (O_27,N_2846,N_2877);
nand UO_28 (O_28,N_2917,N_2970);
or UO_29 (O_29,N_2804,N_2860);
or UO_30 (O_30,N_2933,N_2998);
and UO_31 (O_31,N_2939,N_2829);
nor UO_32 (O_32,N_2922,N_2898);
nand UO_33 (O_33,N_2837,N_2871);
and UO_34 (O_34,N_2878,N_2818);
nor UO_35 (O_35,N_2913,N_2955);
and UO_36 (O_36,N_2918,N_2856);
and UO_37 (O_37,N_2951,N_2889);
nor UO_38 (O_38,N_2971,N_2831);
or UO_39 (O_39,N_2944,N_2835);
or UO_40 (O_40,N_2975,N_2806);
and UO_41 (O_41,N_2808,N_2991);
nand UO_42 (O_42,N_2914,N_2881);
nand UO_43 (O_43,N_2839,N_2852);
nand UO_44 (O_44,N_2894,N_2995);
nand UO_45 (O_45,N_2807,N_2962);
nor UO_46 (O_46,N_2946,N_2897);
nor UO_47 (O_47,N_2925,N_2805);
nor UO_48 (O_48,N_2921,N_2874);
or UO_49 (O_49,N_2900,N_2936);
or UO_50 (O_50,N_2819,N_2961);
nor UO_51 (O_51,N_2916,N_2893);
and UO_52 (O_52,N_2847,N_2960);
nand UO_53 (O_53,N_2923,N_2963);
nor UO_54 (O_54,N_2978,N_2976);
or UO_55 (O_55,N_2990,N_2822);
nor UO_56 (O_56,N_2872,N_2989);
nor UO_57 (O_57,N_2908,N_2836);
nor UO_58 (O_58,N_2828,N_2904);
nor UO_59 (O_59,N_2958,N_2882);
or UO_60 (O_60,N_2974,N_2838);
nor UO_61 (O_61,N_2834,N_2935);
or UO_62 (O_62,N_2920,N_2994);
or UO_63 (O_63,N_2842,N_2919);
nand UO_64 (O_64,N_2940,N_2832);
nand UO_65 (O_65,N_2941,N_2830);
nand UO_66 (O_66,N_2848,N_2858);
and UO_67 (O_67,N_2902,N_2820);
nor UO_68 (O_68,N_2930,N_2886);
nand UO_69 (O_69,N_2968,N_2880);
and UO_70 (O_70,N_2993,N_2884);
nor UO_71 (O_71,N_2977,N_2979);
or UO_72 (O_72,N_2883,N_2906);
and UO_73 (O_73,N_2868,N_2851);
and UO_74 (O_74,N_2855,N_2827);
and UO_75 (O_75,N_2987,N_2988);
or UO_76 (O_76,N_2865,N_2899);
or UO_77 (O_77,N_2814,N_2945);
nand UO_78 (O_78,N_2911,N_2907);
or UO_79 (O_79,N_2901,N_2844);
and UO_80 (O_80,N_2943,N_2867);
nand UO_81 (O_81,N_2811,N_2862);
nand UO_82 (O_82,N_2876,N_2992);
or UO_83 (O_83,N_2850,N_2809);
nand UO_84 (O_84,N_2859,N_2821);
nand UO_85 (O_85,N_2857,N_2890);
and UO_86 (O_86,N_2948,N_2982);
or UO_87 (O_87,N_2801,N_2891);
and UO_88 (O_88,N_2864,N_2909);
nand UO_89 (O_89,N_2927,N_2879);
nand UO_90 (O_90,N_2964,N_2892);
or UO_91 (O_91,N_2895,N_2812);
and UO_92 (O_92,N_2973,N_2981);
nor UO_93 (O_93,N_2924,N_2861);
or UO_94 (O_94,N_2980,N_2802);
and UO_95 (O_95,N_2896,N_2903);
and UO_96 (O_96,N_2853,N_2942);
or UO_97 (O_97,N_2969,N_2929);
nor UO_98 (O_98,N_2938,N_2997);
nand UO_99 (O_99,N_2952,N_2932);
nor UO_100 (O_100,N_2805,N_2851);
nand UO_101 (O_101,N_2879,N_2965);
and UO_102 (O_102,N_2920,N_2889);
nor UO_103 (O_103,N_2914,N_2964);
or UO_104 (O_104,N_2963,N_2999);
nor UO_105 (O_105,N_2814,N_2813);
or UO_106 (O_106,N_2882,N_2987);
nor UO_107 (O_107,N_2909,N_2942);
nor UO_108 (O_108,N_2983,N_2842);
nand UO_109 (O_109,N_2808,N_2823);
nor UO_110 (O_110,N_2854,N_2898);
nand UO_111 (O_111,N_2907,N_2818);
nor UO_112 (O_112,N_2937,N_2895);
or UO_113 (O_113,N_2884,N_2914);
nor UO_114 (O_114,N_2863,N_2898);
or UO_115 (O_115,N_2991,N_2969);
and UO_116 (O_116,N_2895,N_2936);
and UO_117 (O_117,N_2832,N_2914);
or UO_118 (O_118,N_2967,N_2996);
and UO_119 (O_119,N_2879,N_2816);
nor UO_120 (O_120,N_2946,N_2829);
nor UO_121 (O_121,N_2910,N_2854);
nand UO_122 (O_122,N_2869,N_2998);
nor UO_123 (O_123,N_2816,N_2971);
or UO_124 (O_124,N_2942,N_2994);
nor UO_125 (O_125,N_2913,N_2820);
nand UO_126 (O_126,N_2934,N_2875);
or UO_127 (O_127,N_2816,N_2924);
and UO_128 (O_128,N_2951,N_2882);
or UO_129 (O_129,N_2815,N_2801);
nand UO_130 (O_130,N_2848,N_2977);
or UO_131 (O_131,N_2913,N_2878);
or UO_132 (O_132,N_2854,N_2870);
nor UO_133 (O_133,N_2927,N_2874);
or UO_134 (O_134,N_2846,N_2864);
and UO_135 (O_135,N_2907,N_2859);
nor UO_136 (O_136,N_2898,N_2938);
or UO_137 (O_137,N_2951,N_2911);
and UO_138 (O_138,N_2946,N_2833);
or UO_139 (O_139,N_2965,N_2927);
or UO_140 (O_140,N_2882,N_2807);
nor UO_141 (O_141,N_2991,N_2966);
and UO_142 (O_142,N_2936,N_2969);
and UO_143 (O_143,N_2887,N_2940);
and UO_144 (O_144,N_2999,N_2862);
and UO_145 (O_145,N_2931,N_2806);
or UO_146 (O_146,N_2980,N_2807);
nand UO_147 (O_147,N_2892,N_2811);
nand UO_148 (O_148,N_2816,N_2934);
and UO_149 (O_149,N_2961,N_2878);
and UO_150 (O_150,N_2871,N_2942);
nand UO_151 (O_151,N_2948,N_2996);
or UO_152 (O_152,N_2819,N_2816);
or UO_153 (O_153,N_2851,N_2948);
and UO_154 (O_154,N_2856,N_2812);
nand UO_155 (O_155,N_2898,N_2951);
nand UO_156 (O_156,N_2891,N_2959);
and UO_157 (O_157,N_2878,N_2989);
nand UO_158 (O_158,N_2932,N_2958);
and UO_159 (O_159,N_2912,N_2822);
and UO_160 (O_160,N_2905,N_2807);
or UO_161 (O_161,N_2960,N_2856);
nor UO_162 (O_162,N_2827,N_2838);
nor UO_163 (O_163,N_2846,N_2889);
or UO_164 (O_164,N_2904,N_2901);
or UO_165 (O_165,N_2999,N_2948);
xnor UO_166 (O_166,N_2895,N_2848);
and UO_167 (O_167,N_2893,N_2845);
or UO_168 (O_168,N_2898,N_2916);
and UO_169 (O_169,N_2898,N_2892);
and UO_170 (O_170,N_2862,N_2997);
nor UO_171 (O_171,N_2967,N_2907);
and UO_172 (O_172,N_2809,N_2987);
and UO_173 (O_173,N_2969,N_2813);
and UO_174 (O_174,N_2814,N_2870);
or UO_175 (O_175,N_2993,N_2967);
or UO_176 (O_176,N_2805,N_2910);
nor UO_177 (O_177,N_2907,N_2993);
or UO_178 (O_178,N_2960,N_2902);
nor UO_179 (O_179,N_2857,N_2959);
nor UO_180 (O_180,N_2992,N_2965);
and UO_181 (O_181,N_2876,N_2939);
nor UO_182 (O_182,N_2919,N_2867);
or UO_183 (O_183,N_2841,N_2854);
nand UO_184 (O_184,N_2989,N_2856);
and UO_185 (O_185,N_2927,N_2979);
and UO_186 (O_186,N_2944,N_2837);
or UO_187 (O_187,N_2913,N_2943);
nand UO_188 (O_188,N_2863,N_2976);
nand UO_189 (O_189,N_2942,N_2968);
or UO_190 (O_190,N_2985,N_2973);
nand UO_191 (O_191,N_2856,N_2888);
or UO_192 (O_192,N_2892,N_2954);
nand UO_193 (O_193,N_2964,N_2869);
nor UO_194 (O_194,N_2851,N_2939);
and UO_195 (O_195,N_2802,N_2915);
nand UO_196 (O_196,N_2922,N_2962);
nor UO_197 (O_197,N_2948,N_2990);
nor UO_198 (O_198,N_2901,N_2810);
nand UO_199 (O_199,N_2910,N_2997);
nor UO_200 (O_200,N_2998,N_2913);
or UO_201 (O_201,N_2805,N_2868);
nand UO_202 (O_202,N_2996,N_2874);
or UO_203 (O_203,N_2980,N_2895);
nand UO_204 (O_204,N_2972,N_2841);
or UO_205 (O_205,N_2918,N_2928);
nor UO_206 (O_206,N_2905,N_2922);
nor UO_207 (O_207,N_2980,N_2846);
nand UO_208 (O_208,N_2829,N_2854);
and UO_209 (O_209,N_2946,N_2817);
nor UO_210 (O_210,N_2829,N_2983);
nor UO_211 (O_211,N_2976,N_2815);
or UO_212 (O_212,N_2931,N_2948);
nor UO_213 (O_213,N_2979,N_2880);
nor UO_214 (O_214,N_2894,N_2974);
nand UO_215 (O_215,N_2902,N_2913);
and UO_216 (O_216,N_2800,N_2945);
and UO_217 (O_217,N_2841,N_2923);
and UO_218 (O_218,N_2889,N_2973);
or UO_219 (O_219,N_2853,N_2988);
nor UO_220 (O_220,N_2877,N_2929);
nand UO_221 (O_221,N_2926,N_2853);
or UO_222 (O_222,N_2802,N_2975);
nor UO_223 (O_223,N_2814,N_2970);
nor UO_224 (O_224,N_2948,N_2904);
xnor UO_225 (O_225,N_2866,N_2995);
nor UO_226 (O_226,N_2899,N_2844);
or UO_227 (O_227,N_2800,N_2802);
and UO_228 (O_228,N_2872,N_2888);
nor UO_229 (O_229,N_2997,N_2845);
nand UO_230 (O_230,N_2976,N_2870);
and UO_231 (O_231,N_2847,N_2875);
and UO_232 (O_232,N_2971,N_2920);
nor UO_233 (O_233,N_2873,N_2917);
or UO_234 (O_234,N_2973,N_2824);
nor UO_235 (O_235,N_2841,N_2956);
nor UO_236 (O_236,N_2962,N_2933);
or UO_237 (O_237,N_2880,N_2868);
and UO_238 (O_238,N_2908,N_2851);
or UO_239 (O_239,N_2886,N_2828);
and UO_240 (O_240,N_2864,N_2930);
nor UO_241 (O_241,N_2871,N_2838);
nor UO_242 (O_242,N_2932,N_2812);
nor UO_243 (O_243,N_2912,N_2978);
nor UO_244 (O_244,N_2989,N_2827);
nor UO_245 (O_245,N_2840,N_2965);
and UO_246 (O_246,N_2934,N_2865);
or UO_247 (O_247,N_2994,N_2988);
and UO_248 (O_248,N_2974,N_2977);
and UO_249 (O_249,N_2851,N_2850);
nor UO_250 (O_250,N_2910,N_2818);
or UO_251 (O_251,N_2938,N_2950);
nand UO_252 (O_252,N_2898,N_2877);
nor UO_253 (O_253,N_2996,N_2977);
nand UO_254 (O_254,N_2806,N_2903);
or UO_255 (O_255,N_2889,N_2959);
nand UO_256 (O_256,N_2858,N_2966);
or UO_257 (O_257,N_2841,N_2992);
nand UO_258 (O_258,N_2856,N_2870);
xor UO_259 (O_259,N_2824,N_2965);
nor UO_260 (O_260,N_2834,N_2978);
nor UO_261 (O_261,N_2897,N_2985);
nand UO_262 (O_262,N_2953,N_2905);
or UO_263 (O_263,N_2940,N_2918);
and UO_264 (O_264,N_2812,N_2914);
nor UO_265 (O_265,N_2996,N_2941);
nand UO_266 (O_266,N_2803,N_2890);
or UO_267 (O_267,N_2958,N_2862);
or UO_268 (O_268,N_2858,N_2884);
nor UO_269 (O_269,N_2981,N_2877);
nand UO_270 (O_270,N_2934,N_2881);
or UO_271 (O_271,N_2842,N_2896);
and UO_272 (O_272,N_2924,N_2856);
nor UO_273 (O_273,N_2886,N_2960);
nor UO_274 (O_274,N_2921,N_2977);
nand UO_275 (O_275,N_2802,N_2901);
or UO_276 (O_276,N_2959,N_2962);
nor UO_277 (O_277,N_2814,N_2855);
or UO_278 (O_278,N_2976,N_2889);
or UO_279 (O_279,N_2992,N_2912);
nand UO_280 (O_280,N_2847,N_2989);
and UO_281 (O_281,N_2912,N_2996);
nor UO_282 (O_282,N_2904,N_2910);
nand UO_283 (O_283,N_2813,N_2858);
nand UO_284 (O_284,N_2817,N_2986);
nor UO_285 (O_285,N_2841,N_2981);
nand UO_286 (O_286,N_2941,N_2925);
nor UO_287 (O_287,N_2929,N_2837);
and UO_288 (O_288,N_2910,N_2918);
nor UO_289 (O_289,N_2858,N_2839);
nor UO_290 (O_290,N_2915,N_2868);
or UO_291 (O_291,N_2846,N_2817);
or UO_292 (O_292,N_2960,N_2948);
and UO_293 (O_293,N_2889,N_2867);
or UO_294 (O_294,N_2908,N_2872);
nor UO_295 (O_295,N_2872,N_2868);
nor UO_296 (O_296,N_2948,N_2834);
and UO_297 (O_297,N_2887,N_2872);
or UO_298 (O_298,N_2919,N_2822);
and UO_299 (O_299,N_2891,N_2936);
nand UO_300 (O_300,N_2884,N_2910);
nor UO_301 (O_301,N_2951,N_2944);
and UO_302 (O_302,N_2865,N_2946);
nor UO_303 (O_303,N_2848,N_2999);
nand UO_304 (O_304,N_2959,N_2856);
and UO_305 (O_305,N_2870,N_2855);
nor UO_306 (O_306,N_2971,N_2863);
nor UO_307 (O_307,N_2814,N_2869);
nand UO_308 (O_308,N_2978,N_2839);
nand UO_309 (O_309,N_2869,N_2812);
nand UO_310 (O_310,N_2931,N_2989);
nor UO_311 (O_311,N_2930,N_2820);
nor UO_312 (O_312,N_2802,N_2811);
and UO_313 (O_313,N_2835,N_2910);
nor UO_314 (O_314,N_2887,N_2867);
nand UO_315 (O_315,N_2909,N_2938);
and UO_316 (O_316,N_2813,N_2901);
or UO_317 (O_317,N_2843,N_2900);
nor UO_318 (O_318,N_2936,N_2857);
nand UO_319 (O_319,N_2894,N_2998);
or UO_320 (O_320,N_2865,N_2973);
and UO_321 (O_321,N_2983,N_2950);
nand UO_322 (O_322,N_2820,N_2994);
and UO_323 (O_323,N_2953,N_2980);
or UO_324 (O_324,N_2978,N_2911);
nand UO_325 (O_325,N_2808,N_2873);
xor UO_326 (O_326,N_2999,N_2942);
nor UO_327 (O_327,N_2836,N_2991);
nand UO_328 (O_328,N_2807,N_2982);
nand UO_329 (O_329,N_2851,N_2888);
or UO_330 (O_330,N_2912,N_2977);
nand UO_331 (O_331,N_2847,N_2899);
nor UO_332 (O_332,N_2836,N_2976);
nor UO_333 (O_333,N_2980,N_2848);
and UO_334 (O_334,N_2910,N_2868);
nor UO_335 (O_335,N_2880,N_2903);
and UO_336 (O_336,N_2810,N_2904);
or UO_337 (O_337,N_2930,N_2813);
or UO_338 (O_338,N_2926,N_2813);
and UO_339 (O_339,N_2863,N_2979);
and UO_340 (O_340,N_2945,N_2907);
nand UO_341 (O_341,N_2837,N_2935);
nor UO_342 (O_342,N_2998,N_2995);
or UO_343 (O_343,N_2918,N_2820);
and UO_344 (O_344,N_2947,N_2831);
or UO_345 (O_345,N_2979,N_2941);
or UO_346 (O_346,N_2810,N_2802);
and UO_347 (O_347,N_2846,N_2935);
and UO_348 (O_348,N_2952,N_2866);
nor UO_349 (O_349,N_2909,N_2971);
nor UO_350 (O_350,N_2920,N_2977);
nand UO_351 (O_351,N_2841,N_2905);
or UO_352 (O_352,N_2944,N_2840);
or UO_353 (O_353,N_2815,N_2802);
nor UO_354 (O_354,N_2918,N_2970);
nor UO_355 (O_355,N_2839,N_2933);
and UO_356 (O_356,N_2960,N_2868);
nand UO_357 (O_357,N_2851,N_2926);
and UO_358 (O_358,N_2821,N_2974);
nor UO_359 (O_359,N_2976,N_2921);
and UO_360 (O_360,N_2948,N_2837);
nor UO_361 (O_361,N_2928,N_2910);
or UO_362 (O_362,N_2871,N_2888);
and UO_363 (O_363,N_2812,N_2994);
xnor UO_364 (O_364,N_2893,N_2968);
or UO_365 (O_365,N_2901,N_2865);
or UO_366 (O_366,N_2835,N_2862);
nand UO_367 (O_367,N_2995,N_2898);
or UO_368 (O_368,N_2827,N_2836);
and UO_369 (O_369,N_2897,N_2962);
and UO_370 (O_370,N_2967,N_2974);
nor UO_371 (O_371,N_2856,N_2895);
and UO_372 (O_372,N_2962,N_2916);
xor UO_373 (O_373,N_2897,N_2981);
or UO_374 (O_374,N_2999,N_2975);
nor UO_375 (O_375,N_2946,N_2886);
nor UO_376 (O_376,N_2921,N_2901);
nor UO_377 (O_377,N_2923,N_2898);
nor UO_378 (O_378,N_2803,N_2946);
nor UO_379 (O_379,N_2842,N_2985);
nand UO_380 (O_380,N_2916,N_2829);
nor UO_381 (O_381,N_2983,N_2852);
nor UO_382 (O_382,N_2976,N_2959);
or UO_383 (O_383,N_2968,N_2904);
and UO_384 (O_384,N_2872,N_2856);
nand UO_385 (O_385,N_2983,N_2810);
nand UO_386 (O_386,N_2809,N_2965);
xnor UO_387 (O_387,N_2988,N_2873);
nand UO_388 (O_388,N_2992,N_2888);
or UO_389 (O_389,N_2886,N_2881);
nor UO_390 (O_390,N_2819,N_2900);
and UO_391 (O_391,N_2953,N_2931);
nor UO_392 (O_392,N_2853,N_2880);
and UO_393 (O_393,N_2862,N_2894);
and UO_394 (O_394,N_2881,N_2977);
and UO_395 (O_395,N_2992,N_2971);
or UO_396 (O_396,N_2957,N_2945);
or UO_397 (O_397,N_2971,N_2819);
nor UO_398 (O_398,N_2948,N_2890);
and UO_399 (O_399,N_2875,N_2949);
and UO_400 (O_400,N_2975,N_2974);
or UO_401 (O_401,N_2896,N_2897);
and UO_402 (O_402,N_2954,N_2957);
nand UO_403 (O_403,N_2970,N_2890);
or UO_404 (O_404,N_2817,N_2839);
and UO_405 (O_405,N_2974,N_2949);
nand UO_406 (O_406,N_2955,N_2886);
and UO_407 (O_407,N_2830,N_2869);
and UO_408 (O_408,N_2929,N_2945);
nand UO_409 (O_409,N_2805,N_2963);
and UO_410 (O_410,N_2829,N_2868);
nand UO_411 (O_411,N_2965,N_2898);
nand UO_412 (O_412,N_2801,N_2925);
or UO_413 (O_413,N_2874,N_2809);
nand UO_414 (O_414,N_2950,N_2880);
nand UO_415 (O_415,N_2852,N_2876);
nor UO_416 (O_416,N_2908,N_2964);
nand UO_417 (O_417,N_2974,N_2871);
and UO_418 (O_418,N_2931,N_2908);
and UO_419 (O_419,N_2987,N_2877);
or UO_420 (O_420,N_2829,N_2974);
nor UO_421 (O_421,N_2831,N_2824);
or UO_422 (O_422,N_2927,N_2897);
nand UO_423 (O_423,N_2962,N_2927);
nor UO_424 (O_424,N_2950,N_2820);
nor UO_425 (O_425,N_2944,N_2816);
or UO_426 (O_426,N_2974,N_2999);
nor UO_427 (O_427,N_2976,N_2967);
and UO_428 (O_428,N_2844,N_2828);
and UO_429 (O_429,N_2939,N_2964);
or UO_430 (O_430,N_2869,N_2805);
nor UO_431 (O_431,N_2849,N_2901);
nand UO_432 (O_432,N_2900,N_2944);
and UO_433 (O_433,N_2947,N_2818);
or UO_434 (O_434,N_2922,N_2812);
or UO_435 (O_435,N_2896,N_2893);
or UO_436 (O_436,N_2980,N_2925);
or UO_437 (O_437,N_2888,N_2821);
and UO_438 (O_438,N_2901,N_2897);
or UO_439 (O_439,N_2966,N_2853);
nand UO_440 (O_440,N_2838,N_2923);
and UO_441 (O_441,N_2991,N_2951);
or UO_442 (O_442,N_2804,N_2940);
and UO_443 (O_443,N_2877,N_2856);
or UO_444 (O_444,N_2838,N_2927);
nor UO_445 (O_445,N_2938,N_2925);
nand UO_446 (O_446,N_2848,N_2954);
or UO_447 (O_447,N_2969,N_2985);
and UO_448 (O_448,N_2924,N_2869);
and UO_449 (O_449,N_2988,N_2891);
or UO_450 (O_450,N_2839,N_2895);
xnor UO_451 (O_451,N_2806,N_2820);
nor UO_452 (O_452,N_2972,N_2836);
nand UO_453 (O_453,N_2959,N_2921);
and UO_454 (O_454,N_2897,N_2850);
or UO_455 (O_455,N_2950,N_2835);
nor UO_456 (O_456,N_2977,N_2844);
or UO_457 (O_457,N_2954,N_2829);
or UO_458 (O_458,N_2815,N_2975);
nand UO_459 (O_459,N_2911,N_2891);
nand UO_460 (O_460,N_2913,N_2824);
and UO_461 (O_461,N_2887,N_2821);
or UO_462 (O_462,N_2859,N_2815);
nand UO_463 (O_463,N_2919,N_2838);
nand UO_464 (O_464,N_2962,N_2949);
or UO_465 (O_465,N_2809,N_2972);
or UO_466 (O_466,N_2881,N_2923);
nor UO_467 (O_467,N_2971,N_2883);
nand UO_468 (O_468,N_2938,N_2844);
or UO_469 (O_469,N_2976,N_2990);
nand UO_470 (O_470,N_2937,N_2946);
or UO_471 (O_471,N_2874,N_2871);
or UO_472 (O_472,N_2805,N_2945);
nor UO_473 (O_473,N_2950,N_2854);
nand UO_474 (O_474,N_2890,N_2935);
and UO_475 (O_475,N_2891,N_2895);
nand UO_476 (O_476,N_2806,N_2817);
nand UO_477 (O_477,N_2806,N_2899);
and UO_478 (O_478,N_2964,N_2901);
or UO_479 (O_479,N_2816,N_2932);
nor UO_480 (O_480,N_2841,N_2940);
or UO_481 (O_481,N_2993,N_2991);
and UO_482 (O_482,N_2835,N_2831);
or UO_483 (O_483,N_2814,N_2878);
nor UO_484 (O_484,N_2811,N_2969);
or UO_485 (O_485,N_2817,N_2811);
or UO_486 (O_486,N_2904,N_2820);
and UO_487 (O_487,N_2914,N_2998);
or UO_488 (O_488,N_2927,N_2884);
nand UO_489 (O_489,N_2906,N_2932);
nor UO_490 (O_490,N_2986,N_2867);
nand UO_491 (O_491,N_2920,N_2936);
or UO_492 (O_492,N_2840,N_2849);
and UO_493 (O_493,N_2875,N_2884);
nand UO_494 (O_494,N_2950,N_2984);
nor UO_495 (O_495,N_2903,N_2878);
nand UO_496 (O_496,N_2844,N_2987);
or UO_497 (O_497,N_2933,N_2808);
nor UO_498 (O_498,N_2834,N_2992);
xnor UO_499 (O_499,N_2823,N_2887);
endmodule