module basic_2000_20000_2500_125_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1588,In_1142);
and U1 (N_1,In_1636,In_1444);
xor U2 (N_2,In_1420,In_256);
nor U3 (N_3,In_656,In_1885);
or U4 (N_4,In_1982,In_311);
nand U5 (N_5,In_1764,In_1572);
nor U6 (N_6,In_419,In_1864);
nand U7 (N_7,In_258,In_423);
nand U8 (N_8,In_1274,In_39);
xnor U9 (N_9,In_370,In_1539);
nor U10 (N_10,In_1030,In_1309);
or U11 (N_11,In_9,In_1072);
or U12 (N_12,In_1580,In_797);
nor U13 (N_13,In_587,In_88);
and U14 (N_14,In_1323,In_1753);
and U15 (N_15,In_801,In_457);
nand U16 (N_16,In_1369,In_774);
nor U17 (N_17,In_545,In_23);
nor U18 (N_18,In_873,In_721);
xor U19 (N_19,In_818,In_572);
nor U20 (N_20,In_1029,In_1766);
xor U21 (N_21,In_672,In_487);
nor U22 (N_22,In_1715,In_1961);
or U23 (N_23,In_593,In_1952);
and U24 (N_24,In_1288,In_1617);
xnor U25 (N_25,In_1640,In_289);
nor U26 (N_26,In_1631,In_697);
nor U27 (N_27,In_984,In_1249);
xnor U28 (N_28,In_1095,In_249);
and U29 (N_29,In_1910,In_1165);
nand U30 (N_30,In_1209,In_1226);
or U31 (N_31,In_817,In_956);
xnor U32 (N_32,In_518,In_1166);
and U33 (N_33,In_1360,In_3);
xnor U34 (N_34,In_1125,In_1990);
nand U35 (N_35,In_946,In_1428);
or U36 (N_36,In_563,In_1007);
and U37 (N_37,In_1219,In_385);
nand U38 (N_38,In_1550,In_47);
xnor U39 (N_39,In_1692,In_627);
and U40 (N_40,In_1293,In_1198);
nand U41 (N_41,In_283,In_1423);
and U42 (N_42,In_1737,In_1892);
nand U43 (N_43,In_1181,In_1683);
or U44 (N_44,In_867,In_1571);
nor U45 (N_45,In_1242,In_1739);
or U46 (N_46,In_471,In_167);
xnor U47 (N_47,In_55,In_323);
nor U48 (N_48,In_706,In_241);
nand U49 (N_49,In_796,In_1611);
xnor U50 (N_50,In_1337,In_1303);
nor U51 (N_51,In_699,In_1380);
nor U52 (N_52,In_1156,In_855);
xor U53 (N_53,In_1078,In_1121);
xor U54 (N_54,In_287,In_787);
or U55 (N_55,In_1493,In_888);
or U56 (N_56,In_1336,In_1314);
xor U57 (N_57,In_1447,In_621);
nand U58 (N_58,In_381,In_640);
nand U59 (N_59,In_402,In_1793);
nor U60 (N_60,In_333,In_397);
or U61 (N_61,In_53,In_253);
and U62 (N_62,In_1042,In_29);
nand U63 (N_63,In_553,In_1625);
or U64 (N_64,In_490,In_16);
nand U65 (N_65,In_1205,In_305);
xor U66 (N_66,In_1025,In_1708);
nand U67 (N_67,In_754,In_1772);
and U68 (N_68,In_1321,In_775);
nor U69 (N_69,In_1926,In_11);
nand U70 (N_70,In_613,In_739);
nor U71 (N_71,In_332,In_319);
and U72 (N_72,In_840,In_1964);
and U73 (N_73,In_1476,In_1191);
nor U74 (N_74,In_226,In_1341);
xnor U75 (N_75,In_1002,In_164);
or U76 (N_76,In_1752,In_811);
or U77 (N_77,In_1847,In_159);
xor U78 (N_78,In_222,In_1193);
nand U79 (N_79,In_1399,In_1070);
xnor U80 (N_80,In_48,In_1499);
nand U81 (N_81,In_276,In_326);
xor U82 (N_82,In_299,In_990);
xor U83 (N_83,In_106,In_86);
xor U84 (N_84,In_1254,In_433);
xor U85 (N_85,In_71,In_362);
xor U86 (N_86,In_440,In_1626);
and U87 (N_87,In_1100,In_1711);
xnor U88 (N_88,In_995,In_655);
xor U89 (N_89,In_600,In_1650);
and U90 (N_90,In_1895,In_230);
or U91 (N_91,In_1491,In_589);
and U92 (N_92,In_453,In_1412);
xor U93 (N_93,In_1365,In_268);
and U94 (N_94,In_443,In_891);
or U95 (N_95,In_1857,In_1023);
xor U96 (N_96,In_296,In_714);
or U97 (N_97,In_523,In_291);
xnor U98 (N_98,In_1284,In_1803);
and U99 (N_99,In_417,In_665);
nand U100 (N_100,In_1081,In_993);
and U101 (N_101,In_951,In_1881);
nand U102 (N_102,In_547,In_124);
xnor U103 (N_103,In_548,In_1995);
xor U104 (N_104,In_981,In_1467);
nor U105 (N_105,In_1388,In_947);
and U106 (N_106,In_400,In_1109);
or U107 (N_107,In_5,In_1343);
nand U108 (N_108,In_1169,In_1945);
nor U109 (N_109,In_156,In_494);
or U110 (N_110,In_411,In_1807);
xnor U111 (N_111,In_782,In_30);
nor U112 (N_112,In_997,In_1912);
nor U113 (N_113,In_41,In_1747);
and U114 (N_114,In_1258,In_1765);
nor U115 (N_115,In_1163,In_645);
and U116 (N_116,In_1784,In_936);
nor U117 (N_117,In_684,In_1659);
nor U118 (N_118,In_1852,In_246);
or U119 (N_119,In_76,In_602);
nand U120 (N_120,In_1186,In_282);
nand U121 (N_121,In_242,In_452);
nand U122 (N_122,In_649,In_22);
or U123 (N_123,In_123,In_901);
nor U124 (N_124,In_15,In_524);
nand U125 (N_125,In_1728,In_1800);
or U126 (N_126,In_828,In_969);
xnor U127 (N_127,In_1841,In_1662);
nor U128 (N_128,In_890,In_132);
xnor U129 (N_129,In_101,In_506);
nand U130 (N_130,In_339,In_1730);
xor U131 (N_131,In_1347,In_989);
nand U132 (N_132,In_792,In_1830);
nor U133 (N_133,In_1538,In_795);
xor U134 (N_134,In_647,In_130);
nor U135 (N_135,In_975,In_1971);
xnor U136 (N_136,In_1957,In_1200);
nand U137 (N_137,In_442,In_698);
and U138 (N_138,In_1367,In_648);
nand U139 (N_139,In_1415,In_152);
xor U140 (N_140,In_1429,In_131);
nand U141 (N_141,In_1475,In_1522);
and U142 (N_142,In_183,In_467);
nor U143 (N_143,In_195,In_24);
and U144 (N_144,In_1403,In_1265);
xor U145 (N_145,In_1682,In_91);
nor U146 (N_146,In_592,In_1566);
nor U147 (N_147,In_646,In_1699);
nor U148 (N_148,In_1490,In_617);
nand U149 (N_149,In_505,In_1796);
and U150 (N_150,In_1871,In_1727);
or U151 (N_151,In_1328,In_267);
or U152 (N_152,In_1066,In_212);
or U153 (N_153,In_1189,In_743);
nand U154 (N_154,In_1307,In_1177);
nor U155 (N_155,In_1914,In_320);
nand U156 (N_156,In_1985,In_856);
xor U157 (N_157,In_1126,In_193);
and U158 (N_158,In_1050,In_712);
nand U159 (N_159,In_709,In_596);
or U160 (N_160,N_56,In_89);
nand U161 (N_161,In_1221,In_412);
xnor U162 (N_162,In_229,In_175);
xnor U163 (N_163,N_49,In_1676);
and U164 (N_164,In_1808,In_742);
nand U165 (N_165,In_850,In_463);
nand U166 (N_166,In_454,In_704);
nand U167 (N_167,In_1599,In_1921);
xnor U168 (N_168,In_1709,In_1164);
nor U169 (N_169,N_154,In_1695);
xnor U170 (N_170,In_1837,In_1339);
xnor U171 (N_171,In_542,N_19);
nand U172 (N_172,In_1963,In_934);
nor U173 (N_173,In_1667,In_1668);
nor U174 (N_174,In_1589,In_1535);
nand U175 (N_175,In_546,In_1021);
or U176 (N_176,In_1119,In_1696);
nand U177 (N_177,In_1058,In_1247);
and U178 (N_178,In_1489,In_1494);
xor U179 (N_179,In_1865,In_384);
or U180 (N_180,In_1064,In_1915);
nand U181 (N_181,In_474,In_275);
xor U182 (N_182,In_809,In_1679);
xnor U183 (N_183,In_552,In_1459);
nand U184 (N_184,In_1556,In_434);
nor U185 (N_185,In_1455,In_1387);
and U186 (N_186,N_77,In_919);
or U187 (N_187,In_337,In_914);
and U188 (N_188,In_1740,In_466);
nor U189 (N_189,In_1462,In_1889);
and U190 (N_190,N_0,In_1998);
xor U191 (N_191,In_986,In_1931);
nand U192 (N_192,In_168,In_1694);
or U193 (N_193,In_1394,In_1554);
nand U194 (N_194,In_521,In_943);
nand U195 (N_195,In_940,In_972);
or U196 (N_196,In_1612,In_1422);
nand U197 (N_197,In_439,In_315);
and U198 (N_198,In_1601,In_344);
or U199 (N_199,In_1530,In_1630);
nand U200 (N_200,In_1154,In_1065);
xor U201 (N_201,In_302,In_1346);
xor U202 (N_202,In_1144,In_556);
or U203 (N_203,In_982,In_765);
nor U204 (N_204,In_771,In_747);
and U205 (N_205,In_404,In_108);
nand U206 (N_206,In_176,In_752);
and U207 (N_207,In_1128,In_522);
and U208 (N_208,In_1897,In_451);
nor U209 (N_209,In_1812,In_1213);
xor U210 (N_210,In_162,In_582);
xnor U211 (N_211,In_1176,In_626);
or U212 (N_212,In_918,In_1433);
xnor U213 (N_213,In_403,In_1587);
nor U214 (N_214,In_1435,In_762);
nor U215 (N_215,In_1823,In_1940);
and U216 (N_216,In_405,In_1819);
nor U217 (N_217,In_146,In_933);
or U218 (N_218,In_831,In_985);
and U219 (N_219,In_1246,In_670);
and U220 (N_220,In_84,In_863);
or U221 (N_221,In_1120,In_1424);
and U222 (N_222,In_1875,In_331);
nand U223 (N_223,In_1825,In_477);
and U224 (N_224,In_674,In_1335);
and U225 (N_225,In_1295,In_1628);
and U226 (N_226,In_1464,In_727);
nand U227 (N_227,In_508,In_1685);
or U228 (N_228,In_1506,In_830);
nand U229 (N_229,In_1614,In_630);
or U230 (N_230,N_153,In_1018);
nor U231 (N_231,In_1312,In_1319);
or U232 (N_232,In_1267,In_83);
nor U233 (N_233,In_1118,In_500);
xnor U234 (N_234,In_424,In_1206);
and U235 (N_235,In_1868,In_1397);
and U236 (N_236,In_300,In_1517);
and U237 (N_237,In_1561,In_586);
nor U238 (N_238,In_1473,In_346);
or U239 (N_239,In_580,In_749);
and U240 (N_240,In_696,In_1419);
xor U241 (N_241,In_1789,In_1648);
and U242 (N_242,In_756,In_564);
and U243 (N_243,In_929,N_83);
xnor U244 (N_244,In_1974,In_1401);
nand U245 (N_245,In_551,In_18);
nand U246 (N_246,In_1416,In_155);
nand U247 (N_247,In_325,In_1240);
or U248 (N_248,In_1185,In_119);
nor U249 (N_249,In_1542,In_224);
nand U250 (N_250,In_661,In_889);
or U251 (N_251,In_776,In_393);
or U252 (N_252,In_181,In_126);
or U253 (N_253,In_14,In_1389);
nor U254 (N_254,In_1305,In_1618);
or U255 (N_255,In_116,In_838);
nor U256 (N_256,In_875,N_138);
xor U257 (N_257,N_155,N_76);
xor U258 (N_258,In_810,In_893);
or U259 (N_259,In_94,In_1697);
nand U260 (N_260,In_713,In_388);
nand U261 (N_261,In_272,In_1507);
and U262 (N_262,In_1075,In_1463);
nand U263 (N_263,N_64,In_632);
and U264 (N_264,N_135,N_150);
nand U265 (N_265,N_44,In_1508);
nand U266 (N_266,In_171,In_1290);
nand U267 (N_267,In_857,In_1671);
nand U268 (N_268,In_1735,In_172);
nand U269 (N_269,In_912,In_769);
or U270 (N_270,In_571,In_711);
xnor U271 (N_271,In_82,In_1529);
and U272 (N_272,In_1398,In_217);
or U273 (N_273,In_531,In_1393);
nand U274 (N_274,In_1638,In_816);
nand U275 (N_275,N_131,N_108);
nor U276 (N_276,In_1532,In_1955);
xnor U277 (N_277,In_958,In_1215);
or U278 (N_278,In_1190,In_733);
nand U279 (N_279,In_1024,In_363);
and U280 (N_280,In_1904,In_565);
nor U281 (N_281,In_638,In_1076);
nand U282 (N_282,In_1705,In_1280);
nor U283 (N_283,N_118,In_1045);
nor U284 (N_284,In_1570,In_1605);
xor U285 (N_285,In_1101,In_1818);
or U286 (N_286,In_1345,In_504);
or U287 (N_287,In_906,In_703);
xnor U288 (N_288,In_1687,In_915);
nor U289 (N_289,In_110,In_1888);
or U290 (N_290,In_1229,In_96);
or U291 (N_291,In_1324,In_573);
nand U292 (N_292,N_98,In_375);
nor U293 (N_293,In_1408,N_88);
nor U294 (N_294,In_1020,In_1062);
xor U295 (N_295,N_3,N_40);
and U296 (N_296,In_1738,In_1783);
nand U297 (N_297,In_355,In_1568);
nand U298 (N_298,In_664,In_1103);
xnor U299 (N_299,In_1799,In_1311);
and U300 (N_300,In_812,In_1356);
nor U301 (N_301,In_923,In_200);
xnor U302 (N_302,In_390,In_1214);
nor U303 (N_303,In_1653,In_444);
xnor U304 (N_304,In_1677,In_996);
or U305 (N_305,In_1927,In_408);
xor U306 (N_306,In_1850,In_858);
and U307 (N_307,In_42,In_67);
xor U308 (N_308,In_113,In_1551);
nor U309 (N_309,In_689,In_1781);
nand U310 (N_310,In_1460,N_99);
nor U311 (N_311,In_209,In_435);
or U312 (N_312,In_841,N_107);
nor U313 (N_313,In_784,In_140);
nor U314 (N_314,In_1593,N_71);
and U315 (N_315,N_89,In_1012);
xnor U316 (N_316,In_379,In_239);
nand U317 (N_317,In_663,In_1947);
and U318 (N_318,In_1647,In_960);
and U319 (N_319,N_103,In_681);
xor U320 (N_320,In_1344,In_1374);
or U321 (N_321,In_161,In_1669);
nand U322 (N_322,N_109,In_1834);
and U323 (N_323,In_562,In_252);
and U324 (N_324,N_115,In_667);
xor U325 (N_325,N_142,In_1057);
or U326 (N_326,In_372,In_852);
and U327 (N_327,N_207,N_173);
xor U328 (N_328,In_1741,In_312);
nor U329 (N_329,In_1479,N_289);
nor U330 (N_330,In_265,In_1941);
and U331 (N_331,In_376,N_245);
or U332 (N_332,In_770,In_848);
nand U333 (N_333,In_1792,In_666);
nand U334 (N_334,In_1543,In_1302);
and U335 (N_335,In_99,In_1813);
or U336 (N_336,In_620,In_753);
or U337 (N_337,In_1005,In_1821);
nor U338 (N_338,In_716,In_987);
nand U339 (N_339,In_1632,In_886);
nor U340 (N_340,In_1202,In_308);
nand U341 (N_341,In_240,In_93);
nor U342 (N_342,In_1775,In_1684);
or U343 (N_343,In_639,N_263);
nor U344 (N_344,In_529,In_1504);
nor U345 (N_345,N_267,N_284);
nand U346 (N_346,N_9,N_181);
or U347 (N_347,In_1851,N_111);
and U348 (N_348,In_1035,In_208);
nor U349 (N_349,In_1658,In_1273);
or U350 (N_350,In_1935,In_207);
nand U351 (N_351,In_1651,In_1438);
nand U352 (N_352,N_220,In_1782);
xnor U353 (N_353,In_928,In_1849);
and U354 (N_354,In_406,In_27);
nand U355 (N_355,In_307,In_422);
nand U356 (N_356,In_1716,In_1009);
nor U357 (N_357,In_109,In_1513);
or U358 (N_358,N_189,N_45);
nor U359 (N_359,In_881,In_1182);
nor U360 (N_360,In_897,In_1037);
and U361 (N_361,N_105,In_1725);
or U362 (N_362,N_200,In_705);
and U363 (N_363,N_168,In_1856);
nor U364 (N_364,N_274,In_1184);
nor U365 (N_365,In_826,N_170);
nor U366 (N_366,In_1285,N_300);
nand U367 (N_367,In_1440,In_60);
nor U368 (N_368,In_1983,In_780);
nor U369 (N_369,In_1261,In_927);
xnor U370 (N_370,In_1137,In_948);
xnor U371 (N_371,In_717,In_410);
nor U372 (N_372,In_1358,In_1721);
nand U373 (N_373,In_389,In_427);
nor U374 (N_374,In_1903,In_1748);
and U375 (N_375,In_374,In_206);
nor U376 (N_376,In_660,In_1592);
nand U377 (N_377,In_1873,In_693);
nand U378 (N_378,N_141,In_236);
nor U379 (N_379,In_821,In_1316);
nand U380 (N_380,In_1481,In_33);
nor U381 (N_381,In_1731,In_694);
xor U382 (N_382,In_781,In_65);
xor U383 (N_383,In_1286,In_1384);
nor U384 (N_384,N_36,In_437);
nor U385 (N_385,In_270,In_382);
or U386 (N_386,In_1804,In_1641);
and U387 (N_387,In_803,In_583);
and U388 (N_388,N_11,In_1576);
or U389 (N_389,In_849,N_117);
nor U390 (N_390,In_1854,In_1994);
or U391 (N_391,In_965,In_1734);
and U392 (N_392,In_480,In_368);
nor U393 (N_393,In_166,In_227);
nor U394 (N_394,In_1902,N_226);
or U395 (N_395,N_235,N_86);
or U396 (N_396,In_1046,In_1516);
nand U397 (N_397,In_794,In_43);
xnor U398 (N_398,In_1984,In_1067);
xnor U399 (N_399,In_1501,In_1331);
nor U400 (N_400,N_158,N_13);
xnor U401 (N_401,In_277,In_1704);
nor U402 (N_402,In_526,In_854);
or U403 (N_403,In_1729,In_1124);
and U404 (N_404,In_767,In_201);
nor U405 (N_405,In_438,N_84);
and U406 (N_406,In_658,In_1439);
and U407 (N_407,N_249,In_1839);
nor U408 (N_408,N_227,In_654);
or U409 (N_409,N_240,In_677);
and U410 (N_410,N_149,In_691);
nand U411 (N_411,In_1376,In_259);
and U412 (N_412,N_41,In_248);
nand U413 (N_413,In_1750,N_6);
or U414 (N_414,In_1564,In_1713);
xnor U415 (N_415,In_528,In_1524);
nor U416 (N_416,In_1622,In_1060);
nand U417 (N_417,In_1703,In_896);
xnor U418 (N_418,In_1301,In_1000);
and U419 (N_419,In_1271,In_924);
nand U420 (N_420,In_1351,In_662);
and U421 (N_421,In_834,In_428);
and U422 (N_422,In_1448,In_324);
nor U423 (N_423,In_185,In_1071);
or U424 (N_424,In_760,In_497);
or U425 (N_425,In_604,In_481);
and U426 (N_426,In_1038,In_949);
and U427 (N_427,In_824,In_238);
xor U428 (N_428,In_1111,N_57);
and U429 (N_429,In_902,In_1959);
nand U430 (N_430,N_33,In_1672);
xor U431 (N_431,In_1225,In_1342);
and U432 (N_432,In_1364,N_301);
xnor U433 (N_433,In_688,In_1456);
nand U434 (N_434,In_687,In_735);
xor U435 (N_435,In_544,In_846);
nor U436 (N_436,N_85,In_1272);
nand U437 (N_437,In_921,In_58);
or U438 (N_438,In_1405,In_1531);
nor U439 (N_439,N_268,In_1130);
xor U440 (N_440,In_499,In_1196);
and U441 (N_441,In_188,In_1809);
or U442 (N_442,In_154,In_1920);
xor U443 (N_443,In_1275,In_377);
nand U444 (N_444,N_260,In_651);
nor U445 (N_445,In_953,In_429);
and U446 (N_446,In_876,In_578);
or U447 (N_447,N_184,In_907);
xor U448 (N_448,In_1352,In_585);
or U449 (N_449,In_1372,In_1427);
nand U450 (N_450,In_1145,In_1512);
or U451 (N_451,In_1172,In_1743);
nor U452 (N_452,In_880,In_722);
and U453 (N_453,In_501,N_237);
and U454 (N_454,In_1890,In_1033);
and U455 (N_455,In_799,In_720);
and U456 (N_456,In_100,In_1510);
and U457 (N_457,In_910,In_251);
xnor U458 (N_458,In_1744,In_779);
or U459 (N_459,In_1924,In_926);
nor U460 (N_460,In_8,In_823);
nor U461 (N_461,In_335,In_133);
nand U462 (N_462,In_1977,In_1980);
nor U463 (N_463,In_729,In_44);
or U464 (N_464,In_1733,In_1901);
nand U465 (N_465,In_761,In_1786);
and U466 (N_466,In_570,In_1742);
nand U467 (N_467,In_866,In_1844);
xnor U468 (N_468,In_539,In_1546);
xor U469 (N_469,In_1523,N_228);
and U470 (N_470,In_1526,In_1222);
xnor U471 (N_471,In_945,In_347);
nand U472 (N_472,In_470,In_1718);
xor U473 (N_473,N_156,In_1822);
xor U474 (N_474,In_634,N_106);
xor U475 (N_475,In_1159,In_174);
xnor U476 (N_476,N_299,In_724);
nand U477 (N_477,In_1426,In_978);
xnor U478 (N_478,In_746,In_205);
and U479 (N_479,In_455,In_147);
and U480 (N_480,In_612,In_1719);
nand U481 (N_481,In_1537,N_182);
or U482 (N_482,In_75,In_961);
and U483 (N_483,N_464,In_788);
nor U484 (N_484,N_175,In_1905);
nor U485 (N_485,In_1997,N_318);
and U486 (N_486,In_1432,In_723);
or U487 (N_487,In_870,N_157);
xor U488 (N_488,N_321,In_105);
nor U489 (N_489,In_513,In_255);
or U490 (N_490,N_239,In_1223);
or U491 (N_491,In_1886,In_992);
xnor U492 (N_492,In_19,In_1579);
nand U493 (N_493,In_138,N_357);
xor U494 (N_494,N_59,In_637);
xnor U495 (N_495,In_1008,In_568);
xor U496 (N_496,N_96,In_1845);
nor U497 (N_497,In_1698,N_102);
nor U498 (N_498,In_1754,In_950);
xnor U499 (N_499,N_431,In_316);
nand U500 (N_500,N_418,In_1720);
and U501 (N_501,In_1069,N_119);
and U502 (N_502,In_1244,In_744);
nand U503 (N_503,In_804,N_12);
xor U504 (N_504,N_195,In_1);
xor U505 (N_505,N_139,N_162);
nor U506 (N_506,In_1413,N_114);
nor U507 (N_507,In_472,In_77);
xor U508 (N_508,N_215,In_790);
or U509 (N_509,In_925,N_333);
xor U510 (N_510,In_1236,In_1366);
nand U511 (N_511,N_426,In_1661);
and U512 (N_512,In_616,N_63);
and U513 (N_513,In_117,N_259);
nor U514 (N_514,In_1104,In_1266);
nand U515 (N_515,N_397,N_62);
nor U516 (N_516,In_872,In_671);
nand U517 (N_517,In_813,In_519);
nor U518 (N_518,In_1540,N_187);
or U519 (N_519,N_20,In_1179);
and U520 (N_520,In_1835,In_401);
or U521 (N_521,In_345,In_1520);
and U522 (N_522,In_511,In_1094);
xnor U523 (N_523,N_196,In_575);
xnor U524 (N_524,In_1291,In_730);
nor U525 (N_525,N_445,In_213);
nand U526 (N_526,N_309,In_629);
nand U527 (N_527,In_1122,In_286);
and U528 (N_528,In_458,In_1639);
or U529 (N_529,N_330,In_1949);
or U530 (N_530,In_330,N_478);
nand U531 (N_531,In_1906,In_777);
xor U532 (N_532,N_446,N_14);
or U533 (N_533,In_1425,In_0);
xnor U534 (N_534,In_7,In_127);
or U535 (N_535,N_415,In_1884);
nand U536 (N_536,In_1417,In_1279);
or U537 (N_537,N_176,In_1093);
nand U538 (N_538,In_614,N_16);
nand U539 (N_539,In_1157,In_348);
xnor U540 (N_540,In_998,In_40);
nor U541 (N_541,In_461,In_1485);
and U542 (N_542,In_1817,In_789);
nand U543 (N_543,In_1511,In_1978);
xor U544 (N_544,In_1292,In_31);
and U545 (N_545,N_38,In_659);
nand U546 (N_546,In_151,In_1999);
and U547 (N_547,N_315,In_584);
nand U548 (N_548,N_317,In_64);
or U549 (N_549,N_417,In_1624);
nor U550 (N_550,In_418,In_1797);
xnor U551 (N_551,N_230,In_1942);
and U552 (N_552,In_1400,In_882);
xor U553 (N_553,N_476,In_1363);
xnor U554 (N_554,In_1536,In_1114);
and U555 (N_555,In_734,In_68);
xnor U556 (N_556,In_37,N_334);
nor U557 (N_557,In_827,N_474);
or U558 (N_558,In_1357,N_337);
and U559 (N_559,In_835,In_642);
xnor U560 (N_560,In_1987,N_163);
nand U561 (N_561,In_383,In_317);
xnor U562 (N_562,In_653,In_606);
nand U563 (N_563,N_241,In_954);
and U564 (N_564,N_132,N_144);
and U565 (N_565,In_1552,In_1518);
xor U566 (N_566,In_1814,N_375);
xnor U567 (N_567,In_967,In_1635);
or U568 (N_568,In_509,In_1049);
xnor U569 (N_569,N_281,In_1218);
xor U570 (N_570,In_1270,In_57);
nand U571 (N_571,N_223,In_1951);
xor U572 (N_572,N_242,In_701);
and U573 (N_573,In_1268,In_899);
nor U574 (N_574,In_1194,In_1846);
or U575 (N_575,N_219,In_738);
xnor U576 (N_576,In_1168,In_567);
and U577 (N_577,In_1368,N_15);
nand U578 (N_578,In_1210,In_865);
nand U579 (N_579,In_1106,In_399);
or U580 (N_580,In_766,N_75);
nor U581 (N_581,In_1478,N_204);
nor U582 (N_582,N_438,N_25);
xor U583 (N_583,N_116,In_898);
nor U584 (N_584,In_1700,In_98);
or U585 (N_585,In_137,In_737);
or U586 (N_586,N_43,N_414);
and U587 (N_587,N_133,In_558);
nand U588 (N_588,In_1161,In_482);
xnor U589 (N_589,In_1619,N_402);
xor U590 (N_590,In_877,In_917);
and U591 (N_591,N_244,In_1970);
nand U592 (N_592,In_868,In_668);
nand U593 (N_593,In_631,In_1480);
and U594 (N_594,In_581,In_1004);
xnor U595 (N_595,In_1960,In_847);
nand U596 (N_596,N_353,In_1160);
or U597 (N_597,In_1458,In_52);
and U598 (N_598,N_7,In_1633);
nand U599 (N_599,In_1498,In_392);
or U600 (N_600,N_58,In_1252);
or U601 (N_601,In_750,In_469);
or U602 (N_602,In_36,In_719);
xor U603 (N_603,In_1829,N_411);
and U604 (N_604,In_1197,In_1304);
or U605 (N_605,In_129,In_190);
nor U606 (N_606,In_261,N_53);
xnor U607 (N_607,In_1395,N_48);
and U608 (N_608,N_238,In_1787);
xnor U609 (N_609,In_142,In_1032);
nand U610 (N_610,In_941,In_843);
and U611 (N_611,N_35,In_844);
nor U612 (N_612,In_1629,In_233);
xnor U613 (N_613,In_204,In_266);
nor U614 (N_614,In_1801,In_695);
and U615 (N_615,N_91,In_622);
xnor U616 (N_616,In_1877,In_1515);
nand U617 (N_617,N_405,In_1195);
xnor U618 (N_618,In_1031,N_341);
xnor U619 (N_619,N_127,In_1863);
nand U620 (N_620,In_1113,In_1598);
xor U621 (N_621,In_1690,In_512);
xor U622 (N_622,In_1991,In_1088);
nand U623 (N_623,In_1681,In_1880);
nand U624 (N_624,In_1061,In_728);
and U625 (N_625,N_233,In_1264);
nor U626 (N_626,In_430,In_557);
and U627 (N_627,In_878,In_1836);
nor U628 (N_628,In_561,In_1497);
nor U629 (N_629,In_1472,N_5);
xor U630 (N_630,N_390,In_1019);
and U631 (N_631,N_39,In_179);
or U632 (N_632,In_1442,In_1673);
nor U633 (N_633,In_431,In_1872);
nand U634 (N_634,N_213,In_1131);
xnor U635 (N_635,In_25,In_514);
and U636 (N_636,In_1022,In_1678);
xor U637 (N_637,In_1457,N_412);
nand U638 (N_638,In_1874,In_1918);
nand U639 (N_639,In_80,In_1390);
nor U640 (N_640,N_273,In_1928);
nand U641 (N_641,N_78,N_23);
and U642 (N_642,In_869,In_853);
xor U643 (N_643,In_517,In_971);
nand U644 (N_644,In_1477,N_350);
xnor U645 (N_645,In_1139,N_499);
and U646 (N_646,In_153,In_1603);
nor U647 (N_647,In_1027,N_462);
xnor U648 (N_648,N_618,N_466);
nor U649 (N_649,In_135,In_682);
xor U650 (N_650,In_970,N_342);
xor U651 (N_651,In_173,In_1263);
nand U652 (N_652,In_51,N_447);
xor U653 (N_653,In_1574,N_264);
xnor U654 (N_654,In_1333,N_253);
or U655 (N_655,In_1199,In_550);
or U656 (N_656,In_535,In_1108);
or U657 (N_657,N_594,In_409);
nor U658 (N_658,In_1930,In_1495);
nor U659 (N_659,N_450,N_512);
nand U660 (N_660,N_24,N_93);
and U661 (N_661,In_1349,In_21);
or U662 (N_662,In_1565,N_592);
xnor U663 (N_663,N_420,In_1257);
nor U664 (N_664,In_942,N_61);
nor U665 (N_665,N_535,N_169);
and U666 (N_666,In_1028,In_758);
or U667 (N_667,In_1203,In_1860);
nand U668 (N_668,In_257,In_446);
nand U669 (N_669,N_113,In_686);
xor U670 (N_670,N_82,In_1656);
and U671 (N_671,N_18,In_566);
nand U672 (N_672,In_624,In_72);
nand U673 (N_673,In_1474,In_1870);
nor U674 (N_674,In_364,N_632);
and U675 (N_675,N_449,In_465);
nor U676 (N_676,In_1496,N_212);
or U677 (N_677,In_643,In_1544);
nor U678 (N_678,N_540,In_595);
xor U679 (N_679,In_1348,In_1878);
nand U680 (N_680,In_1869,In_1967);
nor U681 (N_681,In_549,N_174);
or U682 (N_682,In_1117,In_180);
xor U683 (N_683,In_1123,In_70);
nand U684 (N_684,In_1717,N_305);
or U685 (N_685,In_1909,In_974);
or U686 (N_686,In_905,In_732);
nor U687 (N_687,In_61,In_973);
nor U688 (N_688,N_101,In_1664);
nand U689 (N_689,In_1127,In_448);
xnor U690 (N_690,In_244,N_564);
nand U691 (N_691,In_1778,In_184);
nand U692 (N_692,In_725,N_605);
nor U693 (N_693,In_1248,N_319);
or U694 (N_694,In_46,In_1581);
and U695 (N_695,In_591,In_533);
nand U696 (N_696,N_256,In_959);
nand U697 (N_697,In_85,In_79);
nand U698 (N_698,N_328,N_516);
or U699 (N_699,N_287,In_1609);
or U700 (N_700,In_1450,In_1443);
nand U701 (N_701,N_247,In_1505);
nand U702 (N_702,In_1298,In_1824);
xor U703 (N_703,In_81,In_294);
xnor U704 (N_704,In_1675,In_1569);
xnor U705 (N_705,In_1143,In_598);
or U706 (N_706,In_1893,N_303);
nand U707 (N_707,In_475,N_60);
nor U708 (N_708,In_768,N_282);
and U709 (N_709,In_609,In_1171);
nand U710 (N_710,N_608,In_1899);
and U711 (N_711,N_294,In_1162);
nor U712 (N_712,N_391,In_1674);
xnor U713 (N_713,N_302,N_612);
xor U714 (N_714,In_1192,In_887);
and U715 (N_715,N_97,In_280);
nand U716 (N_716,N_203,In_628);
xnor U717 (N_717,In_63,N_123);
xor U718 (N_718,In_118,In_590);
xor U719 (N_719,N_498,N_148);
xor U720 (N_720,In_650,In_1404);
nand U721 (N_721,N_639,N_246);
and U722 (N_722,In_976,N_121);
or U723 (N_723,In_211,In_1958);
and U724 (N_724,In_1158,In_1548);
xor U725 (N_725,N_520,N_311);
nand U726 (N_726,N_279,N_584);
and U727 (N_727,In_1660,In_1047);
or U728 (N_728,In_1769,N_210);
and U729 (N_729,N_419,In_820);
nand U730 (N_730,In_218,In_1557);
and U731 (N_731,In_20,In_95);
nand U732 (N_732,N_340,In_641);
and U733 (N_733,In_413,N_546);
xnor U734 (N_734,In_502,N_252);
or U735 (N_735,In_1966,N_143);
nand U736 (N_736,In_503,In_220);
and U737 (N_737,N_270,In_525);
nor U738 (N_738,In_1041,N_532);
or U739 (N_739,N_527,N_295);
nor U740 (N_740,In_1465,N_261);
xnor U741 (N_741,In_807,N_248);
nand U742 (N_742,N_271,In_66);
xnor U743 (N_743,In_73,In_264);
and U744 (N_744,In_186,In_395);
nor U745 (N_745,In_1187,In_107);
and U746 (N_746,In_1112,In_1549);
and U747 (N_747,N_363,In_1151);
xor U748 (N_748,In_1383,In_38);
nand U749 (N_749,In_1585,N_541);
or U750 (N_750,N_413,N_377);
nand U751 (N_751,In_1141,N_556);
or U752 (N_752,In_1533,N_492);
nor U753 (N_753,In_1116,In_1418);
or U754 (N_754,In_492,N_437);
and U755 (N_755,In_702,In_1917);
and U756 (N_756,N_46,In_1712);
and U757 (N_757,N_112,In_1327);
nor U758 (N_758,In_1770,In_879);
and U759 (N_759,In_785,In_864);
and U760 (N_760,In_1780,N_202);
or U761 (N_761,N_278,N_425);
or U762 (N_762,In_1663,In_764);
or U763 (N_763,In_1810,In_1794);
nand U764 (N_764,N_487,In_1528);
and U765 (N_765,N_179,In_2);
xor U766 (N_766,N_549,N_367);
nor U767 (N_767,In_13,In_197);
or U768 (N_768,In_6,In_1665);
or U769 (N_769,In_1649,N_382);
and U770 (N_770,In_489,In_707);
and U771 (N_771,N_381,N_455);
and U772 (N_772,In_1382,N_262);
nor U773 (N_773,In_1680,In_538);
xor U774 (N_774,In_1634,In_1354);
and U775 (N_775,N_358,N_288);
nand U776 (N_776,In_216,In_1250);
and U777 (N_777,In_74,In_387);
or U778 (N_778,N_436,In_269);
xor U779 (N_779,In_1446,In_1231);
xor U780 (N_780,N_552,In_1582);
or U781 (N_781,N_623,In_1256);
nand U782 (N_782,N_368,In_1381);
xnor U783 (N_783,In_736,N_622);
and U784 (N_784,In_1211,In_1183);
or U785 (N_785,In_1297,In_652);
or U786 (N_786,In_351,In_394);
and U787 (N_787,In_908,N_534);
nor U788 (N_788,In_939,In_1670);
nand U789 (N_789,N_70,In_1414);
or U790 (N_790,In_496,In_1749);
nor U791 (N_791,In_1968,In_488);
and U792 (N_792,In_182,In_369);
and U793 (N_793,In_802,In_1876);
or U794 (N_794,N_54,N_308);
and U795 (N_795,N_167,In_555);
xnor U796 (N_796,In_1392,N_255);
nor U797 (N_797,N_559,In_169);
and U798 (N_798,In_1362,In_1326);
nor U799 (N_799,In_1437,In_1805);
or U800 (N_800,In_1320,In_342);
nor U801 (N_801,N_519,In_1627);
nor U802 (N_802,In_1132,In_1938);
or U803 (N_803,In_726,In_755);
nand U804 (N_804,N_234,N_286);
or U805 (N_805,N_501,In_1451);
nand U806 (N_806,N_205,In_1806);
xor U807 (N_807,In_1167,In_1798);
nor U808 (N_808,In_304,In_1726);
or U809 (N_809,In_745,In_1149);
and U810 (N_810,In_1916,N_485);
nand U811 (N_811,In_783,In_1153);
nor U812 (N_812,N_50,In_1937);
and U813 (N_813,In_1562,In_1488);
or U814 (N_814,N_147,In_1514);
nor U815 (N_815,In_214,N_715);
nor U816 (N_816,N_719,N_316);
nand U817 (N_817,N_706,N_723);
nor U818 (N_818,In_1560,In_1948);
xor U819 (N_819,In_415,N_250);
nand U820 (N_820,In_1843,In_223);
or U821 (N_821,In_1950,In_285);
xor U822 (N_822,In_1016,In_1584);
or U823 (N_823,N_566,In_292);
nor U824 (N_824,N_726,In_1773);
nand U825 (N_825,N_544,N_640);
xnor U826 (N_826,N_514,In_516);
xnor U827 (N_827,In_1449,N_633);
or U828 (N_828,N_789,In_930);
and U829 (N_829,N_129,In_1006);
nand U830 (N_830,In_1943,N_243);
nand U831 (N_831,N_593,In_1701);
and U832 (N_832,N_677,In_97);
and U833 (N_833,In_1466,N_643);
nor U834 (N_834,In_1643,N_481);
nand U835 (N_835,N_699,In_577);
nand U836 (N_836,N_225,In_1586);
and U837 (N_837,N_296,N_349);
and U838 (N_838,N_757,N_392);
and U839 (N_839,N_52,In_198);
and U840 (N_840,In_1155,N_550);
or U841 (N_841,N_191,N_380);
and U842 (N_842,N_596,In_1616);
nor U843 (N_843,N_467,In_1862);
and U844 (N_844,In_1235,In_1954);
or U845 (N_845,In_1391,In_1646);
xnor U846 (N_846,In_284,In_1578);
nor U847 (N_847,N_310,In_194);
xnor U848 (N_848,N_406,N_641);
nand U849 (N_849,In_260,In_420);
nor U850 (N_850,In_636,In_690);
or U851 (N_851,In_1003,In_839);
xnor U852 (N_852,In_1107,In_120);
nand U853 (N_853,In_1525,N_10);
and U854 (N_854,N_638,N_495);
or U855 (N_855,N_702,In_825);
xor U856 (N_856,In_1688,N_490);
or U857 (N_857,N_166,In_569);
nand U858 (N_858,N_538,N_429);
and U859 (N_859,In_1642,N_343);
nor U860 (N_860,N_275,N_339);
nor U861 (N_861,In_1325,N_606);
nor U862 (N_862,N_222,In_669);
or U863 (N_863,In_1502,N_194);
or U864 (N_864,N_389,In_1096);
or U865 (N_865,N_488,In_607);
xor U866 (N_866,In_158,N_456);
nand U867 (N_867,In_1953,In_1555);
nor U868 (N_868,N_662,In_498);
nand U869 (N_869,In_1500,N_562);
nor U870 (N_870,In_1073,In_1483);
or U871 (N_871,In_45,N_430);
xnor U872 (N_872,In_904,In_1409);
nand U873 (N_873,N_421,N_509);
xor U874 (N_874,N_457,In_1056);
nand U875 (N_875,In_170,In_1894);
xnor U876 (N_876,N_461,N_697);
and U877 (N_877,In_579,In_1436);
nor U878 (N_878,In_527,N_454);
or U879 (N_879,In_938,In_1595);
and U880 (N_880,In_859,In_806);
nor U881 (N_881,In_983,N_775);
nor U882 (N_882,In_115,In_1224);
or U883 (N_883,N_451,N_529);
and U884 (N_884,In_962,In_618);
or U885 (N_885,N_433,In_143);
nand U886 (N_886,N_722,In_1406);
nand U887 (N_887,N_724,In_883);
and U888 (N_888,N_399,N_764);
nor U889 (N_889,In_1097,In_1234);
xnor U890 (N_890,N_404,N_30);
and U891 (N_891,N_580,In_832);
or U892 (N_892,N_735,In_1939);
nor U893 (N_893,N_561,In_1802);
or U894 (N_894,In_1962,N_620);
xor U895 (N_895,In_1017,In_1993);
nand U896 (N_896,In_1001,N_134);
or U897 (N_897,In_1361,N_428);
nor U898 (N_898,In_1691,In_1484);
nor U899 (N_899,In_1866,N_221);
nand U900 (N_900,In_1559,N_69);
or U901 (N_901,In_1283,In_1152);
or U902 (N_902,In_1136,In_1091);
nand U903 (N_903,In_1492,In_148);
xnor U904 (N_904,N_734,N_713);
xnor U905 (N_905,N_463,In_441);
nor U906 (N_906,N_647,N_403);
and U907 (N_907,In_1329,In_772);
xor U908 (N_908,N_482,N_676);
nor U909 (N_909,In_603,N_422);
or U910 (N_910,N_423,N_555);
and U911 (N_911,In_165,In_610);
xor U912 (N_912,N_768,In_931);
xnor U913 (N_913,In_1220,N_31);
xnor U914 (N_914,N_771,N_769);
or U915 (N_915,N_424,N_796);
and U916 (N_916,In_274,N_2);
and U917 (N_917,In_1026,In_599);
nand U918 (N_918,N_4,N_201);
and U919 (N_919,In_1907,N_335);
or U920 (N_920,N_721,N_68);
nand U921 (N_921,N_55,N_329);
and U922 (N_922,In_1887,In_1573);
or U923 (N_923,N_183,N_743);
or U924 (N_924,N_125,In_462);
xor U925 (N_925,In_1310,N_434);
or U926 (N_926,In_69,In_1842);
xnor U927 (N_927,N_224,N_345);
and U928 (N_928,N_477,N_563);
nor U929 (N_929,In_290,In_386);
nor U930 (N_930,In_1761,N_293);
and U931 (N_931,N_503,In_968);
nor U932 (N_932,N_621,In_1083);
nand U933 (N_933,N_217,In_1757);
or U934 (N_934,N_689,In_1521);
and U935 (N_935,In_1932,N_231);
xnor U936 (N_936,In_778,In_483);
or U937 (N_937,N_551,In_139);
or U938 (N_938,In_221,In_1861);
and U939 (N_939,In_1180,In_228);
nand U940 (N_940,In_1922,In_1133);
and U941 (N_941,In_903,In_1706);
xor U942 (N_942,In_1969,In_871);
or U943 (N_943,N_581,In_378);
or U944 (N_944,In_861,N_648);
xnor U945 (N_945,N_790,In_793);
nor U946 (N_946,N_727,In_837);
or U947 (N_947,N_718,N_486);
nor U948 (N_948,N_442,In_862);
or U949 (N_949,N_646,N_777);
nand U950 (N_950,In_1919,N_439);
nand U951 (N_951,In_1077,N_649);
or U952 (N_952,In_62,In_920);
and U953 (N_953,In_1375,In_1883);
or U954 (N_954,N_94,N_122);
nand U955 (N_955,N_704,In_1756);
or U956 (N_956,N_409,In_191);
nand U957 (N_957,In_700,N_258);
nor U958 (N_958,In_576,In_1989);
and U959 (N_959,In_464,In_1430);
nor U960 (N_960,N_749,In_1838);
nand U961 (N_961,In_1359,N_773);
nand U962 (N_962,In_1355,In_104);
nor U963 (N_963,N_506,In_980);
and U964 (N_964,In_247,In_1099);
xor U965 (N_965,In_944,In_1134);
nor U966 (N_966,In_1431,In_327);
nand U967 (N_967,N_690,In_1212);
or U968 (N_968,N_452,In_1241);
nor U969 (N_969,In_1992,N_867);
and U970 (N_970,N_277,In_396);
xor U971 (N_971,In_192,N_843);
or U972 (N_972,N_955,N_824);
xor U973 (N_973,N_354,In_1452);
or U974 (N_974,In_608,In_1644);
or U975 (N_975,In_1294,In_28);
nor U976 (N_976,In_574,N_692);
and U977 (N_977,In_1386,In_1453);
or U978 (N_978,N_891,N_513);
xor U979 (N_979,N_199,N_628);
and U980 (N_980,In_17,In_520);
or U981 (N_981,In_1853,N_922);
nor U982 (N_982,In_1087,N_806);
nor U983 (N_983,N_809,N_489);
or U984 (N_984,In_1201,N_95);
and U985 (N_985,In_1115,In_1170);
or U986 (N_986,In_1245,In_1996);
and U987 (N_987,In_1085,In_262);
xor U988 (N_988,N_679,In_360);
nand U989 (N_989,N_37,In_484);
and U990 (N_990,In_1820,In_1840);
nor U991 (N_991,In_1828,N_185);
nor U992 (N_992,N_930,N_795);
and U993 (N_993,N_331,In_1322);
and U994 (N_994,In_1082,In_1575);
and U995 (N_995,N_547,In_773);
nor U996 (N_996,In_1929,In_685);
and U997 (N_997,N_578,In_1600);
or U998 (N_998,In_366,N_627);
or U999 (N_999,N_887,N_568);
nor U1000 (N_1000,N_355,In_234);
nor U1001 (N_1001,N_379,In_1795);
nand U1002 (N_1002,In_1896,In_675);
nor U1003 (N_1003,N_291,N_161);
nor U1004 (N_1004,In_935,N_361);
nor U1005 (N_1005,In_122,In_800);
xnor U1006 (N_1006,N_745,In_1173);
and U1007 (N_1007,In_1287,In_1074);
nand U1008 (N_1008,In_1299,N_292);
or U1009 (N_1009,In_1762,N_894);
xnor U1010 (N_1010,N_177,N_822);
xor U1011 (N_1011,N_208,In_1068);
or U1012 (N_1012,N_818,In_1655);
nor U1013 (N_1013,N_821,In_808);
nor U1014 (N_1014,N_304,N_472);
nor U1015 (N_1015,N_666,N_663);
or U1016 (N_1016,N_152,N_800);
or U1017 (N_1017,N_609,In_243);
xor U1018 (N_1018,In_1208,In_1411);
nand U1019 (N_1019,N_783,In_1278);
nor U1020 (N_1020,N_918,N_453);
and U1021 (N_1021,N_826,In_1378);
and U1022 (N_1022,In_1237,In_1956);
xor U1023 (N_1023,N_813,N_832);
or U1024 (N_1024,N_910,N_760);
or U1025 (N_1025,In_900,N_524);
nor U1026 (N_1026,In_751,N_901);
or U1027 (N_1027,In_1751,N_767);
nor U1028 (N_1028,N_794,In_1092);
or U1029 (N_1029,In_1296,N_165);
nor U1030 (N_1030,N_508,In_144);
nand U1031 (N_1031,In_957,In_1965);
and U1032 (N_1032,In_537,N_542);
xnor U1033 (N_1033,N_731,In_1471);
xnor U1034 (N_1034,N_528,N_837);
xor U1035 (N_1035,N_576,N_870);
nand U1036 (N_1036,In_842,N_322);
xor U1037 (N_1037,In_1988,N_372);
or U1038 (N_1038,N_686,N_886);
nor U1039 (N_1039,N_752,N_29);
or U1040 (N_1040,N_709,N_511);
xnor U1041 (N_1041,In_1925,In_1541);
or U1042 (N_1042,In_1138,In_1933);
nor U1043 (N_1043,In_1317,In_1707);
nand U1044 (N_1044,N_332,N_536);
xor U1045 (N_1045,N_920,N_951);
nor U1046 (N_1046,N_674,N_680);
and U1047 (N_1047,In_1882,N_616);
or U1048 (N_1048,N_617,N_385);
and U1049 (N_1049,N_87,In_298);
and U1050 (N_1050,In_215,In_254);
xor U1051 (N_1051,N_313,N_804);
xor U1052 (N_1052,N_925,In_1059);
nor U1053 (N_1053,In_310,N_159);
nor U1054 (N_1054,In_1011,In_1216);
and U1055 (N_1055,N_386,In_1445);
and U1056 (N_1056,In_1308,In_1666);
nand U1057 (N_1057,N_651,N_805);
and U1058 (N_1058,N_599,In_353);
nand U1059 (N_1059,N_73,N_480);
nor U1060 (N_1060,N_665,In_763);
nand U1061 (N_1061,In_1340,N_336);
nor U1062 (N_1062,In_1407,N_776);
nand U1063 (N_1063,N_770,In_1613);
and U1064 (N_1064,In_605,N_861);
nand U1065 (N_1065,N_197,N_604);
xor U1066 (N_1066,In_314,N_742);
nand U1067 (N_1067,In_476,In_103);
and U1068 (N_1068,N_808,N_793);
nand U1069 (N_1069,In_10,N_128);
xnor U1070 (N_1070,In_601,In_673);
and U1071 (N_1071,N_774,N_823);
nor U1072 (N_1072,N_725,N_654);
xnor U1073 (N_1073,N_470,N_946);
or U1074 (N_1074,In_1204,N_954);
and U1075 (N_1075,In_354,N_801);
nand U1076 (N_1076,In_1934,N_410);
nand U1077 (N_1077,In_321,In_350);
and U1078 (N_1078,In_623,N_265);
xor U1079 (N_1079,N_935,In_1689);
or U1080 (N_1080,N_845,In_786);
and U1081 (N_1081,N_67,In_1015);
nor U1082 (N_1082,N_846,N_691);
and U1083 (N_1083,In_1867,N_522);
xor U1084 (N_1084,In_1140,N_517);
and U1085 (N_1085,N_802,N_673);
or U1086 (N_1086,N_587,In_338);
and U1087 (N_1087,In_473,In_819);
nor U1088 (N_1088,N_137,N_577);
and U1089 (N_1089,In_1972,N_530);
nor U1090 (N_1090,N_484,In_748);
and U1091 (N_1091,In_1723,In_1746);
nor U1092 (N_1092,In_1944,N_502);
nand U1093 (N_1093,In_237,N_280);
xor U1094 (N_1094,N_537,In_680);
nand U1095 (N_1095,N_327,N_216);
or U1096 (N_1096,N_500,N_448);
xor U1097 (N_1097,In_1519,N_860);
nor U1098 (N_1098,In_1686,In_49);
nor U1099 (N_1099,In_1315,N_732);
nand U1100 (N_1100,In_1621,In_1657);
nand U1101 (N_1101,In_1080,N_607);
nor U1102 (N_1102,N_518,In_994);
or U1103 (N_1103,N_590,N_394);
xnor U1104 (N_1104,In_1300,N_919);
and U1105 (N_1105,N_254,In_273);
xnor U1106 (N_1106,N_830,In_911);
or U1107 (N_1107,N_748,N_567);
and U1108 (N_1108,N_707,N_746);
or U1109 (N_1109,N_803,N_110);
and U1110 (N_1110,N_570,N_714);
or U1111 (N_1111,N_521,N_700);
nor U1112 (N_1112,In_594,N_615);
and U1113 (N_1113,N_276,In_884);
nor U1114 (N_1114,In_232,N_22);
xnor U1115 (N_1115,N_160,N_814);
or U1116 (N_1116,N_737,N_759);
nor U1117 (N_1117,N_874,In_125);
or U1118 (N_1118,N_408,N_407);
nor U1119 (N_1119,In_507,N_579);
nor U1120 (N_1120,In_1606,N_923);
and U1121 (N_1121,N_781,In_1567);
nor U1122 (N_1122,In_1788,In_149);
or U1123 (N_1123,In_1053,N_172);
nand U1124 (N_1124,N_92,In_515);
nand U1125 (N_1125,N_346,N_882);
nand U1126 (N_1126,In_1238,N_895);
xor U1127 (N_1127,N_1028,N_670);
or U1128 (N_1128,N_1017,In_425);
or U1129 (N_1129,N_523,N_873);
nor U1130 (N_1130,In_798,In_1900);
or U1131 (N_1131,In_1832,N_188);
xor U1132 (N_1132,In_491,In_678);
nor U1133 (N_1133,In_1702,N_842);
or U1134 (N_1134,In_1693,N_469);
nand U1135 (N_1135,In_111,In_187);
nand U1136 (N_1136,In_1610,In_851);
or U1137 (N_1137,In_913,N_650);
and U1138 (N_1138,In_297,In_1563);
nand U1139 (N_1139,N_956,N_320);
nand U1140 (N_1140,N_366,N_325);
nand U1141 (N_1141,N_778,In_845);
nand U1142 (N_1142,N_1088,In_1973);
nor U1143 (N_1143,In_1148,N_947);
and U1144 (N_1144,In_1232,N_1062);
or U1145 (N_1145,N_1038,N_999);
and U1146 (N_1146,In_313,N_669);
nor U1147 (N_1147,N_817,N_851);
xor U1148 (N_1148,In_1898,N_820);
nor U1149 (N_1149,In_543,In_373);
or U1150 (N_1150,N_1048,N_611);
and U1151 (N_1151,N_298,N_1083);
xor U1152 (N_1152,In_1831,In_478);
xor U1153 (N_1153,In_1785,In_416);
nor U1154 (N_1154,In_1986,N_772);
nor U1155 (N_1155,In_1859,N_819);
nand U1156 (N_1156,N_1027,N_465);
nor U1157 (N_1157,In_1276,In_1911);
nor U1158 (N_1158,In_963,In_625);
and U1159 (N_1159,N_1036,N_1029);
xor U1160 (N_1160,In_203,N_683);
nor U1161 (N_1161,N_427,In_874);
nand U1162 (N_1162,N_1016,N_696);
and U1163 (N_1163,N_90,In_1110);
or U1164 (N_1164,In_1790,In_1421);
nor U1165 (N_1165,In_1768,N_573);
or U1166 (N_1166,N_645,N_1002);
or U1167 (N_1167,In_1558,N_678);
and U1168 (N_1168,In_26,In_1338);
or U1169 (N_1169,In_1503,N_980);
or U1170 (N_1170,N_81,In_1936);
or U1171 (N_1171,N_398,N_1082);
nor U1172 (N_1172,N_926,N_991);
xor U1173 (N_1173,N_812,In_1089);
and U1174 (N_1174,N_1011,N_939);
nand U1175 (N_1175,N_1116,In_909);
and U1176 (N_1176,In_309,In_1174);
and U1177 (N_1177,N_493,In_1239);
nand U1178 (N_1178,N_356,N_740);
or U1179 (N_1179,N_993,In_357);
nor U1180 (N_1180,N_1078,N_1111);
nand U1181 (N_1181,In_1410,N_862);
or U1182 (N_1182,In_1441,In_1623);
nand U1183 (N_1183,N_1044,N_1091);
nor U1184 (N_1184,N_936,N_312);
nand U1185 (N_1185,N_140,N_74);
and U1186 (N_1186,N_848,N_900);
and U1187 (N_1187,N_880,N_186);
xnor U1188 (N_1188,N_825,N_602);
xnor U1189 (N_1189,N_192,In_199);
nor U1190 (N_1190,In_1908,In_356);
and U1191 (N_1191,N_973,N_972);
and U1192 (N_1192,In_189,In_1602);
nand U1193 (N_1193,N_51,In_1745);
nand U1194 (N_1194,In_468,N_682);
nor U1195 (N_1195,N_913,In_1777);
nand U1196 (N_1196,N_218,In_833);
or U1197 (N_1197,N_553,In_718);
nor U1198 (N_1198,N_1037,In_365);
nor U1199 (N_1199,N_1104,In_741);
and U1200 (N_1200,N_883,In_1645);
xor U1201 (N_1201,N_698,N_65);
or U1202 (N_1202,N_473,N_675);
nor U1203 (N_1203,In_536,N_872);
or U1204 (N_1204,In_414,N_924);
nand U1205 (N_1205,N_751,N_1058);
or U1206 (N_1206,N_708,In_1855);
or U1207 (N_1207,In_1637,In_1402);
and U1208 (N_1208,In_250,In_1779);
or U1209 (N_1209,N_1117,N_717);
or U1210 (N_1210,N_613,N_889);
and U1211 (N_1211,N_785,In_1079);
or U1212 (N_1212,N_1024,In_56);
xor U1213 (N_1213,N_938,N_750);
nor U1214 (N_1214,In_1318,N_965);
and U1215 (N_1215,In_676,N_744);
or U1216 (N_1216,In_615,N_811);
or U1217 (N_1217,In_1147,In_1253);
and U1218 (N_1218,N_875,In_1233);
or U1219 (N_1219,In_1759,N_815);
nor U1220 (N_1220,In_336,In_486);
xor U1221 (N_1221,In_1370,In_1048);
xor U1222 (N_1222,N_857,In_916);
and U1223 (N_1223,N_976,In_715);
or U1224 (N_1224,N_876,N_841);
xnor U1225 (N_1225,N_952,In_1732);
xor U1226 (N_1226,In_1013,In_1848);
xor U1227 (N_1227,In_178,In_295);
nand U1228 (N_1228,N_1092,In_895);
or U1229 (N_1229,In_1827,In_1306);
xor U1230 (N_1230,In_988,In_456);
nor U1231 (N_1231,N_440,In_759);
nand U1232 (N_1232,N_211,In_1039);
nor U1233 (N_1233,N_927,N_507);
nor U1234 (N_1234,N_903,In_692);
and U1235 (N_1235,N_884,N_1043);
xnor U1236 (N_1236,N_899,N_687);
xnor U1237 (N_1237,In_479,In_1434);
nand U1238 (N_1238,In_163,In_1313);
nor U1239 (N_1239,In_740,In_829);
nand U1240 (N_1240,N_352,In_235);
nor U1241 (N_1241,N_251,In_1468);
and U1242 (N_1242,N_164,In_1654);
or U1243 (N_1243,In_380,N_1021);
or U1244 (N_1244,N_214,N_784);
xnor U1245 (N_1245,In_964,In_436);
or U1246 (N_1246,N_657,N_990);
xor U1247 (N_1247,N_269,N_761);
or U1248 (N_1248,In_421,N_543);
or U1249 (N_1249,N_655,N_780);
xnor U1250 (N_1250,In_1396,N_944);
nor U1251 (N_1251,In_1652,N_1086);
xor U1252 (N_1252,In_407,N_72);
nand U1253 (N_1253,N_1041,N_855);
nand U1254 (N_1254,N_885,In_271);
and U1255 (N_1255,N_987,N_992);
or U1256 (N_1256,N_370,N_949);
and U1257 (N_1257,In_1334,N_736);
and U1258 (N_1258,N_104,N_878);
or U1259 (N_1259,N_574,N_1001);
xor U1260 (N_1260,In_731,In_966);
nand U1261 (N_1261,N_986,In_1188);
xnor U1262 (N_1262,N_1022,N_786);
or U1263 (N_1263,In_952,N_971);
nor U1264 (N_1264,In_1332,N_1030);
nand U1265 (N_1265,N_190,N_728);
or U1266 (N_1266,In_59,In_1879);
nor U1267 (N_1267,N_583,N_844);
xnor U1268 (N_1268,In_708,N_942);
xor U1269 (N_1269,N_871,N_347);
xor U1270 (N_1270,N_652,N_828);
or U1271 (N_1271,In_1724,N_753);
xnor U1272 (N_1272,N_911,In_1102);
and U1273 (N_1273,N_634,N_307);
and U1274 (N_1274,N_1063,In_54);
nor U1275 (N_1275,N_272,In_134);
xor U1276 (N_1276,N_136,N_401);
or U1277 (N_1277,N_934,N_126);
nor U1278 (N_1278,In_219,N_1073);
nor U1279 (N_1279,N_545,N_362);
xnor U1280 (N_1280,In_303,N_829);
xor U1281 (N_1281,In_1034,N_1031);
xor U1282 (N_1282,N_1267,N_585);
nor U1283 (N_1283,N_754,In_318);
or U1284 (N_1284,N_989,In_1547);
and U1285 (N_1285,N_571,N_1141);
xnor U1286 (N_1286,N_653,N_859);
or U1287 (N_1287,In_1596,N_1278);
and U1288 (N_1288,N_589,N_1171);
or U1289 (N_1289,In_245,N_1165);
and U1290 (N_1290,N_917,In_1923);
nand U1291 (N_1291,In_683,N_1145);
nand U1292 (N_1292,N_684,N_1178);
or U1293 (N_1293,N_787,N_1059);
and U1294 (N_1294,N_100,N_957);
or U1295 (N_1295,N_1241,In_1353);
xor U1296 (N_1296,N_387,In_588);
nor U1297 (N_1297,N_1245,N_1157);
nor U1298 (N_1298,N_969,N_854);
xnor U1299 (N_1299,N_916,N_853);
and U1300 (N_1300,N_1142,In_1736);
nand U1301 (N_1301,N_1110,N_960);
nand U1302 (N_1302,N_1052,N_720);
or U1303 (N_1303,N_635,N_1003);
nor U1304 (N_1304,N_1182,In_50);
nor U1305 (N_1305,In_1330,N_626);
nor U1306 (N_1306,N_1026,N_525);
xor U1307 (N_1307,N_1231,In_278);
xor U1308 (N_1308,N_180,In_710);
and U1309 (N_1309,N_1061,N_1097);
nor U1310 (N_1310,In_1175,N_1009);
nand U1311 (N_1311,N_701,N_257);
or U1312 (N_1312,N_1232,N_359);
or U1313 (N_1313,N_283,In_145);
and U1314 (N_1314,N_1257,N_914);
nand U1315 (N_1315,In_150,N_1225);
xnor U1316 (N_1316,N_1103,N_970);
nor U1317 (N_1317,In_1379,In_34);
nor U1318 (N_1318,In_1098,N_1057);
nor U1319 (N_1319,N_1084,In_540);
xor U1320 (N_1320,In_459,In_293);
nand U1321 (N_1321,N_1266,In_1255);
nand U1322 (N_1322,N_1270,N_1269);
and U1323 (N_1323,N_1107,N_1047);
and U1324 (N_1324,In_114,N_1089);
xor U1325 (N_1325,N_1253,N_974);
or U1326 (N_1326,N_1210,N_1094);
and U1327 (N_1327,N_711,N_1223);
nor U1328 (N_1328,In_32,In_359);
xor U1329 (N_1329,In_885,N_730);
and U1330 (N_1330,N_912,In_485);
or U1331 (N_1331,N_565,N_1261);
nand U1332 (N_1332,In_1615,N_1258);
or U1333 (N_1333,N_1175,In_1527);
or U1334 (N_1334,N_338,N_610);
nand U1335 (N_1335,N_598,In_635);
xor U1336 (N_1336,N_1000,N_1197);
and U1337 (N_1337,N_1069,In_493);
nand U1338 (N_1338,N_1272,N_733);
or U1339 (N_1339,N_351,In_1767);
nor U1340 (N_1340,In_136,N_444);
xor U1341 (N_1341,N_1226,N_755);
or U1342 (N_1342,N_659,N_1176);
xnor U1343 (N_1343,N_1208,N_1077);
nand U1344 (N_1344,In_955,N_1147);
nand U1345 (N_1345,N_1139,N_953);
or U1346 (N_1346,In_1105,N_799);
nand U1347 (N_1347,In_1590,In_814);
or U1348 (N_1348,N_1050,N_1192);
xnor U1349 (N_1349,N_1096,N_1168);
or U1350 (N_1350,N_1010,In_352);
nor U1351 (N_1351,N_834,N_1170);
xor U1352 (N_1352,N_597,N_937);
xor U1353 (N_1353,N_344,N_782);
nor U1354 (N_1354,N_124,N_491);
xor U1355 (N_1355,N_779,N_1040);
xnor U1356 (N_1356,N_1230,In_1771);
or U1357 (N_1357,N_80,N_383);
and U1358 (N_1358,N_1006,N_416);
nand U1359 (N_1359,In_1084,N_1033);
or U1360 (N_1360,N_306,In_1608);
nand U1361 (N_1361,N_1229,N_667);
and U1362 (N_1362,N_1177,In_329);
or U1363 (N_1363,N_558,N_1138);
nor U1364 (N_1364,N_1248,N_629);
nor U1365 (N_1365,In_371,In_892);
or U1366 (N_1366,In_78,In_1981);
xnor U1367 (N_1367,N_388,In_1054);
nor U1368 (N_1368,In_860,In_460);
xnor U1369 (N_1369,N_1108,N_603);
xor U1370 (N_1370,N_1167,In_679);
and U1371 (N_1371,N_908,In_1858);
or U1372 (N_1372,N_614,N_747);
xnor U1373 (N_1373,N_994,N_664);
nor U1374 (N_1374,In_432,In_757);
xnor U1375 (N_1375,N_1046,N_1246);
nor U1376 (N_1376,N_1185,N_1095);
and U1377 (N_1377,N_1079,N_1206);
or U1378 (N_1378,N_393,N_661);
and U1379 (N_1379,N_849,N_1242);
and U1380 (N_1380,N_852,N_1150);
and U1381 (N_1381,N_631,N_1237);
and U1382 (N_1382,N_198,In_1055);
nand U1383 (N_1383,N_1072,N_1216);
or U1384 (N_1384,N_554,In_263);
xnor U1385 (N_1385,N_950,N_637);
or U1386 (N_1386,N_1,In_937);
nand U1387 (N_1387,N_966,In_791);
or U1388 (N_1388,N_79,N_1125);
xnor U1389 (N_1389,In_141,In_619);
xor U1390 (N_1390,N_178,N_326);
nand U1391 (N_1391,N_688,N_1251);
and U1392 (N_1392,N_1068,In_1289);
xor U1393 (N_1393,N_1066,N_1075);
or U1394 (N_1394,N_879,In_447);
and U1395 (N_1395,N_1212,N_560);
and U1396 (N_1396,N_1099,N_600);
and U1397 (N_1397,N_232,In_334);
or U1398 (N_1398,N_1121,N_1060);
xnor U1399 (N_1399,N_1156,In_1385);
nor U1400 (N_1400,N_869,N_17);
and U1401 (N_1401,In_1010,N_1112);
or U1402 (N_1402,N_1128,N_569);
or U1403 (N_1403,N_1114,N_1155);
xnor U1404 (N_1404,In_1946,N_671);
nor U1405 (N_1405,In_196,N_933);
and U1406 (N_1406,In_92,In_991);
nor U1407 (N_1407,N_1268,In_1482);
nor U1408 (N_1408,In_450,In_1040);
or U1409 (N_1409,In_815,In_398);
or U1410 (N_1410,N_1163,N_1218);
nand U1411 (N_1411,In_1534,N_1023);
xor U1412 (N_1412,In_611,N_229);
and U1413 (N_1413,N_1227,N_694);
xnor U1414 (N_1414,N_892,N_236);
nand U1415 (N_1415,N_681,N_1090);
xnor U1416 (N_1416,N_1173,N_1109);
nor U1417 (N_1417,N_904,N_984);
or U1418 (N_1418,In_160,N_798);
or U1419 (N_1419,In_922,N_1064);
and U1420 (N_1420,In_979,N_1042);
nand U1421 (N_1421,In_449,N_868);
xor U1422 (N_1422,In_1150,N_1127);
nand U1423 (N_1423,In_1760,In_836);
and U1424 (N_1424,N_1153,In_361);
and U1425 (N_1425,N_373,N_763);
and U1426 (N_1426,N_1049,In_367);
or U1427 (N_1427,In_1891,N_384);
nand U1428 (N_1428,In_1604,N_1126);
nor U1429 (N_1429,N_526,N_977);
and U1430 (N_1430,N_1039,In_1594);
xor U1431 (N_1431,N_371,N_1207);
and U1432 (N_1432,In_1607,N_963);
nor U1433 (N_1433,N_758,In_1260);
xnor U1434 (N_1434,N_1113,N_548);
and U1435 (N_1435,In_90,In_1509);
nor U1436 (N_1436,N_575,N_1236);
nor U1437 (N_1437,In_1014,In_1282);
nor U1438 (N_1438,In_1227,In_1051);
and U1439 (N_1439,N_601,N_1193);
nand U1440 (N_1440,N_1195,In_1350);
and U1441 (N_1441,In_12,N_656);
nand U1442 (N_1442,N_1312,N_840);
xor U1443 (N_1443,In_445,N_928);
nor U1444 (N_1444,N_1374,N_1239);
xnor U1445 (N_1445,N_998,In_1976);
nor U1446 (N_1446,N_1341,N_856);
nor U1447 (N_1447,N_1395,N_958);
nor U1448 (N_1448,N_1323,N_1340);
or U1449 (N_1449,N_360,N_376);
nor U1450 (N_1450,N_1262,N_1406);
nor U1451 (N_1451,N_941,N_130);
or U1452 (N_1452,N_1234,N_1200);
xnor U1453 (N_1453,In_1469,In_1553);
or U1454 (N_1454,N_1336,N_1403);
nor U1455 (N_1455,N_1035,N_1302);
or U1456 (N_1456,In_1052,N_1123);
and U1457 (N_1457,In_1207,N_1339);
and U1458 (N_1458,In_1259,N_1390);
or U1459 (N_1459,N_1160,N_1008);
or U1460 (N_1460,In_1826,N_1131);
xnor U1461 (N_1461,N_1414,N_582);
and U1462 (N_1462,N_1219,In_932);
nor U1463 (N_1463,N_1005,N_34);
nand U1464 (N_1464,N_1282,N_1405);
or U1465 (N_1465,N_1315,N_888);
and U1466 (N_1466,N_1430,N_374);
or U1467 (N_1467,N_1361,N_1265);
or U1468 (N_1468,N_1217,N_1379);
nand U1469 (N_1469,In_1470,N_1007);
nand U1470 (N_1470,N_1398,N_171);
or U1471 (N_1471,N_1065,N_395);
xor U1472 (N_1472,N_964,N_1277);
xor U1473 (N_1473,N_1119,N_365);
xnor U1474 (N_1474,N_968,N_893);
or U1475 (N_1475,N_1364,In_510);
nand U1476 (N_1476,N_1295,N_959);
or U1477 (N_1477,N_1373,N_1369);
and U1478 (N_1478,In_1583,N_1205);
and U1479 (N_1479,N_660,N_1399);
and U1480 (N_1480,N_1321,N_1151);
nor U1481 (N_1481,N_1215,N_756);
xnor U1482 (N_1482,N_1174,N_1427);
or U1483 (N_1483,N_378,N_572);
or U1484 (N_1484,In_1486,N_1129);
or U1485 (N_1485,N_1134,N_1018);
or U1486 (N_1486,N_1318,N_531);
or U1487 (N_1487,In_1228,N_1306);
and U1488 (N_1488,N_1409,N_1169);
or U1489 (N_1489,N_1204,N_1357);
xor U1490 (N_1490,N_1106,N_1328);
xor U1491 (N_1491,N_1102,N_1137);
nor U1492 (N_1492,N_967,In_341);
nand U1493 (N_1493,N_931,N_206);
nor U1494 (N_1494,N_400,N_1428);
nand U1495 (N_1495,N_1201,N_1093);
nand U1496 (N_1496,N_625,N_1196);
xnor U1497 (N_1497,N_1412,N_1019);
nand U1498 (N_1498,N_1235,N_151);
nor U1499 (N_1499,N_738,N_1152);
xor U1500 (N_1500,N_1180,N_847);
nand U1501 (N_1501,N_1311,N_1280);
nand U1502 (N_1502,N_1162,N_1331);
or U1503 (N_1503,N_1419,N_1285);
xor U1504 (N_1504,N_1329,N_1291);
nor U1505 (N_1505,N_792,In_391);
and U1506 (N_1506,N_929,In_894);
xor U1507 (N_1507,N_1190,N_863);
xnor U1508 (N_1508,N_1045,N_1015);
xnor U1509 (N_1509,N_1353,In_1262);
or U1510 (N_1510,N_1377,N_1136);
nand U1511 (N_1511,In_1811,N_1299);
and U1512 (N_1512,N_369,N_1432);
nor U1513 (N_1513,N_658,N_741);
xor U1514 (N_1514,N_1186,In_530);
nor U1515 (N_1515,N_1159,In_225);
nor U1516 (N_1516,N_1307,N_1382);
nand U1517 (N_1517,N_810,N_42);
and U1518 (N_1518,In_1044,N_1238);
nor U1519 (N_1519,N_905,N_906);
nand U1520 (N_1520,N_1025,N_1327);
xnor U1521 (N_1521,In_35,N_297);
nand U1522 (N_1522,N_458,N_866);
nor U1523 (N_1523,N_1279,N_979);
nor U1524 (N_1524,N_838,N_945);
nor U1525 (N_1525,In_560,N_1271);
nand U1526 (N_1526,In_597,N_996);
and U1527 (N_1527,N_588,N_1256);
nand U1528 (N_1528,N_21,N_1014);
nor U1529 (N_1529,N_1352,In_1251);
nand U1530 (N_1530,N_1325,In_343);
xor U1531 (N_1531,N_1020,In_306);
xnor U1532 (N_1532,N_1166,N_475);
or U1533 (N_1533,N_66,N_1334);
nand U1534 (N_1534,N_396,N_710);
nor U1535 (N_1535,N_797,In_532);
or U1536 (N_1536,N_510,N_1202);
xor U1537 (N_1537,N_982,N_1400);
nor U1538 (N_1538,N_1289,N_1431);
nor U1539 (N_1539,N_1316,N_1402);
xnor U1540 (N_1540,N_1244,N_1408);
nand U1541 (N_1541,N_1013,In_426);
or U1542 (N_1542,N_479,In_288);
nor U1543 (N_1543,N_1345,In_1269);
nor U1544 (N_1544,N_1080,N_1397);
or U1545 (N_1545,N_712,N_1228);
nor U1546 (N_1546,N_1296,N_1273);
xnor U1547 (N_1547,N_807,N_1343);
nor U1548 (N_1548,N_1385,N_1146);
nand U1549 (N_1549,N_850,N_1250);
or U1550 (N_1550,N_739,N_985);
or U1551 (N_1551,N_435,N_1143);
and U1552 (N_1552,In_1036,N_494);
nor U1553 (N_1553,In_644,N_1300);
xnor U1554 (N_1554,N_1209,N_1211);
and U1555 (N_1555,N_1100,N_1337);
nand U1556 (N_1556,N_975,N_1132);
nor U1557 (N_1557,N_1338,N_1181);
xor U1558 (N_1558,N_858,N_1281);
and U1559 (N_1559,In_1979,In_534);
nor U1560 (N_1560,N_1144,N_1422);
nor U1561 (N_1561,N_1087,N_1333);
and U1562 (N_1562,In_1487,N_890);
nand U1563 (N_1563,N_1194,N_983);
or U1564 (N_1564,N_1384,N_1425);
or U1565 (N_1565,N_940,N_1351);
or U1566 (N_1566,N_8,N_586);
nor U1567 (N_1567,In_1791,N_668);
nand U1568 (N_1568,N_515,N_978);
nor U1569 (N_1569,N_765,N_644);
xnor U1570 (N_1570,In_541,N_1342);
xnor U1571 (N_1571,In_657,N_898);
xor U1572 (N_1572,N_839,N_1298);
xor U1573 (N_1573,N_1393,N_1292);
or U1574 (N_1574,N_1247,N_1284);
xor U1575 (N_1575,N_1240,N_1404);
nor U1576 (N_1576,In_4,In_1577);
nor U1577 (N_1577,N_988,N_1388);
nand U1578 (N_1578,N_897,N_1378);
nor U1579 (N_1579,N_120,N_1263);
and U1580 (N_1580,N_323,N_1101);
or U1581 (N_1581,In_1373,N_1347);
and U1582 (N_1582,N_1254,N_1115);
and U1583 (N_1583,N_1274,N_471);
nand U1584 (N_1584,In_1277,N_1376);
or U1585 (N_1585,N_1350,N_595);
nand U1586 (N_1586,N_827,N_1359);
and U1587 (N_1587,N_1314,N_1118);
and U1588 (N_1588,N_831,N_1283);
xor U1589 (N_1589,N_907,N_1122);
and U1590 (N_1590,N_1070,N_685);
and U1591 (N_1591,N_1133,N_1415);
and U1592 (N_1592,N_1416,N_1294);
and U1593 (N_1593,N_816,N_1335);
nor U1594 (N_1594,N_1012,N_1310);
xor U1595 (N_1595,N_1383,N_1366);
xnor U1596 (N_1596,In_1146,In_1243);
xor U1597 (N_1597,In_1816,N_1330);
or U1598 (N_1598,N_833,N_1426);
nor U1599 (N_1599,In_281,N_1420);
nand U1600 (N_1600,N_1054,N_1411);
xor U1601 (N_1601,N_1124,N_1386);
or U1602 (N_1602,N_1507,N_1407);
or U1603 (N_1603,In_1086,N_642);
and U1604 (N_1604,N_1452,N_1387);
and U1605 (N_1605,N_1221,N_1290);
xnor U1606 (N_1606,N_630,N_1589);
or U1607 (N_1607,In_1063,In_1281);
nand U1608 (N_1608,N_1004,N_1593);
and U1609 (N_1609,N_1488,N_1472);
and U1610 (N_1610,N_1582,N_1332);
xnor U1611 (N_1611,In_1597,N_1297);
and U1612 (N_1612,N_1497,N_1276);
nor U1613 (N_1613,N_1449,In_1755);
and U1614 (N_1614,N_1566,N_1367);
and U1615 (N_1615,N_1511,N_1220);
and U1616 (N_1616,In_1090,N_1564);
nand U1617 (N_1617,N_788,N_1499);
and U1618 (N_1618,N_881,N_209);
or U1619 (N_1619,N_1465,N_1293);
or U1620 (N_1620,N_1462,N_877);
nand U1621 (N_1621,N_1368,N_1439);
xor U1622 (N_1622,In_495,N_1528);
and U1623 (N_1623,N_1471,N_1509);
and U1624 (N_1624,N_1389,N_1222);
and U1625 (N_1625,N_1464,N_1362);
and U1626 (N_1626,N_1322,N_1067);
or U1627 (N_1627,N_441,N_1555);
and U1628 (N_1628,In_805,N_32);
or U1629 (N_1629,N_193,N_981);
nand U1630 (N_1630,N_1356,N_1287);
xnor U1631 (N_1631,N_1529,N_1392);
xnor U1632 (N_1632,N_1554,N_1568);
nor U1633 (N_1633,N_1578,N_497);
nor U1634 (N_1634,N_1255,N_695);
or U1635 (N_1635,N_1494,N_1493);
nand U1636 (N_1636,In_1710,N_460);
nor U1637 (N_1637,N_1130,N_1518);
nand U1638 (N_1638,N_1490,In_1620);
nor U1639 (N_1639,N_1417,N_1520);
xnor U1640 (N_1640,N_1410,N_591);
nor U1641 (N_1641,N_1451,N_624);
or U1642 (N_1642,N_1433,N_1508);
nor U1643 (N_1643,N_1461,N_1148);
nor U1644 (N_1644,N_1436,N_1538);
nor U1645 (N_1645,N_1561,In_202);
and U1646 (N_1646,N_1442,N_1260);
nand U1647 (N_1647,N_1503,N_1288);
xor U1648 (N_1648,N_1319,N_1598);
xnor U1649 (N_1649,N_1523,N_729);
or U1650 (N_1650,N_1394,N_1303);
nor U1651 (N_1651,N_619,N_1453);
xor U1652 (N_1652,N_314,N_1324);
and U1653 (N_1653,N_1548,In_1129);
xor U1654 (N_1654,N_1135,N_1081);
or U1655 (N_1655,N_1463,N_1381);
nor U1656 (N_1656,N_1543,N_1571);
and U1657 (N_1657,N_1535,N_432);
xor U1658 (N_1658,N_1501,N_1446);
nand U1659 (N_1659,N_1559,In_322);
nor U1660 (N_1660,N_1071,N_1372);
and U1661 (N_1661,N_146,N_1203);
or U1662 (N_1662,In_1763,N_1456);
and U1663 (N_1663,N_539,N_1541);
nor U1664 (N_1664,N_1551,N_1443);
and U1665 (N_1665,N_1348,N_1585);
xnor U1666 (N_1666,N_1224,N_1521);
nor U1667 (N_1667,N_1252,N_1179);
nand U1668 (N_1668,N_1172,In_1833);
nand U1669 (N_1669,N_1587,N_1475);
or U1670 (N_1670,N_835,N_865);
and U1671 (N_1671,N_1592,N_962);
nand U1672 (N_1672,N_1154,N_1478);
nor U1673 (N_1673,In_554,In_1758);
or U1674 (N_1674,N_1574,N_1560);
nor U1675 (N_1675,N_1575,In_1776);
nor U1676 (N_1676,N_1098,N_1309);
nor U1677 (N_1677,N_1085,In_1454);
or U1678 (N_1678,N_1375,In_177);
xor U1679 (N_1679,N_1448,N_1579);
and U1680 (N_1680,N_1477,N_995);
nor U1681 (N_1681,N_1599,N_705);
nor U1682 (N_1682,In_1135,N_703);
or U1683 (N_1683,N_1187,N_1570);
nand U1684 (N_1684,N_1308,N_1542);
or U1685 (N_1685,In_1913,N_1161);
or U1686 (N_1686,N_1074,N_1565);
nand U1687 (N_1687,N_1435,In_822);
and U1688 (N_1688,N_1346,N_557);
and U1689 (N_1689,N_1572,N_1577);
nand U1690 (N_1690,N_1301,N_1441);
nor U1691 (N_1691,N_716,N_1522);
nor U1692 (N_1692,N_1076,N_1259);
or U1693 (N_1693,N_27,N_1583);
nand U1694 (N_1694,In_231,N_1320);
xor U1695 (N_1695,N_1532,N_1105);
nand U1696 (N_1696,N_1495,N_1549);
nor U1697 (N_1697,N_364,N_26);
xor U1698 (N_1698,N_1370,N_1531);
and U1699 (N_1699,N_1595,N_902);
or U1700 (N_1700,N_1539,N_1454);
and U1701 (N_1701,N_1199,N_290);
and U1702 (N_1702,N_1496,N_1483);
and U1703 (N_1703,N_1358,N_1498);
or U1704 (N_1704,N_948,N_1249);
nand U1705 (N_1705,In_358,N_1326);
nand U1706 (N_1706,N_1537,In_87);
or U1707 (N_1707,N_324,N_791);
nor U1708 (N_1708,N_1188,N_1502);
or U1709 (N_1709,In_301,N_1547);
nor U1710 (N_1710,N_1524,In_1975);
nor U1711 (N_1711,N_1457,N_1233);
xnor U1712 (N_1712,In_328,N_1213);
and U1713 (N_1713,N_762,N_1164);
nand U1714 (N_1714,N_1149,N_1032);
and U1715 (N_1715,N_997,N_1487);
nor U1716 (N_1716,N_1525,In_1178);
or U1717 (N_1717,N_1505,N_1344);
or U1718 (N_1718,N_1591,N_1473);
nor U1719 (N_1719,N_921,N_483);
xnor U1720 (N_1720,In_102,N_1482);
nand U1721 (N_1721,N_1467,N_1401);
nand U1722 (N_1722,N_1527,N_693);
or U1723 (N_1723,N_1396,N_1275);
xnor U1724 (N_1724,In_1545,N_1510);
and U1725 (N_1725,N_1540,In_1230);
nand U1726 (N_1726,N_1474,N_1513);
xor U1727 (N_1727,N_47,N_1580);
nand U1728 (N_1728,N_1429,N_1317);
nor U1729 (N_1729,N_672,In_279);
and U1730 (N_1730,N_505,N_961);
nand U1731 (N_1731,N_932,N_1184);
nand U1732 (N_1732,N_468,In_112);
nor U1733 (N_1733,N_1470,N_1056);
and U1734 (N_1734,In_1591,N_1536);
and U1735 (N_1735,N_1380,In_1371);
nor U1736 (N_1736,N_1545,In_977);
xnor U1737 (N_1737,N_1034,N_1469);
and U1738 (N_1738,N_1476,N_1597);
nand U1739 (N_1739,N_1576,N_1051);
xnor U1740 (N_1740,N_1437,N_1588);
nand U1741 (N_1741,N_1486,In_559);
nor U1742 (N_1742,N_1550,N_1460);
xor U1743 (N_1743,N_1447,N_1492);
xnor U1744 (N_1744,N_1444,N_1544);
nand U1745 (N_1745,In_157,N_1371);
or U1746 (N_1746,N_1556,N_1466);
or U1747 (N_1747,N_1354,N_836);
nand U1748 (N_1748,N_1530,N_1055);
nor U1749 (N_1749,N_533,In_633);
or U1750 (N_1750,N_1557,N_1264);
and U1751 (N_1751,N_1590,N_459);
nand U1752 (N_1752,N_1479,N_1519);
nor U1753 (N_1753,N_1573,N_1581);
and U1754 (N_1754,N_1365,In_1774);
nor U1755 (N_1755,In_1043,N_1491);
nor U1756 (N_1756,N_1418,In_340);
xor U1757 (N_1757,N_1434,N_1198);
and U1758 (N_1758,N_285,N_496);
nor U1759 (N_1759,N_1489,N_1313);
nand U1760 (N_1760,N_1742,N_943);
or U1761 (N_1761,N_1614,N_1727);
and U1762 (N_1762,N_1753,N_1423);
or U1763 (N_1763,N_1512,N_1676);
or U1764 (N_1764,N_1748,N_1745);
xor U1765 (N_1765,N_1673,N_1684);
or U1766 (N_1766,N_1715,N_1305);
nand U1767 (N_1767,N_1705,N_1629);
nor U1768 (N_1768,N_1526,N_443);
nor U1769 (N_1769,N_909,N_145);
nor U1770 (N_1770,N_1702,In_210);
nor U1771 (N_1771,N_1634,N_1558);
nor U1772 (N_1772,N_1623,N_1140);
and U1773 (N_1773,N_1601,N_1438);
or U1774 (N_1774,N_1756,N_1650);
nand U1775 (N_1775,N_1594,N_1613);
or U1776 (N_1776,N_1720,N_1724);
nand U1777 (N_1777,N_1214,N_1692);
nor U1778 (N_1778,N_1567,N_1605);
or U1779 (N_1779,N_1730,N_1363);
nand U1780 (N_1780,N_1743,N_1749);
xor U1781 (N_1781,N_1183,N_1754);
nor U1782 (N_1782,N_1620,N_1744);
nor U1783 (N_1783,N_1391,N_1455);
nor U1784 (N_1784,N_1637,N_1612);
nand U1785 (N_1785,N_1717,N_1678);
xor U1786 (N_1786,N_1671,N_28);
or U1787 (N_1787,N_1450,N_1304);
and U1788 (N_1788,N_1189,In_1217);
or U1789 (N_1789,N_1716,N_1533);
nand U1790 (N_1790,N_1711,N_1627);
or U1791 (N_1791,N_1752,N_1685);
xnor U1792 (N_1792,N_1642,N_1706);
and U1793 (N_1793,N_1710,N_1751);
nor U1794 (N_1794,N_1718,N_1622);
nor U1795 (N_1795,N_1586,N_1640);
xnor U1796 (N_1796,N_1611,N_1514);
nor U1797 (N_1797,N_1500,N_1757);
xor U1798 (N_1798,N_1158,N_1602);
or U1799 (N_1799,N_1696,N_1421);
or U1800 (N_1800,N_1355,N_1700);
or U1801 (N_1801,N_1726,N_1680);
nor U1802 (N_1802,N_1615,N_1660);
nor U1803 (N_1803,N_1458,N_1610);
nor U1804 (N_1804,N_1662,N_1504);
nand U1805 (N_1805,N_864,N_896);
and U1806 (N_1806,N_1728,N_1643);
xnor U1807 (N_1807,N_1506,N_504);
or U1808 (N_1808,N_1714,N_1731);
xnor U1809 (N_1809,N_1534,N_1546);
and U1810 (N_1810,N_1651,In_128);
and U1811 (N_1811,In_121,N_1600);
or U1812 (N_1812,N_1687,N_1695);
and U1813 (N_1813,N_1635,N_1563);
nor U1814 (N_1814,N_1698,N_1517);
and U1815 (N_1815,N_1704,N_1670);
and U1816 (N_1816,N_1424,N_1693);
and U1817 (N_1817,N_1658,N_1481);
or U1818 (N_1818,N_1569,N_1739);
xnor U1819 (N_1819,N_1633,N_1689);
xnor U1820 (N_1820,N_1562,N_1120);
nor U1821 (N_1821,In_999,N_1707);
xor U1822 (N_1822,N_1652,N_1674);
xnor U1823 (N_1823,N_1584,N_1661);
nand U1824 (N_1824,N_1683,In_1815);
xnor U1825 (N_1825,N_1734,N_1459);
xor U1826 (N_1826,N_1606,N_1759);
nand U1827 (N_1827,N_1733,N_266);
or U1828 (N_1828,N_1413,N_1618);
nand U1829 (N_1829,N_1675,N_1750);
xnor U1830 (N_1830,N_1626,N_1735);
xor U1831 (N_1831,N_1485,N_1516);
nand U1832 (N_1832,N_1639,N_1657);
and U1833 (N_1833,N_1758,N_1740);
xor U1834 (N_1834,N_1668,N_1607);
nor U1835 (N_1835,N_1723,N_1349);
xor U1836 (N_1836,N_1691,N_1712);
and U1837 (N_1837,N_1737,N_1608);
and U1838 (N_1838,N_1672,N_1624);
nor U1839 (N_1839,N_1641,N_1738);
nand U1840 (N_1840,N_1682,N_1664);
nand U1841 (N_1841,N_1690,N_1552);
nor U1842 (N_1842,N_1677,N_1713);
nor U1843 (N_1843,N_1708,In_349);
nor U1844 (N_1844,N_1515,N_1694);
or U1845 (N_1845,N_1646,N_1663);
nor U1846 (N_1846,N_1621,N_1604);
and U1847 (N_1847,N_1736,N_1647);
xnor U1848 (N_1848,N_1679,N_1699);
nor U1849 (N_1849,N_1648,N_1617);
nor U1850 (N_1850,N_1709,N_1653);
nand U1851 (N_1851,N_1286,N_766);
or U1852 (N_1852,N_1632,N_1619);
and U1853 (N_1853,N_1725,N_1649);
nand U1854 (N_1854,N_1630,N_1360);
or U1855 (N_1855,N_1645,N_915);
nand U1856 (N_1856,N_1681,N_1654);
nor U1857 (N_1857,N_1484,N_1747);
xnor U1858 (N_1858,N_1721,N_1666);
nor U1859 (N_1859,N_1703,N_1722);
and U1860 (N_1860,In_1377,N_1746);
nor U1861 (N_1861,N_1729,N_1732);
nand U1862 (N_1862,N_1445,N_1440);
nand U1863 (N_1863,In_1461,N_1697);
and U1864 (N_1864,N_1686,N_1638);
and U1865 (N_1865,N_1603,N_1665);
and U1866 (N_1866,N_1741,N_1701);
nor U1867 (N_1867,N_1719,N_1616);
or U1868 (N_1868,In_1714,N_1596);
nand U1869 (N_1869,N_1656,N_1625);
and U1870 (N_1870,N_1669,N_1636);
xnor U1871 (N_1871,N_1655,N_1659);
or U1872 (N_1872,N_348,N_1553);
nor U1873 (N_1873,N_1191,N_1688);
nand U1874 (N_1874,N_1480,N_1609);
nand U1875 (N_1875,N_1053,N_636);
nand U1876 (N_1876,N_1631,N_1644);
nor U1877 (N_1877,N_1755,In_1722);
nor U1878 (N_1878,N_1628,N_1667);
nor U1879 (N_1879,N_1468,N_1243);
xor U1880 (N_1880,N_1514,N_1603);
xnor U1881 (N_1881,In_1217,N_1600);
nand U1882 (N_1882,In_1714,N_1445);
and U1883 (N_1883,N_1676,N_1612);
nor U1884 (N_1884,N_1740,N_1697);
and U1885 (N_1885,N_1445,N_1504);
nor U1886 (N_1886,N_1485,In_1815);
xnor U1887 (N_1887,N_1649,N_1440);
nand U1888 (N_1888,N_1747,N_1634);
nand U1889 (N_1889,N_1684,N_1459);
or U1890 (N_1890,N_1671,N_1707);
or U1891 (N_1891,N_1653,N_1723);
nand U1892 (N_1892,N_1756,N_1725);
xnor U1893 (N_1893,N_1632,N_636);
nor U1894 (N_1894,N_1752,N_1712);
and U1895 (N_1895,N_1711,N_1740);
and U1896 (N_1896,N_1655,N_1652);
or U1897 (N_1897,N_1664,N_1660);
nor U1898 (N_1898,N_1700,N_1716);
xor U1899 (N_1899,N_1610,N_1667);
nand U1900 (N_1900,N_1654,N_1183);
nor U1901 (N_1901,N_1608,N_864);
or U1902 (N_1902,N_1642,N_1656);
and U1903 (N_1903,N_1722,N_1678);
nor U1904 (N_1904,N_1733,N_1709);
nand U1905 (N_1905,N_1504,N_1750);
xnor U1906 (N_1906,N_1628,N_1607);
nand U1907 (N_1907,N_1619,N_1666);
nor U1908 (N_1908,N_1243,N_1700);
and U1909 (N_1909,In_121,N_1553);
or U1910 (N_1910,N_1625,N_1603);
xnor U1911 (N_1911,N_1558,In_1377);
nor U1912 (N_1912,In_1461,N_1363);
and U1913 (N_1913,N_1755,N_1711);
or U1914 (N_1914,N_1615,N_1481);
nor U1915 (N_1915,N_1667,N_1708);
xor U1916 (N_1916,N_1754,N_1413);
xnor U1917 (N_1917,N_1744,N_1714);
or U1918 (N_1918,N_1191,N_1605);
or U1919 (N_1919,N_1647,In_1815);
nand U1920 (N_1920,N_1870,N_1874);
or U1921 (N_1921,N_1797,N_1902);
and U1922 (N_1922,N_1798,N_1833);
or U1923 (N_1923,N_1796,N_1762);
or U1924 (N_1924,N_1832,N_1851);
and U1925 (N_1925,N_1800,N_1914);
nand U1926 (N_1926,N_1845,N_1811);
and U1927 (N_1927,N_1881,N_1769);
or U1928 (N_1928,N_1831,N_1862);
or U1929 (N_1929,N_1784,N_1778);
or U1930 (N_1930,N_1821,N_1764);
or U1931 (N_1931,N_1918,N_1846);
xnor U1932 (N_1932,N_1901,N_1850);
nand U1933 (N_1933,N_1854,N_1788);
nand U1934 (N_1934,N_1865,N_1875);
xnor U1935 (N_1935,N_1820,N_1791);
xor U1936 (N_1936,N_1799,N_1830);
or U1937 (N_1937,N_1853,N_1899);
xor U1938 (N_1938,N_1896,N_1891);
xor U1939 (N_1939,N_1824,N_1837);
nand U1940 (N_1940,N_1781,N_1804);
and U1941 (N_1941,N_1916,N_1790);
xnor U1942 (N_1942,N_1774,N_1841);
xnor U1943 (N_1943,N_1909,N_1763);
and U1944 (N_1944,N_1783,N_1908);
xnor U1945 (N_1945,N_1767,N_1879);
or U1946 (N_1946,N_1882,N_1813);
xor U1947 (N_1947,N_1911,N_1838);
and U1948 (N_1948,N_1885,N_1906);
or U1949 (N_1949,N_1771,N_1856);
nand U1950 (N_1950,N_1892,N_1807);
or U1951 (N_1951,N_1768,N_1872);
and U1952 (N_1952,N_1852,N_1910);
nand U1953 (N_1953,N_1913,N_1795);
or U1954 (N_1954,N_1818,N_1794);
or U1955 (N_1955,N_1775,N_1786);
nand U1956 (N_1956,N_1883,N_1772);
or U1957 (N_1957,N_1888,N_1871);
or U1958 (N_1958,N_1808,N_1844);
and U1959 (N_1959,N_1822,N_1919);
nand U1960 (N_1960,N_1836,N_1825);
or U1961 (N_1961,N_1840,N_1814);
or U1962 (N_1962,N_1770,N_1864);
nor U1963 (N_1963,N_1868,N_1785);
nand U1964 (N_1964,N_1760,N_1895);
nand U1965 (N_1965,N_1866,N_1863);
nand U1966 (N_1966,N_1827,N_1878);
xor U1967 (N_1967,N_1861,N_1803);
nand U1968 (N_1968,N_1907,N_1806);
and U1969 (N_1969,N_1773,N_1904);
nand U1970 (N_1970,N_1843,N_1887);
xnor U1971 (N_1971,N_1761,N_1873);
nor U1972 (N_1972,N_1826,N_1877);
nor U1973 (N_1973,N_1823,N_1859);
xor U1974 (N_1974,N_1917,N_1809);
and U1975 (N_1975,N_1793,N_1839);
and U1976 (N_1976,N_1815,N_1812);
and U1977 (N_1977,N_1912,N_1886);
xor U1978 (N_1978,N_1816,N_1894);
nand U1979 (N_1979,N_1858,N_1869);
nand U1980 (N_1980,N_1819,N_1787);
nor U1981 (N_1981,N_1765,N_1889);
nand U1982 (N_1982,N_1893,N_1860);
nand U1983 (N_1983,N_1780,N_1849);
nand U1984 (N_1984,N_1777,N_1801);
nand U1985 (N_1985,N_1805,N_1857);
nand U1986 (N_1986,N_1915,N_1880);
nor U1987 (N_1987,N_1829,N_1782);
nor U1988 (N_1988,N_1817,N_1903);
or U1989 (N_1989,N_1792,N_1900);
nor U1990 (N_1990,N_1789,N_1835);
nor U1991 (N_1991,N_1905,N_1766);
nor U1992 (N_1992,N_1898,N_1867);
or U1993 (N_1993,N_1828,N_1776);
or U1994 (N_1994,N_1848,N_1834);
nand U1995 (N_1995,N_1842,N_1884);
xnor U1996 (N_1996,N_1779,N_1876);
xnor U1997 (N_1997,N_1855,N_1897);
or U1998 (N_1998,N_1802,N_1847);
and U1999 (N_1999,N_1810,N_1890);
xor U2000 (N_2000,N_1785,N_1871);
xor U2001 (N_2001,N_1914,N_1843);
or U2002 (N_2002,N_1866,N_1857);
or U2003 (N_2003,N_1908,N_1897);
nand U2004 (N_2004,N_1761,N_1760);
nor U2005 (N_2005,N_1884,N_1869);
nor U2006 (N_2006,N_1779,N_1843);
nand U2007 (N_2007,N_1761,N_1874);
or U2008 (N_2008,N_1852,N_1906);
nand U2009 (N_2009,N_1815,N_1833);
or U2010 (N_2010,N_1849,N_1785);
nand U2011 (N_2011,N_1904,N_1801);
nand U2012 (N_2012,N_1912,N_1895);
and U2013 (N_2013,N_1845,N_1896);
or U2014 (N_2014,N_1870,N_1784);
nor U2015 (N_2015,N_1814,N_1765);
and U2016 (N_2016,N_1766,N_1783);
and U2017 (N_2017,N_1839,N_1789);
nor U2018 (N_2018,N_1834,N_1899);
or U2019 (N_2019,N_1857,N_1771);
or U2020 (N_2020,N_1855,N_1761);
xor U2021 (N_2021,N_1874,N_1815);
or U2022 (N_2022,N_1780,N_1802);
and U2023 (N_2023,N_1911,N_1806);
nand U2024 (N_2024,N_1878,N_1862);
or U2025 (N_2025,N_1810,N_1898);
nand U2026 (N_2026,N_1802,N_1841);
or U2027 (N_2027,N_1916,N_1765);
and U2028 (N_2028,N_1917,N_1803);
nor U2029 (N_2029,N_1911,N_1809);
xor U2030 (N_2030,N_1890,N_1859);
and U2031 (N_2031,N_1827,N_1776);
and U2032 (N_2032,N_1823,N_1878);
nand U2033 (N_2033,N_1814,N_1808);
nand U2034 (N_2034,N_1867,N_1802);
nor U2035 (N_2035,N_1766,N_1822);
nand U2036 (N_2036,N_1905,N_1893);
or U2037 (N_2037,N_1916,N_1811);
nor U2038 (N_2038,N_1767,N_1820);
and U2039 (N_2039,N_1777,N_1886);
xnor U2040 (N_2040,N_1855,N_1862);
nor U2041 (N_2041,N_1770,N_1781);
nand U2042 (N_2042,N_1824,N_1762);
nor U2043 (N_2043,N_1897,N_1866);
and U2044 (N_2044,N_1786,N_1801);
nand U2045 (N_2045,N_1815,N_1777);
nand U2046 (N_2046,N_1833,N_1840);
xnor U2047 (N_2047,N_1856,N_1875);
and U2048 (N_2048,N_1856,N_1794);
nand U2049 (N_2049,N_1833,N_1907);
and U2050 (N_2050,N_1898,N_1767);
and U2051 (N_2051,N_1794,N_1863);
and U2052 (N_2052,N_1899,N_1763);
nor U2053 (N_2053,N_1899,N_1788);
nand U2054 (N_2054,N_1771,N_1891);
nor U2055 (N_2055,N_1912,N_1766);
xnor U2056 (N_2056,N_1919,N_1785);
nand U2057 (N_2057,N_1831,N_1841);
nand U2058 (N_2058,N_1884,N_1760);
nand U2059 (N_2059,N_1785,N_1783);
and U2060 (N_2060,N_1886,N_1893);
or U2061 (N_2061,N_1837,N_1788);
nand U2062 (N_2062,N_1842,N_1907);
and U2063 (N_2063,N_1807,N_1897);
nand U2064 (N_2064,N_1836,N_1889);
or U2065 (N_2065,N_1873,N_1836);
nand U2066 (N_2066,N_1874,N_1812);
or U2067 (N_2067,N_1806,N_1791);
and U2068 (N_2068,N_1846,N_1866);
or U2069 (N_2069,N_1824,N_1850);
xnor U2070 (N_2070,N_1783,N_1919);
nor U2071 (N_2071,N_1820,N_1808);
and U2072 (N_2072,N_1826,N_1851);
and U2073 (N_2073,N_1817,N_1809);
or U2074 (N_2074,N_1767,N_1899);
xnor U2075 (N_2075,N_1891,N_1801);
nor U2076 (N_2076,N_1774,N_1825);
or U2077 (N_2077,N_1850,N_1813);
nor U2078 (N_2078,N_1779,N_1883);
xnor U2079 (N_2079,N_1785,N_1800);
or U2080 (N_2080,N_1975,N_2069);
nand U2081 (N_2081,N_1927,N_2045);
and U2082 (N_2082,N_2047,N_1996);
and U2083 (N_2083,N_1925,N_2048);
nand U2084 (N_2084,N_2010,N_1974);
or U2085 (N_2085,N_2022,N_2038);
or U2086 (N_2086,N_2056,N_2067);
nand U2087 (N_2087,N_1958,N_1960);
and U2088 (N_2088,N_1934,N_2000);
nand U2089 (N_2089,N_1994,N_1935);
nand U2090 (N_2090,N_2009,N_1998);
or U2091 (N_2091,N_1968,N_2029);
nand U2092 (N_2092,N_2071,N_2033);
and U2093 (N_2093,N_1963,N_1976);
nand U2094 (N_2094,N_1982,N_1947);
and U2095 (N_2095,N_2065,N_2060);
xor U2096 (N_2096,N_2053,N_1950);
and U2097 (N_2097,N_2030,N_2079);
xor U2098 (N_2098,N_1999,N_1940);
xor U2099 (N_2099,N_1990,N_2021);
and U2100 (N_2100,N_1929,N_1964);
xor U2101 (N_2101,N_2017,N_1933);
xor U2102 (N_2102,N_1983,N_1961);
and U2103 (N_2103,N_2051,N_1920);
xor U2104 (N_2104,N_1944,N_2059);
and U2105 (N_2105,N_2003,N_1997);
nand U2106 (N_2106,N_2011,N_2004);
xnor U2107 (N_2107,N_1995,N_2024);
nand U2108 (N_2108,N_1943,N_2001);
nor U2109 (N_2109,N_2007,N_1993);
nand U2110 (N_2110,N_1985,N_2023);
or U2111 (N_2111,N_1955,N_2002);
nand U2112 (N_2112,N_2037,N_1932);
nor U2113 (N_2113,N_2014,N_1967);
nor U2114 (N_2114,N_2061,N_1965);
xor U2115 (N_2115,N_2031,N_2042);
nand U2116 (N_2116,N_1991,N_2040);
xor U2117 (N_2117,N_2054,N_2027);
nand U2118 (N_2118,N_2066,N_1977);
xor U2119 (N_2119,N_2063,N_2025);
and U2120 (N_2120,N_1941,N_1948);
xor U2121 (N_2121,N_2028,N_2020);
xnor U2122 (N_2122,N_2046,N_2043);
xor U2123 (N_2123,N_2052,N_2013);
nand U2124 (N_2124,N_1954,N_1969);
nor U2125 (N_2125,N_2068,N_2026);
xnor U2126 (N_2126,N_1989,N_1937);
xor U2127 (N_2127,N_2012,N_1942);
nand U2128 (N_2128,N_1946,N_1981);
or U2129 (N_2129,N_2070,N_1986);
xnor U2130 (N_2130,N_2015,N_2058);
nand U2131 (N_2131,N_2074,N_2032);
and U2132 (N_2132,N_1957,N_1921);
nor U2133 (N_2133,N_1980,N_1962);
nor U2134 (N_2134,N_1928,N_1987);
nor U2135 (N_2135,N_2072,N_2064);
xor U2136 (N_2136,N_1971,N_2036);
nand U2137 (N_2137,N_2049,N_2057);
nor U2138 (N_2138,N_1992,N_2077);
and U2139 (N_2139,N_2073,N_2019);
nor U2140 (N_2140,N_1923,N_1938);
or U2141 (N_2141,N_1924,N_2055);
and U2142 (N_2142,N_2076,N_1931);
xor U2143 (N_2143,N_1951,N_1945);
nand U2144 (N_2144,N_1939,N_2008);
and U2145 (N_2145,N_2006,N_2041);
or U2146 (N_2146,N_1984,N_1953);
or U2147 (N_2147,N_2039,N_1936);
nor U2148 (N_2148,N_2075,N_1978);
and U2149 (N_2149,N_1956,N_2005);
or U2150 (N_2150,N_1959,N_1970);
and U2151 (N_2151,N_1973,N_1922);
and U2152 (N_2152,N_2034,N_1930);
nor U2153 (N_2153,N_1972,N_1949);
nor U2154 (N_2154,N_2044,N_1979);
nor U2155 (N_2155,N_1926,N_2062);
xor U2156 (N_2156,N_2050,N_2035);
nor U2157 (N_2157,N_2078,N_1988);
nor U2158 (N_2158,N_2018,N_1966);
nand U2159 (N_2159,N_2016,N_1952);
nand U2160 (N_2160,N_1965,N_2013);
and U2161 (N_2161,N_1964,N_2055);
nor U2162 (N_2162,N_2020,N_2042);
and U2163 (N_2163,N_2050,N_1922);
or U2164 (N_2164,N_1928,N_1977);
and U2165 (N_2165,N_2002,N_2007);
or U2166 (N_2166,N_1923,N_1936);
nor U2167 (N_2167,N_2051,N_1936);
or U2168 (N_2168,N_2043,N_2021);
xor U2169 (N_2169,N_2048,N_2076);
xnor U2170 (N_2170,N_2048,N_1938);
nand U2171 (N_2171,N_2010,N_2032);
and U2172 (N_2172,N_2047,N_2041);
nand U2173 (N_2173,N_2055,N_1993);
or U2174 (N_2174,N_1990,N_2009);
nor U2175 (N_2175,N_1932,N_2077);
nand U2176 (N_2176,N_1950,N_2072);
and U2177 (N_2177,N_2040,N_2011);
xnor U2178 (N_2178,N_1960,N_2061);
nand U2179 (N_2179,N_1967,N_1990);
nand U2180 (N_2180,N_2060,N_2048);
or U2181 (N_2181,N_2031,N_1954);
and U2182 (N_2182,N_1988,N_1921);
nor U2183 (N_2183,N_2045,N_2002);
and U2184 (N_2184,N_1928,N_2047);
or U2185 (N_2185,N_1972,N_2061);
xnor U2186 (N_2186,N_2006,N_2007);
nor U2187 (N_2187,N_1998,N_2074);
nor U2188 (N_2188,N_1973,N_1933);
or U2189 (N_2189,N_1940,N_1991);
or U2190 (N_2190,N_2015,N_2052);
nor U2191 (N_2191,N_2051,N_1957);
and U2192 (N_2192,N_1994,N_2039);
and U2193 (N_2193,N_2060,N_1939);
or U2194 (N_2194,N_2062,N_2007);
nand U2195 (N_2195,N_2032,N_1970);
or U2196 (N_2196,N_2040,N_1983);
or U2197 (N_2197,N_2060,N_2030);
nand U2198 (N_2198,N_2060,N_1927);
nand U2199 (N_2199,N_1991,N_1921);
nor U2200 (N_2200,N_2044,N_2047);
nand U2201 (N_2201,N_2043,N_2031);
and U2202 (N_2202,N_2009,N_2049);
nand U2203 (N_2203,N_2079,N_2002);
nor U2204 (N_2204,N_1931,N_2022);
or U2205 (N_2205,N_1938,N_2039);
nand U2206 (N_2206,N_2004,N_2048);
xor U2207 (N_2207,N_1950,N_1998);
and U2208 (N_2208,N_1970,N_1932);
or U2209 (N_2209,N_1951,N_2072);
or U2210 (N_2210,N_2046,N_2005);
nand U2211 (N_2211,N_1952,N_2028);
and U2212 (N_2212,N_2051,N_1932);
xor U2213 (N_2213,N_2065,N_2046);
and U2214 (N_2214,N_1958,N_2063);
and U2215 (N_2215,N_1995,N_1948);
or U2216 (N_2216,N_1942,N_1967);
or U2217 (N_2217,N_1963,N_2068);
or U2218 (N_2218,N_1960,N_1956);
and U2219 (N_2219,N_1962,N_2025);
or U2220 (N_2220,N_1980,N_1928);
or U2221 (N_2221,N_1967,N_1977);
nor U2222 (N_2222,N_1956,N_2045);
and U2223 (N_2223,N_1960,N_1973);
xnor U2224 (N_2224,N_2042,N_1969);
nand U2225 (N_2225,N_2047,N_2061);
nor U2226 (N_2226,N_2056,N_2029);
nand U2227 (N_2227,N_2019,N_1988);
xnor U2228 (N_2228,N_2015,N_2041);
and U2229 (N_2229,N_1966,N_1938);
nand U2230 (N_2230,N_1968,N_1979);
nand U2231 (N_2231,N_1946,N_1940);
or U2232 (N_2232,N_2052,N_2076);
nor U2233 (N_2233,N_2071,N_1974);
xnor U2234 (N_2234,N_2041,N_2035);
nor U2235 (N_2235,N_1970,N_2002);
nor U2236 (N_2236,N_1962,N_1996);
nand U2237 (N_2237,N_1939,N_1950);
xnor U2238 (N_2238,N_2076,N_1990);
xor U2239 (N_2239,N_1960,N_1924);
or U2240 (N_2240,N_2198,N_2122);
xor U2241 (N_2241,N_2140,N_2084);
nand U2242 (N_2242,N_2116,N_2189);
and U2243 (N_2243,N_2109,N_2102);
xor U2244 (N_2244,N_2225,N_2186);
xnor U2245 (N_2245,N_2211,N_2143);
nor U2246 (N_2246,N_2185,N_2086);
and U2247 (N_2247,N_2098,N_2137);
and U2248 (N_2248,N_2081,N_2239);
xor U2249 (N_2249,N_2136,N_2206);
xnor U2250 (N_2250,N_2147,N_2133);
nor U2251 (N_2251,N_2144,N_2105);
or U2252 (N_2252,N_2181,N_2167);
and U2253 (N_2253,N_2123,N_2155);
nor U2254 (N_2254,N_2236,N_2171);
or U2255 (N_2255,N_2210,N_2127);
nand U2256 (N_2256,N_2183,N_2232);
and U2257 (N_2257,N_2209,N_2174);
xor U2258 (N_2258,N_2219,N_2104);
and U2259 (N_2259,N_2132,N_2100);
nand U2260 (N_2260,N_2165,N_2159);
nor U2261 (N_2261,N_2138,N_2180);
or U2262 (N_2262,N_2222,N_2148);
or U2263 (N_2263,N_2226,N_2141);
nand U2264 (N_2264,N_2094,N_2107);
xor U2265 (N_2265,N_2119,N_2182);
or U2266 (N_2266,N_2217,N_2135);
nor U2267 (N_2267,N_2233,N_2164);
nand U2268 (N_2268,N_2205,N_2082);
nand U2269 (N_2269,N_2090,N_2175);
nand U2270 (N_2270,N_2163,N_2190);
nor U2271 (N_2271,N_2128,N_2150);
nand U2272 (N_2272,N_2202,N_2207);
nor U2273 (N_2273,N_2224,N_2199);
nand U2274 (N_2274,N_2214,N_2237);
or U2275 (N_2275,N_2112,N_2231);
and U2276 (N_2276,N_2161,N_2216);
nor U2277 (N_2277,N_2125,N_2177);
nor U2278 (N_2278,N_2153,N_2166);
xnor U2279 (N_2279,N_2184,N_2091);
or U2280 (N_2280,N_2126,N_2194);
or U2281 (N_2281,N_2187,N_2218);
and U2282 (N_2282,N_2156,N_2117);
or U2283 (N_2283,N_2221,N_2162);
nor U2284 (N_2284,N_2213,N_2191);
xor U2285 (N_2285,N_2192,N_2201);
xor U2286 (N_2286,N_2193,N_2106);
xnor U2287 (N_2287,N_2121,N_2124);
or U2288 (N_2288,N_2089,N_2080);
or U2289 (N_2289,N_2134,N_2092);
or U2290 (N_2290,N_2230,N_2095);
nor U2291 (N_2291,N_2085,N_2170);
xor U2292 (N_2292,N_2168,N_2154);
nand U2293 (N_2293,N_2139,N_2160);
nor U2294 (N_2294,N_2173,N_2195);
nand U2295 (N_2295,N_2097,N_2130);
nand U2296 (N_2296,N_2197,N_2235);
and U2297 (N_2297,N_2227,N_2101);
xnor U2298 (N_2298,N_2113,N_2200);
xor U2299 (N_2299,N_2169,N_2203);
or U2300 (N_2300,N_2196,N_2103);
or U2301 (N_2301,N_2099,N_2151);
nor U2302 (N_2302,N_2176,N_2131);
xor U2303 (N_2303,N_2145,N_2146);
and U2304 (N_2304,N_2157,N_2087);
or U2305 (N_2305,N_2114,N_2118);
and U2306 (N_2306,N_2220,N_2204);
nor U2307 (N_2307,N_2188,N_2234);
nor U2308 (N_2308,N_2093,N_2152);
xor U2309 (N_2309,N_2228,N_2238);
or U2310 (N_2310,N_2120,N_2172);
or U2311 (N_2311,N_2088,N_2108);
nor U2312 (N_2312,N_2129,N_2142);
xor U2313 (N_2313,N_2149,N_2096);
xnor U2314 (N_2314,N_2223,N_2083);
nor U2315 (N_2315,N_2158,N_2208);
and U2316 (N_2316,N_2215,N_2179);
xnor U2317 (N_2317,N_2212,N_2111);
nand U2318 (N_2318,N_2229,N_2178);
or U2319 (N_2319,N_2115,N_2110);
and U2320 (N_2320,N_2086,N_2084);
and U2321 (N_2321,N_2148,N_2107);
and U2322 (N_2322,N_2231,N_2098);
nor U2323 (N_2323,N_2215,N_2204);
nand U2324 (N_2324,N_2147,N_2193);
xnor U2325 (N_2325,N_2157,N_2129);
or U2326 (N_2326,N_2143,N_2085);
or U2327 (N_2327,N_2141,N_2207);
xor U2328 (N_2328,N_2119,N_2199);
or U2329 (N_2329,N_2222,N_2154);
nor U2330 (N_2330,N_2101,N_2239);
and U2331 (N_2331,N_2220,N_2155);
or U2332 (N_2332,N_2170,N_2099);
nor U2333 (N_2333,N_2133,N_2212);
nand U2334 (N_2334,N_2225,N_2115);
or U2335 (N_2335,N_2236,N_2113);
nor U2336 (N_2336,N_2207,N_2218);
nor U2337 (N_2337,N_2180,N_2122);
xnor U2338 (N_2338,N_2100,N_2102);
xnor U2339 (N_2339,N_2125,N_2110);
or U2340 (N_2340,N_2226,N_2208);
xor U2341 (N_2341,N_2192,N_2145);
and U2342 (N_2342,N_2149,N_2113);
nand U2343 (N_2343,N_2112,N_2237);
or U2344 (N_2344,N_2221,N_2223);
or U2345 (N_2345,N_2126,N_2231);
nor U2346 (N_2346,N_2146,N_2150);
and U2347 (N_2347,N_2211,N_2123);
nand U2348 (N_2348,N_2207,N_2100);
and U2349 (N_2349,N_2226,N_2162);
nor U2350 (N_2350,N_2210,N_2082);
xnor U2351 (N_2351,N_2083,N_2222);
and U2352 (N_2352,N_2080,N_2159);
nand U2353 (N_2353,N_2087,N_2127);
and U2354 (N_2354,N_2232,N_2130);
and U2355 (N_2355,N_2232,N_2196);
nor U2356 (N_2356,N_2097,N_2225);
and U2357 (N_2357,N_2128,N_2236);
nand U2358 (N_2358,N_2207,N_2122);
nand U2359 (N_2359,N_2081,N_2180);
or U2360 (N_2360,N_2172,N_2087);
nand U2361 (N_2361,N_2140,N_2142);
xor U2362 (N_2362,N_2217,N_2232);
nor U2363 (N_2363,N_2225,N_2100);
nand U2364 (N_2364,N_2187,N_2113);
or U2365 (N_2365,N_2102,N_2224);
nand U2366 (N_2366,N_2088,N_2133);
and U2367 (N_2367,N_2111,N_2165);
or U2368 (N_2368,N_2169,N_2222);
xor U2369 (N_2369,N_2168,N_2175);
nor U2370 (N_2370,N_2087,N_2219);
or U2371 (N_2371,N_2179,N_2182);
and U2372 (N_2372,N_2236,N_2197);
nor U2373 (N_2373,N_2089,N_2152);
nor U2374 (N_2374,N_2165,N_2214);
nand U2375 (N_2375,N_2096,N_2136);
xor U2376 (N_2376,N_2166,N_2178);
or U2377 (N_2377,N_2080,N_2148);
xnor U2378 (N_2378,N_2167,N_2199);
xnor U2379 (N_2379,N_2176,N_2103);
and U2380 (N_2380,N_2188,N_2217);
and U2381 (N_2381,N_2199,N_2210);
or U2382 (N_2382,N_2116,N_2171);
nor U2383 (N_2383,N_2149,N_2214);
and U2384 (N_2384,N_2222,N_2239);
or U2385 (N_2385,N_2120,N_2173);
nand U2386 (N_2386,N_2176,N_2193);
or U2387 (N_2387,N_2139,N_2206);
xnor U2388 (N_2388,N_2100,N_2111);
nor U2389 (N_2389,N_2219,N_2209);
nor U2390 (N_2390,N_2226,N_2185);
xnor U2391 (N_2391,N_2098,N_2136);
or U2392 (N_2392,N_2134,N_2159);
nand U2393 (N_2393,N_2173,N_2204);
xor U2394 (N_2394,N_2189,N_2152);
nor U2395 (N_2395,N_2232,N_2233);
and U2396 (N_2396,N_2204,N_2196);
and U2397 (N_2397,N_2132,N_2164);
and U2398 (N_2398,N_2187,N_2177);
or U2399 (N_2399,N_2167,N_2154);
nor U2400 (N_2400,N_2261,N_2283);
and U2401 (N_2401,N_2343,N_2332);
nor U2402 (N_2402,N_2337,N_2340);
or U2403 (N_2403,N_2313,N_2255);
or U2404 (N_2404,N_2336,N_2399);
nor U2405 (N_2405,N_2366,N_2338);
and U2406 (N_2406,N_2325,N_2354);
or U2407 (N_2407,N_2330,N_2265);
or U2408 (N_2408,N_2248,N_2384);
and U2409 (N_2409,N_2281,N_2379);
nand U2410 (N_2410,N_2351,N_2364);
nor U2411 (N_2411,N_2381,N_2365);
and U2412 (N_2412,N_2382,N_2249);
nor U2413 (N_2413,N_2356,N_2246);
or U2414 (N_2414,N_2329,N_2275);
and U2415 (N_2415,N_2323,N_2298);
nor U2416 (N_2416,N_2314,N_2308);
or U2417 (N_2417,N_2335,N_2363);
nand U2418 (N_2418,N_2357,N_2374);
xor U2419 (N_2419,N_2282,N_2259);
xor U2420 (N_2420,N_2303,N_2274);
and U2421 (N_2421,N_2291,N_2254);
or U2422 (N_2422,N_2373,N_2258);
xor U2423 (N_2423,N_2344,N_2348);
nor U2424 (N_2424,N_2306,N_2369);
xnor U2425 (N_2425,N_2243,N_2304);
xnor U2426 (N_2426,N_2375,N_2268);
xnor U2427 (N_2427,N_2285,N_2267);
or U2428 (N_2428,N_2288,N_2321);
or U2429 (N_2429,N_2262,N_2392);
nor U2430 (N_2430,N_2253,N_2318);
or U2431 (N_2431,N_2279,N_2386);
and U2432 (N_2432,N_2264,N_2353);
or U2433 (N_2433,N_2331,N_2397);
nor U2434 (N_2434,N_2247,N_2250);
xor U2435 (N_2435,N_2266,N_2293);
and U2436 (N_2436,N_2311,N_2347);
nand U2437 (N_2437,N_2342,N_2297);
nand U2438 (N_2438,N_2257,N_2387);
or U2439 (N_2439,N_2320,N_2395);
xor U2440 (N_2440,N_2241,N_2371);
xnor U2441 (N_2441,N_2358,N_2292);
or U2442 (N_2442,N_2385,N_2276);
and U2443 (N_2443,N_2240,N_2339);
nand U2444 (N_2444,N_2345,N_2301);
nand U2445 (N_2445,N_2256,N_2355);
and U2446 (N_2446,N_2307,N_2360);
nand U2447 (N_2447,N_2300,N_2380);
and U2448 (N_2448,N_2287,N_2328);
nand U2449 (N_2449,N_2396,N_2327);
nand U2450 (N_2450,N_2389,N_2388);
xnor U2451 (N_2451,N_2309,N_2290);
xnor U2452 (N_2452,N_2263,N_2322);
and U2453 (N_2453,N_2361,N_2277);
and U2454 (N_2454,N_2296,N_2284);
nand U2455 (N_2455,N_2359,N_2350);
and U2456 (N_2456,N_2295,N_2333);
nand U2457 (N_2457,N_2251,N_2310);
and U2458 (N_2458,N_2390,N_2362);
nand U2459 (N_2459,N_2370,N_2305);
and U2460 (N_2460,N_2299,N_2245);
nand U2461 (N_2461,N_2289,N_2352);
and U2462 (N_2462,N_2242,N_2341);
nor U2463 (N_2463,N_2286,N_2317);
or U2464 (N_2464,N_2272,N_2324);
and U2465 (N_2465,N_2398,N_2315);
nand U2466 (N_2466,N_2394,N_2378);
or U2467 (N_2467,N_2312,N_2368);
or U2468 (N_2468,N_2319,N_2326);
nor U2469 (N_2469,N_2376,N_2391);
nand U2470 (N_2470,N_2294,N_2302);
or U2471 (N_2471,N_2260,N_2393);
or U2472 (N_2472,N_2244,N_2383);
nand U2473 (N_2473,N_2252,N_2269);
or U2474 (N_2474,N_2349,N_2278);
and U2475 (N_2475,N_2377,N_2270);
nor U2476 (N_2476,N_2334,N_2271);
nor U2477 (N_2477,N_2367,N_2280);
nor U2478 (N_2478,N_2372,N_2346);
xor U2479 (N_2479,N_2273,N_2316);
nor U2480 (N_2480,N_2271,N_2241);
or U2481 (N_2481,N_2367,N_2369);
nand U2482 (N_2482,N_2263,N_2333);
and U2483 (N_2483,N_2305,N_2294);
xor U2484 (N_2484,N_2338,N_2260);
nor U2485 (N_2485,N_2252,N_2317);
nand U2486 (N_2486,N_2335,N_2266);
or U2487 (N_2487,N_2301,N_2330);
or U2488 (N_2488,N_2288,N_2342);
nand U2489 (N_2489,N_2262,N_2378);
xnor U2490 (N_2490,N_2248,N_2253);
nand U2491 (N_2491,N_2370,N_2343);
nand U2492 (N_2492,N_2384,N_2265);
nand U2493 (N_2493,N_2305,N_2333);
nand U2494 (N_2494,N_2305,N_2241);
and U2495 (N_2495,N_2268,N_2371);
or U2496 (N_2496,N_2390,N_2294);
xnor U2497 (N_2497,N_2353,N_2317);
nand U2498 (N_2498,N_2271,N_2319);
and U2499 (N_2499,N_2304,N_2282);
xor U2500 (N_2500,N_2285,N_2244);
and U2501 (N_2501,N_2245,N_2268);
nor U2502 (N_2502,N_2316,N_2248);
nand U2503 (N_2503,N_2255,N_2382);
nor U2504 (N_2504,N_2392,N_2304);
or U2505 (N_2505,N_2306,N_2292);
or U2506 (N_2506,N_2328,N_2240);
nor U2507 (N_2507,N_2325,N_2355);
xor U2508 (N_2508,N_2383,N_2297);
nor U2509 (N_2509,N_2312,N_2247);
nand U2510 (N_2510,N_2266,N_2257);
xnor U2511 (N_2511,N_2276,N_2344);
xnor U2512 (N_2512,N_2302,N_2319);
xor U2513 (N_2513,N_2348,N_2304);
and U2514 (N_2514,N_2249,N_2384);
xnor U2515 (N_2515,N_2330,N_2324);
xor U2516 (N_2516,N_2297,N_2287);
or U2517 (N_2517,N_2286,N_2333);
and U2518 (N_2518,N_2281,N_2255);
nand U2519 (N_2519,N_2362,N_2307);
and U2520 (N_2520,N_2276,N_2289);
and U2521 (N_2521,N_2326,N_2332);
or U2522 (N_2522,N_2322,N_2241);
or U2523 (N_2523,N_2315,N_2332);
nor U2524 (N_2524,N_2381,N_2371);
nand U2525 (N_2525,N_2346,N_2378);
nor U2526 (N_2526,N_2271,N_2308);
nand U2527 (N_2527,N_2247,N_2273);
xnor U2528 (N_2528,N_2336,N_2388);
nor U2529 (N_2529,N_2384,N_2307);
nand U2530 (N_2530,N_2349,N_2246);
nor U2531 (N_2531,N_2310,N_2366);
nor U2532 (N_2532,N_2307,N_2306);
and U2533 (N_2533,N_2270,N_2337);
nor U2534 (N_2534,N_2354,N_2368);
nand U2535 (N_2535,N_2394,N_2253);
or U2536 (N_2536,N_2350,N_2384);
and U2537 (N_2537,N_2261,N_2290);
nand U2538 (N_2538,N_2326,N_2362);
nor U2539 (N_2539,N_2261,N_2293);
nor U2540 (N_2540,N_2253,N_2279);
or U2541 (N_2541,N_2392,N_2385);
nand U2542 (N_2542,N_2273,N_2266);
and U2543 (N_2543,N_2311,N_2315);
xor U2544 (N_2544,N_2259,N_2357);
nand U2545 (N_2545,N_2376,N_2313);
nor U2546 (N_2546,N_2304,N_2281);
nand U2547 (N_2547,N_2257,N_2370);
and U2548 (N_2548,N_2277,N_2374);
xnor U2549 (N_2549,N_2269,N_2264);
nor U2550 (N_2550,N_2299,N_2272);
nand U2551 (N_2551,N_2242,N_2356);
nor U2552 (N_2552,N_2300,N_2367);
and U2553 (N_2553,N_2355,N_2339);
nand U2554 (N_2554,N_2317,N_2287);
or U2555 (N_2555,N_2390,N_2287);
nand U2556 (N_2556,N_2354,N_2348);
xor U2557 (N_2557,N_2334,N_2260);
xor U2558 (N_2558,N_2269,N_2265);
xnor U2559 (N_2559,N_2308,N_2340);
xor U2560 (N_2560,N_2450,N_2541);
and U2561 (N_2561,N_2402,N_2547);
or U2562 (N_2562,N_2471,N_2473);
or U2563 (N_2563,N_2453,N_2407);
and U2564 (N_2564,N_2431,N_2486);
xnor U2565 (N_2565,N_2554,N_2558);
nand U2566 (N_2566,N_2434,N_2521);
or U2567 (N_2567,N_2439,N_2442);
nand U2568 (N_2568,N_2451,N_2514);
xnor U2569 (N_2569,N_2529,N_2504);
nor U2570 (N_2570,N_2538,N_2530);
and U2571 (N_2571,N_2446,N_2524);
and U2572 (N_2572,N_2411,N_2458);
nand U2573 (N_2573,N_2447,N_2444);
or U2574 (N_2574,N_2469,N_2443);
and U2575 (N_2575,N_2499,N_2415);
nor U2576 (N_2576,N_2548,N_2491);
and U2577 (N_2577,N_2476,N_2463);
xor U2578 (N_2578,N_2494,N_2408);
xnor U2579 (N_2579,N_2527,N_2557);
or U2580 (N_2580,N_2428,N_2474);
and U2581 (N_2581,N_2424,N_2401);
and U2582 (N_2582,N_2542,N_2472);
or U2583 (N_2583,N_2420,N_2533);
xnor U2584 (N_2584,N_2440,N_2412);
nor U2585 (N_2585,N_2449,N_2427);
or U2586 (N_2586,N_2510,N_2478);
or U2587 (N_2587,N_2556,N_2459);
xnor U2588 (N_2588,N_2438,N_2468);
nand U2589 (N_2589,N_2559,N_2500);
nor U2590 (N_2590,N_2534,N_2454);
nand U2591 (N_2591,N_2508,N_2421);
and U2592 (N_2592,N_2553,N_2543);
xor U2593 (N_2593,N_2516,N_2522);
xnor U2594 (N_2594,N_2502,N_2496);
nor U2595 (N_2595,N_2495,N_2461);
nand U2596 (N_2596,N_2416,N_2513);
nor U2597 (N_2597,N_2544,N_2436);
and U2598 (N_2598,N_2422,N_2519);
or U2599 (N_2599,N_2426,N_2456);
or U2600 (N_2600,N_2549,N_2413);
nor U2601 (N_2601,N_2492,N_2403);
xor U2602 (N_2602,N_2405,N_2525);
nand U2603 (N_2603,N_2505,N_2455);
nand U2604 (N_2604,N_2441,N_2515);
or U2605 (N_2605,N_2552,N_2539);
and U2606 (N_2606,N_2437,N_2483);
nor U2607 (N_2607,N_2400,N_2546);
or U2608 (N_2608,N_2445,N_2410);
and U2609 (N_2609,N_2462,N_2485);
nand U2610 (N_2610,N_2452,N_2520);
or U2611 (N_2611,N_2435,N_2404);
nor U2612 (N_2612,N_2503,N_2497);
xnor U2613 (N_2613,N_2512,N_2409);
nor U2614 (N_2614,N_2550,N_2406);
or U2615 (N_2615,N_2531,N_2423);
nand U2616 (N_2616,N_2506,N_2419);
and U2617 (N_2617,N_2532,N_2414);
xnor U2618 (N_2618,N_2457,N_2460);
nand U2619 (N_2619,N_2432,N_2535);
or U2620 (N_2620,N_2498,N_2448);
and U2621 (N_2621,N_2475,N_2466);
and U2622 (N_2622,N_2523,N_2488);
or U2623 (N_2623,N_2477,N_2490);
or U2624 (N_2624,N_2482,N_2417);
nand U2625 (N_2625,N_2507,N_2465);
and U2626 (N_2626,N_2481,N_2493);
or U2627 (N_2627,N_2425,N_2517);
nand U2628 (N_2628,N_2551,N_2540);
nor U2629 (N_2629,N_2537,N_2555);
and U2630 (N_2630,N_2487,N_2470);
or U2631 (N_2631,N_2418,N_2518);
or U2632 (N_2632,N_2480,N_2545);
and U2633 (N_2633,N_2511,N_2484);
xnor U2634 (N_2634,N_2526,N_2536);
xor U2635 (N_2635,N_2467,N_2528);
nor U2636 (N_2636,N_2429,N_2489);
nand U2637 (N_2637,N_2430,N_2501);
nand U2638 (N_2638,N_2464,N_2509);
or U2639 (N_2639,N_2433,N_2479);
and U2640 (N_2640,N_2458,N_2548);
nor U2641 (N_2641,N_2529,N_2462);
nor U2642 (N_2642,N_2552,N_2444);
or U2643 (N_2643,N_2534,N_2455);
and U2644 (N_2644,N_2493,N_2462);
nand U2645 (N_2645,N_2499,N_2432);
xor U2646 (N_2646,N_2553,N_2469);
xor U2647 (N_2647,N_2472,N_2405);
and U2648 (N_2648,N_2437,N_2403);
and U2649 (N_2649,N_2526,N_2416);
or U2650 (N_2650,N_2485,N_2435);
or U2651 (N_2651,N_2545,N_2488);
nor U2652 (N_2652,N_2534,N_2461);
nand U2653 (N_2653,N_2483,N_2548);
nand U2654 (N_2654,N_2558,N_2469);
xor U2655 (N_2655,N_2501,N_2545);
nand U2656 (N_2656,N_2416,N_2431);
xnor U2657 (N_2657,N_2456,N_2545);
and U2658 (N_2658,N_2429,N_2452);
nor U2659 (N_2659,N_2405,N_2420);
nor U2660 (N_2660,N_2554,N_2518);
and U2661 (N_2661,N_2539,N_2509);
nand U2662 (N_2662,N_2474,N_2496);
nor U2663 (N_2663,N_2453,N_2552);
nor U2664 (N_2664,N_2510,N_2533);
xnor U2665 (N_2665,N_2530,N_2500);
nor U2666 (N_2666,N_2486,N_2509);
nand U2667 (N_2667,N_2485,N_2530);
xor U2668 (N_2668,N_2496,N_2499);
xor U2669 (N_2669,N_2504,N_2406);
or U2670 (N_2670,N_2542,N_2424);
and U2671 (N_2671,N_2498,N_2526);
xnor U2672 (N_2672,N_2528,N_2479);
and U2673 (N_2673,N_2429,N_2528);
or U2674 (N_2674,N_2526,N_2463);
or U2675 (N_2675,N_2498,N_2461);
and U2676 (N_2676,N_2484,N_2431);
or U2677 (N_2677,N_2457,N_2511);
nor U2678 (N_2678,N_2444,N_2449);
nor U2679 (N_2679,N_2455,N_2530);
nor U2680 (N_2680,N_2462,N_2428);
nor U2681 (N_2681,N_2490,N_2426);
xnor U2682 (N_2682,N_2494,N_2446);
xor U2683 (N_2683,N_2453,N_2436);
nor U2684 (N_2684,N_2455,N_2432);
nor U2685 (N_2685,N_2424,N_2534);
nand U2686 (N_2686,N_2532,N_2519);
or U2687 (N_2687,N_2444,N_2471);
nand U2688 (N_2688,N_2550,N_2465);
and U2689 (N_2689,N_2541,N_2481);
xor U2690 (N_2690,N_2435,N_2440);
or U2691 (N_2691,N_2553,N_2421);
nor U2692 (N_2692,N_2548,N_2539);
and U2693 (N_2693,N_2499,N_2444);
or U2694 (N_2694,N_2503,N_2439);
nand U2695 (N_2695,N_2487,N_2559);
xor U2696 (N_2696,N_2489,N_2438);
and U2697 (N_2697,N_2485,N_2495);
or U2698 (N_2698,N_2493,N_2402);
or U2699 (N_2699,N_2497,N_2469);
or U2700 (N_2700,N_2483,N_2420);
or U2701 (N_2701,N_2495,N_2491);
and U2702 (N_2702,N_2520,N_2518);
nand U2703 (N_2703,N_2486,N_2502);
nor U2704 (N_2704,N_2452,N_2502);
xor U2705 (N_2705,N_2504,N_2494);
and U2706 (N_2706,N_2529,N_2505);
xnor U2707 (N_2707,N_2548,N_2446);
nor U2708 (N_2708,N_2422,N_2450);
nor U2709 (N_2709,N_2447,N_2479);
nand U2710 (N_2710,N_2483,N_2537);
or U2711 (N_2711,N_2448,N_2540);
nand U2712 (N_2712,N_2474,N_2470);
xnor U2713 (N_2713,N_2559,N_2408);
nor U2714 (N_2714,N_2544,N_2556);
nor U2715 (N_2715,N_2507,N_2532);
nand U2716 (N_2716,N_2434,N_2509);
xor U2717 (N_2717,N_2436,N_2400);
nor U2718 (N_2718,N_2439,N_2507);
nand U2719 (N_2719,N_2523,N_2408);
nand U2720 (N_2720,N_2686,N_2690);
nand U2721 (N_2721,N_2683,N_2673);
nor U2722 (N_2722,N_2696,N_2681);
nor U2723 (N_2723,N_2614,N_2568);
nor U2724 (N_2724,N_2573,N_2689);
and U2725 (N_2725,N_2648,N_2662);
or U2726 (N_2726,N_2678,N_2562);
nor U2727 (N_2727,N_2659,N_2709);
xnor U2728 (N_2728,N_2637,N_2591);
nor U2729 (N_2729,N_2569,N_2605);
or U2730 (N_2730,N_2666,N_2704);
xnor U2731 (N_2731,N_2688,N_2649);
and U2732 (N_2732,N_2589,N_2584);
and U2733 (N_2733,N_2616,N_2611);
or U2734 (N_2734,N_2622,N_2707);
and U2735 (N_2735,N_2585,N_2667);
and U2736 (N_2736,N_2596,N_2634);
and U2737 (N_2737,N_2620,N_2638);
and U2738 (N_2738,N_2685,N_2706);
nand U2739 (N_2739,N_2576,N_2699);
and U2740 (N_2740,N_2618,N_2711);
or U2741 (N_2741,N_2660,N_2714);
and U2742 (N_2742,N_2646,N_2564);
xor U2743 (N_2743,N_2587,N_2623);
nor U2744 (N_2744,N_2694,N_2679);
nor U2745 (N_2745,N_2599,N_2684);
nand U2746 (N_2746,N_2570,N_2644);
and U2747 (N_2747,N_2626,N_2639);
xor U2748 (N_2748,N_2652,N_2574);
xnor U2749 (N_2749,N_2687,N_2635);
xnor U2750 (N_2750,N_2661,N_2641);
nand U2751 (N_2751,N_2566,N_2705);
nand U2752 (N_2752,N_2600,N_2668);
nand U2753 (N_2753,N_2563,N_2653);
and U2754 (N_2754,N_2593,N_2636);
and U2755 (N_2755,N_2565,N_2633);
nor U2756 (N_2756,N_2663,N_2700);
and U2757 (N_2757,N_2671,N_2619);
nor U2758 (N_2758,N_2571,N_2680);
and U2759 (N_2759,N_2695,N_2627);
nand U2760 (N_2760,N_2655,N_2613);
or U2761 (N_2761,N_2604,N_2672);
nor U2762 (N_2762,N_2677,N_2590);
and U2763 (N_2763,N_2597,N_2598);
nand U2764 (N_2764,N_2628,N_2643);
or U2765 (N_2765,N_2609,N_2612);
and U2766 (N_2766,N_2601,N_2697);
nor U2767 (N_2767,N_2716,N_2703);
nor U2768 (N_2768,N_2698,N_2664);
and U2769 (N_2769,N_2581,N_2645);
xnor U2770 (N_2770,N_2674,N_2629);
and U2771 (N_2771,N_2650,N_2602);
or U2772 (N_2772,N_2670,N_2665);
or U2773 (N_2773,N_2594,N_2572);
and U2774 (N_2774,N_2608,N_2583);
nor U2775 (N_2775,N_2640,N_2647);
xnor U2776 (N_2776,N_2715,N_2610);
or U2777 (N_2777,N_2606,N_2607);
nor U2778 (N_2778,N_2682,N_2701);
nor U2779 (N_2779,N_2713,N_2708);
or U2780 (N_2780,N_2691,N_2718);
or U2781 (N_2781,N_2561,N_2632);
xnor U2782 (N_2782,N_2582,N_2669);
nor U2783 (N_2783,N_2656,N_2615);
nor U2784 (N_2784,N_2630,N_2575);
and U2785 (N_2785,N_2675,N_2658);
or U2786 (N_2786,N_2617,N_2651);
or U2787 (N_2787,N_2567,N_2624);
or U2788 (N_2788,N_2693,N_2631);
and U2789 (N_2789,N_2595,N_2692);
xnor U2790 (N_2790,N_2642,N_2719);
nor U2791 (N_2791,N_2603,N_2592);
nor U2792 (N_2792,N_2621,N_2654);
or U2793 (N_2793,N_2560,N_2588);
nand U2794 (N_2794,N_2579,N_2702);
xor U2795 (N_2795,N_2578,N_2586);
nand U2796 (N_2796,N_2717,N_2625);
nor U2797 (N_2797,N_2657,N_2676);
or U2798 (N_2798,N_2580,N_2712);
and U2799 (N_2799,N_2710,N_2577);
or U2800 (N_2800,N_2585,N_2659);
nor U2801 (N_2801,N_2623,N_2698);
xor U2802 (N_2802,N_2662,N_2602);
nor U2803 (N_2803,N_2672,N_2610);
and U2804 (N_2804,N_2666,N_2579);
nand U2805 (N_2805,N_2619,N_2604);
nand U2806 (N_2806,N_2614,N_2705);
nand U2807 (N_2807,N_2652,N_2713);
or U2808 (N_2808,N_2711,N_2676);
or U2809 (N_2809,N_2652,N_2616);
or U2810 (N_2810,N_2690,N_2590);
nor U2811 (N_2811,N_2594,N_2662);
and U2812 (N_2812,N_2618,N_2703);
and U2813 (N_2813,N_2641,N_2624);
nand U2814 (N_2814,N_2654,N_2573);
nand U2815 (N_2815,N_2654,N_2648);
and U2816 (N_2816,N_2690,N_2703);
or U2817 (N_2817,N_2643,N_2635);
and U2818 (N_2818,N_2618,N_2648);
or U2819 (N_2819,N_2568,N_2694);
nor U2820 (N_2820,N_2639,N_2670);
and U2821 (N_2821,N_2611,N_2641);
nor U2822 (N_2822,N_2624,N_2709);
and U2823 (N_2823,N_2649,N_2626);
nand U2824 (N_2824,N_2577,N_2617);
xor U2825 (N_2825,N_2613,N_2569);
nand U2826 (N_2826,N_2592,N_2585);
and U2827 (N_2827,N_2650,N_2627);
nor U2828 (N_2828,N_2627,N_2618);
and U2829 (N_2829,N_2607,N_2624);
nor U2830 (N_2830,N_2592,N_2608);
and U2831 (N_2831,N_2597,N_2574);
or U2832 (N_2832,N_2690,N_2580);
xor U2833 (N_2833,N_2640,N_2670);
xnor U2834 (N_2834,N_2662,N_2633);
xnor U2835 (N_2835,N_2678,N_2623);
or U2836 (N_2836,N_2708,N_2613);
and U2837 (N_2837,N_2642,N_2563);
nand U2838 (N_2838,N_2595,N_2654);
and U2839 (N_2839,N_2703,N_2568);
xor U2840 (N_2840,N_2680,N_2703);
nand U2841 (N_2841,N_2612,N_2611);
or U2842 (N_2842,N_2584,N_2594);
or U2843 (N_2843,N_2709,N_2655);
nor U2844 (N_2844,N_2572,N_2591);
nor U2845 (N_2845,N_2581,N_2597);
or U2846 (N_2846,N_2646,N_2707);
xnor U2847 (N_2847,N_2688,N_2718);
nor U2848 (N_2848,N_2675,N_2711);
nor U2849 (N_2849,N_2666,N_2625);
and U2850 (N_2850,N_2645,N_2601);
and U2851 (N_2851,N_2719,N_2701);
xor U2852 (N_2852,N_2646,N_2706);
nand U2853 (N_2853,N_2674,N_2581);
or U2854 (N_2854,N_2566,N_2702);
and U2855 (N_2855,N_2672,N_2680);
and U2856 (N_2856,N_2668,N_2630);
xnor U2857 (N_2857,N_2577,N_2637);
or U2858 (N_2858,N_2670,N_2646);
nand U2859 (N_2859,N_2672,N_2595);
nor U2860 (N_2860,N_2617,N_2565);
or U2861 (N_2861,N_2689,N_2639);
xnor U2862 (N_2862,N_2703,N_2714);
xnor U2863 (N_2863,N_2703,N_2702);
xnor U2864 (N_2864,N_2682,N_2581);
or U2865 (N_2865,N_2713,N_2705);
nor U2866 (N_2866,N_2637,N_2574);
xnor U2867 (N_2867,N_2592,N_2568);
nand U2868 (N_2868,N_2577,N_2588);
and U2869 (N_2869,N_2696,N_2597);
and U2870 (N_2870,N_2588,N_2631);
nand U2871 (N_2871,N_2608,N_2640);
or U2872 (N_2872,N_2609,N_2577);
or U2873 (N_2873,N_2585,N_2663);
nand U2874 (N_2874,N_2671,N_2711);
nand U2875 (N_2875,N_2681,N_2666);
or U2876 (N_2876,N_2715,N_2567);
nor U2877 (N_2877,N_2669,N_2683);
or U2878 (N_2878,N_2666,N_2608);
xor U2879 (N_2879,N_2701,N_2593);
nand U2880 (N_2880,N_2830,N_2814);
nor U2881 (N_2881,N_2865,N_2825);
or U2882 (N_2882,N_2745,N_2743);
xor U2883 (N_2883,N_2862,N_2760);
and U2884 (N_2884,N_2779,N_2818);
xor U2885 (N_2885,N_2799,N_2874);
or U2886 (N_2886,N_2741,N_2769);
and U2887 (N_2887,N_2785,N_2790);
or U2888 (N_2888,N_2746,N_2750);
xnor U2889 (N_2889,N_2756,N_2762);
or U2890 (N_2890,N_2798,N_2723);
or U2891 (N_2891,N_2774,N_2752);
and U2892 (N_2892,N_2801,N_2808);
and U2893 (N_2893,N_2813,N_2787);
nand U2894 (N_2894,N_2852,N_2740);
xor U2895 (N_2895,N_2731,N_2747);
nand U2896 (N_2896,N_2835,N_2796);
xnor U2897 (N_2897,N_2828,N_2758);
and U2898 (N_2898,N_2850,N_2856);
nand U2899 (N_2899,N_2800,N_2821);
nor U2900 (N_2900,N_2749,N_2786);
xnor U2901 (N_2901,N_2840,N_2775);
xnor U2902 (N_2902,N_2875,N_2791);
nor U2903 (N_2903,N_2795,N_2869);
and U2904 (N_2904,N_2807,N_2757);
nor U2905 (N_2905,N_2824,N_2725);
nor U2906 (N_2906,N_2811,N_2861);
xor U2907 (N_2907,N_2817,N_2763);
nand U2908 (N_2908,N_2794,N_2803);
and U2909 (N_2909,N_2772,N_2777);
nor U2910 (N_2910,N_2753,N_2768);
nand U2911 (N_2911,N_2735,N_2759);
nand U2912 (N_2912,N_2806,N_2739);
and U2913 (N_2913,N_2802,N_2726);
nor U2914 (N_2914,N_2871,N_2848);
nand U2915 (N_2915,N_2847,N_2822);
nand U2916 (N_2916,N_2858,N_2863);
xnor U2917 (N_2917,N_2866,N_2730);
nor U2918 (N_2918,N_2832,N_2810);
xor U2919 (N_2919,N_2827,N_2805);
and U2920 (N_2920,N_2771,N_2845);
nor U2921 (N_2921,N_2733,N_2837);
xor U2922 (N_2922,N_2857,N_2844);
nand U2923 (N_2923,N_2838,N_2833);
nor U2924 (N_2924,N_2784,N_2843);
nor U2925 (N_2925,N_2778,N_2776);
xnor U2926 (N_2926,N_2873,N_2721);
or U2927 (N_2927,N_2834,N_2789);
xnor U2928 (N_2928,N_2860,N_2732);
and U2929 (N_2929,N_2878,N_2734);
or U2930 (N_2930,N_2783,N_2727);
nand U2931 (N_2931,N_2754,N_2766);
and U2932 (N_2932,N_2842,N_2742);
xor U2933 (N_2933,N_2764,N_2851);
and U2934 (N_2934,N_2782,N_2836);
nand U2935 (N_2935,N_2815,N_2770);
and U2936 (N_2936,N_2767,N_2872);
xnor U2937 (N_2937,N_2781,N_2792);
xnor U2938 (N_2938,N_2839,N_2864);
nand U2939 (N_2939,N_2870,N_2720);
and U2940 (N_2940,N_2829,N_2823);
nand U2941 (N_2941,N_2736,N_2728);
or U2942 (N_2942,N_2868,N_2812);
or U2943 (N_2943,N_2737,N_2820);
or U2944 (N_2944,N_2816,N_2724);
nor U2945 (N_2945,N_2744,N_2867);
or U2946 (N_2946,N_2780,N_2722);
and U2947 (N_2947,N_2804,N_2855);
nor U2948 (N_2948,N_2793,N_2859);
xor U2949 (N_2949,N_2819,N_2761);
and U2950 (N_2950,N_2729,N_2841);
nor U2951 (N_2951,N_2788,N_2877);
or U2952 (N_2952,N_2773,N_2809);
or U2953 (N_2953,N_2876,N_2738);
nor U2954 (N_2954,N_2797,N_2846);
xnor U2955 (N_2955,N_2755,N_2879);
or U2956 (N_2956,N_2748,N_2831);
nor U2957 (N_2957,N_2849,N_2853);
and U2958 (N_2958,N_2765,N_2854);
nor U2959 (N_2959,N_2826,N_2751);
nand U2960 (N_2960,N_2853,N_2730);
or U2961 (N_2961,N_2838,N_2792);
xnor U2962 (N_2962,N_2768,N_2794);
and U2963 (N_2963,N_2789,N_2871);
or U2964 (N_2964,N_2786,N_2852);
xnor U2965 (N_2965,N_2878,N_2721);
and U2966 (N_2966,N_2865,N_2831);
and U2967 (N_2967,N_2818,N_2769);
nor U2968 (N_2968,N_2861,N_2828);
nand U2969 (N_2969,N_2851,N_2799);
nor U2970 (N_2970,N_2777,N_2786);
nor U2971 (N_2971,N_2744,N_2791);
and U2972 (N_2972,N_2730,N_2862);
nor U2973 (N_2973,N_2809,N_2799);
or U2974 (N_2974,N_2732,N_2783);
or U2975 (N_2975,N_2794,N_2770);
nand U2976 (N_2976,N_2752,N_2794);
nor U2977 (N_2977,N_2777,N_2720);
xnor U2978 (N_2978,N_2749,N_2797);
xnor U2979 (N_2979,N_2833,N_2770);
xor U2980 (N_2980,N_2865,N_2857);
xor U2981 (N_2981,N_2872,N_2789);
and U2982 (N_2982,N_2781,N_2755);
or U2983 (N_2983,N_2797,N_2814);
nor U2984 (N_2984,N_2797,N_2858);
or U2985 (N_2985,N_2776,N_2774);
nor U2986 (N_2986,N_2748,N_2735);
or U2987 (N_2987,N_2781,N_2826);
nand U2988 (N_2988,N_2731,N_2778);
and U2989 (N_2989,N_2756,N_2823);
nor U2990 (N_2990,N_2752,N_2754);
or U2991 (N_2991,N_2844,N_2835);
and U2992 (N_2992,N_2860,N_2743);
nand U2993 (N_2993,N_2743,N_2722);
and U2994 (N_2994,N_2825,N_2759);
nor U2995 (N_2995,N_2839,N_2757);
and U2996 (N_2996,N_2872,N_2841);
nand U2997 (N_2997,N_2855,N_2748);
nand U2998 (N_2998,N_2815,N_2733);
and U2999 (N_2999,N_2736,N_2795);
nand U3000 (N_3000,N_2777,N_2861);
and U3001 (N_3001,N_2787,N_2805);
and U3002 (N_3002,N_2788,N_2832);
and U3003 (N_3003,N_2753,N_2844);
nand U3004 (N_3004,N_2874,N_2831);
or U3005 (N_3005,N_2845,N_2859);
or U3006 (N_3006,N_2803,N_2753);
or U3007 (N_3007,N_2810,N_2875);
nand U3008 (N_3008,N_2741,N_2785);
xnor U3009 (N_3009,N_2819,N_2782);
nand U3010 (N_3010,N_2814,N_2808);
and U3011 (N_3011,N_2874,N_2817);
and U3012 (N_3012,N_2877,N_2727);
or U3013 (N_3013,N_2772,N_2824);
xnor U3014 (N_3014,N_2734,N_2732);
xor U3015 (N_3015,N_2782,N_2807);
xnor U3016 (N_3016,N_2720,N_2737);
or U3017 (N_3017,N_2758,N_2814);
or U3018 (N_3018,N_2854,N_2800);
xnor U3019 (N_3019,N_2776,N_2801);
or U3020 (N_3020,N_2832,N_2793);
nor U3021 (N_3021,N_2876,N_2762);
nor U3022 (N_3022,N_2852,N_2723);
nor U3023 (N_3023,N_2780,N_2865);
and U3024 (N_3024,N_2782,N_2777);
xnor U3025 (N_3025,N_2879,N_2822);
xor U3026 (N_3026,N_2789,N_2809);
or U3027 (N_3027,N_2865,N_2855);
xnor U3028 (N_3028,N_2822,N_2726);
or U3029 (N_3029,N_2820,N_2865);
nor U3030 (N_3030,N_2789,N_2870);
and U3031 (N_3031,N_2823,N_2773);
xor U3032 (N_3032,N_2873,N_2769);
nand U3033 (N_3033,N_2745,N_2728);
nand U3034 (N_3034,N_2758,N_2845);
nand U3035 (N_3035,N_2822,N_2805);
nand U3036 (N_3036,N_2749,N_2839);
xor U3037 (N_3037,N_2728,N_2840);
xor U3038 (N_3038,N_2757,N_2833);
nor U3039 (N_3039,N_2823,N_2759);
nor U3040 (N_3040,N_2937,N_2924);
or U3041 (N_3041,N_2986,N_2992);
and U3042 (N_3042,N_2906,N_2916);
nor U3043 (N_3043,N_2907,N_2985);
and U3044 (N_3044,N_2982,N_2917);
nand U3045 (N_3045,N_3007,N_3034);
and U3046 (N_3046,N_3006,N_2911);
nor U3047 (N_3047,N_2957,N_3029);
or U3048 (N_3048,N_2961,N_3013);
nand U3049 (N_3049,N_2970,N_2981);
and U3050 (N_3050,N_3010,N_2974);
nand U3051 (N_3051,N_2882,N_2969);
nor U3052 (N_3052,N_2884,N_2929);
or U3053 (N_3053,N_2909,N_2895);
xnor U3054 (N_3054,N_3032,N_3022);
nand U3055 (N_3055,N_2944,N_2931);
nand U3056 (N_3056,N_2989,N_2902);
and U3057 (N_3057,N_2993,N_3026);
xor U3058 (N_3058,N_2978,N_2891);
nand U3059 (N_3059,N_3025,N_2959);
nand U3060 (N_3060,N_2976,N_2960);
xor U3061 (N_3061,N_3015,N_2933);
xnor U3062 (N_3062,N_2942,N_3036);
or U3063 (N_3063,N_2893,N_2897);
nand U3064 (N_3064,N_2980,N_2964);
xnor U3065 (N_3065,N_2997,N_2988);
xor U3066 (N_3066,N_2887,N_2925);
nand U3067 (N_3067,N_2936,N_2896);
xor U3068 (N_3068,N_2881,N_2910);
and U3069 (N_3069,N_3002,N_2935);
nand U3070 (N_3070,N_2927,N_2938);
nor U3071 (N_3071,N_2901,N_2940);
nand U3072 (N_3072,N_3005,N_2955);
xnor U3073 (N_3073,N_3018,N_3028);
nor U3074 (N_3074,N_3016,N_2903);
and U3075 (N_3075,N_2979,N_3027);
xor U3076 (N_3076,N_3000,N_2920);
nor U3077 (N_3077,N_2971,N_2922);
xnor U3078 (N_3078,N_2888,N_2990);
and U3079 (N_3079,N_2965,N_2880);
or U3080 (N_3080,N_2983,N_2967);
and U3081 (N_3081,N_2943,N_2899);
xnor U3082 (N_3082,N_2975,N_3037);
or U3083 (N_3083,N_2928,N_2894);
or U3084 (N_3084,N_2908,N_2890);
xor U3085 (N_3085,N_2954,N_2995);
nand U3086 (N_3086,N_2972,N_3004);
and U3087 (N_3087,N_2921,N_2958);
and U3088 (N_3088,N_2926,N_2956);
and U3089 (N_3089,N_3003,N_2951);
xor U3090 (N_3090,N_2952,N_2945);
nor U3091 (N_3091,N_2968,N_2950);
xnor U3092 (N_3092,N_2991,N_2977);
and U3093 (N_3093,N_2930,N_2905);
nor U3094 (N_3094,N_2947,N_2889);
xnor U3095 (N_3095,N_3001,N_3012);
xnor U3096 (N_3096,N_2996,N_2913);
and U3097 (N_3097,N_2934,N_2998);
nor U3098 (N_3098,N_2885,N_2923);
or U3099 (N_3099,N_2994,N_3017);
and U3100 (N_3100,N_3030,N_2999);
and U3101 (N_3101,N_2963,N_2984);
or U3102 (N_3102,N_3035,N_2914);
and U3103 (N_3103,N_3014,N_2948);
and U3104 (N_3104,N_2915,N_3024);
and U3105 (N_3105,N_3021,N_3019);
or U3106 (N_3106,N_2892,N_3023);
nor U3107 (N_3107,N_2886,N_3033);
nand U3108 (N_3108,N_3031,N_2900);
nor U3109 (N_3109,N_2941,N_2966);
nor U3110 (N_3110,N_2949,N_2932);
xor U3111 (N_3111,N_2904,N_2953);
or U3112 (N_3112,N_2919,N_3039);
or U3113 (N_3113,N_2898,N_2973);
nor U3114 (N_3114,N_3009,N_2987);
or U3115 (N_3115,N_2939,N_2883);
xor U3116 (N_3116,N_3038,N_3020);
or U3117 (N_3117,N_2918,N_2962);
nand U3118 (N_3118,N_3011,N_2946);
xnor U3119 (N_3119,N_3008,N_2912);
nor U3120 (N_3120,N_2987,N_2929);
nand U3121 (N_3121,N_2900,N_2968);
and U3122 (N_3122,N_2918,N_2968);
and U3123 (N_3123,N_2956,N_2999);
nor U3124 (N_3124,N_2990,N_2906);
xor U3125 (N_3125,N_2901,N_2992);
xor U3126 (N_3126,N_2906,N_2936);
or U3127 (N_3127,N_2927,N_2926);
or U3128 (N_3128,N_2882,N_2919);
xnor U3129 (N_3129,N_2968,N_3003);
or U3130 (N_3130,N_2904,N_3030);
nand U3131 (N_3131,N_2880,N_2901);
or U3132 (N_3132,N_3037,N_2963);
nand U3133 (N_3133,N_2969,N_2952);
nand U3134 (N_3134,N_2882,N_2982);
xor U3135 (N_3135,N_3006,N_2921);
or U3136 (N_3136,N_2941,N_2891);
or U3137 (N_3137,N_2919,N_3028);
and U3138 (N_3138,N_3004,N_3021);
and U3139 (N_3139,N_2921,N_2927);
xor U3140 (N_3140,N_2903,N_2990);
nand U3141 (N_3141,N_2904,N_2888);
and U3142 (N_3142,N_3021,N_2889);
or U3143 (N_3143,N_2939,N_2929);
xnor U3144 (N_3144,N_2987,N_2953);
nand U3145 (N_3145,N_2942,N_2881);
xnor U3146 (N_3146,N_2963,N_2988);
or U3147 (N_3147,N_3014,N_3030);
nand U3148 (N_3148,N_2910,N_2996);
and U3149 (N_3149,N_2880,N_2975);
xor U3150 (N_3150,N_2906,N_2953);
nand U3151 (N_3151,N_3031,N_2908);
nor U3152 (N_3152,N_2921,N_2891);
xnor U3153 (N_3153,N_2932,N_2953);
nor U3154 (N_3154,N_2892,N_2943);
nor U3155 (N_3155,N_3015,N_3029);
or U3156 (N_3156,N_3005,N_2967);
nand U3157 (N_3157,N_2880,N_2946);
xor U3158 (N_3158,N_2917,N_3034);
or U3159 (N_3159,N_2902,N_2892);
nor U3160 (N_3160,N_3022,N_2966);
nor U3161 (N_3161,N_2956,N_3035);
and U3162 (N_3162,N_3037,N_2940);
nor U3163 (N_3163,N_2942,N_2993);
and U3164 (N_3164,N_2886,N_2980);
nor U3165 (N_3165,N_2909,N_3036);
and U3166 (N_3166,N_3006,N_2900);
nand U3167 (N_3167,N_2935,N_3006);
xor U3168 (N_3168,N_2906,N_3009);
nand U3169 (N_3169,N_2924,N_2946);
or U3170 (N_3170,N_3030,N_2997);
or U3171 (N_3171,N_3014,N_3010);
and U3172 (N_3172,N_2935,N_2981);
xnor U3173 (N_3173,N_2955,N_2884);
nand U3174 (N_3174,N_3026,N_2998);
or U3175 (N_3175,N_2908,N_2949);
nand U3176 (N_3176,N_2963,N_2995);
nor U3177 (N_3177,N_2963,N_2896);
nor U3178 (N_3178,N_2928,N_2986);
nand U3179 (N_3179,N_3026,N_2984);
nand U3180 (N_3180,N_2953,N_2897);
or U3181 (N_3181,N_3001,N_3022);
or U3182 (N_3182,N_2969,N_2922);
nor U3183 (N_3183,N_2981,N_2923);
or U3184 (N_3184,N_3018,N_3023);
nor U3185 (N_3185,N_3035,N_2911);
nand U3186 (N_3186,N_3039,N_3028);
or U3187 (N_3187,N_3008,N_2956);
and U3188 (N_3188,N_2954,N_2941);
or U3189 (N_3189,N_2940,N_3006);
nor U3190 (N_3190,N_2964,N_3019);
and U3191 (N_3191,N_2922,N_2895);
nand U3192 (N_3192,N_2984,N_2955);
nand U3193 (N_3193,N_2897,N_2998);
or U3194 (N_3194,N_3039,N_3021);
or U3195 (N_3195,N_2955,N_3011);
or U3196 (N_3196,N_2964,N_2988);
or U3197 (N_3197,N_3034,N_2971);
and U3198 (N_3198,N_2903,N_3033);
nand U3199 (N_3199,N_2917,N_2990);
or U3200 (N_3200,N_3180,N_3056);
nor U3201 (N_3201,N_3081,N_3112);
and U3202 (N_3202,N_3074,N_3143);
xor U3203 (N_3203,N_3150,N_3170);
and U3204 (N_3204,N_3192,N_3189);
or U3205 (N_3205,N_3120,N_3127);
xnor U3206 (N_3206,N_3132,N_3063);
xnor U3207 (N_3207,N_3092,N_3146);
nand U3208 (N_3208,N_3142,N_3116);
and U3209 (N_3209,N_3085,N_3161);
or U3210 (N_3210,N_3131,N_3094);
or U3211 (N_3211,N_3055,N_3100);
xnor U3212 (N_3212,N_3171,N_3096);
and U3213 (N_3213,N_3086,N_3190);
or U3214 (N_3214,N_3174,N_3137);
and U3215 (N_3215,N_3159,N_3105);
xor U3216 (N_3216,N_3156,N_3070);
xnor U3217 (N_3217,N_3153,N_3110);
and U3218 (N_3218,N_3123,N_3117);
and U3219 (N_3219,N_3182,N_3148);
or U3220 (N_3220,N_3169,N_3175);
or U3221 (N_3221,N_3128,N_3193);
xor U3222 (N_3222,N_3125,N_3065);
xor U3223 (N_3223,N_3139,N_3178);
and U3224 (N_3224,N_3099,N_3091);
nand U3225 (N_3225,N_3163,N_3162);
nand U3226 (N_3226,N_3060,N_3167);
nor U3227 (N_3227,N_3145,N_3053);
xnor U3228 (N_3228,N_3149,N_3165);
nand U3229 (N_3229,N_3047,N_3090);
and U3230 (N_3230,N_3183,N_3118);
nor U3231 (N_3231,N_3124,N_3064);
xor U3232 (N_3232,N_3135,N_3134);
or U3233 (N_3233,N_3059,N_3164);
or U3234 (N_3234,N_3046,N_3122);
nor U3235 (N_3235,N_3185,N_3166);
or U3236 (N_3236,N_3154,N_3084);
and U3237 (N_3237,N_3126,N_3066);
or U3238 (N_3238,N_3089,N_3101);
nand U3239 (N_3239,N_3079,N_3103);
or U3240 (N_3240,N_3196,N_3058);
and U3241 (N_3241,N_3144,N_3195);
and U3242 (N_3242,N_3088,N_3114);
nor U3243 (N_3243,N_3051,N_3129);
xor U3244 (N_3244,N_3057,N_3157);
xnor U3245 (N_3245,N_3152,N_3198);
nand U3246 (N_3246,N_3173,N_3177);
nand U3247 (N_3247,N_3176,N_3199);
or U3248 (N_3248,N_3188,N_3141);
xor U3249 (N_3249,N_3158,N_3111);
and U3250 (N_3250,N_3187,N_3045);
nor U3251 (N_3251,N_3044,N_3049);
or U3252 (N_3252,N_3077,N_3184);
or U3253 (N_3253,N_3071,N_3078);
and U3254 (N_3254,N_3107,N_3042);
or U3255 (N_3255,N_3043,N_3073);
or U3256 (N_3256,N_3113,N_3061);
xor U3257 (N_3257,N_3041,N_3069);
nor U3258 (N_3258,N_3121,N_3062);
or U3259 (N_3259,N_3181,N_3080);
nor U3260 (N_3260,N_3095,N_3104);
nand U3261 (N_3261,N_3130,N_3197);
or U3262 (N_3262,N_3179,N_3172);
xor U3263 (N_3263,N_3054,N_3082);
nand U3264 (N_3264,N_3106,N_3140);
nand U3265 (N_3265,N_3068,N_3133);
nor U3266 (N_3266,N_3075,N_3147);
nand U3267 (N_3267,N_3098,N_3050);
nand U3268 (N_3268,N_3155,N_3115);
xor U3269 (N_3269,N_3108,N_3067);
nor U3270 (N_3270,N_3119,N_3072);
xnor U3271 (N_3271,N_3151,N_3040);
nor U3272 (N_3272,N_3093,N_3186);
xor U3273 (N_3273,N_3138,N_3097);
xnor U3274 (N_3274,N_3102,N_3136);
and U3275 (N_3275,N_3052,N_3048);
and U3276 (N_3276,N_3083,N_3076);
nor U3277 (N_3277,N_3168,N_3191);
and U3278 (N_3278,N_3194,N_3087);
and U3279 (N_3279,N_3109,N_3160);
nor U3280 (N_3280,N_3142,N_3175);
or U3281 (N_3281,N_3094,N_3141);
nor U3282 (N_3282,N_3167,N_3116);
xor U3283 (N_3283,N_3058,N_3193);
xor U3284 (N_3284,N_3150,N_3098);
nand U3285 (N_3285,N_3086,N_3169);
or U3286 (N_3286,N_3161,N_3133);
nor U3287 (N_3287,N_3081,N_3095);
xor U3288 (N_3288,N_3088,N_3080);
and U3289 (N_3289,N_3108,N_3154);
nand U3290 (N_3290,N_3085,N_3050);
xnor U3291 (N_3291,N_3156,N_3068);
and U3292 (N_3292,N_3090,N_3155);
nor U3293 (N_3293,N_3179,N_3150);
nand U3294 (N_3294,N_3145,N_3131);
nand U3295 (N_3295,N_3134,N_3068);
nor U3296 (N_3296,N_3042,N_3044);
or U3297 (N_3297,N_3145,N_3147);
and U3298 (N_3298,N_3167,N_3111);
nor U3299 (N_3299,N_3120,N_3052);
and U3300 (N_3300,N_3091,N_3104);
nor U3301 (N_3301,N_3132,N_3184);
and U3302 (N_3302,N_3197,N_3092);
or U3303 (N_3303,N_3104,N_3111);
nand U3304 (N_3304,N_3097,N_3114);
or U3305 (N_3305,N_3120,N_3093);
or U3306 (N_3306,N_3078,N_3062);
nand U3307 (N_3307,N_3095,N_3194);
nand U3308 (N_3308,N_3182,N_3187);
nand U3309 (N_3309,N_3077,N_3110);
nand U3310 (N_3310,N_3048,N_3132);
nand U3311 (N_3311,N_3096,N_3054);
and U3312 (N_3312,N_3144,N_3103);
xor U3313 (N_3313,N_3192,N_3046);
xnor U3314 (N_3314,N_3125,N_3101);
and U3315 (N_3315,N_3162,N_3121);
xor U3316 (N_3316,N_3176,N_3146);
nand U3317 (N_3317,N_3057,N_3137);
or U3318 (N_3318,N_3182,N_3057);
or U3319 (N_3319,N_3188,N_3171);
or U3320 (N_3320,N_3194,N_3065);
nor U3321 (N_3321,N_3067,N_3153);
or U3322 (N_3322,N_3186,N_3196);
and U3323 (N_3323,N_3122,N_3102);
nand U3324 (N_3324,N_3064,N_3135);
nor U3325 (N_3325,N_3109,N_3166);
or U3326 (N_3326,N_3149,N_3198);
xor U3327 (N_3327,N_3188,N_3156);
xor U3328 (N_3328,N_3048,N_3044);
and U3329 (N_3329,N_3160,N_3059);
xor U3330 (N_3330,N_3090,N_3183);
and U3331 (N_3331,N_3139,N_3172);
or U3332 (N_3332,N_3103,N_3114);
nor U3333 (N_3333,N_3084,N_3129);
and U3334 (N_3334,N_3149,N_3174);
nor U3335 (N_3335,N_3067,N_3096);
or U3336 (N_3336,N_3125,N_3072);
and U3337 (N_3337,N_3164,N_3136);
nor U3338 (N_3338,N_3171,N_3095);
nand U3339 (N_3339,N_3194,N_3088);
or U3340 (N_3340,N_3122,N_3172);
xnor U3341 (N_3341,N_3042,N_3062);
nor U3342 (N_3342,N_3197,N_3132);
nand U3343 (N_3343,N_3153,N_3122);
xnor U3344 (N_3344,N_3198,N_3133);
and U3345 (N_3345,N_3097,N_3127);
nand U3346 (N_3346,N_3126,N_3087);
nand U3347 (N_3347,N_3157,N_3167);
nand U3348 (N_3348,N_3152,N_3168);
nor U3349 (N_3349,N_3119,N_3096);
or U3350 (N_3350,N_3115,N_3088);
or U3351 (N_3351,N_3123,N_3064);
xnor U3352 (N_3352,N_3159,N_3075);
nor U3353 (N_3353,N_3181,N_3051);
nand U3354 (N_3354,N_3124,N_3137);
and U3355 (N_3355,N_3173,N_3199);
nand U3356 (N_3356,N_3171,N_3144);
and U3357 (N_3357,N_3187,N_3122);
nand U3358 (N_3358,N_3196,N_3136);
xnor U3359 (N_3359,N_3085,N_3131);
xnor U3360 (N_3360,N_3274,N_3264);
or U3361 (N_3361,N_3344,N_3216);
xor U3362 (N_3362,N_3279,N_3266);
or U3363 (N_3363,N_3288,N_3290);
xor U3364 (N_3364,N_3254,N_3356);
xor U3365 (N_3365,N_3257,N_3323);
or U3366 (N_3366,N_3305,N_3289);
nor U3367 (N_3367,N_3241,N_3222);
or U3368 (N_3368,N_3238,N_3276);
nor U3369 (N_3369,N_3286,N_3228);
nor U3370 (N_3370,N_3233,N_3340);
or U3371 (N_3371,N_3236,N_3255);
and U3372 (N_3372,N_3339,N_3333);
nand U3373 (N_3373,N_3329,N_3327);
xnor U3374 (N_3374,N_3309,N_3250);
or U3375 (N_3375,N_3318,N_3297);
or U3376 (N_3376,N_3225,N_3253);
nand U3377 (N_3377,N_3211,N_3310);
or U3378 (N_3378,N_3212,N_3335);
and U3379 (N_3379,N_3240,N_3322);
xor U3380 (N_3380,N_3204,N_3226);
and U3381 (N_3381,N_3292,N_3353);
or U3382 (N_3382,N_3312,N_3351);
nor U3383 (N_3383,N_3301,N_3205);
xor U3384 (N_3384,N_3298,N_3268);
nand U3385 (N_3385,N_3251,N_3300);
nand U3386 (N_3386,N_3302,N_3352);
and U3387 (N_3387,N_3252,N_3337);
xor U3388 (N_3388,N_3330,N_3317);
and U3389 (N_3389,N_3345,N_3206);
or U3390 (N_3390,N_3332,N_3359);
nor U3391 (N_3391,N_3324,N_3307);
or U3392 (N_3392,N_3336,N_3275);
nand U3393 (N_3393,N_3350,N_3315);
nand U3394 (N_3394,N_3278,N_3280);
or U3395 (N_3395,N_3210,N_3334);
nor U3396 (N_3396,N_3273,N_3218);
nand U3397 (N_3397,N_3270,N_3220);
nand U3398 (N_3398,N_3328,N_3263);
nor U3399 (N_3399,N_3295,N_3316);
nand U3400 (N_3400,N_3311,N_3281);
nor U3401 (N_3401,N_3314,N_3239);
or U3402 (N_3402,N_3200,N_3213);
xor U3403 (N_3403,N_3320,N_3261);
nand U3404 (N_3404,N_3247,N_3357);
and U3405 (N_3405,N_3231,N_3269);
or U3406 (N_3406,N_3230,N_3223);
nand U3407 (N_3407,N_3272,N_3342);
nor U3408 (N_3408,N_3293,N_3237);
nand U3409 (N_3409,N_3294,N_3326);
xor U3410 (N_3410,N_3265,N_3347);
or U3411 (N_3411,N_3209,N_3341);
and U3412 (N_3412,N_3343,N_3271);
and U3413 (N_3413,N_3277,N_3313);
and U3414 (N_3414,N_3321,N_3202);
nor U3415 (N_3415,N_3207,N_3215);
nand U3416 (N_3416,N_3214,N_3259);
nor U3417 (N_3417,N_3245,N_3304);
xor U3418 (N_3418,N_3258,N_3287);
nor U3419 (N_3419,N_3244,N_3355);
and U3420 (N_3420,N_3296,N_3303);
and U3421 (N_3421,N_3346,N_3354);
or U3422 (N_3422,N_3234,N_3284);
or U3423 (N_3423,N_3282,N_3267);
and U3424 (N_3424,N_3256,N_3217);
or U3425 (N_3425,N_3201,N_3348);
and U3426 (N_3426,N_3285,N_3358);
xnor U3427 (N_3427,N_3227,N_3325);
or U3428 (N_3428,N_3248,N_3338);
or U3429 (N_3429,N_3221,N_3306);
or U3430 (N_3430,N_3331,N_3262);
and U3431 (N_3431,N_3319,N_3291);
xor U3432 (N_3432,N_3249,N_3299);
xnor U3433 (N_3433,N_3229,N_3283);
nor U3434 (N_3434,N_3246,N_3208);
and U3435 (N_3435,N_3219,N_3242);
or U3436 (N_3436,N_3243,N_3260);
and U3437 (N_3437,N_3232,N_3224);
nor U3438 (N_3438,N_3235,N_3349);
or U3439 (N_3439,N_3308,N_3203);
or U3440 (N_3440,N_3232,N_3282);
nor U3441 (N_3441,N_3295,N_3290);
xor U3442 (N_3442,N_3342,N_3310);
xnor U3443 (N_3443,N_3239,N_3201);
xnor U3444 (N_3444,N_3260,N_3209);
or U3445 (N_3445,N_3248,N_3267);
or U3446 (N_3446,N_3211,N_3292);
or U3447 (N_3447,N_3213,N_3226);
nand U3448 (N_3448,N_3336,N_3224);
or U3449 (N_3449,N_3346,N_3253);
or U3450 (N_3450,N_3261,N_3359);
xnor U3451 (N_3451,N_3265,N_3276);
xnor U3452 (N_3452,N_3334,N_3289);
and U3453 (N_3453,N_3264,N_3263);
or U3454 (N_3454,N_3319,N_3354);
and U3455 (N_3455,N_3240,N_3213);
nand U3456 (N_3456,N_3261,N_3293);
nor U3457 (N_3457,N_3268,N_3314);
xor U3458 (N_3458,N_3329,N_3322);
and U3459 (N_3459,N_3246,N_3206);
or U3460 (N_3460,N_3313,N_3340);
nor U3461 (N_3461,N_3346,N_3310);
xnor U3462 (N_3462,N_3356,N_3292);
nand U3463 (N_3463,N_3336,N_3318);
or U3464 (N_3464,N_3204,N_3301);
nor U3465 (N_3465,N_3296,N_3339);
or U3466 (N_3466,N_3268,N_3245);
nand U3467 (N_3467,N_3236,N_3215);
nor U3468 (N_3468,N_3237,N_3243);
nand U3469 (N_3469,N_3310,N_3358);
nor U3470 (N_3470,N_3236,N_3321);
nand U3471 (N_3471,N_3217,N_3214);
nand U3472 (N_3472,N_3306,N_3340);
and U3473 (N_3473,N_3225,N_3287);
or U3474 (N_3474,N_3340,N_3274);
and U3475 (N_3475,N_3268,N_3278);
or U3476 (N_3476,N_3251,N_3321);
nand U3477 (N_3477,N_3233,N_3244);
nand U3478 (N_3478,N_3315,N_3202);
or U3479 (N_3479,N_3322,N_3313);
nand U3480 (N_3480,N_3258,N_3230);
and U3481 (N_3481,N_3267,N_3230);
or U3482 (N_3482,N_3295,N_3274);
nand U3483 (N_3483,N_3307,N_3332);
xor U3484 (N_3484,N_3262,N_3247);
nor U3485 (N_3485,N_3230,N_3242);
nor U3486 (N_3486,N_3346,N_3270);
nor U3487 (N_3487,N_3232,N_3264);
nor U3488 (N_3488,N_3200,N_3245);
and U3489 (N_3489,N_3279,N_3336);
nand U3490 (N_3490,N_3324,N_3343);
nor U3491 (N_3491,N_3235,N_3211);
nand U3492 (N_3492,N_3353,N_3297);
and U3493 (N_3493,N_3334,N_3301);
or U3494 (N_3494,N_3243,N_3235);
nor U3495 (N_3495,N_3236,N_3306);
xnor U3496 (N_3496,N_3290,N_3226);
and U3497 (N_3497,N_3321,N_3338);
and U3498 (N_3498,N_3239,N_3209);
nand U3499 (N_3499,N_3349,N_3359);
or U3500 (N_3500,N_3213,N_3277);
nand U3501 (N_3501,N_3213,N_3353);
xor U3502 (N_3502,N_3269,N_3346);
xnor U3503 (N_3503,N_3259,N_3249);
and U3504 (N_3504,N_3328,N_3226);
nand U3505 (N_3505,N_3331,N_3200);
nand U3506 (N_3506,N_3214,N_3289);
xnor U3507 (N_3507,N_3204,N_3294);
and U3508 (N_3508,N_3269,N_3336);
nor U3509 (N_3509,N_3359,N_3348);
and U3510 (N_3510,N_3256,N_3282);
nand U3511 (N_3511,N_3241,N_3323);
nor U3512 (N_3512,N_3336,N_3316);
nand U3513 (N_3513,N_3321,N_3359);
xnor U3514 (N_3514,N_3318,N_3356);
nand U3515 (N_3515,N_3206,N_3330);
xnor U3516 (N_3516,N_3210,N_3254);
or U3517 (N_3517,N_3308,N_3333);
nand U3518 (N_3518,N_3335,N_3253);
xor U3519 (N_3519,N_3283,N_3264);
nor U3520 (N_3520,N_3437,N_3457);
and U3521 (N_3521,N_3503,N_3409);
nand U3522 (N_3522,N_3417,N_3464);
nor U3523 (N_3523,N_3515,N_3364);
and U3524 (N_3524,N_3443,N_3453);
or U3525 (N_3525,N_3402,N_3423);
nand U3526 (N_3526,N_3381,N_3411);
xor U3527 (N_3527,N_3518,N_3498);
nor U3528 (N_3528,N_3444,N_3425);
xnor U3529 (N_3529,N_3413,N_3490);
nand U3530 (N_3530,N_3394,N_3400);
or U3531 (N_3531,N_3482,N_3382);
nand U3532 (N_3532,N_3408,N_3493);
and U3533 (N_3533,N_3511,N_3412);
xor U3534 (N_3534,N_3448,N_3474);
and U3535 (N_3535,N_3508,N_3505);
and U3536 (N_3536,N_3513,N_3407);
nor U3537 (N_3537,N_3377,N_3432);
and U3538 (N_3538,N_3429,N_3371);
xor U3539 (N_3539,N_3439,N_3370);
or U3540 (N_3540,N_3486,N_3395);
and U3541 (N_3541,N_3450,N_3468);
or U3542 (N_3542,N_3398,N_3435);
and U3543 (N_3543,N_3452,N_3436);
nand U3544 (N_3544,N_3475,N_3496);
nand U3545 (N_3545,N_3424,N_3454);
nor U3546 (N_3546,N_3441,N_3451);
xor U3547 (N_3547,N_3494,N_3438);
nand U3548 (N_3548,N_3492,N_3368);
and U3549 (N_3549,N_3445,N_3366);
nand U3550 (N_3550,N_3491,N_3419);
or U3551 (N_3551,N_3447,N_3405);
or U3552 (N_3552,N_3479,N_3433);
and U3553 (N_3553,N_3465,N_3485);
or U3554 (N_3554,N_3361,N_3516);
and U3555 (N_3555,N_3387,N_3509);
and U3556 (N_3556,N_3471,N_3415);
xor U3557 (N_3557,N_3507,N_3495);
nand U3558 (N_3558,N_3463,N_3484);
nor U3559 (N_3559,N_3460,N_3519);
and U3560 (N_3560,N_3386,N_3363);
nand U3561 (N_3561,N_3430,N_3442);
and U3562 (N_3562,N_3477,N_3389);
and U3563 (N_3563,N_3388,N_3514);
or U3564 (N_3564,N_3421,N_3478);
nand U3565 (N_3565,N_3502,N_3431);
and U3566 (N_3566,N_3397,N_3367);
and U3567 (N_3567,N_3362,N_3497);
and U3568 (N_3568,N_3365,N_3480);
and U3569 (N_3569,N_3376,N_3420);
and U3570 (N_3570,N_3458,N_3383);
or U3571 (N_3571,N_3440,N_3427);
or U3572 (N_3572,N_3373,N_3476);
xnor U3573 (N_3573,N_3517,N_3360);
and U3574 (N_3574,N_3428,N_3456);
or U3575 (N_3575,N_3391,N_3390);
nor U3576 (N_3576,N_3470,N_3385);
or U3577 (N_3577,N_3467,N_3375);
or U3578 (N_3578,N_3506,N_3481);
nand U3579 (N_3579,N_3449,N_3501);
and U3580 (N_3580,N_3401,N_3510);
or U3581 (N_3581,N_3483,N_3500);
and U3582 (N_3582,N_3403,N_3462);
nor U3583 (N_3583,N_3499,N_3384);
xnor U3584 (N_3584,N_3469,N_3410);
and U3585 (N_3585,N_3473,N_3416);
or U3586 (N_3586,N_3472,N_3489);
xor U3587 (N_3587,N_3512,N_3406);
xnor U3588 (N_3588,N_3434,N_3372);
or U3589 (N_3589,N_3393,N_3418);
nand U3590 (N_3590,N_3392,N_3455);
and U3591 (N_3591,N_3422,N_3396);
nor U3592 (N_3592,N_3380,N_3504);
xor U3593 (N_3593,N_3378,N_3404);
or U3594 (N_3594,N_3466,N_3459);
and U3595 (N_3595,N_3446,N_3379);
nand U3596 (N_3596,N_3399,N_3461);
nand U3597 (N_3597,N_3487,N_3414);
nor U3598 (N_3598,N_3374,N_3488);
or U3599 (N_3599,N_3369,N_3426);
nand U3600 (N_3600,N_3384,N_3398);
xnor U3601 (N_3601,N_3464,N_3389);
or U3602 (N_3602,N_3479,N_3435);
and U3603 (N_3603,N_3383,N_3360);
or U3604 (N_3604,N_3382,N_3431);
nor U3605 (N_3605,N_3495,N_3399);
and U3606 (N_3606,N_3499,N_3478);
or U3607 (N_3607,N_3401,N_3416);
nand U3608 (N_3608,N_3368,N_3490);
nor U3609 (N_3609,N_3494,N_3460);
or U3610 (N_3610,N_3519,N_3500);
or U3611 (N_3611,N_3460,N_3418);
nand U3612 (N_3612,N_3409,N_3495);
nand U3613 (N_3613,N_3515,N_3488);
xnor U3614 (N_3614,N_3398,N_3378);
xor U3615 (N_3615,N_3461,N_3430);
nor U3616 (N_3616,N_3457,N_3416);
nand U3617 (N_3617,N_3506,N_3416);
and U3618 (N_3618,N_3468,N_3505);
and U3619 (N_3619,N_3363,N_3429);
or U3620 (N_3620,N_3402,N_3404);
nor U3621 (N_3621,N_3378,N_3459);
and U3622 (N_3622,N_3464,N_3374);
nand U3623 (N_3623,N_3472,N_3452);
nand U3624 (N_3624,N_3444,N_3361);
nand U3625 (N_3625,N_3462,N_3455);
and U3626 (N_3626,N_3449,N_3500);
nand U3627 (N_3627,N_3501,N_3416);
or U3628 (N_3628,N_3453,N_3444);
nand U3629 (N_3629,N_3370,N_3501);
or U3630 (N_3630,N_3409,N_3440);
and U3631 (N_3631,N_3362,N_3377);
and U3632 (N_3632,N_3453,N_3427);
nor U3633 (N_3633,N_3371,N_3372);
nor U3634 (N_3634,N_3421,N_3403);
and U3635 (N_3635,N_3481,N_3367);
or U3636 (N_3636,N_3454,N_3453);
xnor U3637 (N_3637,N_3460,N_3363);
xor U3638 (N_3638,N_3376,N_3386);
and U3639 (N_3639,N_3467,N_3470);
or U3640 (N_3640,N_3403,N_3396);
nand U3641 (N_3641,N_3397,N_3482);
or U3642 (N_3642,N_3376,N_3501);
nand U3643 (N_3643,N_3383,N_3467);
and U3644 (N_3644,N_3470,N_3371);
or U3645 (N_3645,N_3416,N_3466);
nor U3646 (N_3646,N_3403,N_3493);
and U3647 (N_3647,N_3374,N_3487);
and U3648 (N_3648,N_3362,N_3378);
or U3649 (N_3649,N_3426,N_3486);
and U3650 (N_3650,N_3429,N_3517);
xnor U3651 (N_3651,N_3361,N_3392);
nand U3652 (N_3652,N_3383,N_3435);
and U3653 (N_3653,N_3439,N_3448);
nand U3654 (N_3654,N_3366,N_3506);
nand U3655 (N_3655,N_3495,N_3435);
nor U3656 (N_3656,N_3446,N_3502);
xor U3657 (N_3657,N_3457,N_3405);
nor U3658 (N_3658,N_3376,N_3488);
nand U3659 (N_3659,N_3461,N_3478);
xor U3660 (N_3660,N_3381,N_3490);
nand U3661 (N_3661,N_3419,N_3437);
nor U3662 (N_3662,N_3399,N_3481);
xnor U3663 (N_3663,N_3428,N_3503);
nand U3664 (N_3664,N_3379,N_3410);
and U3665 (N_3665,N_3431,N_3516);
xnor U3666 (N_3666,N_3447,N_3401);
or U3667 (N_3667,N_3402,N_3446);
nor U3668 (N_3668,N_3464,N_3444);
and U3669 (N_3669,N_3375,N_3381);
and U3670 (N_3670,N_3458,N_3480);
nand U3671 (N_3671,N_3436,N_3478);
and U3672 (N_3672,N_3394,N_3368);
xnor U3673 (N_3673,N_3383,N_3457);
nand U3674 (N_3674,N_3382,N_3407);
or U3675 (N_3675,N_3477,N_3453);
nor U3676 (N_3676,N_3386,N_3379);
nand U3677 (N_3677,N_3416,N_3442);
and U3678 (N_3678,N_3380,N_3415);
nand U3679 (N_3679,N_3415,N_3482);
nand U3680 (N_3680,N_3586,N_3583);
xor U3681 (N_3681,N_3614,N_3632);
xor U3682 (N_3682,N_3557,N_3587);
nand U3683 (N_3683,N_3677,N_3618);
nand U3684 (N_3684,N_3604,N_3643);
nor U3685 (N_3685,N_3592,N_3554);
or U3686 (N_3686,N_3619,N_3631);
nor U3687 (N_3687,N_3527,N_3674);
xnor U3688 (N_3688,N_3542,N_3574);
xor U3689 (N_3689,N_3546,N_3679);
nor U3690 (N_3690,N_3622,N_3522);
or U3691 (N_3691,N_3573,N_3575);
or U3692 (N_3692,N_3629,N_3598);
xnor U3693 (N_3693,N_3625,N_3675);
nand U3694 (N_3694,N_3596,N_3676);
xnor U3695 (N_3695,N_3637,N_3539);
nor U3696 (N_3696,N_3562,N_3566);
xor U3697 (N_3697,N_3582,N_3572);
and U3698 (N_3698,N_3535,N_3634);
nand U3699 (N_3699,N_3594,N_3523);
and U3700 (N_3700,N_3659,N_3662);
or U3701 (N_3701,N_3521,N_3644);
or U3702 (N_3702,N_3646,N_3548);
or U3703 (N_3703,N_3612,N_3616);
xnor U3704 (N_3704,N_3669,N_3597);
nor U3705 (N_3705,N_3623,N_3526);
nand U3706 (N_3706,N_3638,N_3652);
xnor U3707 (N_3707,N_3569,N_3571);
xnor U3708 (N_3708,N_3590,N_3593);
and U3709 (N_3709,N_3529,N_3520);
nor U3710 (N_3710,N_3530,N_3670);
nand U3711 (N_3711,N_3615,N_3556);
and U3712 (N_3712,N_3552,N_3567);
xor U3713 (N_3713,N_3544,N_3600);
xor U3714 (N_3714,N_3601,N_3649);
xnor U3715 (N_3715,N_3621,N_3578);
xnor U3716 (N_3716,N_3534,N_3543);
xor U3717 (N_3717,N_3609,N_3541);
xnor U3718 (N_3718,N_3560,N_3606);
nand U3719 (N_3719,N_3536,N_3651);
and U3720 (N_3720,N_3605,N_3627);
or U3721 (N_3721,N_3610,N_3540);
nor U3722 (N_3722,N_3673,N_3648);
nor U3723 (N_3723,N_3570,N_3666);
nor U3724 (N_3724,N_3663,N_3549);
nor U3725 (N_3725,N_3568,N_3672);
or U3726 (N_3726,N_3640,N_3550);
or U3727 (N_3727,N_3668,N_3532);
nor U3728 (N_3728,N_3559,N_3645);
xor U3729 (N_3729,N_3664,N_3531);
or U3730 (N_3730,N_3551,N_3564);
or U3731 (N_3731,N_3528,N_3657);
nor U3732 (N_3732,N_3555,N_3577);
and U3733 (N_3733,N_3613,N_3576);
xnor U3734 (N_3734,N_3620,N_3642);
nand U3735 (N_3735,N_3547,N_3563);
or U3736 (N_3736,N_3584,N_3628);
or U3737 (N_3737,N_3658,N_3537);
nand U3738 (N_3738,N_3653,N_3639);
xor U3739 (N_3739,N_3595,N_3671);
or U3740 (N_3740,N_3553,N_3588);
nand U3741 (N_3741,N_3533,N_3635);
xnor U3742 (N_3742,N_3589,N_3585);
nor U3743 (N_3743,N_3558,N_3580);
or U3744 (N_3744,N_3607,N_3665);
and U3745 (N_3745,N_3565,N_3611);
or U3746 (N_3746,N_3579,N_3603);
nor U3747 (N_3747,N_3654,N_3581);
xor U3748 (N_3748,N_3525,N_3626);
nor U3749 (N_3749,N_3678,N_3656);
nand U3750 (N_3750,N_3667,N_3650);
xnor U3751 (N_3751,N_3545,N_3624);
and U3752 (N_3752,N_3641,N_3636);
or U3753 (N_3753,N_3602,N_3538);
nor U3754 (N_3754,N_3608,N_3660);
xor U3755 (N_3755,N_3599,N_3591);
nand U3756 (N_3756,N_3617,N_3561);
or U3757 (N_3757,N_3524,N_3655);
and U3758 (N_3758,N_3633,N_3647);
xor U3759 (N_3759,N_3661,N_3630);
and U3760 (N_3760,N_3590,N_3553);
and U3761 (N_3761,N_3620,N_3606);
and U3762 (N_3762,N_3657,N_3627);
or U3763 (N_3763,N_3630,N_3526);
or U3764 (N_3764,N_3678,N_3535);
xnor U3765 (N_3765,N_3567,N_3647);
or U3766 (N_3766,N_3525,N_3675);
and U3767 (N_3767,N_3674,N_3679);
or U3768 (N_3768,N_3546,N_3597);
nand U3769 (N_3769,N_3525,N_3602);
nor U3770 (N_3770,N_3604,N_3588);
nand U3771 (N_3771,N_3633,N_3549);
and U3772 (N_3772,N_3665,N_3520);
and U3773 (N_3773,N_3618,N_3662);
xnor U3774 (N_3774,N_3529,N_3580);
and U3775 (N_3775,N_3632,N_3675);
xnor U3776 (N_3776,N_3546,N_3654);
nand U3777 (N_3777,N_3526,N_3569);
and U3778 (N_3778,N_3560,N_3548);
nand U3779 (N_3779,N_3579,N_3663);
xnor U3780 (N_3780,N_3552,N_3619);
and U3781 (N_3781,N_3667,N_3563);
or U3782 (N_3782,N_3568,N_3647);
nor U3783 (N_3783,N_3637,N_3526);
nor U3784 (N_3784,N_3591,N_3555);
nor U3785 (N_3785,N_3547,N_3568);
or U3786 (N_3786,N_3605,N_3677);
nor U3787 (N_3787,N_3533,N_3658);
or U3788 (N_3788,N_3551,N_3671);
xnor U3789 (N_3789,N_3651,N_3598);
xnor U3790 (N_3790,N_3536,N_3650);
nand U3791 (N_3791,N_3650,N_3551);
xor U3792 (N_3792,N_3532,N_3599);
and U3793 (N_3793,N_3614,N_3642);
nand U3794 (N_3794,N_3549,N_3604);
nor U3795 (N_3795,N_3640,N_3650);
and U3796 (N_3796,N_3550,N_3644);
nor U3797 (N_3797,N_3664,N_3595);
nor U3798 (N_3798,N_3653,N_3534);
xnor U3799 (N_3799,N_3604,N_3614);
nor U3800 (N_3800,N_3599,N_3623);
xnor U3801 (N_3801,N_3527,N_3585);
or U3802 (N_3802,N_3528,N_3542);
or U3803 (N_3803,N_3612,N_3657);
nand U3804 (N_3804,N_3651,N_3678);
xor U3805 (N_3805,N_3533,N_3604);
xor U3806 (N_3806,N_3643,N_3618);
xor U3807 (N_3807,N_3631,N_3559);
nor U3808 (N_3808,N_3608,N_3568);
nand U3809 (N_3809,N_3609,N_3669);
nand U3810 (N_3810,N_3641,N_3656);
and U3811 (N_3811,N_3621,N_3640);
nand U3812 (N_3812,N_3520,N_3620);
xor U3813 (N_3813,N_3555,N_3581);
nand U3814 (N_3814,N_3639,N_3593);
nand U3815 (N_3815,N_3654,N_3636);
xor U3816 (N_3816,N_3585,N_3676);
and U3817 (N_3817,N_3633,N_3590);
and U3818 (N_3818,N_3583,N_3610);
nand U3819 (N_3819,N_3538,N_3667);
nor U3820 (N_3820,N_3624,N_3653);
or U3821 (N_3821,N_3539,N_3580);
or U3822 (N_3822,N_3648,N_3570);
nand U3823 (N_3823,N_3568,N_3651);
nor U3824 (N_3824,N_3583,N_3580);
nor U3825 (N_3825,N_3547,N_3536);
nor U3826 (N_3826,N_3605,N_3524);
nor U3827 (N_3827,N_3608,N_3620);
nor U3828 (N_3828,N_3613,N_3617);
xor U3829 (N_3829,N_3654,N_3660);
nor U3830 (N_3830,N_3632,N_3592);
nor U3831 (N_3831,N_3636,N_3593);
nand U3832 (N_3832,N_3554,N_3556);
or U3833 (N_3833,N_3546,N_3643);
nor U3834 (N_3834,N_3557,N_3564);
nor U3835 (N_3835,N_3520,N_3558);
xnor U3836 (N_3836,N_3522,N_3545);
nand U3837 (N_3837,N_3576,N_3555);
nand U3838 (N_3838,N_3646,N_3594);
and U3839 (N_3839,N_3590,N_3559);
and U3840 (N_3840,N_3719,N_3772);
and U3841 (N_3841,N_3798,N_3702);
and U3842 (N_3842,N_3818,N_3721);
and U3843 (N_3843,N_3807,N_3788);
and U3844 (N_3844,N_3715,N_3824);
and U3845 (N_3845,N_3685,N_3720);
or U3846 (N_3846,N_3749,N_3794);
xor U3847 (N_3847,N_3727,N_3823);
xor U3848 (N_3848,N_3746,N_3802);
xnor U3849 (N_3849,N_3728,N_3690);
nand U3850 (N_3850,N_3747,N_3765);
or U3851 (N_3851,N_3808,N_3785);
or U3852 (N_3852,N_3726,N_3713);
nor U3853 (N_3853,N_3722,N_3832);
or U3854 (N_3854,N_3680,N_3683);
nor U3855 (N_3855,N_3835,N_3793);
nor U3856 (N_3856,N_3718,N_3745);
and U3857 (N_3857,N_3767,N_3730);
nor U3858 (N_3858,N_3742,N_3790);
or U3859 (N_3859,N_3812,N_3725);
xor U3860 (N_3860,N_3731,N_3744);
xnor U3861 (N_3861,N_3752,N_3831);
nand U3862 (N_3862,N_3733,N_3696);
nor U3863 (N_3863,N_3710,N_3756);
and U3864 (N_3864,N_3754,N_3780);
and U3865 (N_3865,N_3688,N_3819);
nand U3866 (N_3866,N_3748,N_3682);
nand U3867 (N_3867,N_3829,N_3757);
and U3868 (N_3868,N_3777,N_3801);
nand U3869 (N_3869,N_3769,N_3751);
xnor U3870 (N_3870,N_3741,N_3686);
nand U3871 (N_3871,N_3701,N_3714);
nor U3872 (N_3872,N_3833,N_3804);
nor U3873 (N_3873,N_3740,N_3707);
nand U3874 (N_3874,N_3732,N_3792);
and U3875 (N_3875,N_3779,N_3813);
nand U3876 (N_3876,N_3783,N_3787);
or U3877 (N_3877,N_3753,N_3768);
nand U3878 (N_3878,N_3795,N_3805);
nor U3879 (N_3879,N_3723,N_3729);
or U3880 (N_3880,N_3814,N_3828);
or U3881 (N_3881,N_3736,N_3773);
or U3882 (N_3882,N_3758,N_3698);
xnor U3883 (N_3883,N_3826,N_3761);
nor U3884 (N_3884,N_3684,N_3735);
and U3885 (N_3885,N_3820,N_3778);
nor U3886 (N_3886,N_3709,N_3763);
or U3887 (N_3887,N_3695,N_3734);
or U3888 (N_3888,N_3704,N_3737);
and U3889 (N_3889,N_3810,N_3760);
and U3890 (N_3890,N_3822,N_3782);
nand U3891 (N_3891,N_3681,N_3799);
xor U3892 (N_3892,N_3774,N_3706);
xor U3893 (N_3893,N_3750,N_3691);
nor U3894 (N_3894,N_3837,N_3711);
and U3895 (N_3895,N_3825,N_3775);
xnor U3896 (N_3896,N_3806,N_3781);
nor U3897 (N_3897,N_3743,N_3700);
and U3898 (N_3898,N_3803,N_3703);
nand U3899 (N_3899,N_3789,N_3739);
and U3900 (N_3900,N_3817,N_3776);
nor U3901 (N_3901,N_3821,N_3809);
and U3902 (N_3902,N_3764,N_3770);
xnor U3903 (N_3903,N_3811,N_3830);
nor U3904 (N_3904,N_3692,N_3712);
nand U3905 (N_3905,N_3816,N_3716);
xor U3906 (N_3906,N_3708,N_3836);
xor U3907 (N_3907,N_3689,N_3834);
nand U3908 (N_3908,N_3800,N_3838);
nor U3909 (N_3909,N_3762,N_3738);
and U3910 (N_3910,N_3784,N_3697);
or U3911 (N_3911,N_3791,N_3796);
or U3912 (N_3912,N_3699,N_3797);
xor U3913 (N_3913,N_3815,N_3693);
nand U3914 (N_3914,N_3724,N_3705);
nor U3915 (N_3915,N_3755,N_3786);
nor U3916 (N_3916,N_3717,N_3766);
nor U3917 (N_3917,N_3687,N_3759);
and U3918 (N_3918,N_3839,N_3827);
or U3919 (N_3919,N_3694,N_3771);
xor U3920 (N_3920,N_3809,N_3830);
or U3921 (N_3921,N_3789,N_3773);
and U3922 (N_3922,N_3767,N_3710);
and U3923 (N_3923,N_3720,N_3818);
and U3924 (N_3924,N_3695,N_3781);
and U3925 (N_3925,N_3699,N_3716);
or U3926 (N_3926,N_3684,N_3731);
xnor U3927 (N_3927,N_3811,N_3686);
nand U3928 (N_3928,N_3720,N_3694);
nor U3929 (N_3929,N_3829,N_3792);
or U3930 (N_3930,N_3715,N_3688);
nand U3931 (N_3931,N_3788,N_3690);
and U3932 (N_3932,N_3761,N_3760);
nand U3933 (N_3933,N_3788,N_3735);
xor U3934 (N_3934,N_3753,N_3750);
or U3935 (N_3935,N_3684,N_3738);
xnor U3936 (N_3936,N_3745,N_3813);
or U3937 (N_3937,N_3839,N_3809);
xor U3938 (N_3938,N_3766,N_3774);
and U3939 (N_3939,N_3728,N_3783);
xnor U3940 (N_3940,N_3769,N_3746);
nand U3941 (N_3941,N_3746,N_3784);
or U3942 (N_3942,N_3688,N_3759);
nand U3943 (N_3943,N_3797,N_3821);
nand U3944 (N_3944,N_3766,N_3684);
xor U3945 (N_3945,N_3728,N_3697);
nor U3946 (N_3946,N_3685,N_3760);
nand U3947 (N_3947,N_3802,N_3796);
nand U3948 (N_3948,N_3836,N_3775);
xor U3949 (N_3949,N_3814,N_3707);
and U3950 (N_3950,N_3721,N_3771);
nand U3951 (N_3951,N_3741,N_3732);
xnor U3952 (N_3952,N_3831,N_3785);
nor U3953 (N_3953,N_3710,N_3785);
nand U3954 (N_3954,N_3691,N_3762);
and U3955 (N_3955,N_3787,N_3704);
and U3956 (N_3956,N_3751,N_3796);
nor U3957 (N_3957,N_3822,N_3687);
and U3958 (N_3958,N_3804,N_3752);
xnor U3959 (N_3959,N_3730,N_3825);
nand U3960 (N_3960,N_3725,N_3717);
and U3961 (N_3961,N_3764,N_3798);
and U3962 (N_3962,N_3837,N_3805);
xor U3963 (N_3963,N_3789,N_3711);
and U3964 (N_3964,N_3685,N_3684);
xnor U3965 (N_3965,N_3799,N_3791);
xnor U3966 (N_3966,N_3690,N_3836);
or U3967 (N_3967,N_3802,N_3728);
or U3968 (N_3968,N_3793,N_3766);
nand U3969 (N_3969,N_3729,N_3728);
nor U3970 (N_3970,N_3740,N_3692);
nor U3971 (N_3971,N_3746,N_3708);
and U3972 (N_3972,N_3725,N_3727);
and U3973 (N_3973,N_3707,N_3684);
nand U3974 (N_3974,N_3774,N_3763);
or U3975 (N_3975,N_3774,N_3745);
nand U3976 (N_3976,N_3723,N_3818);
and U3977 (N_3977,N_3681,N_3721);
nand U3978 (N_3978,N_3689,N_3806);
xor U3979 (N_3979,N_3719,N_3705);
xor U3980 (N_3980,N_3766,N_3812);
or U3981 (N_3981,N_3702,N_3734);
xor U3982 (N_3982,N_3747,N_3792);
and U3983 (N_3983,N_3761,N_3694);
nand U3984 (N_3984,N_3683,N_3836);
or U3985 (N_3985,N_3753,N_3814);
xor U3986 (N_3986,N_3690,N_3744);
or U3987 (N_3987,N_3789,N_3811);
or U3988 (N_3988,N_3823,N_3701);
and U3989 (N_3989,N_3768,N_3718);
nor U3990 (N_3990,N_3697,N_3814);
and U3991 (N_3991,N_3812,N_3694);
nor U3992 (N_3992,N_3794,N_3696);
xor U3993 (N_3993,N_3803,N_3760);
nand U3994 (N_3994,N_3715,N_3800);
xnor U3995 (N_3995,N_3836,N_3730);
or U3996 (N_3996,N_3839,N_3784);
nand U3997 (N_3997,N_3797,N_3755);
or U3998 (N_3998,N_3792,N_3775);
or U3999 (N_3999,N_3838,N_3697);
nor U4000 (N_4000,N_3974,N_3868);
nand U4001 (N_4001,N_3958,N_3897);
nand U4002 (N_4002,N_3875,N_3845);
or U4003 (N_4003,N_3883,N_3996);
nor U4004 (N_4004,N_3862,N_3870);
or U4005 (N_4005,N_3983,N_3926);
or U4006 (N_4006,N_3960,N_3962);
or U4007 (N_4007,N_3850,N_3898);
or U4008 (N_4008,N_3994,N_3989);
nor U4009 (N_4009,N_3855,N_3890);
nor U4010 (N_4010,N_3916,N_3904);
or U4011 (N_4011,N_3886,N_3967);
nor U4012 (N_4012,N_3963,N_3876);
nor U4013 (N_4013,N_3976,N_3851);
nand U4014 (N_4014,N_3881,N_3987);
xnor U4015 (N_4015,N_3867,N_3884);
or U4016 (N_4016,N_3859,N_3921);
xnor U4017 (N_4017,N_3912,N_3950);
xor U4018 (N_4018,N_3937,N_3847);
and U4019 (N_4019,N_3914,N_3968);
nand U4020 (N_4020,N_3892,N_3879);
xor U4021 (N_4021,N_3894,N_3938);
or U4022 (N_4022,N_3840,N_3857);
nor U4023 (N_4023,N_3891,N_3854);
xor U4024 (N_4024,N_3978,N_3952);
nand U4025 (N_4025,N_3911,N_3947);
nand U4026 (N_4026,N_3972,N_3988);
or U4027 (N_4027,N_3946,N_3929);
and U4028 (N_4028,N_3858,N_3910);
nor U4029 (N_4029,N_3917,N_3882);
xor U4030 (N_4030,N_3990,N_3860);
nand U4031 (N_4031,N_3841,N_3955);
or U4032 (N_4032,N_3942,N_3901);
and U4033 (N_4033,N_3985,N_3940);
nor U4034 (N_4034,N_3930,N_3935);
or U4035 (N_4035,N_3915,N_3872);
or U4036 (N_4036,N_3948,N_3936);
and U4037 (N_4037,N_3856,N_3895);
nor U4038 (N_4038,N_3893,N_3975);
nand U4039 (N_4039,N_3969,N_3902);
or U4040 (N_4040,N_3995,N_3887);
or U4041 (N_4041,N_3924,N_3889);
nor U4042 (N_4042,N_3923,N_3964);
xor U4043 (N_4043,N_3998,N_3866);
nor U4044 (N_4044,N_3843,N_3844);
nor U4045 (N_4045,N_3846,N_3900);
nor U4046 (N_4046,N_3931,N_3909);
or U4047 (N_4047,N_3874,N_3849);
xor U4048 (N_4048,N_3943,N_3906);
nand U4049 (N_4049,N_3878,N_3918);
nor U4050 (N_4050,N_3956,N_3944);
xor U4051 (N_4051,N_3853,N_3899);
and U4052 (N_4052,N_3903,N_3980);
xnor U4053 (N_4053,N_3939,N_3984);
and U4054 (N_4054,N_3966,N_3873);
nor U4055 (N_4055,N_3869,N_3864);
and U4056 (N_4056,N_3877,N_3919);
and U4057 (N_4057,N_3885,N_3953);
nor U4058 (N_4058,N_3888,N_3973);
xor U4059 (N_4059,N_3992,N_3954);
or U4060 (N_4060,N_3908,N_3951);
nand U4061 (N_4061,N_3991,N_3945);
and U4062 (N_4062,N_3863,N_3965);
or U4063 (N_4063,N_3928,N_3957);
or U4064 (N_4064,N_3852,N_3922);
nor U4065 (N_4065,N_3979,N_3871);
or U4066 (N_4066,N_3932,N_3842);
or U4067 (N_4067,N_3977,N_3993);
xnor U4068 (N_4068,N_3920,N_3880);
nand U4069 (N_4069,N_3848,N_3971);
nand U4070 (N_4070,N_3949,N_3861);
nand U4071 (N_4071,N_3905,N_3997);
or U4072 (N_4072,N_3927,N_3913);
nor U4073 (N_4073,N_3986,N_3865);
or U4074 (N_4074,N_3999,N_3907);
or U4075 (N_4075,N_3933,N_3934);
nor U4076 (N_4076,N_3961,N_3896);
xnor U4077 (N_4077,N_3981,N_3970);
and U4078 (N_4078,N_3982,N_3925);
or U4079 (N_4079,N_3941,N_3959);
xor U4080 (N_4080,N_3937,N_3939);
and U4081 (N_4081,N_3871,N_3875);
or U4082 (N_4082,N_3856,N_3878);
or U4083 (N_4083,N_3861,N_3923);
nor U4084 (N_4084,N_3946,N_3901);
nor U4085 (N_4085,N_3988,N_3925);
xor U4086 (N_4086,N_3992,N_3908);
nand U4087 (N_4087,N_3924,N_3896);
xor U4088 (N_4088,N_3989,N_3864);
nand U4089 (N_4089,N_3969,N_3924);
and U4090 (N_4090,N_3924,N_3891);
and U4091 (N_4091,N_3913,N_3848);
and U4092 (N_4092,N_3949,N_3862);
nand U4093 (N_4093,N_3875,N_3987);
and U4094 (N_4094,N_3939,N_3987);
and U4095 (N_4095,N_3968,N_3864);
nor U4096 (N_4096,N_3953,N_3978);
xor U4097 (N_4097,N_3926,N_3995);
nand U4098 (N_4098,N_3915,N_3916);
and U4099 (N_4099,N_3873,N_3994);
or U4100 (N_4100,N_3987,N_3904);
and U4101 (N_4101,N_3918,N_3949);
nor U4102 (N_4102,N_3999,N_3943);
and U4103 (N_4103,N_3880,N_3939);
and U4104 (N_4104,N_3840,N_3910);
or U4105 (N_4105,N_3874,N_3913);
xor U4106 (N_4106,N_3980,N_3956);
or U4107 (N_4107,N_3948,N_3937);
nor U4108 (N_4108,N_3935,N_3964);
or U4109 (N_4109,N_3960,N_3917);
and U4110 (N_4110,N_3894,N_3988);
xnor U4111 (N_4111,N_3955,N_3979);
or U4112 (N_4112,N_3883,N_3887);
xnor U4113 (N_4113,N_3854,N_3973);
nand U4114 (N_4114,N_3903,N_3894);
nor U4115 (N_4115,N_3863,N_3984);
and U4116 (N_4116,N_3922,N_3935);
nand U4117 (N_4117,N_3967,N_3854);
and U4118 (N_4118,N_3911,N_3926);
nand U4119 (N_4119,N_3841,N_3944);
nor U4120 (N_4120,N_3941,N_3886);
or U4121 (N_4121,N_3858,N_3979);
and U4122 (N_4122,N_3912,N_3952);
or U4123 (N_4123,N_3961,N_3992);
and U4124 (N_4124,N_3900,N_3896);
and U4125 (N_4125,N_3990,N_3887);
and U4126 (N_4126,N_3886,N_3865);
nor U4127 (N_4127,N_3869,N_3969);
and U4128 (N_4128,N_3949,N_3972);
and U4129 (N_4129,N_3859,N_3933);
xor U4130 (N_4130,N_3953,N_3918);
nand U4131 (N_4131,N_3904,N_3871);
xnor U4132 (N_4132,N_3987,N_3982);
xor U4133 (N_4133,N_3887,N_3889);
xor U4134 (N_4134,N_3951,N_3891);
and U4135 (N_4135,N_3945,N_3926);
and U4136 (N_4136,N_3927,N_3921);
xor U4137 (N_4137,N_3942,N_3978);
nor U4138 (N_4138,N_3919,N_3841);
or U4139 (N_4139,N_3852,N_3863);
nand U4140 (N_4140,N_3930,N_3931);
and U4141 (N_4141,N_3857,N_3937);
or U4142 (N_4142,N_3959,N_3957);
nand U4143 (N_4143,N_3963,N_3858);
xor U4144 (N_4144,N_3971,N_3886);
nor U4145 (N_4145,N_3861,N_3895);
nand U4146 (N_4146,N_3901,N_3875);
xor U4147 (N_4147,N_3941,N_3868);
nor U4148 (N_4148,N_3845,N_3854);
or U4149 (N_4149,N_3927,N_3876);
and U4150 (N_4150,N_3897,N_3925);
xnor U4151 (N_4151,N_3962,N_3868);
nor U4152 (N_4152,N_3914,N_3845);
nand U4153 (N_4153,N_3885,N_3861);
nor U4154 (N_4154,N_3936,N_3905);
nand U4155 (N_4155,N_3918,N_3929);
nor U4156 (N_4156,N_3859,N_3858);
or U4157 (N_4157,N_3878,N_3971);
and U4158 (N_4158,N_3903,N_3921);
or U4159 (N_4159,N_3986,N_3967);
nor U4160 (N_4160,N_4017,N_4043);
or U4161 (N_4161,N_4128,N_4025);
or U4162 (N_4162,N_4086,N_4116);
and U4163 (N_4163,N_4014,N_4133);
nor U4164 (N_4164,N_4042,N_4099);
and U4165 (N_4165,N_4089,N_4144);
and U4166 (N_4166,N_4120,N_4040);
or U4167 (N_4167,N_4131,N_4072);
nand U4168 (N_4168,N_4057,N_4065);
and U4169 (N_4169,N_4005,N_4092);
and U4170 (N_4170,N_4064,N_4037);
nor U4171 (N_4171,N_4002,N_4053);
or U4172 (N_4172,N_4032,N_4123);
xor U4173 (N_4173,N_4115,N_4126);
nand U4174 (N_4174,N_4117,N_4024);
or U4175 (N_4175,N_4157,N_4097);
and U4176 (N_4176,N_4104,N_4114);
nand U4177 (N_4177,N_4008,N_4134);
nor U4178 (N_4178,N_4041,N_4074);
nand U4179 (N_4179,N_4029,N_4085);
and U4180 (N_4180,N_4052,N_4150);
and U4181 (N_4181,N_4106,N_4012);
xnor U4182 (N_4182,N_4075,N_4094);
or U4183 (N_4183,N_4050,N_4101);
xor U4184 (N_4184,N_4118,N_4148);
xnor U4185 (N_4185,N_4078,N_4054);
or U4186 (N_4186,N_4132,N_4135);
xnor U4187 (N_4187,N_4142,N_4080);
nor U4188 (N_4188,N_4045,N_4098);
nand U4189 (N_4189,N_4143,N_4141);
xor U4190 (N_4190,N_4076,N_4107);
xnor U4191 (N_4191,N_4071,N_4011);
xor U4192 (N_4192,N_4060,N_4129);
nor U4193 (N_4193,N_4103,N_4146);
xnor U4194 (N_4194,N_4038,N_4009);
xnor U4195 (N_4195,N_4001,N_4051);
xor U4196 (N_4196,N_4034,N_4109);
nor U4197 (N_4197,N_4046,N_4010);
and U4198 (N_4198,N_4121,N_4159);
nor U4199 (N_4199,N_4073,N_4026);
and U4200 (N_4200,N_4136,N_4039);
or U4201 (N_4201,N_4059,N_4091);
and U4202 (N_4202,N_4055,N_4048);
or U4203 (N_4203,N_4147,N_4061);
nor U4204 (N_4204,N_4003,N_4058);
nand U4205 (N_4205,N_4068,N_4093);
and U4206 (N_4206,N_4000,N_4006);
and U4207 (N_4207,N_4139,N_4067);
or U4208 (N_4208,N_4082,N_4021);
and U4209 (N_4209,N_4140,N_4130);
nor U4210 (N_4210,N_4063,N_4004);
and U4211 (N_4211,N_4020,N_4007);
and U4212 (N_4212,N_4028,N_4111);
xor U4213 (N_4213,N_4122,N_4138);
nand U4214 (N_4214,N_4018,N_4022);
nand U4215 (N_4215,N_4090,N_4105);
or U4216 (N_4216,N_4031,N_4016);
or U4217 (N_4217,N_4044,N_4013);
xnor U4218 (N_4218,N_4108,N_4027);
nand U4219 (N_4219,N_4096,N_4056);
nor U4220 (N_4220,N_4088,N_4047);
and U4221 (N_4221,N_4087,N_4095);
nor U4222 (N_4222,N_4153,N_4079);
or U4223 (N_4223,N_4149,N_4036);
xnor U4224 (N_4224,N_4081,N_4033);
xnor U4225 (N_4225,N_4030,N_4112);
xnor U4226 (N_4226,N_4102,N_4066);
nand U4227 (N_4227,N_4049,N_4035);
and U4228 (N_4228,N_4083,N_4070);
xnor U4229 (N_4229,N_4015,N_4110);
and U4230 (N_4230,N_4127,N_4019);
nor U4231 (N_4231,N_4152,N_4158);
xnor U4232 (N_4232,N_4151,N_4100);
nor U4233 (N_4233,N_4145,N_4137);
xor U4234 (N_4234,N_4155,N_4084);
nand U4235 (N_4235,N_4062,N_4124);
and U4236 (N_4236,N_4119,N_4154);
nand U4237 (N_4237,N_4077,N_4125);
and U4238 (N_4238,N_4113,N_4023);
nand U4239 (N_4239,N_4069,N_4156);
xnor U4240 (N_4240,N_4087,N_4004);
nand U4241 (N_4241,N_4101,N_4013);
or U4242 (N_4242,N_4134,N_4147);
nor U4243 (N_4243,N_4098,N_4050);
and U4244 (N_4244,N_4089,N_4079);
nor U4245 (N_4245,N_4033,N_4120);
nand U4246 (N_4246,N_4003,N_4089);
and U4247 (N_4247,N_4010,N_4089);
and U4248 (N_4248,N_4145,N_4149);
and U4249 (N_4249,N_4088,N_4010);
and U4250 (N_4250,N_4111,N_4122);
and U4251 (N_4251,N_4006,N_4126);
or U4252 (N_4252,N_4056,N_4097);
and U4253 (N_4253,N_4045,N_4005);
or U4254 (N_4254,N_4101,N_4109);
nand U4255 (N_4255,N_4141,N_4064);
nor U4256 (N_4256,N_4105,N_4127);
nor U4257 (N_4257,N_4122,N_4113);
or U4258 (N_4258,N_4103,N_4085);
nor U4259 (N_4259,N_4139,N_4025);
xor U4260 (N_4260,N_4132,N_4016);
xnor U4261 (N_4261,N_4018,N_4068);
or U4262 (N_4262,N_4123,N_4000);
or U4263 (N_4263,N_4065,N_4046);
nor U4264 (N_4264,N_4066,N_4083);
xnor U4265 (N_4265,N_4131,N_4158);
xnor U4266 (N_4266,N_4110,N_4044);
nor U4267 (N_4267,N_4096,N_4020);
or U4268 (N_4268,N_4028,N_4070);
xnor U4269 (N_4269,N_4027,N_4153);
or U4270 (N_4270,N_4063,N_4127);
xnor U4271 (N_4271,N_4043,N_4106);
and U4272 (N_4272,N_4087,N_4106);
or U4273 (N_4273,N_4051,N_4078);
xor U4274 (N_4274,N_4138,N_4099);
nand U4275 (N_4275,N_4084,N_4136);
or U4276 (N_4276,N_4092,N_4070);
and U4277 (N_4277,N_4013,N_4047);
and U4278 (N_4278,N_4072,N_4099);
xnor U4279 (N_4279,N_4078,N_4124);
nor U4280 (N_4280,N_4024,N_4010);
xor U4281 (N_4281,N_4071,N_4047);
or U4282 (N_4282,N_4121,N_4046);
or U4283 (N_4283,N_4107,N_4036);
nand U4284 (N_4284,N_4138,N_4139);
nor U4285 (N_4285,N_4051,N_4149);
or U4286 (N_4286,N_4082,N_4022);
nor U4287 (N_4287,N_4135,N_4078);
nor U4288 (N_4288,N_4066,N_4112);
and U4289 (N_4289,N_4069,N_4118);
nand U4290 (N_4290,N_4125,N_4028);
or U4291 (N_4291,N_4008,N_4011);
or U4292 (N_4292,N_4063,N_4075);
and U4293 (N_4293,N_4123,N_4112);
nand U4294 (N_4294,N_4016,N_4095);
or U4295 (N_4295,N_4059,N_4124);
nand U4296 (N_4296,N_4028,N_4077);
nor U4297 (N_4297,N_4093,N_4009);
xnor U4298 (N_4298,N_4103,N_4070);
and U4299 (N_4299,N_4124,N_4145);
xor U4300 (N_4300,N_4099,N_4057);
xnor U4301 (N_4301,N_4143,N_4050);
or U4302 (N_4302,N_4076,N_4142);
xor U4303 (N_4303,N_4116,N_4051);
nand U4304 (N_4304,N_4112,N_4127);
xnor U4305 (N_4305,N_4146,N_4029);
nand U4306 (N_4306,N_4029,N_4159);
and U4307 (N_4307,N_4121,N_4035);
or U4308 (N_4308,N_4053,N_4137);
nor U4309 (N_4309,N_4137,N_4022);
and U4310 (N_4310,N_4012,N_4022);
nor U4311 (N_4311,N_4138,N_4061);
or U4312 (N_4312,N_4041,N_4129);
and U4313 (N_4313,N_4037,N_4002);
nor U4314 (N_4314,N_4128,N_4082);
and U4315 (N_4315,N_4005,N_4113);
nand U4316 (N_4316,N_4069,N_4145);
nand U4317 (N_4317,N_4005,N_4019);
xor U4318 (N_4318,N_4109,N_4141);
or U4319 (N_4319,N_4057,N_4009);
or U4320 (N_4320,N_4308,N_4204);
xor U4321 (N_4321,N_4261,N_4276);
nand U4322 (N_4322,N_4298,N_4221);
xor U4323 (N_4323,N_4263,N_4246);
or U4324 (N_4324,N_4272,N_4288);
and U4325 (N_4325,N_4319,N_4220);
nor U4326 (N_4326,N_4181,N_4300);
xnor U4327 (N_4327,N_4294,N_4282);
nand U4328 (N_4328,N_4219,N_4213);
nor U4329 (N_4329,N_4257,N_4193);
or U4330 (N_4330,N_4250,N_4232);
and U4331 (N_4331,N_4208,N_4160);
nand U4332 (N_4332,N_4316,N_4200);
xor U4333 (N_4333,N_4217,N_4179);
and U4334 (N_4334,N_4206,N_4191);
and U4335 (N_4335,N_4172,N_4162);
nor U4336 (N_4336,N_4266,N_4182);
or U4337 (N_4337,N_4164,N_4210);
or U4338 (N_4338,N_4203,N_4198);
nor U4339 (N_4339,N_4174,N_4199);
or U4340 (N_4340,N_4166,N_4314);
nor U4341 (N_4341,N_4167,N_4242);
nand U4342 (N_4342,N_4177,N_4241);
nand U4343 (N_4343,N_4201,N_4194);
and U4344 (N_4344,N_4259,N_4280);
and U4345 (N_4345,N_4278,N_4161);
and U4346 (N_4346,N_4163,N_4183);
or U4347 (N_4347,N_4315,N_4192);
nor U4348 (N_4348,N_4229,N_4239);
nor U4349 (N_4349,N_4245,N_4189);
and U4350 (N_4350,N_4311,N_4313);
or U4351 (N_4351,N_4253,N_4236);
or U4352 (N_4352,N_4240,N_4297);
nor U4353 (N_4353,N_4234,N_4281);
or U4354 (N_4354,N_4291,N_4285);
or U4355 (N_4355,N_4265,N_4279);
nor U4356 (N_4356,N_4283,N_4214);
xnor U4357 (N_4357,N_4271,N_4277);
nor U4358 (N_4358,N_4286,N_4270);
nor U4359 (N_4359,N_4223,N_4317);
or U4360 (N_4360,N_4244,N_4168);
or U4361 (N_4361,N_4267,N_4258);
nand U4362 (N_4362,N_4195,N_4231);
and U4363 (N_4363,N_4218,N_4260);
nand U4364 (N_4364,N_4228,N_4180);
xnor U4365 (N_4365,N_4310,N_4301);
and U4366 (N_4366,N_4309,N_4268);
or U4367 (N_4367,N_4171,N_4293);
and U4368 (N_4368,N_4185,N_4275);
nor U4369 (N_4369,N_4237,N_4256);
xor U4370 (N_4370,N_4186,N_4227);
nand U4371 (N_4371,N_4305,N_4207);
xor U4372 (N_4372,N_4302,N_4307);
nor U4373 (N_4373,N_4304,N_4295);
nor U4374 (N_4374,N_4178,N_4205);
or U4375 (N_4375,N_4209,N_4296);
xnor U4376 (N_4376,N_4292,N_4238);
xor U4377 (N_4377,N_4269,N_4252);
nor U4378 (N_4378,N_4169,N_4224);
or U4379 (N_4379,N_4289,N_4235);
nor U4380 (N_4380,N_4262,N_4173);
xor U4381 (N_4381,N_4312,N_4197);
nand U4382 (N_4382,N_4165,N_4190);
nor U4383 (N_4383,N_4170,N_4254);
nor U4384 (N_4384,N_4287,N_4255);
nor U4385 (N_4385,N_4196,N_4216);
nand U4386 (N_4386,N_4175,N_4233);
and U4387 (N_4387,N_4249,N_4222);
or U4388 (N_4388,N_4211,N_4184);
nor U4389 (N_4389,N_4176,N_4187);
xnor U4390 (N_4390,N_4274,N_4248);
nand U4391 (N_4391,N_4290,N_4264);
xnor U4392 (N_4392,N_4251,N_4225);
and U4393 (N_4393,N_4247,N_4230);
and U4394 (N_4394,N_4188,N_4318);
or U4395 (N_4395,N_4243,N_4202);
or U4396 (N_4396,N_4299,N_4215);
and U4397 (N_4397,N_4212,N_4303);
xor U4398 (N_4398,N_4273,N_4284);
and U4399 (N_4399,N_4226,N_4306);
and U4400 (N_4400,N_4288,N_4228);
nor U4401 (N_4401,N_4294,N_4192);
and U4402 (N_4402,N_4244,N_4245);
or U4403 (N_4403,N_4232,N_4171);
or U4404 (N_4404,N_4210,N_4296);
or U4405 (N_4405,N_4169,N_4251);
or U4406 (N_4406,N_4208,N_4174);
and U4407 (N_4407,N_4200,N_4218);
and U4408 (N_4408,N_4296,N_4280);
nand U4409 (N_4409,N_4191,N_4281);
or U4410 (N_4410,N_4251,N_4189);
xor U4411 (N_4411,N_4200,N_4209);
xnor U4412 (N_4412,N_4242,N_4169);
or U4413 (N_4413,N_4198,N_4246);
and U4414 (N_4414,N_4239,N_4179);
or U4415 (N_4415,N_4314,N_4308);
xnor U4416 (N_4416,N_4257,N_4211);
and U4417 (N_4417,N_4184,N_4267);
nand U4418 (N_4418,N_4228,N_4213);
and U4419 (N_4419,N_4229,N_4197);
or U4420 (N_4420,N_4195,N_4309);
xor U4421 (N_4421,N_4168,N_4208);
or U4422 (N_4422,N_4273,N_4261);
and U4423 (N_4423,N_4244,N_4257);
nor U4424 (N_4424,N_4161,N_4276);
xor U4425 (N_4425,N_4199,N_4300);
nand U4426 (N_4426,N_4266,N_4180);
or U4427 (N_4427,N_4182,N_4160);
or U4428 (N_4428,N_4235,N_4265);
xor U4429 (N_4429,N_4240,N_4209);
and U4430 (N_4430,N_4209,N_4197);
and U4431 (N_4431,N_4311,N_4305);
nor U4432 (N_4432,N_4265,N_4266);
or U4433 (N_4433,N_4310,N_4172);
or U4434 (N_4434,N_4286,N_4304);
or U4435 (N_4435,N_4228,N_4273);
xor U4436 (N_4436,N_4222,N_4250);
nor U4437 (N_4437,N_4248,N_4262);
xor U4438 (N_4438,N_4269,N_4280);
nor U4439 (N_4439,N_4281,N_4168);
or U4440 (N_4440,N_4267,N_4238);
nand U4441 (N_4441,N_4177,N_4208);
nand U4442 (N_4442,N_4209,N_4251);
nand U4443 (N_4443,N_4308,N_4189);
and U4444 (N_4444,N_4288,N_4238);
xnor U4445 (N_4445,N_4229,N_4271);
and U4446 (N_4446,N_4294,N_4296);
xnor U4447 (N_4447,N_4306,N_4165);
and U4448 (N_4448,N_4168,N_4279);
and U4449 (N_4449,N_4200,N_4168);
nand U4450 (N_4450,N_4279,N_4253);
and U4451 (N_4451,N_4287,N_4186);
nor U4452 (N_4452,N_4279,N_4237);
and U4453 (N_4453,N_4206,N_4213);
nor U4454 (N_4454,N_4186,N_4174);
nor U4455 (N_4455,N_4280,N_4193);
and U4456 (N_4456,N_4182,N_4186);
or U4457 (N_4457,N_4300,N_4257);
xnor U4458 (N_4458,N_4206,N_4291);
nor U4459 (N_4459,N_4217,N_4220);
or U4460 (N_4460,N_4234,N_4161);
or U4461 (N_4461,N_4317,N_4316);
nand U4462 (N_4462,N_4309,N_4252);
nand U4463 (N_4463,N_4186,N_4254);
or U4464 (N_4464,N_4264,N_4257);
nor U4465 (N_4465,N_4255,N_4276);
xor U4466 (N_4466,N_4302,N_4264);
nand U4467 (N_4467,N_4297,N_4260);
and U4468 (N_4468,N_4319,N_4243);
nor U4469 (N_4469,N_4309,N_4303);
or U4470 (N_4470,N_4283,N_4278);
nand U4471 (N_4471,N_4224,N_4304);
and U4472 (N_4472,N_4237,N_4287);
or U4473 (N_4473,N_4249,N_4319);
and U4474 (N_4474,N_4171,N_4202);
nand U4475 (N_4475,N_4301,N_4304);
nand U4476 (N_4476,N_4208,N_4265);
or U4477 (N_4477,N_4304,N_4275);
or U4478 (N_4478,N_4315,N_4168);
and U4479 (N_4479,N_4280,N_4263);
and U4480 (N_4480,N_4406,N_4368);
or U4481 (N_4481,N_4373,N_4418);
xor U4482 (N_4482,N_4407,N_4336);
nor U4483 (N_4483,N_4411,N_4396);
or U4484 (N_4484,N_4459,N_4466);
nand U4485 (N_4485,N_4405,N_4323);
and U4486 (N_4486,N_4453,N_4380);
and U4487 (N_4487,N_4346,N_4369);
and U4488 (N_4488,N_4385,N_4342);
or U4489 (N_4489,N_4364,N_4402);
or U4490 (N_4490,N_4353,N_4470);
and U4491 (N_4491,N_4362,N_4479);
xor U4492 (N_4492,N_4413,N_4387);
nand U4493 (N_4493,N_4360,N_4448);
and U4494 (N_4494,N_4356,N_4465);
nor U4495 (N_4495,N_4374,N_4442);
or U4496 (N_4496,N_4439,N_4367);
or U4497 (N_4497,N_4386,N_4460);
xor U4498 (N_4498,N_4434,N_4392);
nor U4499 (N_4499,N_4348,N_4471);
or U4500 (N_4500,N_4416,N_4433);
nand U4501 (N_4501,N_4330,N_4436);
nor U4502 (N_4502,N_4426,N_4437);
or U4503 (N_4503,N_4452,N_4320);
xnor U4504 (N_4504,N_4444,N_4422);
nand U4505 (N_4505,N_4420,N_4352);
nand U4506 (N_4506,N_4450,N_4438);
nor U4507 (N_4507,N_4399,N_4335);
or U4508 (N_4508,N_4337,N_4446);
nand U4509 (N_4509,N_4325,N_4350);
nor U4510 (N_4510,N_4467,N_4324);
and U4511 (N_4511,N_4358,N_4400);
xor U4512 (N_4512,N_4344,N_4351);
or U4513 (N_4513,N_4375,N_4359);
and U4514 (N_4514,N_4469,N_4449);
and U4515 (N_4515,N_4334,N_4332);
nor U4516 (N_4516,N_4461,N_4428);
nand U4517 (N_4517,N_4365,N_4409);
nor U4518 (N_4518,N_4427,N_4455);
xor U4519 (N_4519,N_4322,N_4424);
nand U4520 (N_4520,N_4475,N_4363);
or U4521 (N_4521,N_4457,N_4458);
nor U4522 (N_4522,N_4435,N_4329);
nor U4523 (N_4523,N_4404,N_4349);
or U4524 (N_4524,N_4454,N_4445);
xor U4525 (N_4525,N_4378,N_4476);
and U4526 (N_4526,N_4463,N_4401);
or U4527 (N_4527,N_4340,N_4390);
xnor U4528 (N_4528,N_4403,N_4414);
xor U4529 (N_4529,N_4474,N_4394);
or U4530 (N_4530,N_4377,N_4477);
nand U4531 (N_4531,N_4347,N_4472);
nand U4532 (N_4532,N_4361,N_4328);
nor U4533 (N_4533,N_4425,N_4397);
nand U4534 (N_4534,N_4423,N_4379);
nand U4535 (N_4535,N_4381,N_4410);
and U4536 (N_4536,N_4395,N_4354);
or U4537 (N_4537,N_4341,N_4326);
and U4538 (N_4538,N_4333,N_4331);
and U4539 (N_4539,N_4393,N_4451);
nand U4540 (N_4540,N_4355,N_4408);
and U4541 (N_4541,N_4376,N_4398);
and U4542 (N_4542,N_4343,N_4388);
nand U4543 (N_4543,N_4345,N_4464);
and U4544 (N_4544,N_4383,N_4447);
xnor U4545 (N_4545,N_4370,N_4432);
nor U4546 (N_4546,N_4431,N_4443);
and U4547 (N_4547,N_4372,N_4419);
or U4548 (N_4548,N_4389,N_4441);
and U4549 (N_4549,N_4456,N_4468);
or U4550 (N_4550,N_4421,N_4412);
or U4551 (N_4551,N_4429,N_4430);
nand U4552 (N_4552,N_4339,N_4391);
or U4553 (N_4553,N_4417,N_4371);
xor U4554 (N_4554,N_4366,N_4382);
xor U4555 (N_4555,N_4473,N_4415);
xnor U4556 (N_4556,N_4462,N_4440);
nor U4557 (N_4557,N_4384,N_4357);
and U4558 (N_4558,N_4478,N_4327);
xor U4559 (N_4559,N_4338,N_4321);
xor U4560 (N_4560,N_4406,N_4345);
xnor U4561 (N_4561,N_4442,N_4435);
or U4562 (N_4562,N_4331,N_4366);
and U4563 (N_4563,N_4409,N_4423);
or U4564 (N_4564,N_4389,N_4329);
nor U4565 (N_4565,N_4445,N_4344);
nor U4566 (N_4566,N_4438,N_4390);
and U4567 (N_4567,N_4447,N_4432);
or U4568 (N_4568,N_4468,N_4358);
nand U4569 (N_4569,N_4434,N_4406);
nand U4570 (N_4570,N_4321,N_4392);
xnor U4571 (N_4571,N_4376,N_4358);
nor U4572 (N_4572,N_4419,N_4325);
nor U4573 (N_4573,N_4365,N_4441);
nor U4574 (N_4574,N_4387,N_4384);
or U4575 (N_4575,N_4329,N_4373);
nand U4576 (N_4576,N_4372,N_4466);
or U4577 (N_4577,N_4470,N_4361);
or U4578 (N_4578,N_4369,N_4325);
and U4579 (N_4579,N_4444,N_4383);
and U4580 (N_4580,N_4433,N_4419);
xor U4581 (N_4581,N_4429,N_4406);
nor U4582 (N_4582,N_4450,N_4399);
nand U4583 (N_4583,N_4394,N_4455);
nand U4584 (N_4584,N_4326,N_4373);
and U4585 (N_4585,N_4479,N_4463);
nor U4586 (N_4586,N_4393,N_4366);
and U4587 (N_4587,N_4357,N_4447);
xor U4588 (N_4588,N_4344,N_4396);
nand U4589 (N_4589,N_4444,N_4457);
xnor U4590 (N_4590,N_4434,N_4449);
or U4591 (N_4591,N_4421,N_4322);
xnor U4592 (N_4592,N_4331,N_4450);
nand U4593 (N_4593,N_4439,N_4420);
nor U4594 (N_4594,N_4377,N_4328);
xor U4595 (N_4595,N_4326,N_4426);
xor U4596 (N_4596,N_4381,N_4454);
nand U4597 (N_4597,N_4378,N_4432);
xnor U4598 (N_4598,N_4384,N_4360);
xor U4599 (N_4599,N_4461,N_4478);
nand U4600 (N_4600,N_4440,N_4338);
and U4601 (N_4601,N_4336,N_4415);
or U4602 (N_4602,N_4353,N_4437);
or U4603 (N_4603,N_4470,N_4432);
and U4604 (N_4604,N_4443,N_4395);
or U4605 (N_4605,N_4416,N_4367);
nand U4606 (N_4606,N_4391,N_4412);
and U4607 (N_4607,N_4459,N_4469);
xor U4608 (N_4608,N_4324,N_4339);
and U4609 (N_4609,N_4415,N_4325);
nor U4610 (N_4610,N_4368,N_4446);
nor U4611 (N_4611,N_4447,N_4412);
nand U4612 (N_4612,N_4466,N_4360);
or U4613 (N_4613,N_4365,N_4341);
xor U4614 (N_4614,N_4437,N_4367);
xor U4615 (N_4615,N_4372,N_4377);
or U4616 (N_4616,N_4460,N_4346);
xor U4617 (N_4617,N_4461,N_4358);
or U4618 (N_4618,N_4343,N_4432);
xor U4619 (N_4619,N_4330,N_4418);
xor U4620 (N_4620,N_4430,N_4328);
nor U4621 (N_4621,N_4433,N_4430);
or U4622 (N_4622,N_4463,N_4373);
nand U4623 (N_4623,N_4380,N_4446);
nor U4624 (N_4624,N_4417,N_4344);
and U4625 (N_4625,N_4366,N_4380);
nor U4626 (N_4626,N_4404,N_4445);
nand U4627 (N_4627,N_4417,N_4369);
xnor U4628 (N_4628,N_4404,N_4476);
and U4629 (N_4629,N_4457,N_4361);
nand U4630 (N_4630,N_4446,N_4451);
nor U4631 (N_4631,N_4391,N_4363);
or U4632 (N_4632,N_4383,N_4398);
or U4633 (N_4633,N_4406,N_4346);
and U4634 (N_4634,N_4359,N_4332);
or U4635 (N_4635,N_4466,N_4348);
xnor U4636 (N_4636,N_4447,N_4394);
or U4637 (N_4637,N_4399,N_4395);
xnor U4638 (N_4638,N_4457,N_4455);
nor U4639 (N_4639,N_4426,N_4451);
nor U4640 (N_4640,N_4547,N_4639);
and U4641 (N_4641,N_4582,N_4631);
or U4642 (N_4642,N_4554,N_4617);
nand U4643 (N_4643,N_4605,N_4561);
xor U4644 (N_4644,N_4579,N_4533);
and U4645 (N_4645,N_4520,N_4516);
nand U4646 (N_4646,N_4552,N_4538);
or U4647 (N_4647,N_4513,N_4614);
nor U4648 (N_4648,N_4600,N_4522);
nand U4649 (N_4649,N_4498,N_4621);
and U4650 (N_4650,N_4595,N_4620);
nand U4651 (N_4651,N_4574,N_4573);
xnor U4652 (N_4652,N_4481,N_4637);
or U4653 (N_4653,N_4628,N_4511);
or U4654 (N_4654,N_4506,N_4613);
nor U4655 (N_4655,N_4603,N_4592);
nand U4656 (N_4656,N_4581,N_4590);
or U4657 (N_4657,N_4508,N_4524);
or U4658 (N_4658,N_4487,N_4504);
nand U4659 (N_4659,N_4505,N_4619);
or U4660 (N_4660,N_4594,N_4517);
nor U4661 (N_4661,N_4486,N_4583);
or U4662 (N_4662,N_4612,N_4559);
and U4663 (N_4663,N_4503,N_4586);
nand U4664 (N_4664,N_4591,N_4537);
nor U4665 (N_4665,N_4609,N_4615);
nor U4666 (N_4666,N_4575,N_4518);
and U4667 (N_4667,N_4497,N_4555);
nor U4668 (N_4668,N_4560,N_4512);
and U4669 (N_4669,N_4489,N_4588);
or U4670 (N_4670,N_4550,N_4568);
and U4671 (N_4671,N_4601,N_4584);
nand U4672 (N_4672,N_4545,N_4526);
and U4673 (N_4673,N_4523,N_4565);
nor U4674 (N_4674,N_4585,N_4548);
and U4675 (N_4675,N_4540,N_4627);
and U4676 (N_4676,N_4490,N_4536);
nand U4677 (N_4677,N_4485,N_4598);
nor U4678 (N_4678,N_4571,N_4535);
nor U4679 (N_4679,N_4567,N_4578);
xnor U4680 (N_4680,N_4521,N_4558);
and U4681 (N_4681,N_4610,N_4563);
xor U4682 (N_4682,N_4564,N_4514);
nand U4683 (N_4683,N_4624,N_4556);
xor U4684 (N_4684,N_4569,N_4611);
or U4685 (N_4685,N_4562,N_4492);
nand U4686 (N_4686,N_4551,N_4572);
and U4687 (N_4687,N_4634,N_4606);
xor U4688 (N_4688,N_4488,N_4608);
and U4689 (N_4689,N_4502,N_4553);
nor U4690 (N_4690,N_4597,N_4638);
or U4691 (N_4691,N_4494,N_4480);
nor U4692 (N_4692,N_4530,N_4529);
nand U4693 (N_4693,N_4629,N_4499);
or U4694 (N_4694,N_4630,N_4618);
or U4695 (N_4695,N_4576,N_4607);
nand U4696 (N_4696,N_4566,N_4636);
xor U4697 (N_4697,N_4483,N_4577);
and U4698 (N_4698,N_4635,N_4507);
xnor U4699 (N_4699,N_4542,N_4549);
nand U4700 (N_4700,N_4633,N_4599);
nor U4701 (N_4701,N_4509,N_4510);
or U4702 (N_4702,N_4625,N_4589);
xnor U4703 (N_4703,N_4501,N_4534);
nand U4704 (N_4704,N_4616,N_4580);
nor U4705 (N_4705,N_4626,N_4484);
or U4706 (N_4706,N_4532,N_4557);
or U4707 (N_4707,N_4544,N_4519);
xnor U4708 (N_4708,N_4528,N_4632);
and U4709 (N_4709,N_4539,N_4593);
nand U4710 (N_4710,N_4527,N_4541);
or U4711 (N_4711,N_4500,N_4496);
or U4712 (N_4712,N_4515,N_4623);
xor U4713 (N_4713,N_4602,N_4482);
nor U4714 (N_4714,N_4604,N_4570);
nand U4715 (N_4715,N_4531,N_4543);
xnor U4716 (N_4716,N_4495,N_4491);
nand U4717 (N_4717,N_4546,N_4525);
nor U4718 (N_4718,N_4587,N_4622);
and U4719 (N_4719,N_4493,N_4596);
nand U4720 (N_4720,N_4542,N_4521);
or U4721 (N_4721,N_4571,N_4544);
xnor U4722 (N_4722,N_4480,N_4495);
nand U4723 (N_4723,N_4547,N_4509);
nand U4724 (N_4724,N_4632,N_4562);
or U4725 (N_4725,N_4515,N_4513);
or U4726 (N_4726,N_4486,N_4563);
xnor U4727 (N_4727,N_4547,N_4607);
nand U4728 (N_4728,N_4609,N_4563);
or U4729 (N_4729,N_4566,N_4539);
or U4730 (N_4730,N_4578,N_4618);
or U4731 (N_4731,N_4628,N_4590);
and U4732 (N_4732,N_4561,N_4589);
nand U4733 (N_4733,N_4550,N_4558);
nand U4734 (N_4734,N_4503,N_4594);
or U4735 (N_4735,N_4597,N_4494);
and U4736 (N_4736,N_4506,N_4502);
or U4737 (N_4737,N_4637,N_4544);
and U4738 (N_4738,N_4614,N_4624);
nand U4739 (N_4739,N_4484,N_4504);
or U4740 (N_4740,N_4494,N_4516);
nor U4741 (N_4741,N_4624,N_4512);
nor U4742 (N_4742,N_4616,N_4557);
nor U4743 (N_4743,N_4586,N_4528);
nor U4744 (N_4744,N_4622,N_4507);
nand U4745 (N_4745,N_4507,N_4579);
and U4746 (N_4746,N_4568,N_4535);
nand U4747 (N_4747,N_4535,N_4574);
and U4748 (N_4748,N_4586,N_4571);
nor U4749 (N_4749,N_4612,N_4637);
nor U4750 (N_4750,N_4581,N_4607);
nor U4751 (N_4751,N_4606,N_4628);
nor U4752 (N_4752,N_4557,N_4486);
and U4753 (N_4753,N_4532,N_4606);
xor U4754 (N_4754,N_4613,N_4513);
and U4755 (N_4755,N_4562,N_4513);
nand U4756 (N_4756,N_4620,N_4585);
xor U4757 (N_4757,N_4525,N_4520);
or U4758 (N_4758,N_4633,N_4515);
xor U4759 (N_4759,N_4628,N_4595);
nor U4760 (N_4760,N_4501,N_4530);
nor U4761 (N_4761,N_4511,N_4637);
nor U4762 (N_4762,N_4582,N_4513);
xnor U4763 (N_4763,N_4567,N_4535);
nor U4764 (N_4764,N_4523,N_4592);
nor U4765 (N_4765,N_4540,N_4485);
nand U4766 (N_4766,N_4484,N_4603);
or U4767 (N_4767,N_4608,N_4627);
xnor U4768 (N_4768,N_4529,N_4568);
xnor U4769 (N_4769,N_4605,N_4545);
and U4770 (N_4770,N_4615,N_4600);
and U4771 (N_4771,N_4566,N_4531);
or U4772 (N_4772,N_4612,N_4510);
xnor U4773 (N_4773,N_4498,N_4515);
xnor U4774 (N_4774,N_4637,N_4518);
and U4775 (N_4775,N_4559,N_4563);
xor U4776 (N_4776,N_4485,N_4530);
and U4777 (N_4777,N_4553,N_4526);
nor U4778 (N_4778,N_4538,N_4519);
xnor U4779 (N_4779,N_4617,N_4592);
nand U4780 (N_4780,N_4547,N_4631);
or U4781 (N_4781,N_4631,N_4615);
nand U4782 (N_4782,N_4507,N_4489);
and U4783 (N_4783,N_4496,N_4552);
nand U4784 (N_4784,N_4500,N_4628);
xnor U4785 (N_4785,N_4533,N_4566);
or U4786 (N_4786,N_4626,N_4611);
or U4787 (N_4787,N_4560,N_4491);
or U4788 (N_4788,N_4546,N_4578);
nor U4789 (N_4789,N_4507,N_4629);
or U4790 (N_4790,N_4552,N_4635);
nor U4791 (N_4791,N_4533,N_4518);
and U4792 (N_4792,N_4501,N_4546);
nand U4793 (N_4793,N_4524,N_4591);
nand U4794 (N_4794,N_4590,N_4539);
xor U4795 (N_4795,N_4526,N_4635);
xnor U4796 (N_4796,N_4586,N_4537);
xnor U4797 (N_4797,N_4625,N_4592);
nand U4798 (N_4798,N_4582,N_4571);
nor U4799 (N_4799,N_4637,N_4507);
xnor U4800 (N_4800,N_4688,N_4725);
or U4801 (N_4801,N_4647,N_4643);
nor U4802 (N_4802,N_4739,N_4655);
or U4803 (N_4803,N_4715,N_4780);
xnor U4804 (N_4804,N_4767,N_4758);
and U4805 (N_4805,N_4673,N_4703);
and U4806 (N_4806,N_4734,N_4705);
nand U4807 (N_4807,N_4662,N_4669);
nand U4808 (N_4808,N_4752,N_4663);
nor U4809 (N_4809,N_4747,N_4763);
xor U4810 (N_4810,N_4671,N_4736);
xnor U4811 (N_4811,N_4754,N_4790);
nor U4812 (N_4812,N_4724,N_4666);
and U4813 (N_4813,N_4727,N_4690);
nand U4814 (N_4814,N_4784,N_4730);
nor U4815 (N_4815,N_4696,N_4676);
or U4816 (N_4816,N_4685,N_4711);
or U4817 (N_4817,N_4645,N_4772);
and U4818 (N_4818,N_4674,N_4698);
or U4819 (N_4819,N_4721,N_4659);
nand U4820 (N_4820,N_4794,N_4708);
and U4821 (N_4821,N_4755,N_4644);
nor U4822 (N_4822,N_4686,N_4665);
nor U4823 (N_4823,N_4760,N_4661);
nand U4824 (N_4824,N_4751,N_4651);
nor U4825 (N_4825,N_4774,N_4793);
or U4826 (N_4826,N_4726,N_4710);
nand U4827 (N_4827,N_4749,N_4672);
or U4828 (N_4828,N_4741,N_4687);
xnor U4829 (N_4829,N_4795,N_4709);
xnor U4830 (N_4830,N_4762,N_4742);
nor U4831 (N_4831,N_4712,N_4664);
nand U4832 (N_4832,N_4720,N_4729);
xor U4833 (N_4833,N_4768,N_4646);
nor U4834 (N_4834,N_4733,N_4798);
xor U4835 (N_4835,N_4702,N_4738);
nor U4836 (N_4836,N_4693,N_4700);
or U4837 (N_4837,N_4719,N_4797);
nor U4838 (N_4838,N_4704,N_4783);
or U4839 (N_4839,N_4746,N_4640);
nor U4840 (N_4840,N_4678,N_4650);
and U4841 (N_4841,N_4680,N_4670);
or U4842 (N_4842,N_4771,N_4737);
nor U4843 (N_4843,N_4691,N_4744);
and U4844 (N_4844,N_4679,N_4789);
nor U4845 (N_4845,N_4775,N_4735);
nor U4846 (N_4846,N_4718,N_4778);
nor U4847 (N_4847,N_4759,N_4682);
and U4848 (N_4848,N_4648,N_4731);
xnor U4849 (N_4849,N_4799,N_4779);
nand U4850 (N_4850,N_4695,N_4785);
or U4851 (N_4851,N_4641,N_4667);
or U4852 (N_4852,N_4722,N_4786);
or U4853 (N_4853,N_4753,N_4743);
nor U4854 (N_4854,N_4732,N_4713);
xor U4855 (N_4855,N_4728,N_4697);
nor U4856 (N_4856,N_4781,N_4764);
nor U4857 (N_4857,N_4756,N_4675);
nor U4858 (N_4858,N_4692,N_4765);
and U4859 (N_4859,N_4681,N_4654);
nor U4860 (N_4860,N_4694,N_4660);
nor U4861 (N_4861,N_4714,N_4748);
nor U4862 (N_4862,N_4788,N_4657);
nand U4863 (N_4863,N_4750,N_4653);
nor U4864 (N_4864,N_4656,N_4745);
or U4865 (N_4865,N_4787,N_4707);
nand U4866 (N_4866,N_4689,N_4683);
nor U4867 (N_4867,N_4642,N_4677);
nor U4868 (N_4868,N_4770,N_4769);
xor U4869 (N_4869,N_4796,N_4684);
xor U4870 (N_4870,N_4723,N_4777);
and U4871 (N_4871,N_4701,N_4766);
nand U4872 (N_4872,N_4761,N_4792);
nand U4873 (N_4873,N_4740,N_4658);
and U4874 (N_4874,N_4717,N_4699);
and U4875 (N_4875,N_4716,N_4791);
nor U4876 (N_4876,N_4652,N_4649);
xor U4877 (N_4877,N_4757,N_4668);
nor U4878 (N_4878,N_4782,N_4776);
nand U4879 (N_4879,N_4773,N_4706);
nor U4880 (N_4880,N_4789,N_4662);
and U4881 (N_4881,N_4702,N_4706);
nand U4882 (N_4882,N_4684,N_4719);
and U4883 (N_4883,N_4674,N_4775);
nor U4884 (N_4884,N_4746,N_4698);
nand U4885 (N_4885,N_4784,N_4790);
nor U4886 (N_4886,N_4674,N_4778);
and U4887 (N_4887,N_4682,N_4700);
or U4888 (N_4888,N_4695,N_4716);
or U4889 (N_4889,N_4704,N_4782);
xnor U4890 (N_4890,N_4732,N_4731);
nor U4891 (N_4891,N_4720,N_4717);
xor U4892 (N_4892,N_4689,N_4788);
and U4893 (N_4893,N_4672,N_4702);
and U4894 (N_4894,N_4710,N_4760);
xnor U4895 (N_4895,N_4755,N_4777);
nor U4896 (N_4896,N_4710,N_4776);
nand U4897 (N_4897,N_4725,N_4655);
nor U4898 (N_4898,N_4766,N_4774);
nand U4899 (N_4899,N_4709,N_4718);
nor U4900 (N_4900,N_4727,N_4660);
xor U4901 (N_4901,N_4715,N_4777);
nor U4902 (N_4902,N_4672,N_4736);
or U4903 (N_4903,N_4687,N_4790);
nor U4904 (N_4904,N_4714,N_4709);
or U4905 (N_4905,N_4783,N_4752);
and U4906 (N_4906,N_4653,N_4646);
nor U4907 (N_4907,N_4655,N_4768);
or U4908 (N_4908,N_4689,N_4640);
xor U4909 (N_4909,N_4738,N_4765);
xnor U4910 (N_4910,N_4675,N_4703);
and U4911 (N_4911,N_4691,N_4699);
xor U4912 (N_4912,N_4669,N_4794);
xor U4913 (N_4913,N_4752,N_4737);
and U4914 (N_4914,N_4778,N_4689);
nor U4915 (N_4915,N_4766,N_4661);
and U4916 (N_4916,N_4713,N_4741);
nor U4917 (N_4917,N_4671,N_4692);
nor U4918 (N_4918,N_4705,N_4777);
or U4919 (N_4919,N_4728,N_4659);
and U4920 (N_4920,N_4756,N_4667);
or U4921 (N_4921,N_4718,N_4657);
and U4922 (N_4922,N_4692,N_4781);
xnor U4923 (N_4923,N_4686,N_4670);
nor U4924 (N_4924,N_4725,N_4768);
nor U4925 (N_4925,N_4703,N_4658);
and U4926 (N_4926,N_4656,N_4688);
nand U4927 (N_4927,N_4769,N_4644);
nor U4928 (N_4928,N_4782,N_4733);
and U4929 (N_4929,N_4709,N_4759);
nand U4930 (N_4930,N_4686,N_4694);
nand U4931 (N_4931,N_4772,N_4747);
nor U4932 (N_4932,N_4703,N_4727);
nor U4933 (N_4933,N_4650,N_4709);
nand U4934 (N_4934,N_4653,N_4672);
nand U4935 (N_4935,N_4750,N_4640);
xnor U4936 (N_4936,N_4657,N_4770);
nand U4937 (N_4937,N_4760,N_4642);
or U4938 (N_4938,N_4773,N_4686);
or U4939 (N_4939,N_4681,N_4725);
and U4940 (N_4940,N_4672,N_4769);
and U4941 (N_4941,N_4745,N_4703);
xor U4942 (N_4942,N_4656,N_4647);
or U4943 (N_4943,N_4734,N_4686);
xor U4944 (N_4944,N_4764,N_4763);
and U4945 (N_4945,N_4642,N_4764);
or U4946 (N_4946,N_4787,N_4692);
nand U4947 (N_4947,N_4760,N_4781);
nand U4948 (N_4948,N_4764,N_4690);
nor U4949 (N_4949,N_4684,N_4739);
nand U4950 (N_4950,N_4707,N_4738);
xnor U4951 (N_4951,N_4651,N_4739);
nand U4952 (N_4952,N_4757,N_4644);
xnor U4953 (N_4953,N_4687,N_4732);
nor U4954 (N_4954,N_4699,N_4641);
and U4955 (N_4955,N_4709,N_4796);
and U4956 (N_4956,N_4655,N_4670);
or U4957 (N_4957,N_4742,N_4651);
nor U4958 (N_4958,N_4727,N_4699);
xnor U4959 (N_4959,N_4657,N_4645);
and U4960 (N_4960,N_4839,N_4915);
and U4961 (N_4961,N_4892,N_4802);
or U4962 (N_4962,N_4930,N_4810);
or U4963 (N_4963,N_4908,N_4854);
and U4964 (N_4964,N_4806,N_4817);
nand U4965 (N_4965,N_4847,N_4832);
xnor U4966 (N_4966,N_4920,N_4828);
nor U4967 (N_4967,N_4922,N_4870);
nor U4968 (N_4968,N_4884,N_4891);
or U4969 (N_4969,N_4871,N_4883);
or U4970 (N_4970,N_4852,N_4835);
xnor U4971 (N_4971,N_4815,N_4935);
or U4972 (N_4972,N_4803,N_4917);
and U4973 (N_4973,N_4913,N_4840);
and U4974 (N_4974,N_4931,N_4939);
or U4975 (N_4975,N_4907,N_4896);
xor U4976 (N_4976,N_4946,N_4910);
xnor U4977 (N_4977,N_4925,N_4887);
xor U4978 (N_4978,N_4843,N_4873);
and U4979 (N_4979,N_4842,N_4865);
xor U4980 (N_4980,N_4914,N_4808);
nand U4981 (N_4981,N_4837,N_4900);
nor U4982 (N_4982,N_4918,N_4876);
and U4983 (N_4983,N_4814,N_4841);
nand U4984 (N_4984,N_4895,N_4947);
or U4985 (N_4985,N_4937,N_4813);
and U4986 (N_4986,N_4912,N_4861);
nor U4987 (N_4987,N_4903,N_4956);
xnor U4988 (N_4988,N_4822,N_4889);
or U4989 (N_4989,N_4899,N_4885);
nor U4990 (N_4990,N_4825,N_4949);
or U4991 (N_4991,N_4958,N_4834);
nor U4992 (N_4992,N_4936,N_4853);
nor U4993 (N_4993,N_4845,N_4909);
and U4994 (N_4994,N_4880,N_4878);
or U4995 (N_4995,N_4857,N_4951);
xor U4996 (N_4996,N_4906,N_4872);
and U4997 (N_4997,N_4924,N_4945);
and U4998 (N_4998,N_4863,N_4805);
or U4999 (N_4999,N_4849,N_4816);
nor U5000 (N_5000,N_4938,N_4905);
nand U5001 (N_5001,N_4933,N_4953);
nor U5002 (N_5002,N_4859,N_4846);
and U5003 (N_5003,N_4955,N_4902);
xor U5004 (N_5004,N_4940,N_4862);
nand U5005 (N_5005,N_4819,N_4901);
xnor U5006 (N_5006,N_4886,N_4893);
and U5007 (N_5007,N_4875,N_4897);
and U5008 (N_5008,N_4833,N_4809);
nor U5009 (N_5009,N_4820,N_4919);
nand U5010 (N_5010,N_4868,N_4874);
xor U5011 (N_5011,N_4830,N_4812);
or U5012 (N_5012,N_4890,N_4954);
nor U5013 (N_5013,N_4911,N_4826);
nor U5014 (N_5014,N_4927,N_4877);
nand U5015 (N_5015,N_4836,N_4821);
xor U5016 (N_5016,N_4818,N_4898);
or U5017 (N_5017,N_4801,N_4869);
xnor U5018 (N_5018,N_4867,N_4844);
or U5019 (N_5019,N_4824,N_4838);
nor U5020 (N_5020,N_4948,N_4864);
and U5021 (N_5021,N_4941,N_4904);
nor U5022 (N_5022,N_4823,N_4950);
xor U5023 (N_5023,N_4916,N_4921);
nor U5024 (N_5024,N_4943,N_4804);
or U5025 (N_5025,N_4860,N_4952);
xor U5026 (N_5026,N_4858,N_4894);
nor U5027 (N_5027,N_4881,N_4811);
nand U5028 (N_5028,N_4829,N_4855);
nor U5029 (N_5029,N_4928,N_4929);
or U5030 (N_5030,N_4866,N_4848);
nand U5031 (N_5031,N_4800,N_4851);
xor U5032 (N_5032,N_4831,N_4944);
xnor U5033 (N_5033,N_4827,N_4888);
or U5034 (N_5034,N_4942,N_4850);
nand U5035 (N_5035,N_4959,N_4856);
xnor U5036 (N_5036,N_4807,N_4957);
and U5037 (N_5037,N_4926,N_4934);
nor U5038 (N_5038,N_4882,N_4879);
nand U5039 (N_5039,N_4923,N_4932);
xor U5040 (N_5040,N_4826,N_4852);
nand U5041 (N_5041,N_4810,N_4832);
nand U5042 (N_5042,N_4868,N_4837);
and U5043 (N_5043,N_4932,N_4942);
xor U5044 (N_5044,N_4908,N_4871);
nand U5045 (N_5045,N_4932,N_4853);
or U5046 (N_5046,N_4835,N_4802);
or U5047 (N_5047,N_4804,N_4896);
or U5048 (N_5048,N_4864,N_4876);
and U5049 (N_5049,N_4865,N_4944);
nor U5050 (N_5050,N_4898,N_4938);
nor U5051 (N_5051,N_4840,N_4923);
nand U5052 (N_5052,N_4902,N_4922);
xnor U5053 (N_5053,N_4843,N_4807);
or U5054 (N_5054,N_4824,N_4831);
or U5055 (N_5055,N_4959,N_4894);
nand U5056 (N_5056,N_4853,N_4911);
xnor U5057 (N_5057,N_4848,N_4858);
xnor U5058 (N_5058,N_4804,N_4899);
nor U5059 (N_5059,N_4952,N_4825);
nand U5060 (N_5060,N_4956,N_4857);
xor U5061 (N_5061,N_4876,N_4848);
nand U5062 (N_5062,N_4893,N_4840);
nand U5063 (N_5063,N_4927,N_4846);
nor U5064 (N_5064,N_4843,N_4919);
xnor U5065 (N_5065,N_4864,N_4923);
or U5066 (N_5066,N_4886,N_4937);
nor U5067 (N_5067,N_4810,N_4856);
and U5068 (N_5068,N_4842,N_4837);
nand U5069 (N_5069,N_4915,N_4876);
and U5070 (N_5070,N_4848,N_4807);
nand U5071 (N_5071,N_4866,N_4867);
nor U5072 (N_5072,N_4868,N_4877);
nand U5073 (N_5073,N_4806,N_4814);
xnor U5074 (N_5074,N_4823,N_4864);
nand U5075 (N_5075,N_4957,N_4872);
and U5076 (N_5076,N_4939,N_4904);
nor U5077 (N_5077,N_4867,N_4927);
or U5078 (N_5078,N_4879,N_4922);
or U5079 (N_5079,N_4857,N_4821);
xor U5080 (N_5080,N_4809,N_4896);
and U5081 (N_5081,N_4931,N_4947);
nor U5082 (N_5082,N_4844,N_4814);
and U5083 (N_5083,N_4890,N_4948);
or U5084 (N_5084,N_4941,N_4882);
xor U5085 (N_5085,N_4813,N_4858);
xor U5086 (N_5086,N_4959,N_4858);
xnor U5087 (N_5087,N_4850,N_4802);
nand U5088 (N_5088,N_4818,N_4857);
nor U5089 (N_5089,N_4858,N_4924);
or U5090 (N_5090,N_4822,N_4934);
nor U5091 (N_5091,N_4838,N_4813);
or U5092 (N_5092,N_4928,N_4888);
and U5093 (N_5093,N_4831,N_4871);
nand U5094 (N_5094,N_4941,N_4893);
nor U5095 (N_5095,N_4812,N_4822);
nand U5096 (N_5096,N_4874,N_4955);
nor U5097 (N_5097,N_4814,N_4875);
nor U5098 (N_5098,N_4858,N_4871);
and U5099 (N_5099,N_4831,N_4862);
xnor U5100 (N_5100,N_4837,N_4830);
nor U5101 (N_5101,N_4808,N_4917);
xor U5102 (N_5102,N_4853,N_4897);
and U5103 (N_5103,N_4861,N_4848);
or U5104 (N_5104,N_4914,N_4910);
nor U5105 (N_5105,N_4959,N_4814);
or U5106 (N_5106,N_4939,N_4956);
xor U5107 (N_5107,N_4904,N_4871);
nand U5108 (N_5108,N_4903,N_4846);
nand U5109 (N_5109,N_4895,N_4932);
nor U5110 (N_5110,N_4832,N_4898);
nand U5111 (N_5111,N_4859,N_4883);
xnor U5112 (N_5112,N_4936,N_4821);
nor U5113 (N_5113,N_4881,N_4839);
nor U5114 (N_5114,N_4884,N_4938);
nand U5115 (N_5115,N_4941,N_4846);
nand U5116 (N_5116,N_4841,N_4907);
xor U5117 (N_5117,N_4818,N_4868);
nor U5118 (N_5118,N_4820,N_4902);
nand U5119 (N_5119,N_4855,N_4892);
and U5120 (N_5120,N_5048,N_5019);
xnor U5121 (N_5121,N_5026,N_4967);
nand U5122 (N_5122,N_5111,N_5071);
and U5123 (N_5123,N_5015,N_5009);
nand U5124 (N_5124,N_5023,N_5104);
nand U5125 (N_5125,N_4994,N_4970);
nand U5126 (N_5126,N_5018,N_5010);
nand U5127 (N_5127,N_5068,N_5058);
xor U5128 (N_5128,N_5053,N_4964);
or U5129 (N_5129,N_4974,N_5105);
xor U5130 (N_5130,N_5092,N_5093);
nor U5131 (N_5131,N_5021,N_4987);
nand U5132 (N_5132,N_5038,N_5001);
or U5133 (N_5133,N_4984,N_5036);
nand U5134 (N_5134,N_5106,N_5103);
and U5135 (N_5135,N_4996,N_5011);
nor U5136 (N_5136,N_5114,N_5096);
xnor U5137 (N_5137,N_5099,N_4992);
and U5138 (N_5138,N_5008,N_5109);
or U5139 (N_5139,N_5069,N_5100);
and U5140 (N_5140,N_5032,N_5037);
and U5141 (N_5141,N_4961,N_5003);
xnor U5142 (N_5142,N_5033,N_5049);
and U5143 (N_5143,N_5073,N_5085);
nand U5144 (N_5144,N_5004,N_5075);
and U5145 (N_5145,N_5091,N_5112);
nand U5146 (N_5146,N_5059,N_4976);
nor U5147 (N_5147,N_4978,N_5056);
nor U5148 (N_5148,N_4997,N_4983);
nand U5149 (N_5149,N_5086,N_5046);
or U5150 (N_5150,N_4973,N_5024);
nor U5151 (N_5151,N_5110,N_5060);
and U5152 (N_5152,N_4993,N_5084);
nand U5153 (N_5153,N_5057,N_5094);
and U5154 (N_5154,N_4966,N_5020);
nor U5155 (N_5155,N_4968,N_5012);
nand U5156 (N_5156,N_5067,N_5113);
xnor U5157 (N_5157,N_5042,N_5051);
xor U5158 (N_5158,N_5050,N_5089);
and U5159 (N_5159,N_5062,N_5014);
and U5160 (N_5160,N_5115,N_4982);
and U5161 (N_5161,N_5063,N_4975);
nor U5162 (N_5162,N_4969,N_5101);
and U5163 (N_5163,N_5076,N_5066);
or U5164 (N_5164,N_5030,N_5077);
nand U5165 (N_5165,N_4971,N_5095);
or U5166 (N_5166,N_5064,N_5088);
xnor U5167 (N_5167,N_4960,N_5043);
nand U5168 (N_5168,N_5102,N_5098);
xnor U5169 (N_5169,N_5025,N_5029);
or U5170 (N_5170,N_4986,N_5107);
or U5171 (N_5171,N_4963,N_4972);
xnor U5172 (N_5172,N_5000,N_5087);
nor U5173 (N_5173,N_5047,N_5054);
nor U5174 (N_5174,N_5119,N_5039);
and U5175 (N_5175,N_5080,N_5072);
or U5176 (N_5176,N_5005,N_5016);
xnor U5177 (N_5177,N_5006,N_5013);
xnor U5178 (N_5178,N_4988,N_5081);
or U5179 (N_5179,N_5074,N_5065);
or U5180 (N_5180,N_4995,N_5035);
and U5181 (N_5181,N_5017,N_5083);
or U5182 (N_5182,N_5044,N_4999);
nand U5183 (N_5183,N_5034,N_5079);
or U5184 (N_5184,N_4991,N_5040);
nor U5185 (N_5185,N_5108,N_5028);
xor U5186 (N_5186,N_5045,N_5061);
xor U5187 (N_5187,N_5041,N_5052);
or U5188 (N_5188,N_5082,N_4980);
xor U5189 (N_5189,N_5055,N_5117);
nand U5190 (N_5190,N_4989,N_5116);
or U5191 (N_5191,N_5031,N_5118);
or U5192 (N_5192,N_4977,N_4985);
or U5193 (N_5193,N_4981,N_5002);
or U5194 (N_5194,N_5078,N_4965);
and U5195 (N_5195,N_4979,N_5022);
nand U5196 (N_5196,N_5070,N_5097);
nor U5197 (N_5197,N_5027,N_5007);
xnor U5198 (N_5198,N_4962,N_4990);
nand U5199 (N_5199,N_5090,N_4998);
nand U5200 (N_5200,N_5036,N_5046);
and U5201 (N_5201,N_4997,N_4989);
nand U5202 (N_5202,N_4967,N_5078);
nor U5203 (N_5203,N_5029,N_4972);
or U5204 (N_5204,N_5036,N_5019);
and U5205 (N_5205,N_5011,N_5115);
nor U5206 (N_5206,N_4992,N_5033);
xnor U5207 (N_5207,N_5046,N_5112);
nand U5208 (N_5208,N_5031,N_5010);
nand U5209 (N_5209,N_5032,N_5006);
xnor U5210 (N_5210,N_4961,N_4973);
xor U5211 (N_5211,N_4975,N_4973);
nand U5212 (N_5212,N_4978,N_4984);
nand U5213 (N_5213,N_5018,N_4962);
xor U5214 (N_5214,N_5099,N_4961);
or U5215 (N_5215,N_5075,N_5006);
and U5216 (N_5216,N_5056,N_5066);
nand U5217 (N_5217,N_5040,N_5041);
or U5218 (N_5218,N_5009,N_5005);
and U5219 (N_5219,N_5085,N_5045);
nand U5220 (N_5220,N_5031,N_5075);
or U5221 (N_5221,N_5037,N_4969);
and U5222 (N_5222,N_5105,N_5115);
nand U5223 (N_5223,N_4962,N_5073);
or U5224 (N_5224,N_5026,N_5045);
and U5225 (N_5225,N_5062,N_5080);
nand U5226 (N_5226,N_4964,N_5110);
or U5227 (N_5227,N_4976,N_5058);
xor U5228 (N_5228,N_4997,N_5024);
xor U5229 (N_5229,N_5039,N_4997);
and U5230 (N_5230,N_5035,N_5004);
or U5231 (N_5231,N_4995,N_5008);
nand U5232 (N_5232,N_5046,N_5099);
and U5233 (N_5233,N_5117,N_5059);
nand U5234 (N_5234,N_5035,N_5010);
nand U5235 (N_5235,N_5036,N_5045);
nor U5236 (N_5236,N_4999,N_5096);
xor U5237 (N_5237,N_5066,N_5108);
nor U5238 (N_5238,N_4988,N_5110);
nor U5239 (N_5239,N_5108,N_4986);
and U5240 (N_5240,N_5088,N_5018);
nand U5241 (N_5241,N_5104,N_4980);
xor U5242 (N_5242,N_5004,N_4998);
or U5243 (N_5243,N_5097,N_5025);
nand U5244 (N_5244,N_5057,N_4997);
xnor U5245 (N_5245,N_5090,N_5071);
xnor U5246 (N_5246,N_5097,N_4999);
nor U5247 (N_5247,N_5070,N_5065);
nor U5248 (N_5248,N_5008,N_5099);
or U5249 (N_5249,N_5110,N_5080);
nand U5250 (N_5250,N_5088,N_5004);
or U5251 (N_5251,N_5109,N_5061);
xnor U5252 (N_5252,N_4973,N_5081);
or U5253 (N_5253,N_5017,N_4976);
or U5254 (N_5254,N_5091,N_5107);
nand U5255 (N_5255,N_5098,N_4998);
and U5256 (N_5256,N_5068,N_5024);
nor U5257 (N_5257,N_5066,N_5055);
and U5258 (N_5258,N_4991,N_5083);
xnor U5259 (N_5259,N_5067,N_4971);
or U5260 (N_5260,N_5115,N_5047);
or U5261 (N_5261,N_5081,N_4981);
xnor U5262 (N_5262,N_4965,N_4995);
or U5263 (N_5263,N_5089,N_4982);
nor U5264 (N_5264,N_5068,N_5041);
xor U5265 (N_5265,N_4987,N_4975);
xor U5266 (N_5266,N_5069,N_5045);
xnor U5267 (N_5267,N_4991,N_5057);
and U5268 (N_5268,N_5114,N_5050);
or U5269 (N_5269,N_4971,N_4978);
nor U5270 (N_5270,N_4966,N_5106);
or U5271 (N_5271,N_5047,N_5073);
or U5272 (N_5272,N_4974,N_5074);
and U5273 (N_5273,N_4972,N_5059);
xnor U5274 (N_5274,N_4974,N_4987);
nor U5275 (N_5275,N_5025,N_4985);
xnor U5276 (N_5276,N_5012,N_4983);
and U5277 (N_5277,N_5004,N_5100);
nand U5278 (N_5278,N_4980,N_5027);
xor U5279 (N_5279,N_4973,N_4974);
nor U5280 (N_5280,N_5204,N_5164);
nand U5281 (N_5281,N_5225,N_5208);
xnor U5282 (N_5282,N_5128,N_5177);
xnor U5283 (N_5283,N_5277,N_5182);
nand U5284 (N_5284,N_5250,N_5137);
and U5285 (N_5285,N_5210,N_5162);
or U5286 (N_5286,N_5171,N_5256);
nor U5287 (N_5287,N_5197,N_5264);
nor U5288 (N_5288,N_5157,N_5235);
xnor U5289 (N_5289,N_5276,N_5165);
and U5290 (N_5290,N_5124,N_5255);
or U5291 (N_5291,N_5275,N_5237);
or U5292 (N_5292,N_5246,N_5192);
nand U5293 (N_5293,N_5163,N_5205);
xor U5294 (N_5294,N_5198,N_5254);
or U5295 (N_5295,N_5244,N_5174);
or U5296 (N_5296,N_5156,N_5155);
xnor U5297 (N_5297,N_5200,N_5209);
xor U5298 (N_5298,N_5233,N_5228);
nand U5299 (N_5299,N_5271,N_5258);
or U5300 (N_5300,N_5199,N_5261);
xor U5301 (N_5301,N_5146,N_5180);
nand U5302 (N_5302,N_5196,N_5147);
nor U5303 (N_5303,N_5168,N_5179);
nor U5304 (N_5304,N_5176,N_5234);
xnor U5305 (N_5305,N_5215,N_5266);
nand U5306 (N_5306,N_5273,N_5141);
or U5307 (N_5307,N_5207,N_5152);
or U5308 (N_5308,N_5133,N_5189);
or U5309 (N_5309,N_5251,N_5236);
and U5310 (N_5310,N_5263,N_5130);
or U5311 (N_5311,N_5178,N_5184);
or U5312 (N_5312,N_5181,N_5148);
and U5313 (N_5313,N_5153,N_5220);
xor U5314 (N_5314,N_5145,N_5249);
or U5315 (N_5315,N_5190,N_5227);
or U5316 (N_5316,N_5247,N_5239);
nand U5317 (N_5317,N_5195,N_5240);
nand U5318 (N_5318,N_5214,N_5169);
and U5319 (N_5319,N_5172,N_5127);
nand U5320 (N_5320,N_5166,N_5245);
nor U5321 (N_5321,N_5151,N_5229);
or U5322 (N_5322,N_5170,N_5238);
nand U5323 (N_5323,N_5121,N_5120);
nor U5324 (N_5324,N_5202,N_5191);
or U5325 (N_5325,N_5231,N_5134);
or U5326 (N_5326,N_5274,N_5125);
xnor U5327 (N_5327,N_5262,N_5252);
or U5328 (N_5328,N_5267,N_5243);
nor U5329 (N_5329,N_5126,N_5265);
xnor U5330 (N_5330,N_5257,N_5144);
xnor U5331 (N_5331,N_5224,N_5226);
and U5332 (N_5332,N_5136,N_5216);
nor U5333 (N_5333,N_5219,N_5158);
or U5334 (N_5334,N_5278,N_5212);
and U5335 (N_5335,N_5242,N_5135);
or U5336 (N_5336,N_5213,N_5272);
nand U5337 (N_5337,N_5173,N_5221);
xor U5338 (N_5338,N_5222,N_5188);
nand U5339 (N_5339,N_5183,N_5193);
and U5340 (N_5340,N_5260,N_5253);
xor U5341 (N_5341,N_5159,N_5232);
xnor U5342 (N_5342,N_5149,N_5270);
or U5343 (N_5343,N_5218,N_5138);
nor U5344 (N_5344,N_5201,N_5187);
nand U5345 (N_5345,N_5154,N_5132);
and U5346 (N_5346,N_5150,N_5167);
nand U5347 (N_5347,N_5185,N_5160);
nor U5348 (N_5348,N_5139,N_5131);
xnor U5349 (N_5349,N_5122,N_5268);
and U5350 (N_5350,N_5175,N_5279);
xnor U5351 (N_5351,N_5241,N_5129);
nand U5352 (N_5352,N_5186,N_5269);
and U5353 (N_5353,N_5123,N_5194);
nor U5354 (N_5354,N_5223,N_5143);
and U5355 (N_5355,N_5211,N_5142);
nor U5356 (N_5356,N_5217,N_5161);
xor U5357 (N_5357,N_5230,N_5203);
nor U5358 (N_5358,N_5248,N_5206);
xor U5359 (N_5359,N_5259,N_5140);
xnor U5360 (N_5360,N_5191,N_5264);
nor U5361 (N_5361,N_5158,N_5195);
nor U5362 (N_5362,N_5243,N_5175);
nor U5363 (N_5363,N_5125,N_5168);
xor U5364 (N_5364,N_5275,N_5151);
xor U5365 (N_5365,N_5226,N_5125);
and U5366 (N_5366,N_5274,N_5232);
nor U5367 (N_5367,N_5278,N_5204);
nand U5368 (N_5368,N_5139,N_5222);
xnor U5369 (N_5369,N_5250,N_5143);
and U5370 (N_5370,N_5261,N_5256);
or U5371 (N_5371,N_5256,N_5210);
and U5372 (N_5372,N_5192,N_5235);
or U5373 (N_5373,N_5202,N_5169);
and U5374 (N_5374,N_5139,N_5164);
xnor U5375 (N_5375,N_5140,N_5227);
or U5376 (N_5376,N_5154,N_5248);
and U5377 (N_5377,N_5231,N_5270);
and U5378 (N_5378,N_5127,N_5223);
nand U5379 (N_5379,N_5234,N_5208);
and U5380 (N_5380,N_5141,N_5266);
nor U5381 (N_5381,N_5217,N_5187);
nor U5382 (N_5382,N_5196,N_5197);
or U5383 (N_5383,N_5176,N_5154);
nand U5384 (N_5384,N_5180,N_5159);
nor U5385 (N_5385,N_5201,N_5124);
and U5386 (N_5386,N_5176,N_5188);
xnor U5387 (N_5387,N_5243,N_5165);
or U5388 (N_5388,N_5249,N_5174);
or U5389 (N_5389,N_5154,N_5235);
or U5390 (N_5390,N_5162,N_5232);
nor U5391 (N_5391,N_5163,N_5150);
nand U5392 (N_5392,N_5187,N_5153);
nor U5393 (N_5393,N_5237,N_5277);
or U5394 (N_5394,N_5239,N_5268);
and U5395 (N_5395,N_5278,N_5174);
nor U5396 (N_5396,N_5130,N_5129);
and U5397 (N_5397,N_5248,N_5277);
and U5398 (N_5398,N_5126,N_5247);
and U5399 (N_5399,N_5220,N_5157);
nand U5400 (N_5400,N_5162,N_5153);
and U5401 (N_5401,N_5270,N_5207);
and U5402 (N_5402,N_5180,N_5209);
nand U5403 (N_5403,N_5269,N_5223);
xor U5404 (N_5404,N_5206,N_5127);
nand U5405 (N_5405,N_5238,N_5243);
or U5406 (N_5406,N_5164,N_5132);
xnor U5407 (N_5407,N_5152,N_5131);
nand U5408 (N_5408,N_5148,N_5267);
nand U5409 (N_5409,N_5263,N_5121);
nor U5410 (N_5410,N_5203,N_5245);
and U5411 (N_5411,N_5170,N_5245);
and U5412 (N_5412,N_5274,N_5136);
nor U5413 (N_5413,N_5160,N_5141);
xnor U5414 (N_5414,N_5133,N_5126);
nor U5415 (N_5415,N_5211,N_5264);
nand U5416 (N_5416,N_5264,N_5199);
or U5417 (N_5417,N_5239,N_5278);
or U5418 (N_5418,N_5273,N_5231);
nand U5419 (N_5419,N_5181,N_5188);
nor U5420 (N_5420,N_5141,N_5129);
nor U5421 (N_5421,N_5142,N_5173);
and U5422 (N_5422,N_5148,N_5142);
xor U5423 (N_5423,N_5231,N_5129);
or U5424 (N_5424,N_5225,N_5174);
xor U5425 (N_5425,N_5143,N_5199);
or U5426 (N_5426,N_5158,N_5265);
nand U5427 (N_5427,N_5126,N_5207);
and U5428 (N_5428,N_5134,N_5123);
nand U5429 (N_5429,N_5132,N_5231);
nor U5430 (N_5430,N_5141,N_5151);
and U5431 (N_5431,N_5136,N_5212);
nand U5432 (N_5432,N_5130,N_5139);
or U5433 (N_5433,N_5141,N_5261);
and U5434 (N_5434,N_5135,N_5160);
or U5435 (N_5435,N_5180,N_5137);
nor U5436 (N_5436,N_5127,N_5160);
nand U5437 (N_5437,N_5279,N_5209);
xnor U5438 (N_5438,N_5126,N_5166);
and U5439 (N_5439,N_5279,N_5217);
or U5440 (N_5440,N_5291,N_5386);
nand U5441 (N_5441,N_5329,N_5416);
xor U5442 (N_5442,N_5419,N_5427);
and U5443 (N_5443,N_5305,N_5353);
nor U5444 (N_5444,N_5421,N_5319);
nand U5445 (N_5445,N_5412,N_5381);
and U5446 (N_5446,N_5299,N_5298);
or U5447 (N_5447,N_5339,N_5293);
nand U5448 (N_5448,N_5360,N_5334);
nor U5449 (N_5449,N_5436,N_5284);
xnor U5450 (N_5450,N_5430,N_5428);
or U5451 (N_5451,N_5313,N_5337);
and U5452 (N_5452,N_5324,N_5340);
or U5453 (N_5453,N_5431,N_5415);
and U5454 (N_5454,N_5434,N_5349);
xor U5455 (N_5455,N_5378,N_5287);
nor U5456 (N_5456,N_5406,N_5343);
and U5457 (N_5457,N_5317,N_5388);
nor U5458 (N_5458,N_5344,N_5368);
nand U5459 (N_5459,N_5425,N_5411);
nand U5460 (N_5460,N_5373,N_5303);
xor U5461 (N_5461,N_5438,N_5312);
and U5462 (N_5462,N_5409,N_5366);
nand U5463 (N_5463,N_5379,N_5357);
nor U5464 (N_5464,N_5375,N_5398);
and U5465 (N_5465,N_5374,N_5304);
xnor U5466 (N_5466,N_5332,N_5403);
and U5467 (N_5467,N_5439,N_5320);
nand U5468 (N_5468,N_5323,N_5365);
nand U5469 (N_5469,N_5370,N_5372);
or U5470 (N_5470,N_5437,N_5422);
xnor U5471 (N_5471,N_5338,N_5396);
or U5472 (N_5472,N_5347,N_5367);
or U5473 (N_5473,N_5399,N_5327);
or U5474 (N_5474,N_5432,N_5296);
nand U5475 (N_5475,N_5389,N_5341);
xor U5476 (N_5476,N_5363,N_5325);
xnor U5477 (N_5477,N_5306,N_5376);
and U5478 (N_5478,N_5395,N_5391);
nor U5479 (N_5479,N_5429,N_5336);
or U5480 (N_5480,N_5310,N_5316);
nand U5481 (N_5481,N_5286,N_5280);
nor U5482 (N_5482,N_5387,N_5394);
nor U5483 (N_5483,N_5435,N_5326);
or U5484 (N_5484,N_5414,N_5342);
and U5485 (N_5485,N_5315,N_5423);
nor U5486 (N_5486,N_5369,N_5330);
xnor U5487 (N_5487,N_5301,N_5377);
nand U5488 (N_5488,N_5289,N_5358);
or U5489 (N_5489,N_5354,N_5294);
nand U5490 (N_5490,N_5426,N_5346);
nor U5491 (N_5491,N_5401,N_5418);
nor U5492 (N_5492,N_5348,N_5385);
xnor U5493 (N_5493,N_5400,N_5362);
and U5494 (N_5494,N_5382,N_5371);
xnor U5495 (N_5495,N_5420,N_5307);
nand U5496 (N_5496,N_5413,N_5292);
or U5497 (N_5497,N_5333,N_5404);
or U5498 (N_5498,N_5295,N_5433);
or U5499 (N_5499,N_5345,N_5290);
nand U5500 (N_5500,N_5281,N_5300);
xor U5501 (N_5501,N_5380,N_5355);
nor U5502 (N_5502,N_5335,N_5383);
nand U5503 (N_5503,N_5351,N_5417);
or U5504 (N_5504,N_5302,N_5410);
nand U5505 (N_5505,N_5359,N_5314);
nor U5506 (N_5506,N_5408,N_5318);
or U5507 (N_5507,N_5424,N_5288);
nor U5508 (N_5508,N_5350,N_5311);
or U5509 (N_5509,N_5390,N_5308);
nand U5510 (N_5510,N_5352,N_5356);
nand U5511 (N_5511,N_5364,N_5322);
or U5512 (N_5512,N_5309,N_5402);
or U5513 (N_5513,N_5328,N_5285);
or U5514 (N_5514,N_5331,N_5297);
nand U5515 (N_5515,N_5397,N_5282);
nand U5516 (N_5516,N_5407,N_5392);
xnor U5517 (N_5517,N_5361,N_5283);
nor U5518 (N_5518,N_5321,N_5393);
or U5519 (N_5519,N_5405,N_5384);
nor U5520 (N_5520,N_5430,N_5409);
nor U5521 (N_5521,N_5303,N_5366);
and U5522 (N_5522,N_5364,N_5383);
or U5523 (N_5523,N_5300,N_5374);
nand U5524 (N_5524,N_5370,N_5285);
or U5525 (N_5525,N_5396,N_5364);
and U5526 (N_5526,N_5390,N_5367);
nor U5527 (N_5527,N_5341,N_5303);
nor U5528 (N_5528,N_5376,N_5288);
nand U5529 (N_5529,N_5291,N_5340);
nor U5530 (N_5530,N_5388,N_5429);
nand U5531 (N_5531,N_5284,N_5400);
and U5532 (N_5532,N_5398,N_5335);
nand U5533 (N_5533,N_5391,N_5396);
nor U5534 (N_5534,N_5288,N_5418);
nand U5535 (N_5535,N_5325,N_5405);
and U5536 (N_5536,N_5382,N_5297);
xnor U5537 (N_5537,N_5360,N_5353);
nor U5538 (N_5538,N_5387,N_5419);
nand U5539 (N_5539,N_5297,N_5303);
nor U5540 (N_5540,N_5320,N_5297);
nor U5541 (N_5541,N_5413,N_5392);
nor U5542 (N_5542,N_5333,N_5433);
nand U5543 (N_5543,N_5343,N_5433);
and U5544 (N_5544,N_5293,N_5316);
or U5545 (N_5545,N_5400,N_5296);
and U5546 (N_5546,N_5337,N_5346);
xor U5547 (N_5547,N_5348,N_5350);
nand U5548 (N_5548,N_5334,N_5320);
nor U5549 (N_5549,N_5428,N_5427);
nor U5550 (N_5550,N_5351,N_5295);
nand U5551 (N_5551,N_5378,N_5293);
xor U5552 (N_5552,N_5359,N_5328);
xor U5553 (N_5553,N_5319,N_5403);
nor U5554 (N_5554,N_5436,N_5338);
and U5555 (N_5555,N_5429,N_5419);
xor U5556 (N_5556,N_5342,N_5314);
or U5557 (N_5557,N_5302,N_5365);
nor U5558 (N_5558,N_5406,N_5381);
nor U5559 (N_5559,N_5366,N_5296);
xor U5560 (N_5560,N_5396,N_5362);
nand U5561 (N_5561,N_5428,N_5410);
nor U5562 (N_5562,N_5410,N_5303);
and U5563 (N_5563,N_5374,N_5428);
and U5564 (N_5564,N_5351,N_5390);
nor U5565 (N_5565,N_5372,N_5382);
nor U5566 (N_5566,N_5349,N_5336);
nand U5567 (N_5567,N_5420,N_5359);
nand U5568 (N_5568,N_5296,N_5421);
and U5569 (N_5569,N_5298,N_5375);
nand U5570 (N_5570,N_5399,N_5284);
nand U5571 (N_5571,N_5409,N_5367);
and U5572 (N_5572,N_5290,N_5293);
xnor U5573 (N_5573,N_5333,N_5397);
nor U5574 (N_5574,N_5332,N_5370);
xor U5575 (N_5575,N_5281,N_5312);
nor U5576 (N_5576,N_5407,N_5337);
nor U5577 (N_5577,N_5402,N_5376);
or U5578 (N_5578,N_5314,N_5333);
xnor U5579 (N_5579,N_5330,N_5332);
nand U5580 (N_5580,N_5321,N_5428);
nand U5581 (N_5581,N_5385,N_5364);
nor U5582 (N_5582,N_5420,N_5347);
nand U5583 (N_5583,N_5425,N_5433);
xnor U5584 (N_5584,N_5381,N_5281);
nor U5585 (N_5585,N_5323,N_5352);
xnor U5586 (N_5586,N_5412,N_5281);
nand U5587 (N_5587,N_5283,N_5401);
and U5588 (N_5588,N_5303,N_5380);
nand U5589 (N_5589,N_5368,N_5405);
xnor U5590 (N_5590,N_5437,N_5302);
or U5591 (N_5591,N_5384,N_5434);
nand U5592 (N_5592,N_5412,N_5323);
or U5593 (N_5593,N_5286,N_5384);
nand U5594 (N_5594,N_5417,N_5423);
xor U5595 (N_5595,N_5287,N_5292);
xor U5596 (N_5596,N_5312,N_5307);
nand U5597 (N_5597,N_5409,N_5317);
and U5598 (N_5598,N_5389,N_5353);
xnor U5599 (N_5599,N_5284,N_5389);
or U5600 (N_5600,N_5599,N_5505);
xor U5601 (N_5601,N_5516,N_5563);
nor U5602 (N_5602,N_5501,N_5573);
nand U5603 (N_5603,N_5530,N_5535);
and U5604 (N_5604,N_5556,N_5534);
nor U5605 (N_5605,N_5532,N_5497);
or U5606 (N_5606,N_5592,N_5476);
nor U5607 (N_5607,N_5551,N_5565);
xor U5608 (N_5608,N_5538,N_5536);
or U5609 (N_5609,N_5562,N_5455);
nor U5610 (N_5610,N_5579,N_5493);
xor U5611 (N_5611,N_5576,N_5520);
nor U5612 (N_5612,N_5528,N_5555);
nand U5613 (N_5613,N_5442,N_5567);
or U5614 (N_5614,N_5509,N_5450);
and U5615 (N_5615,N_5456,N_5477);
or U5616 (N_5616,N_5572,N_5460);
xor U5617 (N_5617,N_5494,N_5527);
nand U5618 (N_5618,N_5486,N_5480);
nor U5619 (N_5619,N_5447,N_5585);
and U5620 (N_5620,N_5594,N_5503);
or U5621 (N_5621,N_5471,N_5500);
and U5622 (N_5622,N_5513,N_5441);
and U5623 (N_5623,N_5544,N_5479);
nand U5624 (N_5624,N_5444,N_5490);
nand U5625 (N_5625,N_5539,N_5484);
and U5626 (N_5626,N_5537,N_5596);
or U5627 (N_5627,N_5475,N_5577);
nand U5628 (N_5628,N_5468,N_5511);
xnor U5629 (N_5629,N_5558,N_5464);
nand U5630 (N_5630,N_5517,N_5591);
xor U5631 (N_5631,N_5550,N_5514);
or U5632 (N_5632,N_5448,N_5524);
and U5633 (N_5633,N_5459,N_5578);
and U5634 (N_5634,N_5489,N_5512);
xnor U5635 (N_5635,N_5443,N_5481);
nand U5636 (N_5636,N_5546,N_5508);
and U5637 (N_5637,N_5545,N_5483);
xor U5638 (N_5638,N_5465,N_5529);
nand U5639 (N_5639,N_5571,N_5548);
nor U5640 (N_5640,N_5440,N_5589);
and U5641 (N_5641,N_5518,N_5553);
xnor U5642 (N_5642,N_5522,N_5496);
nor U5643 (N_5643,N_5543,N_5510);
xor U5644 (N_5644,N_5474,N_5507);
nor U5645 (N_5645,N_5547,N_5566);
xnor U5646 (N_5646,N_5526,N_5469);
xnor U5647 (N_5647,N_5554,N_5446);
nand U5648 (N_5648,N_5570,N_5597);
xor U5649 (N_5649,N_5541,N_5533);
nor U5650 (N_5650,N_5557,N_5478);
or U5651 (N_5651,N_5466,N_5552);
xnor U5652 (N_5652,N_5467,N_5595);
xnor U5653 (N_5653,N_5568,N_5523);
nand U5654 (N_5654,N_5582,N_5485);
nor U5655 (N_5655,N_5488,N_5525);
xnor U5656 (N_5656,N_5561,N_5491);
nor U5657 (N_5657,N_5495,N_5560);
or U5658 (N_5658,N_5586,N_5593);
and U5659 (N_5659,N_5462,N_5487);
or U5660 (N_5660,N_5519,N_5504);
nand U5661 (N_5661,N_5584,N_5449);
nor U5662 (N_5662,N_5598,N_5506);
and U5663 (N_5663,N_5492,N_5531);
nor U5664 (N_5664,N_5470,N_5458);
or U5665 (N_5665,N_5461,N_5498);
nor U5666 (N_5666,N_5502,N_5587);
or U5667 (N_5667,N_5521,N_5580);
nand U5668 (N_5668,N_5542,N_5463);
and U5669 (N_5669,N_5540,N_5564);
nor U5670 (N_5670,N_5515,N_5454);
nor U5671 (N_5671,N_5581,N_5559);
nor U5672 (N_5672,N_5499,N_5472);
and U5673 (N_5673,N_5451,N_5590);
and U5674 (N_5674,N_5588,N_5452);
nor U5675 (N_5675,N_5575,N_5583);
and U5676 (N_5676,N_5569,N_5453);
and U5677 (N_5677,N_5574,N_5473);
nand U5678 (N_5678,N_5482,N_5445);
xnor U5679 (N_5679,N_5457,N_5549);
nand U5680 (N_5680,N_5591,N_5484);
xor U5681 (N_5681,N_5596,N_5570);
nor U5682 (N_5682,N_5562,N_5480);
xnor U5683 (N_5683,N_5469,N_5462);
xnor U5684 (N_5684,N_5537,N_5574);
and U5685 (N_5685,N_5525,N_5441);
and U5686 (N_5686,N_5530,N_5445);
nand U5687 (N_5687,N_5587,N_5569);
xnor U5688 (N_5688,N_5459,N_5444);
or U5689 (N_5689,N_5514,N_5559);
nand U5690 (N_5690,N_5579,N_5572);
xor U5691 (N_5691,N_5539,N_5522);
nand U5692 (N_5692,N_5456,N_5537);
nor U5693 (N_5693,N_5444,N_5596);
and U5694 (N_5694,N_5533,N_5526);
or U5695 (N_5695,N_5476,N_5472);
nand U5696 (N_5696,N_5496,N_5499);
and U5697 (N_5697,N_5538,N_5564);
nor U5698 (N_5698,N_5511,N_5441);
nor U5699 (N_5699,N_5476,N_5562);
and U5700 (N_5700,N_5441,N_5445);
xor U5701 (N_5701,N_5588,N_5493);
nand U5702 (N_5702,N_5492,N_5484);
nand U5703 (N_5703,N_5516,N_5448);
or U5704 (N_5704,N_5507,N_5520);
and U5705 (N_5705,N_5593,N_5544);
nor U5706 (N_5706,N_5546,N_5554);
or U5707 (N_5707,N_5460,N_5549);
nor U5708 (N_5708,N_5534,N_5586);
nand U5709 (N_5709,N_5512,N_5498);
and U5710 (N_5710,N_5594,N_5549);
xor U5711 (N_5711,N_5542,N_5516);
xor U5712 (N_5712,N_5546,N_5531);
nor U5713 (N_5713,N_5478,N_5463);
or U5714 (N_5714,N_5534,N_5559);
and U5715 (N_5715,N_5535,N_5590);
or U5716 (N_5716,N_5481,N_5489);
and U5717 (N_5717,N_5463,N_5535);
or U5718 (N_5718,N_5447,N_5467);
xor U5719 (N_5719,N_5556,N_5560);
nand U5720 (N_5720,N_5522,N_5469);
and U5721 (N_5721,N_5523,N_5527);
xnor U5722 (N_5722,N_5547,N_5468);
nand U5723 (N_5723,N_5504,N_5547);
nand U5724 (N_5724,N_5461,N_5567);
and U5725 (N_5725,N_5498,N_5484);
or U5726 (N_5726,N_5526,N_5490);
xnor U5727 (N_5727,N_5594,N_5570);
and U5728 (N_5728,N_5495,N_5482);
nor U5729 (N_5729,N_5528,N_5571);
and U5730 (N_5730,N_5532,N_5549);
and U5731 (N_5731,N_5571,N_5590);
and U5732 (N_5732,N_5554,N_5544);
nand U5733 (N_5733,N_5526,N_5472);
nor U5734 (N_5734,N_5499,N_5568);
xor U5735 (N_5735,N_5452,N_5590);
and U5736 (N_5736,N_5456,N_5519);
and U5737 (N_5737,N_5556,N_5490);
nand U5738 (N_5738,N_5451,N_5534);
or U5739 (N_5739,N_5556,N_5456);
xnor U5740 (N_5740,N_5587,N_5582);
xor U5741 (N_5741,N_5521,N_5505);
nand U5742 (N_5742,N_5469,N_5474);
and U5743 (N_5743,N_5449,N_5539);
xnor U5744 (N_5744,N_5569,N_5526);
xor U5745 (N_5745,N_5531,N_5524);
xnor U5746 (N_5746,N_5508,N_5440);
and U5747 (N_5747,N_5527,N_5571);
nor U5748 (N_5748,N_5515,N_5592);
xnor U5749 (N_5749,N_5466,N_5486);
and U5750 (N_5750,N_5448,N_5547);
nand U5751 (N_5751,N_5483,N_5535);
or U5752 (N_5752,N_5545,N_5574);
nor U5753 (N_5753,N_5570,N_5543);
nor U5754 (N_5754,N_5482,N_5516);
nor U5755 (N_5755,N_5446,N_5466);
and U5756 (N_5756,N_5532,N_5526);
nand U5757 (N_5757,N_5551,N_5546);
nand U5758 (N_5758,N_5481,N_5521);
nor U5759 (N_5759,N_5521,N_5542);
nor U5760 (N_5760,N_5688,N_5661);
xor U5761 (N_5761,N_5731,N_5750);
nor U5762 (N_5762,N_5625,N_5659);
or U5763 (N_5763,N_5614,N_5702);
nor U5764 (N_5764,N_5717,N_5678);
nand U5765 (N_5765,N_5752,N_5670);
and U5766 (N_5766,N_5646,N_5756);
nand U5767 (N_5767,N_5738,N_5677);
xor U5768 (N_5768,N_5711,N_5697);
nor U5769 (N_5769,N_5696,N_5732);
and U5770 (N_5770,N_5654,N_5631);
and U5771 (N_5771,N_5716,N_5617);
and U5772 (N_5772,N_5724,N_5603);
xor U5773 (N_5773,N_5753,N_5606);
and U5774 (N_5774,N_5748,N_5723);
xnor U5775 (N_5775,N_5728,N_5747);
or U5776 (N_5776,N_5628,N_5710);
nand U5777 (N_5777,N_5657,N_5726);
or U5778 (N_5778,N_5675,N_5663);
nor U5779 (N_5779,N_5705,N_5658);
nand U5780 (N_5780,N_5609,N_5638);
nand U5781 (N_5781,N_5703,N_5645);
and U5782 (N_5782,N_5686,N_5727);
nor U5783 (N_5783,N_5642,N_5616);
nor U5784 (N_5784,N_5721,N_5665);
xor U5785 (N_5785,N_5698,N_5744);
or U5786 (N_5786,N_5668,N_5713);
or U5787 (N_5787,N_5626,N_5704);
or U5788 (N_5788,N_5734,N_5637);
xor U5789 (N_5789,N_5608,N_5664);
or U5790 (N_5790,N_5630,N_5693);
or U5791 (N_5791,N_5641,N_5676);
or U5792 (N_5792,N_5739,N_5680);
xor U5793 (N_5793,N_5610,N_5699);
nor U5794 (N_5794,N_5619,N_5701);
or U5795 (N_5795,N_5640,N_5743);
nand U5796 (N_5796,N_5687,N_5707);
xnor U5797 (N_5797,N_5751,N_5615);
nand U5798 (N_5798,N_5759,N_5695);
nand U5799 (N_5799,N_5706,N_5655);
nor U5800 (N_5800,N_5666,N_5639);
nor U5801 (N_5801,N_5671,N_5629);
nor U5802 (N_5802,N_5684,N_5644);
and U5803 (N_5803,N_5700,N_5730);
xor U5804 (N_5804,N_5754,N_5736);
nand U5805 (N_5805,N_5689,N_5719);
xnor U5806 (N_5806,N_5712,N_5643);
nor U5807 (N_5807,N_5600,N_5740);
xor U5808 (N_5808,N_5733,N_5656);
or U5809 (N_5809,N_5650,N_5745);
or U5810 (N_5810,N_5691,N_5651);
nor U5811 (N_5811,N_5690,N_5624);
xnor U5812 (N_5812,N_5634,N_5622);
xor U5813 (N_5813,N_5683,N_5714);
xor U5814 (N_5814,N_5737,N_5601);
nor U5815 (N_5815,N_5604,N_5652);
and U5816 (N_5816,N_5648,N_5674);
nor U5817 (N_5817,N_5673,N_5653);
nor U5818 (N_5818,N_5758,N_5709);
nand U5819 (N_5819,N_5605,N_5613);
or U5820 (N_5820,N_5618,N_5669);
and U5821 (N_5821,N_5722,N_5620);
and U5822 (N_5822,N_5647,N_5662);
nor U5823 (N_5823,N_5720,N_5649);
and U5824 (N_5824,N_5621,N_5660);
or U5825 (N_5825,N_5635,N_5685);
xnor U5826 (N_5826,N_5694,N_5632);
and U5827 (N_5827,N_5633,N_5708);
xor U5828 (N_5828,N_5607,N_5612);
or U5829 (N_5829,N_5725,N_5667);
nor U5830 (N_5830,N_5611,N_5692);
nand U5831 (N_5831,N_5755,N_5672);
and U5832 (N_5832,N_5681,N_5746);
and U5833 (N_5833,N_5682,N_5741);
or U5834 (N_5834,N_5718,N_5729);
and U5835 (N_5835,N_5623,N_5636);
xor U5836 (N_5836,N_5749,N_5679);
nand U5837 (N_5837,N_5757,N_5602);
or U5838 (N_5838,N_5627,N_5715);
xor U5839 (N_5839,N_5742,N_5735);
xnor U5840 (N_5840,N_5617,N_5671);
or U5841 (N_5841,N_5661,N_5643);
xor U5842 (N_5842,N_5757,N_5711);
or U5843 (N_5843,N_5733,N_5643);
nand U5844 (N_5844,N_5729,N_5759);
or U5845 (N_5845,N_5719,N_5702);
or U5846 (N_5846,N_5734,N_5722);
nor U5847 (N_5847,N_5693,N_5680);
or U5848 (N_5848,N_5693,N_5712);
xor U5849 (N_5849,N_5725,N_5672);
nor U5850 (N_5850,N_5670,N_5640);
nand U5851 (N_5851,N_5750,N_5709);
nor U5852 (N_5852,N_5634,N_5704);
xnor U5853 (N_5853,N_5712,N_5706);
nand U5854 (N_5854,N_5610,N_5612);
xnor U5855 (N_5855,N_5704,N_5689);
or U5856 (N_5856,N_5752,N_5637);
nand U5857 (N_5857,N_5701,N_5681);
and U5858 (N_5858,N_5757,N_5759);
and U5859 (N_5859,N_5747,N_5681);
nand U5860 (N_5860,N_5728,N_5606);
nor U5861 (N_5861,N_5684,N_5723);
and U5862 (N_5862,N_5726,N_5690);
xor U5863 (N_5863,N_5669,N_5634);
and U5864 (N_5864,N_5712,N_5748);
nor U5865 (N_5865,N_5611,N_5681);
nand U5866 (N_5866,N_5652,N_5730);
nor U5867 (N_5867,N_5693,N_5648);
nor U5868 (N_5868,N_5750,N_5606);
nand U5869 (N_5869,N_5619,N_5660);
xor U5870 (N_5870,N_5623,N_5711);
nand U5871 (N_5871,N_5604,N_5636);
nand U5872 (N_5872,N_5641,N_5757);
or U5873 (N_5873,N_5699,N_5743);
or U5874 (N_5874,N_5610,N_5611);
xor U5875 (N_5875,N_5686,N_5656);
nand U5876 (N_5876,N_5743,N_5696);
nand U5877 (N_5877,N_5738,N_5711);
and U5878 (N_5878,N_5657,N_5607);
and U5879 (N_5879,N_5615,N_5609);
nor U5880 (N_5880,N_5643,N_5726);
and U5881 (N_5881,N_5745,N_5602);
nor U5882 (N_5882,N_5691,N_5663);
nor U5883 (N_5883,N_5726,N_5757);
nand U5884 (N_5884,N_5645,N_5743);
nor U5885 (N_5885,N_5669,N_5673);
or U5886 (N_5886,N_5604,N_5746);
nand U5887 (N_5887,N_5654,N_5614);
nor U5888 (N_5888,N_5719,N_5608);
nand U5889 (N_5889,N_5692,N_5742);
nor U5890 (N_5890,N_5665,N_5609);
and U5891 (N_5891,N_5740,N_5605);
or U5892 (N_5892,N_5684,N_5616);
nor U5893 (N_5893,N_5744,N_5678);
or U5894 (N_5894,N_5721,N_5739);
xnor U5895 (N_5895,N_5715,N_5734);
nor U5896 (N_5896,N_5689,N_5627);
nand U5897 (N_5897,N_5699,N_5650);
or U5898 (N_5898,N_5675,N_5629);
nor U5899 (N_5899,N_5601,N_5744);
and U5900 (N_5900,N_5724,N_5729);
and U5901 (N_5901,N_5648,N_5627);
xnor U5902 (N_5902,N_5658,N_5608);
or U5903 (N_5903,N_5731,N_5619);
and U5904 (N_5904,N_5640,N_5617);
or U5905 (N_5905,N_5700,N_5755);
or U5906 (N_5906,N_5616,N_5693);
xnor U5907 (N_5907,N_5628,N_5687);
nand U5908 (N_5908,N_5673,N_5616);
and U5909 (N_5909,N_5704,N_5665);
nand U5910 (N_5910,N_5604,N_5600);
xnor U5911 (N_5911,N_5649,N_5734);
nor U5912 (N_5912,N_5624,N_5666);
or U5913 (N_5913,N_5677,N_5709);
xnor U5914 (N_5914,N_5736,N_5622);
nor U5915 (N_5915,N_5625,N_5672);
and U5916 (N_5916,N_5705,N_5663);
or U5917 (N_5917,N_5608,N_5614);
xnor U5918 (N_5918,N_5629,N_5600);
and U5919 (N_5919,N_5755,N_5699);
and U5920 (N_5920,N_5915,N_5839);
xnor U5921 (N_5921,N_5826,N_5905);
nor U5922 (N_5922,N_5806,N_5824);
or U5923 (N_5923,N_5810,N_5881);
xor U5924 (N_5924,N_5903,N_5820);
nand U5925 (N_5925,N_5788,N_5893);
and U5926 (N_5926,N_5911,N_5849);
and U5927 (N_5927,N_5880,N_5790);
and U5928 (N_5928,N_5803,N_5845);
xnor U5929 (N_5929,N_5816,N_5888);
and U5930 (N_5930,N_5856,N_5818);
nand U5931 (N_5931,N_5896,N_5857);
nor U5932 (N_5932,N_5798,N_5882);
nor U5933 (N_5933,N_5774,N_5868);
xnor U5934 (N_5934,N_5779,N_5869);
and U5935 (N_5935,N_5815,N_5840);
and U5936 (N_5936,N_5874,N_5791);
and U5937 (N_5937,N_5793,N_5827);
nor U5938 (N_5938,N_5797,N_5764);
and U5939 (N_5939,N_5813,N_5767);
nand U5940 (N_5940,N_5802,N_5783);
nand U5941 (N_5941,N_5873,N_5807);
or U5942 (N_5942,N_5914,N_5789);
nor U5943 (N_5943,N_5808,N_5848);
xnor U5944 (N_5944,N_5835,N_5852);
nand U5945 (N_5945,N_5867,N_5780);
nor U5946 (N_5946,N_5821,N_5823);
xor U5947 (N_5947,N_5918,N_5895);
and U5948 (N_5948,N_5909,N_5865);
xnor U5949 (N_5949,N_5907,N_5838);
or U5950 (N_5950,N_5784,N_5870);
and U5951 (N_5951,N_5825,N_5829);
nor U5952 (N_5952,N_5832,N_5760);
or U5953 (N_5953,N_5777,N_5775);
xor U5954 (N_5954,N_5828,N_5898);
or U5955 (N_5955,N_5805,N_5879);
and U5956 (N_5956,N_5811,N_5906);
xor U5957 (N_5957,N_5843,N_5902);
and U5958 (N_5958,N_5831,N_5875);
nor U5959 (N_5959,N_5772,N_5846);
xor U5960 (N_5960,N_5792,N_5904);
nand U5961 (N_5961,N_5889,N_5769);
nor U5962 (N_5962,N_5916,N_5910);
nand U5963 (N_5963,N_5897,N_5864);
and U5964 (N_5964,N_5883,N_5876);
and U5965 (N_5965,N_5887,N_5833);
and U5966 (N_5966,N_5917,N_5901);
or U5967 (N_5967,N_5795,N_5766);
or U5968 (N_5968,N_5770,N_5855);
nand U5969 (N_5969,N_5830,N_5771);
nor U5970 (N_5970,N_5809,N_5786);
nand U5971 (N_5971,N_5776,N_5894);
and U5972 (N_5972,N_5801,N_5885);
or U5973 (N_5973,N_5900,N_5861);
xor U5974 (N_5974,N_5871,N_5872);
and U5975 (N_5975,N_5853,N_5773);
nand U5976 (N_5976,N_5850,N_5782);
nor U5977 (N_5977,N_5765,N_5858);
nor U5978 (N_5978,N_5817,N_5794);
nor U5979 (N_5979,N_5785,N_5787);
and U5980 (N_5980,N_5866,N_5822);
nand U5981 (N_5981,N_5847,N_5859);
xnor U5982 (N_5982,N_5908,N_5800);
nand U5983 (N_5983,N_5837,N_5854);
xnor U5984 (N_5984,N_5892,N_5814);
nand U5985 (N_5985,N_5844,N_5796);
or U5986 (N_5986,N_5819,N_5842);
nor U5987 (N_5987,N_5913,N_5862);
nand U5988 (N_5988,N_5877,N_5778);
xor U5989 (N_5989,N_5878,N_5890);
nor U5990 (N_5990,N_5860,N_5919);
nor U5991 (N_5991,N_5891,N_5762);
and U5992 (N_5992,N_5851,N_5768);
xnor U5993 (N_5993,N_5841,N_5912);
nand U5994 (N_5994,N_5812,N_5834);
xor U5995 (N_5995,N_5863,N_5836);
xnor U5996 (N_5996,N_5804,N_5799);
xor U5997 (N_5997,N_5763,N_5781);
nor U5998 (N_5998,N_5886,N_5884);
or U5999 (N_5999,N_5899,N_5761);
nor U6000 (N_6000,N_5836,N_5877);
and U6001 (N_6001,N_5854,N_5789);
and U6002 (N_6002,N_5848,N_5899);
nand U6003 (N_6003,N_5869,N_5786);
nor U6004 (N_6004,N_5762,N_5760);
nor U6005 (N_6005,N_5878,N_5876);
xnor U6006 (N_6006,N_5771,N_5819);
xor U6007 (N_6007,N_5856,N_5905);
nor U6008 (N_6008,N_5829,N_5862);
or U6009 (N_6009,N_5799,N_5760);
nand U6010 (N_6010,N_5806,N_5805);
xor U6011 (N_6011,N_5769,N_5864);
nand U6012 (N_6012,N_5771,N_5770);
nor U6013 (N_6013,N_5886,N_5760);
nand U6014 (N_6014,N_5838,N_5769);
nor U6015 (N_6015,N_5859,N_5852);
nor U6016 (N_6016,N_5792,N_5905);
and U6017 (N_6017,N_5916,N_5769);
nand U6018 (N_6018,N_5779,N_5879);
and U6019 (N_6019,N_5895,N_5914);
nand U6020 (N_6020,N_5773,N_5903);
nor U6021 (N_6021,N_5869,N_5794);
xor U6022 (N_6022,N_5801,N_5843);
nand U6023 (N_6023,N_5850,N_5902);
and U6024 (N_6024,N_5854,N_5788);
nor U6025 (N_6025,N_5888,N_5902);
or U6026 (N_6026,N_5768,N_5911);
and U6027 (N_6027,N_5916,N_5779);
xor U6028 (N_6028,N_5831,N_5902);
xor U6029 (N_6029,N_5881,N_5779);
or U6030 (N_6030,N_5846,N_5799);
nor U6031 (N_6031,N_5888,N_5912);
xor U6032 (N_6032,N_5908,N_5819);
and U6033 (N_6033,N_5874,N_5893);
nand U6034 (N_6034,N_5892,N_5786);
or U6035 (N_6035,N_5843,N_5853);
and U6036 (N_6036,N_5841,N_5761);
and U6037 (N_6037,N_5772,N_5880);
or U6038 (N_6038,N_5780,N_5917);
xnor U6039 (N_6039,N_5779,N_5760);
xnor U6040 (N_6040,N_5795,N_5801);
xnor U6041 (N_6041,N_5763,N_5883);
and U6042 (N_6042,N_5871,N_5902);
or U6043 (N_6043,N_5825,N_5819);
nand U6044 (N_6044,N_5896,N_5809);
or U6045 (N_6045,N_5886,N_5856);
and U6046 (N_6046,N_5905,N_5815);
nand U6047 (N_6047,N_5823,N_5869);
or U6048 (N_6048,N_5838,N_5809);
xor U6049 (N_6049,N_5850,N_5790);
or U6050 (N_6050,N_5903,N_5881);
and U6051 (N_6051,N_5856,N_5772);
nor U6052 (N_6052,N_5816,N_5760);
or U6053 (N_6053,N_5818,N_5813);
and U6054 (N_6054,N_5794,N_5905);
xor U6055 (N_6055,N_5817,N_5763);
xor U6056 (N_6056,N_5875,N_5771);
or U6057 (N_6057,N_5913,N_5845);
xor U6058 (N_6058,N_5777,N_5793);
xor U6059 (N_6059,N_5775,N_5854);
nand U6060 (N_6060,N_5818,N_5840);
and U6061 (N_6061,N_5801,N_5828);
xor U6062 (N_6062,N_5900,N_5919);
or U6063 (N_6063,N_5810,N_5912);
or U6064 (N_6064,N_5865,N_5777);
or U6065 (N_6065,N_5839,N_5769);
or U6066 (N_6066,N_5869,N_5829);
or U6067 (N_6067,N_5823,N_5781);
and U6068 (N_6068,N_5825,N_5800);
nand U6069 (N_6069,N_5898,N_5850);
nand U6070 (N_6070,N_5906,N_5860);
or U6071 (N_6071,N_5847,N_5814);
or U6072 (N_6072,N_5847,N_5852);
xnor U6073 (N_6073,N_5917,N_5843);
nand U6074 (N_6074,N_5822,N_5910);
xor U6075 (N_6075,N_5802,N_5835);
or U6076 (N_6076,N_5770,N_5864);
nand U6077 (N_6077,N_5907,N_5798);
and U6078 (N_6078,N_5914,N_5874);
or U6079 (N_6079,N_5868,N_5788);
nor U6080 (N_6080,N_5983,N_5944);
nand U6081 (N_6081,N_6065,N_6011);
or U6082 (N_6082,N_5989,N_5976);
xor U6083 (N_6083,N_6019,N_6010);
nor U6084 (N_6084,N_5921,N_5945);
and U6085 (N_6085,N_5996,N_5965);
or U6086 (N_6086,N_5986,N_6004);
and U6087 (N_6087,N_5990,N_5961);
nor U6088 (N_6088,N_6037,N_5924);
nor U6089 (N_6089,N_5982,N_5954);
xnor U6090 (N_6090,N_6071,N_6053);
xnor U6091 (N_6091,N_5977,N_5966);
nor U6092 (N_6092,N_5967,N_6020);
nand U6093 (N_6093,N_6025,N_5973);
xor U6094 (N_6094,N_5991,N_6076);
and U6095 (N_6095,N_6048,N_5949);
nand U6096 (N_6096,N_6073,N_6044);
nor U6097 (N_6097,N_6066,N_6009);
nor U6098 (N_6098,N_5936,N_5930);
and U6099 (N_6099,N_6036,N_6074);
xor U6100 (N_6100,N_6070,N_6006);
or U6101 (N_6101,N_6024,N_5985);
xnor U6102 (N_6102,N_6014,N_6041);
nand U6103 (N_6103,N_5987,N_6007);
and U6104 (N_6104,N_6028,N_5934);
or U6105 (N_6105,N_6002,N_5953);
nor U6106 (N_6106,N_6077,N_5960);
nand U6107 (N_6107,N_6051,N_6050);
nor U6108 (N_6108,N_5946,N_5963);
nor U6109 (N_6109,N_5931,N_5999);
or U6110 (N_6110,N_5968,N_5964);
xor U6111 (N_6111,N_5984,N_6055);
and U6112 (N_6112,N_5971,N_5951);
nor U6113 (N_6113,N_5988,N_5935);
nand U6114 (N_6114,N_6069,N_5955);
or U6115 (N_6115,N_5938,N_6021);
nand U6116 (N_6116,N_6072,N_6005);
nor U6117 (N_6117,N_6056,N_5942);
nand U6118 (N_6118,N_6047,N_5943);
xnor U6119 (N_6119,N_6060,N_5957);
or U6120 (N_6120,N_6032,N_5970);
and U6121 (N_6121,N_6046,N_6030);
nand U6122 (N_6122,N_5952,N_5920);
nor U6123 (N_6123,N_5993,N_5956);
and U6124 (N_6124,N_6034,N_5925);
nor U6125 (N_6125,N_5997,N_6042);
or U6126 (N_6126,N_6013,N_5981);
nand U6127 (N_6127,N_6000,N_5939);
and U6128 (N_6128,N_6045,N_5950);
xnor U6129 (N_6129,N_5940,N_6026);
nand U6130 (N_6130,N_6067,N_5998);
xnor U6131 (N_6131,N_6079,N_5948);
xnor U6132 (N_6132,N_6039,N_5959);
nand U6133 (N_6133,N_5958,N_6068);
or U6134 (N_6134,N_6078,N_6049);
nor U6135 (N_6135,N_6035,N_6018);
nor U6136 (N_6136,N_5992,N_6001);
xor U6137 (N_6137,N_5978,N_6015);
xor U6138 (N_6138,N_5995,N_6064);
nand U6139 (N_6139,N_5947,N_6063);
and U6140 (N_6140,N_5933,N_6027);
or U6141 (N_6141,N_6057,N_6003);
nor U6142 (N_6142,N_5929,N_6043);
and U6143 (N_6143,N_6058,N_5941);
xor U6144 (N_6144,N_5937,N_5962);
and U6145 (N_6145,N_5975,N_6031);
or U6146 (N_6146,N_5926,N_6017);
nor U6147 (N_6147,N_6054,N_5994);
nand U6148 (N_6148,N_6008,N_6040);
nand U6149 (N_6149,N_6038,N_6016);
xor U6150 (N_6150,N_5974,N_6061);
xor U6151 (N_6151,N_5979,N_5922);
or U6152 (N_6152,N_6062,N_6029);
and U6153 (N_6153,N_6075,N_5969);
or U6154 (N_6154,N_6012,N_5932);
xnor U6155 (N_6155,N_6033,N_5972);
xor U6156 (N_6156,N_5980,N_6023);
nand U6157 (N_6157,N_6022,N_6052);
or U6158 (N_6158,N_5928,N_5927);
xnor U6159 (N_6159,N_5923,N_6059);
xor U6160 (N_6160,N_6071,N_6047);
nand U6161 (N_6161,N_5982,N_5941);
xnor U6162 (N_6162,N_6042,N_5937);
or U6163 (N_6163,N_6034,N_5947);
xnor U6164 (N_6164,N_5996,N_6039);
nor U6165 (N_6165,N_5948,N_6050);
nor U6166 (N_6166,N_6026,N_5946);
nand U6167 (N_6167,N_5966,N_6048);
nand U6168 (N_6168,N_6023,N_5989);
and U6169 (N_6169,N_6025,N_6042);
nand U6170 (N_6170,N_6006,N_5990);
nand U6171 (N_6171,N_6041,N_6076);
nor U6172 (N_6172,N_6058,N_5995);
nand U6173 (N_6173,N_5991,N_6060);
or U6174 (N_6174,N_5964,N_6049);
or U6175 (N_6175,N_6035,N_6064);
or U6176 (N_6176,N_5935,N_6024);
and U6177 (N_6177,N_6044,N_5948);
xnor U6178 (N_6178,N_5944,N_5981);
nor U6179 (N_6179,N_6073,N_5935);
nand U6180 (N_6180,N_6009,N_5927);
xor U6181 (N_6181,N_5968,N_5989);
or U6182 (N_6182,N_5981,N_5972);
and U6183 (N_6183,N_5984,N_6040);
or U6184 (N_6184,N_6016,N_5924);
or U6185 (N_6185,N_6021,N_5976);
and U6186 (N_6186,N_6058,N_6048);
or U6187 (N_6187,N_6068,N_6020);
or U6188 (N_6188,N_5920,N_5991);
nor U6189 (N_6189,N_6031,N_5944);
xor U6190 (N_6190,N_5958,N_5954);
nor U6191 (N_6191,N_6054,N_6019);
xnor U6192 (N_6192,N_5943,N_5923);
nor U6193 (N_6193,N_6022,N_5931);
or U6194 (N_6194,N_6026,N_6033);
nor U6195 (N_6195,N_5986,N_6018);
xnor U6196 (N_6196,N_6001,N_5986);
xnor U6197 (N_6197,N_5967,N_6065);
nor U6198 (N_6198,N_6042,N_5960);
and U6199 (N_6199,N_5968,N_6077);
or U6200 (N_6200,N_5989,N_5961);
nand U6201 (N_6201,N_5927,N_6059);
or U6202 (N_6202,N_6054,N_5999);
nand U6203 (N_6203,N_5943,N_5988);
or U6204 (N_6204,N_5966,N_5934);
or U6205 (N_6205,N_6018,N_6015);
nand U6206 (N_6206,N_5995,N_5941);
and U6207 (N_6207,N_6039,N_5949);
nor U6208 (N_6208,N_5934,N_5991);
nand U6209 (N_6209,N_6020,N_6035);
xor U6210 (N_6210,N_6027,N_6053);
or U6211 (N_6211,N_6004,N_6040);
xor U6212 (N_6212,N_5943,N_5976);
xnor U6213 (N_6213,N_6069,N_6057);
xnor U6214 (N_6214,N_5977,N_6039);
nor U6215 (N_6215,N_6052,N_6059);
and U6216 (N_6216,N_5983,N_5970);
nand U6217 (N_6217,N_5941,N_5935);
nand U6218 (N_6218,N_5962,N_5928);
or U6219 (N_6219,N_6074,N_6043);
nand U6220 (N_6220,N_6054,N_6000);
nand U6221 (N_6221,N_5943,N_5991);
nor U6222 (N_6222,N_6016,N_6052);
and U6223 (N_6223,N_5961,N_6016);
nand U6224 (N_6224,N_5955,N_6070);
or U6225 (N_6225,N_5966,N_5960);
or U6226 (N_6226,N_6003,N_6039);
nor U6227 (N_6227,N_5980,N_6033);
nand U6228 (N_6228,N_6055,N_6030);
nand U6229 (N_6229,N_6062,N_5999);
nand U6230 (N_6230,N_6005,N_6046);
and U6231 (N_6231,N_6057,N_6029);
or U6232 (N_6232,N_6013,N_6014);
xnor U6233 (N_6233,N_6060,N_5967);
nor U6234 (N_6234,N_6039,N_5941);
nand U6235 (N_6235,N_6006,N_5956);
xnor U6236 (N_6236,N_5954,N_6016);
nand U6237 (N_6237,N_5974,N_6026);
nand U6238 (N_6238,N_6028,N_6040);
xnor U6239 (N_6239,N_6052,N_6029);
xor U6240 (N_6240,N_6209,N_6219);
xnor U6241 (N_6241,N_6157,N_6174);
xor U6242 (N_6242,N_6234,N_6135);
xor U6243 (N_6243,N_6111,N_6117);
xor U6244 (N_6244,N_6166,N_6103);
or U6245 (N_6245,N_6092,N_6083);
and U6246 (N_6246,N_6142,N_6105);
or U6247 (N_6247,N_6239,N_6194);
nand U6248 (N_6248,N_6218,N_6152);
xor U6249 (N_6249,N_6133,N_6122);
and U6250 (N_6250,N_6238,N_6099);
and U6251 (N_6251,N_6098,N_6224);
or U6252 (N_6252,N_6195,N_6160);
xnor U6253 (N_6253,N_6106,N_6186);
and U6254 (N_6254,N_6140,N_6197);
nand U6255 (N_6255,N_6205,N_6231);
xor U6256 (N_6256,N_6089,N_6125);
xnor U6257 (N_6257,N_6093,N_6182);
and U6258 (N_6258,N_6136,N_6175);
nor U6259 (N_6259,N_6080,N_6088);
nor U6260 (N_6260,N_6168,N_6236);
and U6261 (N_6261,N_6216,N_6109);
xor U6262 (N_6262,N_6176,N_6147);
nor U6263 (N_6263,N_6091,N_6115);
or U6264 (N_6264,N_6156,N_6127);
nor U6265 (N_6265,N_6131,N_6217);
xor U6266 (N_6266,N_6108,N_6210);
nand U6267 (N_6267,N_6200,N_6207);
nand U6268 (N_6268,N_6188,N_6084);
nand U6269 (N_6269,N_6081,N_6162);
and U6270 (N_6270,N_6094,N_6097);
nor U6271 (N_6271,N_6096,N_6113);
or U6272 (N_6272,N_6235,N_6086);
or U6273 (N_6273,N_6145,N_6149);
nand U6274 (N_6274,N_6110,N_6100);
or U6275 (N_6275,N_6201,N_6163);
nand U6276 (N_6276,N_6198,N_6165);
or U6277 (N_6277,N_6185,N_6114);
nand U6278 (N_6278,N_6112,N_6090);
xnor U6279 (N_6279,N_6126,N_6159);
nor U6280 (N_6280,N_6232,N_6183);
nor U6281 (N_6281,N_6120,N_6085);
or U6282 (N_6282,N_6144,N_6171);
nand U6283 (N_6283,N_6164,N_6208);
nor U6284 (N_6284,N_6203,N_6212);
nand U6285 (N_6285,N_6129,N_6119);
xnor U6286 (N_6286,N_6121,N_6206);
or U6287 (N_6287,N_6204,N_6177);
and U6288 (N_6288,N_6179,N_6237);
nand U6289 (N_6289,N_6101,N_6141);
nand U6290 (N_6290,N_6107,N_6229);
and U6291 (N_6291,N_6199,N_6180);
and U6292 (N_6292,N_6158,N_6102);
or U6293 (N_6293,N_6220,N_6146);
and U6294 (N_6294,N_6172,N_6184);
xor U6295 (N_6295,N_6095,N_6223);
nand U6296 (N_6296,N_6150,N_6190);
nand U6297 (N_6297,N_6118,N_6124);
nor U6298 (N_6298,N_6128,N_6170);
and U6299 (N_6299,N_6167,N_6230);
nand U6300 (N_6300,N_6155,N_6202);
nand U6301 (N_6301,N_6137,N_6151);
or U6302 (N_6302,N_6233,N_6173);
xnor U6303 (N_6303,N_6222,N_6138);
nor U6304 (N_6304,N_6193,N_6123);
xor U6305 (N_6305,N_6187,N_6196);
nor U6306 (N_6306,N_6215,N_6082);
or U6307 (N_6307,N_6192,N_6134);
or U6308 (N_6308,N_6148,N_6161);
nand U6309 (N_6309,N_6227,N_6214);
nand U6310 (N_6310,N_6228,N_6178);
or U6311 (N_6311,N_6226,N_6181);
and U6312 (N_6312,N_6221,N_6169);
nand U6313 (N_6313,N_6104,N_6139);
nand U6314 (N_6314,N_6130,N_6087);
xor U6315 (N_6315,N_6211,N_6154);
and U6316 (N_6316,N_6153,N_6191);
and U6317 (N_6317,N_6225,N_6213);
xor U6318 (N_6318,N_6189,N_6116);
or U6319 (N_6319,N_6143,N_6132);
nor U6320 (N_6320,N_6198,N_6211);
nand U6321 (N_6321,N_6128,N_6120);
xnor U6322 (N_6322,N_6096,N_6207);
and U6323 (N_6323,N_6106,N_6090);
nor U6324 (N_6324,N_6157,N_6127);
or U6325 (N_6325,N_6178,N_6196);
or U6326 (N_6326,N_6095,N_6234);
and U6327 (N_6327,N_6124,N_6108);
or U6328 (N_6328,N_6113,N_6110);
nand U6329 (N_6329,N_6113,N_6158);
nor U6330 (N_6330,N_6157,N_6130);
nor U6331 (N_6331,N_6209,N_6172);
nor U6332 (N_6332,N_6148,N_6197);
or U6333 (N_6333,N_6220,N_6218);
nand U6334 (N_6334,N_6140,N_6206);
and U6335 (N_6335,N_6173,N_6102);
or U6336 (N_6336,N_6170,N_6208);
and U6337 (N_6337,N_6176,N_6198);
nor U6338 (N_6338,N_6143,N_6142);
xor U6339 (N_6339,N_6098,N_6222);
nor U6340 (N_6340,N_6214,N_6119);
xnor U6341 (N_6341,N_6088,N_6159);
and U6342 (N_6342,N_6175,N_6116);
nor U6343 (N_6343,N_6219,N_6213);
or U6344 (N_6344,N_6219,N_6088);
xnor U6345 (N_6345,N_6140,N_6160);
or U6346 (N_6346,N_6184,N_6092);
and U6347 (N_6347,N_6132,N_6163);
xor U6348 (N_6348,N_6135,N_6168);
or U6349 (N_6349,N_6197,N_6208);
nor U6350 (N_6350,N_6215,N_6096);
xor U6351 (N_6351,N_6092,N_6094);
and U6352 (N_6352,N_6237,N_6086);
nor U6353 (N_6353,N_6089,N_6098);
or U6354 (N_6354,N_6110,N_6189);
xor U6355 (N_6355,N_6199,N_6159);
or U6356 (N_6356,N_6216,N_6225);
xnor U6357 (N_6357,N_6131,N_6206);
or U6358 (N_6358,N_6174,N_6085);
or U6359 (N_6359,N_6197,N_6094);
xor U6360 (N_6360,N_6143,N_6167);
nand U6361 (N_6361,N_6235,N_6183);
xor U6362 (N_6362,N_6224,N_6149);
and U6363 (N_6363,N_6123,N_6210);
nand U6364 (N_6364,N_6179,N_6202);
and U6365 (N_6365,N_6153,N_6188);
nand U6366 (N_6366,N_6120,N_6187);
nand U6367 (N_6367,N_6108,N_6155);
or U6368 (N_6368,N_6214,N_6183);
and U6369 (N_6369,N_6227,N_6237);
and U6370 (N_6370,N_6165,N_6200);
xor U6371 (N_6371,N_6094,N_6129);
and U6372 (N_6372,N_6238,N_6134);
nand U6373 (N_6373,N_6086,N_6185);
nor U6374 (N_6374,N_6166,N_6147);
nor U6375 (N_6375,N_6193,N_6104);
nor U6376 (N_6376,N_6119,N_6120);
xnor U6377 (N_6377,N_6084,N_6141);
nand U6378 (N_6378,N_6092,N_6201);
and U6379 (N_6379,N_6135,N_6160);
nand U6380 (N_6380,N_6222,N_6177);
xnor U6381 (N_6381,N_6106,N_6181);
or U6382 (N_6382,N_6111,N_6228);
xor U6383 (N_6383,N_6192,N_6119);
nor U6384 (N_6384,N_6175,N_6199);
nand U6385 (N_6385,N_6236,N_6143);
and U6386 (N_6386,N_6086,N_6138);
or U6387 (N_6387,N_6226,N_6215);
and U6388 (N_6388,N_6238,N_6149);
nor U6389 (N_6389,N_6196,N_6165);
nor U6390 (N_6390,N_6141,N_6212);
nor U6391 (N_6391,N_6187,N_6100);
or U6392 (N_6392,N_6126,N_6086);
nand U6393 (N_6393,N_6112,N_6215);
or U6394 (N_6394,N_6159,N_6146);
or U6395 (N_6395,N_6157,N_6096);
or U6396 (N_6396,N_6220,N_6197);
xnor U6397 (N_6397,N_6211,N_6137);
xnor U6398 (N_6398,N_6118,N_6192);
or U6399 (N_6399,N_6220,N_6081);
or U6400 (N_6400,N_6300,N_6274);
nor U6401 (N_6401,N_6399,N_6299);
nand U6402 (N_6402,N_6367,N_6273);
nand U6403 (N_6403,N_6292,N_6327);
nor U6404 (N_6404,N_6341,N_6352);
or U6405 (N_6405,N_6387,N_6378);
xnor U6406 (N_6406,N_6289,N_6391);
or U6407 (N_6407,N_6381,N_6297);
or U6408 (N_6408,N_6253,N_6397);
nor U6409 (N_6409,N_6247,N_6287);
nor U6410 (N_6410,N_6250,N_6265);
or U6411 (N_6411,N_6376,N_6285);
nand U6412 (N_6412,N_6375,N_6386);
and U6413 (N_6413,N_6304,N_6240);
and U6414 (N_6414,N_6332,N_6363);
nand U6415 (N_6415,N_6358,N_6267);
nor U6416 (N_6416,N_6241,N_6322);
or U6417 (N_6417,N_6349,N_6317);
and U6418 (N_6418,N_6277,N_6283);
xnor U6419 (N_6419,N_6369,N_6345);
nor U6420 (N_6420,N_6294,N_6258);
nand U6421 (N_6421,N_6371,N_6256);
and U6422 (N_6422,N_6337,N_6270);
xnor U6423 (N_6423,N_6260,N_6353);
nand U6424 (N_6424,N_6315,N_6394);
or U6425 (N_6425,N_6343,N_6388);
nand U6426 (N_6426,N_6370,N_6310);
nor U6427 (N_6427,N_6279,N_6336);
nand U6428 (N_6428,N_6246,N_6312);
nor U6429 (N_6429,N_6264,N_6347);
nand U6430 (N_6430,N_6320,N_6362);
nand U6431 (N_6431,N_6281,N_6326);
nand U6432 (N_6432,N_6360,N_6309);
and U6433 (N_6433,N_6251,N_6302);
nor U6434 (N_6434,N_6372,N_6377);
nor U6435 (N_6435,N_6262,N_6321);
nor U6436 (N_6436,N_6252,N_6325);
nor U6437 (N_6437,N_6242,N_6263);
and U6438 (N_6438,N_6269,N_6348);
xnor U6439 (N_6439,N_6293,N_6382);
xnor U6440 (N_6440,N_6318,N_6384);
xor U6441 (N_6441,N_6338,N_6357);
or U6442 (N_6442,N_6314,N_6366);
xnor U6443 (N_6443,N_6261,N_6330);
or U6444 (N_6444,N_6307,N_6385);
xnor U6445 (N_6445,N_6323,N_6266);
xor U6446 (N_6446,N_6329,N_6396);
or U6447 (N_6447,N_6374,N_6259);
or U6448 (N_6448,N_6245,N_6311);
and U6449 (N_6449,N_6303,N_6350);
nand U6450 (N_6450,N_6380,N_6243);
and U6451 (N_6451,N_6255,N_6373);
nand U6452 (N_6452,N_6340,N_6334);
nor U6453 (N_6453,N_6390,N_6324);
xnor U6454 (N_6454,N_6342,N_6248);
xnor U6455 (N_6455,N_6295,N_6286);
or U6456 (N_6456,N_6301,N_6308);
and U6457 (N_6457,N_6288,N_6305);
nor U6458 (N_6458,N_6393,N_6383);
and U6459 (N_6459,N_6339,N_6271);
nand U6460 (N_6460,N_6284,N_6365);
xnor U6461 (N_6461,N_6276,N_6354);
nor U6462 (N_6462,N_6389,N_6333);
nor U6463 (N_6463,N_6280,N_6328);
nand U6464 (N_6464,N_6282,N_6398);
and U6465 (N_6465,N_6268,N_6361);
nand U6466 (N_6466,N_6275,N_6344);
nand U6467 (N_6467,N_6368,N_6249);
nand U6468 (N_6468,N_6244,N_6306);
and U6469 (N_6469,N_6272,N_6316);
nand U6470 (N_6470,N_6331,N_6290);
nand U6471 (N_6471,N_6346,N_6319);
and U6472 (N_6472,N_6254,N_6356);
xnor U6473 (N_6473,N_6335,N_6395);
nand U6474 (N_6474,N_6364,N_6296);
or U6475 (N_6475,N_6313,N_6278);
and U6476 (N_6476,N_6355,N_6257);
or U6477 (N_6477,N_6298,N_6379);
nand U6478 (N_6478,N_6392,N_6291);
or U6479 (N_6479,N_6359,N_6351);
xnor U6480 (N_6480,N_6269,N_6274);
or U6481 (N_6481,N_6290,N_6378);
and U6482 (N_6482,N_6309,N_6291);
nor U6483 (N_6483,N_6301,N_6366);
and U6484 (N_6484,N_6258,N_6317);
and U6485 (N_6485,N_6374,N_6262);
and U6486 (N_6486,N_6394,N_6279);
xor U6487 (N_6487,N_6310,N_6337);
and U6488 (N_6488,N_6372,N_6375);
nand U6489 (N_6489,N_6286,N_6306);
xor U6490 (N_6490,N_6366,N_6249);
and U6491 (N_6491,N_6295,N_6378);
xor U6492 (N_6492,N_6306,N_6292);
nand U6493 (N_6493,N_6297,N_6270);
and U6494 (N_6494,N_6381,N_6258);
nor U6495 (N_6495,N_6264,N_6368);
xor U6496 (N_6496,N_6294,N_6268);
and U6497 (N_6497,N_6306,N_6275);
xor U6498 (N_6498,N_6323,N_6295);
nor U6499 (N_6499,N_6252,N_6370);
xnor U6500 (N_6500,N_6256,N_6333);
nand U6501 (N_6501,N_6376,N_6241);
or U6502 (N_6502,N_6350,N_6278);
xor U6503 (N_6503,N_6392,N_6355);
nand U6504 (N_6504,N_6254,N_6360);
nand U6505 (N_6505,N_6251,N_6310);
and U6506 (N_6506,N_6380,N_6291);
or U6507 (N_6507,N_6332,N_6264);
nor U6508 (N_6508,N_6355,N_6351);
or U6509 (N_6509,N_6296,N_6395);
nand U6510 (N_6510,N_6285,N_6316);
nand U6511 (N_6511,N_6297,N_6394);
and U6512 (N_6512,N_6342,N_6245);
nand U6513 (N_6513,N_6380,N_6346);
and U6514 (N_6514,N_6327,N_6350);
nand U6515 (N_6515,N_6361,N_6380);
nor U6516 (N_6516,N_6338,N_6386);
nand U6517 (N_6517,N_6278,N_6279);
nand U6518 (N_6518,N_6336,N_6392);
xor U6519 (N_6519,N_6308,N_6367);
nand U6520 (N_6520,N_6322,N_6337);
nor U6521 (N_6521,N_6266,N_6291);
or U6522 (N_6522,N_6247,N_6321);
xnor U6523 (N_6523,N_6361,N_6337);
nand U6524 (N_6524,N_6322,N_6302);
and U6525 (N_6525,N_6296,N_6283);
nor U6526 (N_6526,N_6276,N_6267);
and U6527 (N_6527,N_6299,N_6363);
or U6528 (N_6528,N_6289,N_6276);
or U6529 (N_6529,N_6373,N_6388);
xor U6530 (N_6530,N_6344,N_6296);
or U6531 (N_6531,N_6265,N_6283);
and U6532 (N_6532,N_6346,N_6367);
xnor U6533 (N_6533,N_6296,N_6307);
or U6534 (N_6534,N_6395,N_6328);
nor U6535 (N_6535,N_6372,N_6283);
nand U6536 (N_6536,N_6255,N_6337);
nand U6537 (N_6537,N_6287,N_6354);
and U6538 (N_6538,N_6248,N_6259);
nand U6539 (N_6539,N_6343,N_6297);
nand U6540 (N_6540,N_6348,N_6250);
nor U6541 (N_6541,N_6355,N_6364);
nor U6542 (N_6542,N_6383,N_6254);
or U6543 (N_6543,N_6280,N_6379);
xnor U6544 (N_6544,N_6323,N_6268);
and U6545 (N_6545,N_6338,N_6319);
xnor U6546 (N_6546,N_6340,N_6251);
nor U6547 (N_6547,N_6386,N_6302);
nor U6548 (N_6548,N_6387,N_6271);
nand U6549 (N_6549,N_6380,N_6269);
xnor U6550 (N_6550,N_6261,N_6282);
or U6551 (N_6551,N_6264,N_6275);
or U6552 (N_6552,N_6306,N_6340);
nor U6553 (N_6553,N_6383,N_6370);
nand U6554 (N_6554,N_6271,N_6371);
nor U6555 (N_6555,N_6328,N_6282);
xnor U6556 (N_6556,N_6341,N_6278);
nand U6557 (N_6557,N_6399,N_6297);
nand U6558 (N_6558,N_6361,N_6332);
and U6559 (N_6559,N_6317,N_6268);
xor U6560 (N_6560,N_6535,N_6502);
or U6561 (N_6561,N_6423,N_6531);
nand U6562 (N_6562,N_6415,N_6500);
nor U6563 (N_6563,N_6449,N_6419);
nor U6564 (N_6564,N_6430,N_6557);
nand U6565 (N_6565,N_6468,N_6435);
nand U6566 (N_6566,N_6472,N_6559);
or U6567 (N_6567,N_6515,N_6479);
nand U6568 (N_6568,N_6474,N_6407);
nand U6569 (N_6569,N_6495,N_6492);
and U6570 (N_6570,N_6504,N_6544);
xor U6571 (N_6571,N_6409,N_6508);
nor U6572 (N_6572,N_6480,N_6408);
nor U6573 (N_6573,N_6525,N_6401);
nor U6574 (N_6574,N_6510,N_6484);
xnor U6575 (N_6575,N_6477,N_6455);
nor U6576 (N_6576,N_6530,N_6452);
or U6577 (N_6577,N_6436,N_6550);
or U6578 (N_6578,N_6505,N_6469);
xor U6579 (N_6579,N_6555,N_6412);
or U6580 (N_6580,N_6497,N_6417);
xor U6581 (N_6581,N_6503,N_6458);
nor U6582 (N_6582,N_6493,N_6533);
xor U6583 (N_6583,N_6486,N_6459);
or U6584 (N_6584,N_6438,N_6539);
nand U6585 (N_6585,N_6517,N_6463);
nor U6586 (N_6586,N_6487,N_6520);
xnor U6587 (N_6587,N_6519,N_6428);
nor U6588 (N_6588,N_6441,N_6432);
and U6589 (N_6589,N_6478,N_6437);
nand U6590 (N_6590,N_6473,N_6427);
and U6591 (N_6591,N_6498,N_6558);
nand U6592 (N_6592,N_6470,N_6462);
and U6593 (N_6593,N_6461,N_6434);
nor U6594 (N_6594,N_6414,N_6481);
nand U6595 (N_6595,N_6464,N_6451);
nand U6596 (N_6596,N_6526,N_6482);
and U6597 (N_6597,N_6400,N_6460);
or U6598 (N_6598,N_6444,N_6418);
or U6599 (N_6599,N_6507,N_6411);
or U6600 (N_6600,N_6522,N_6521);
nand U6601 (N_6601,N_6466,N_6440);
nor U6602 (N_6602,N_6406,N_6552);
nor U6603 (N_6603,N_6403,N_6532);
and U6604 (N_6604,N_6446,N_6516);
or U6605 (N_6605,N_6404,N_6511);
or U6606 (N_6606,N_6546,N_6524);
and U6607 (N_6607,N_6547,N_6485);
or U6608 (N_6608,N_6410,N_6433);
nand U6609 (N_6609,N_6431,N_6443);
and U6610 (N_6610,N_6529,N_6422);
nand U6611 (N_6611,N_6534,N_6509);
nand U6612 (N_6612,N_6402,N_6556);
and U6613 (N_6613,N_6499,N_6513);
nand U6614 (N_6614,N_6551,N_6537);
and U6615 (N_6615,N_6442,N_6545);
nor U6616 (N_6616,N_6483,N_6501);
xnor U6617 (N_6617,N_6540,N_6439);
nor U6618 (N_6618,N_6506,N_6548);
nor U6619 (N_6619,N_6528,N_6457);
nor U6620 (N_6620,N_6543,N_6518);
nand U6621 (N_6621,N_6512,N_6448);
xnor U6622 (N_6622,N_6514,N_6475);
nor U6623 (N_6623,N_6421,N_6405);
and U6624 (N_6624,N_6496,N_6488);
xor U6625 (N_6625,N_6447,N_6453);
xor U6626 (N_6626,N_6541,N_6527);
nor U6627 (N_6627,N_6420,N_6476);
xor U6628 (N_6628,N_6465,N_6554);
nor U6629 (N_6629,N_6456,N_6549);
or U6630 (N_6630,N_6413,N_6490);
xnor U6631 (N_6631,N_6424,N_6553);
nor U6632 (N_6632,N_6454,N_6467);
and U6633 (N_6633,N_6450,N_6538);
and U6634 (N_6634,N_6489,N_6491);
nand U6635 (N_6635,N_6494,N_6429);
nand U6636 (N_6636,N_6536,N_6445);
xor U6637 (N_6637,N_6425,N_6416);
xnor U6638 (N_6638,N_6426,N_6471);
xor U6639 (N_6639,N_6542,N_6523);
xnor U6640 (N_6640,N_6434,N_6533);
nand U6641 (N_6641,N_6521,N_6420);
xnor U6642 (N_6642,N_6419,N_6464);
and U6643 (N_6643,N_6430,N_6411);
nand U6644 (N_6644,N_6441,N_6525);
or U6645 (N_6645,N_6404,N_6531);
xnor U6646 (N_6646,N_6535,N_6523);
nor U6647 (N_6647,N_6503,N_6525);
xor U6648 (N_6648,N_6475,N_6554);
nor U6649 (N_6649,N_6532,N_6530);
and U6650 (N_6650,N_6460,N_6405);
and U6651 (N_6651,N_6401,N_6454);
nor U6652 (N_6652,N_6485,N_6526);
and U6653 (N_6653,N_6460,N_6434);
or U6654 (N_6654,N_6443,N_6515);
or U6655 (N_6655,N_6552,N_6428);
or U6656 (N_6656,N_6513,N_6557);
xor U6657 (N_6657,N_6554,N_6409);
nand U6658 (N_6658,N_6426,N_6552);
nand U6659 (N_6659,N_6460,N_6556);
nor U6660 (N_6660,N_6456,N_6510);
and U6661 (N_6661,N_6437,N_6454);
nor U6662 (N_6662,N_6424,N_6491);
or U6663 (N_6663,N_6529,N_6501);
or U6664 (N_6664,N_6508,N_6454);
or U6665 (N_6665,N_6553,N_6471);
and U6666 (N_6666,N_6438,N_6517);
nor U6667 (N_6667,N_6447,N_6516);
or U6668 (N_6668,N_6450,N_6462);
nand U6669 (N_6669,N_6476,N_6417);
or U6670 (N_6670,N_6409,N_6513);
or U6671 (N_6671,N_6487,N_6470);
nor U6672 (N_6672,N_6502,N_6459);
xnor U6673 (N_6673,N_6461,N_6553);
nor U6674 (N_6674,N_6410,N_6471);
nor U6675 (N_6675,N_6434,N_6527);
nor U6676 (N_6676,N_6460,N_6517);
and U6677 (N_6677,N_6496,N_6555);
or U6678 (N_6678,N_6544,N_6470);
and U6679 (N_6679,N_6405,N_6428);
nor U6680 (N_6680,N_6468,N_6423);
nor U6681 (N_6681,N_6409,N_6434);
and U6682 (N_6682,N_6405,N_6534);
xnor U6683 (N_6683,N_6548,N_6403);
or U6684 (N_6684,N_6400,N_6409);
nor U6685 (N_6685,N_6468,N_6535);
xor U6686 (N_6686,N_6458,N_6417);
and U6687 (N_6687,N_6524,N_6400);
and U6688 (N_6688,N_6524,N_6443);
or U6689 (N_6689,N_6557,N_6521);
and U6690 (N_6690,N_6547,N_6534);
nor U6691 (N_6691,N_6435,N_6497);
nand U6692 (N_6692,N_6525,N_6522);
or U6693 (N_6693,N_6460,N_6472);
nor U6694 (N_6694,N_6484,N_6534);
nand U6695 (N_6695,N_6507,N_6510);
xor U6696 (N_6696,N_6417,N_6483);
xor U6697 (N_6697,N_6419,N_6478);
nor U6698 (N_6698,N_6460,N_6468);
xnor U6699 (N_6699,N_6494,N_6471);
nor U6700 (N_6700,N_6453,N_6487);
or U6701 (N_6701,N_6485,N_6428);
xnor U6702 (N_6702,N_6436,N_6492);
or U6703 (N_6703,N_6404,N_6549);
and U6704 (N_6704,N_6536,N_6558);
nor U6705 (N_6705,N_6506,N_6424);
xnor U6706 (N_6706,N_6504,N_6401);
xnor U6707 (N_6707,N_6466,N_6443);
or U6708 (N_6708,N_6403,N_6433);
nor U6709 (N_6709,N_6459,N_6420);
nor U6710 (N_6710,N_6530,N_6431);
nand U6711 (N_6711,N_6404,N_6558);
or U6712 (N_6712,N_6490,N_6547);
and U6713 (N_6713,N_6503,N_6427);
and U6714 (N_6714,N_6400,N_6503);
xor U6715 (N_6715,N_6555,N_6413);
xnor U6716 (N_6716,N_6461,N_6474);
and U6717 (N_6717,N_6418,N_6441);
nor U6718 (N_6718,N_6507,N_6485);
nor U6719 (N_6719,N_6552,N_6401);
and U6720 (N_6720,N_6697,N_6662);
nand U6721 (N_6721,N_6702,N_6581);
nor U6722 (N_6722,N_6578,N_6604);
or U6723 (N_6723,N_6677,N_6717);
or U6724 (N_6724,N_6715,N_6563);
or U6725 (N_6725,N_6709,N_6653);
and U6726 (N_6726,N_6634,N_6647);
xor U6727 (N_6727,N_6703,N_6659);
or U6728 (N_6728,N_6620,N_6698);
xor U6729 (N_6729,N_6590,N_6665);
xor U6730 (N_6730,N_6585,N_6638);
or U6731 (N_6731,N_6577,N_6694);
and U6732 (N_6732,N_6627,N_6615);
xnor U6733 (N_6733,N_6716,N_6654);
nand U6734 (N_6734,N_6586,N_6598);
xnor U6735 (N_6735,N_6648,N_6655);
nand U6736 (N_6736,N_6616,N_6688);
and U6737 (N_6737,N_6641,N_6631);
xnor U6738 (N_6738,N_6678,N_6574);
or U6739 (N_6739,N_6672,N_6576);
xor U6740 (N_6740,N_6630,N_6658);
nand U6741 (N_6741,N_6637,N_6711);
nor U6742 (N_6742,N_6568,N_6707);
xor U6743 (N_6743,N_6593,N_6679);
nor U6744 (N_6744,N_6676,N_6691);
nor U6745 (N_6745,N_6583,N_6609);
xnor U6746 (N_6746,N_6696,N_6569);
and U6747 (N_6747,N_6682,N_6644);
xnor U6748 (N_6748,N_6596,N_6700);
or U6749 (N_6749,N_6614,N_6708);
or U6750 (N_6750,N_6610,N_6626);
or U6751 (N_6751,N_6690,N_6680);
nor U6752 (N_6752,N_6719,N_6608);
and U6753 (N_6753,N_6618,N_6589);
nand U6754 (N_6754,N_6623,N_6571);
nor U6755 (N_6755,N_6668,N_6600);
nor U6756 (N_6756,N_6591,N_6612);
and U6757 (N_6757,N_6692,N_6642);
xnor U6758 (N_6758,N_6613,N_6718);
and U6759 (N_6759,N_6663,N_6617);
nand U6760 (N_6760,N_6671,N_6652);
or U6761 (N_6761,N_6628,N_6588);
xor U6762 (N_6762,N_6629,N_6649);
or U6763 (N_6763,N_6584,N_6602);
or U6764 (N_6764,N_6687,N_6689);
and U6765 (N_6765,N_6575,N_6666);
nor U6766 (N_6766,N_6695,N_6566);
and U6767 (N_6767,N_6660,N_6664);
nand U6768 (N_6768,N_6714,N_6639);
nand U6769 (N_6769,N_6673,N_6632);
nand U6770 (N_6770,N_6640,N_6651);
or U6771 (N_6771,N_6636,N_6699);
or U6772 (N_6772,N_6607,N_6560);
nor U6773 (N_6773,N_6624,N_6562);
and U6774 (N_6774,N_6683,N_6580);
and U6775 (N_6775,N_6594,N_6669);
and U6776 (N_6776,N_6592,N_6572);
xnor U6777 (N_6777,N_6643,N_6595);
or U6778 (N_6778,N_6605,N_6667);
nand U6779 (N_6779,N_6701,N_6582);
nor U6780 (N_6780,N_6684,N_6706);
nor U6781 (N_6781,N_6603,N_6599);
or U6782 (N_6782,N_6573,N_6674);
or U6783 (N_6783,N_6681,N_6661);
nor U6784 (N_6784,N_6686,N_6650);
and U6785 (N_6785,N_6635,N_6567);
xnor U6786 (N_6786,N_6633,N_6564);
or U6787 (N_6787,N_6646,N_6685);
xor U6788 (N_6788,N_6579,N_6621);
xor U6789 (N_6789,N_6675,N_6587);
nor U6790 (N_6790,N_6565,N_6645);
and U6791 (N_6791,N_6622,N_6670);
and U6792 (N_6792,N_6597,N_6712);
nor U6793 (N_6793,N_6713,N_6611);
or U6794 (N_6794,N_6625,N_6705);
nand U6795 (N_6795,N_6656,N_6693);
nor U6796 (N_6796,N_6570,N_6561);
xnor U6797 (N_6797,N_6657,N_6710);
and U6798 (N_6798,N_6619,N_6606);
nor U6799 (N_6799,N_6704,N_6601);
nor U6800 (N_6800,N_6711,N_6587);
or U6801 (N_6801,N_6649,N_6576);
nor U6802 (N_6802,N_6687,N_6597);
or U6803 (N_6803,N_6609,N_6594);
and U6804 (N_6804,N_6638,N_6624);
or U6805 (N_6805,N_6704,N_6642);
nand U6806 (N_6806,N_6644,N_6563);
nand U6807 (N_6807,N_6579,N_6612);
nand U6808 (N_6808,N_6619,N_6589);
nor U6809 (N_6809,N_6578,N_6651);
nor U6810 (N_6810,N_6683,N_6622);
and U6811 (N_6811,N_6716,N_6594);
or U6812 (N_6812,N_6698,N_6713);
nand U6813 (N_6813,N_6717,N_6567);
and U6814 (N_6814,N_6670,N_6712);
nand U6815 (N_6815,N_6679,N_6578);
and U6816 (N_6816,N_6672,N_6696);
or U6817 (N_6817,N_6714,N_6679);
nor U6818 (N_6818,N_6699,N_6579);
and U6819 (N_6819,N_6577,N_6573);
nor U6820 (N_6820,N_6651,N_6596);
nand U6821 (N_6821,N_6610,N_6571);
and U6822 (N_6822,N_6716,N_6616);
or U6823 (N_6823,N_6677,N_6574);
and U6824 (N_6824,N_6567,N_6580);
nor U6825 (N_6825,N_6652,N_6567);
xnor U6826 (N_6826,N_6592,N_6631);
and U6827 (N_6827,N_6592,N_6663);
nand U6828 (N_6828,N_6633,N_6662);
and U6829 (N_6829,N_6622,N_6578);
or U6830 (N_6830,N_6598,N_6705);
nand U6831 (N_6831,N_6560,N_6599);
nand U6832 (N_6832,N_6615,N_6569);
nand U6833 (N_6833,N_6582,N_6675);
xor U6834 (N_6834,N_6685,N_6591);
or U6835 (N_6835,N_6715,N_6622);
nor U6836 (N_6836,N_6616,N_6642);
nor U6837 (N_6837,N_6674,N_6591);
and U6838 (N_6838,N_6614,N_6714);
nand U6839 (N_6839,N_6674,N_6669);
xor U6840 (N_6840,N_6637,N_6640);
or U6841 (N_6841,N_6643,N_6565);
nor U6842 (N_6842,N_6623,N_6609);
nand U6843 (N_6843,N_6561,N_6630);
xnor U6844 (N_6844,N_6610,N_6642);
and U6845 (N_6845,N_6686,N_6708);
and U6846 (N_6846,N_6658,N_6674);
nor U6847 (N_6847,N_6699,N_6715);
xor U6848 (N_6848,N_6651,N_6575);
or U6849 (N_6849,N_6709,N_6676);
or U6850 (N_6850,N_6562,N_6697);
and U6851 (N_6851,N_6679,N_6658);
and U6852 (N_6852,N_6591,N_6682);
xor U6853 (N_6853,N_6678,N_6659);
nand U6854 (N_6854,N_6686,N_6628);
or U6855 (N_6855,N_6718,N_6620);
nand U6856 (N_6856,N_6584,N_6714);
or U6857 (N_6857,N_6621,N_6715);
and U6858 (N_6858,N_6697,N_6695);
nand U6859 (N_6859,N_6624,N_6567);
nand U6860 (N_6860,N_6603,N_6676);
xor U6861 (N_6861,N_6598,N_6627);
or U6862 (N_6862,N_6669,N_6617);
nand U6863 (N_6863,N_6681,N_6704);
nand U6864 (N_6864,N_6607,N_6657);
and U6865 (N_6865,N_6595,N_6623);
and U6866 (N_6866,N_6697,N_6593);
and U6867 (N_6867,N_6644,N_6589);
and U6868 (N_6868,N_6646,N_6589);
xnor U6869 (N_6869,N_6609,N_6603);
and U6870 (N_6870,N_6693,N_6718);
nand U6871 (N_6871,N_6682,N_6618);
nor U6872 (N_6872,N_6645,N_6561);
and U6873 (N_6873,N_6613,N_6603);
nor U6874 (N_6874,N_6644,N_6717);
xor U6875 (N_6875,N_6560,N_6626);
nand U6876 (N_6876,N_6644,N_6659);
xnor U6877 (N_6877,N_6595,N_6612);
and U6878 (N_6878,N_6616,N_6675);
xor U6879 (N_6879,N_6593,N_6592);
or U6880 (N_6880,N_6872,N_6794);
xor U6881 (N_6881,N_6727,N_6821);
nand U6882 (N_6882,N_6808,N_6789);
xor U6883 (N_6883,N_6877,N_6744);
xor U6884 (N_6884,N_6871,N_6737);
and U6885 (N_6885,N_6866,N_6743);
and U6886 (N_6886,N_6762,N_6764);
nor U6887 (N_6887,N_6813,N_6878);
xnor U6888 (N_6888,N_6766,N_6859);
and U6889 (N_6889,N_6775,N_6782);
nor U6890 (N_6890,N_6822,N_6779);
nor U6891 (N_6891,N_6752,N_6805);
and U6892 (N_6892,N_6834,N_6863);
or U6893 (N_6893,N_6853,N_6826);
xor U6894 (N_6894,N_6824,N_6765);
xor U6895 (N_6895,N_6786,N_6799);
or U6896 (N_6896,N_6839,N_6759);
nor U6897 (N_6897,N_6725,N_6770);
and U6898 (N_6898,N_6778,N_6795);
xnor U6899 (N_6899,N_6849,N_6723);
nand U6900 (N_6900,N_6784,N_6800);
and U6901 (N_6901,N_6817,N_6865);
nand U6902 (N_6902,N_6857,N_6787);
and U6903 (N_6903,N_6746,N_6769);
and U6904 (N_6904,N_6736,N_6793);
xnor U6905 (N_6905,N_6850,N_6753);
nor U6906 (N_6906,N_6831,N_6829);
nand U6907 (N_6907,N_6875,N_6721);
nor U6908 (N_6908,N_6830,N_6856);
or U6909 (N_6909,N_6855,N_6814);
xnor U6910 (N_6910,N_6873,N_6798);
or U6911 (N_6911,N_6861,N_6760);
nor U6912 (N_6912,N_6734,N_6869);
nand U6913 (N_6913,N_6776,N_6748);
nand U6914 (N_6914,N_6858,N_6722);
nand U6915 (N_6915,N_6728,N_6809);
nor U6916 (N_6916,N_6754,N_6763);
or U6917 (N_6917,N_6772,N_6726);
nor U6918 (N_6918,N_6720,N_6806);
and U6919 (N_6919,N_6832,N_6788);
xor U6920 (N_6920,N_6835,N_6796);
nand U6921 (N_6921,N_6874,N_6774);
xor U6922 (N_6922,N_6843,N_6845);
or U6923 (N_6923,N_6867,N_6815);
or U6924 (N_6924,N_6847,N_6876);
nor U6925 (N_6925,N_6757,N_6783);
xor U6926 (N_6926,N_6724,N_6749);
nand U6927 (N_6927,N_6758,N_6823);
xnor U6928 (N_6928,N_6862,N_6818);
or U6929 (N_6929,N_6739,N_6750);
and U6930 (N_6930,N_6785,N_6828);
nand U6931 (N_6931,N_6846,N_6836);
xor U6932 (N_6932,N_6820,N_6802);
and U6933 (N_6933,N_6860,N_6851);
nand U6934 (N_6934,N_6768,N_6837);
nand U6935 (N_6935,N_6792,N_6740);
or U6936 (N_6936,N_6733,N_6790);
and U6937 (N_6937,N_6825,N_6868);
or U6938 (N_6938,N_6730,N_6747);
and U6939 (N_6939,N_6797,N_6767);
nand U6940 (N_6940,N_6870,N_6780);
or U6941 (N_6941,N_6854,N_6738);
nand U6942 (N_6942,N_6741,N_6755);
nand U6943 (N_6943,N_6864,N_6731);
or U6944 (N_6944,N_6751,N_6841);
nand U6945 (N_6945,N_6807,N_6848);
nor U6946 (N_6946,N_6819,N_6777);
or U6947 (N_6947,N_6742,N_6781);
and U6948 (N_6948,N_6810,N_6801);
nand U6949 (N_6949,N_6804,N_6827);
or U6950 (N_6950,N_6840,N_6852);
and U6951 (N_6951,N_6879,N_6756);
nand U6952 (N_6952,N_6812,N_6745);
nor U6953 (N_6953,N_6735,N_6842);
and U6954 (N_6954,N_6761,N_6732);
or U6955 (N_6955,N_6844,N_6803);
and U6956 (N_6956,N_6816,N_6833);
nand U6957 (N_6957,N_6773,N_6771);
and U6958 (N_6958,N_6838,N_6729);
nand U6959 (N_6959,N_6811,N_6791);
nand U6960 (N_6960,N_6765,N_6796);
nor U6961 (N_6961,N_6844,N_6848);
xor U6962 (N_6962,N_6787,N_6792);
xnor U6963 (N_6963,N_6749,N_6855);
or U6964 (N_6964,N_6723,N_6821);
nand U6965 (N_6965,N_6773,N_6873);
and U6966 (N_6966,N_6864,N_6818);
xor U6967 (N_6967,N_6826,N_6869);
or U6968 (N_6968,N_6751,N_6800);
or U6969 (N_6969,N_6741,N_6810);
nor U6970 (N_6970,N_6724,N_6763);
nand U6971 (N_6971,N_6848,N_6783);
or U6972 (N_6972,N_6720,N_6745);
and U6973 (N_6973,N_6864,N_6754);
and U6974 (N_6974,N_6807,N_6736);
xor U6975 (N_6975,N_6754,N_6866);
nand U6976 (N_6976,N_6871,N_6738);
nand U6977 (N_6977,N_6858,N_6794);
or U6978 (N_6978,N_6772,N_6783);
nor U6979 (N_6979,N_6807,N_6767);
or U6980 (N_6980,N_6727,N_6753);
and U6981 (N_6981,N_6789,N_6778);
or U6982 (N_6982,N_6801,N_6816);
nand U6983 (N_6983,N_6854,N_6856);
or U6984 (N_6984,N_6764,N_6868);
and U6985 (N_6985,N_6857,N_6845);
nor U6986 (N_6986,N_6793,N_6772);
nand U6987 (N_6987,N_6866,N_6863);
nor U6988 (N_6988,N_6835,N_6842);
nor U6989 (N_6989,N_6816,N_6791);
or U6990 (N_6990,N_6813,N_6746);
xor U6991 (N_6991,N_6745,N_6792);
nand U6992 (N_6992,N_6786,N_6751);
and U6993 (N_6993,N_6762,N_6746);
nand U6994 (N_6994,N_6812,N_6818);
and U6995 (N_6995,N_6878,N_6756);
xnor U6996 (N_6996,N_6809,N_6784);
nor U6997 (N_6997,N_6812,N_6848);
nor U6998 (N_6998,N_6782,N_6752);
xor U6999 (N_6999,N_6862,N_6742);
nand U7000 (N_7000,N_6733,N_6846);
or U7001 (N_7001,N_6822,N_6774);
xnor U7002 (N_7002,N_6860,N_6843);
or U7003 (N_7003,N_6823,N_6769);
or U7004 (N_7004,N_6785,N_6846);
xnor U7005 (N_7005,N_6720,N_6812);
nand U7006 (N_7006,N_6874,N_6768);
and U7007 (N_7007,N_6808,N_6752);
or U7008 (N_7008,N_6834,N_6747);
nor U7009 (N_7009,N_6829,N_6810);
nor U7010 (N_7010,N_6769,N_6779);
nand U7011 (N_7011,N_6765,N_6811);
and U7012 (N_7012,N_6842,N_6818);
or U7013 (N_7013,N_6869,N_6857);
nor U7014 (N_7014,N_6749,N_6803);
nand U7015 (N_7015,N_6731,N_6728);
and U7016 (N_7016,N_6852,N_6744);
nand U7017 (N_7017,N_6774,N_6766);
xnor U7018 (N_7018,N_6757,N_6879);
nor U7019 (N_7019,N_6812,N_6838);
nor U7020 (N_7020,N_6756,N_6843);
nor U7021 (N_7021,N_6784,N_6859);
or U7022 (N_7022,N_6770,N_6802);
and U7023 (N_7023,N_6865,N_6748);
and U7024 (N_7024,N_6728,N_6830);
or U7025 (N_7025,N_6788,N_6878);
nor U7026 (N_7026,N_6791,N_6817);
or U7027 (N_7027,N_6863,N_6741);
and U7028 (N_7028,N_6747,N_6736);
xnor U7029 (N_7029,N_6742,N_6739);
or U7030 (N_7030,N_6770,N_6750);
nand U7031 (N_7031,N_6862,N_6775);
xnor U7032 (N_7032,N_6819,N_6807);
or U7033 (N_7033,N_6734,N_6848);
xnor U7034 (N_7034,N_6873,N_6746);
xor U7035 (N_7035,N_6773,N_6865);
nand U7036 (N_7036,N_6843,N_6876);
or U7037 (N_7037,N_6845,N_6725);
nor U7038 (N_7038,N_6849,N_6798);
nand U7039 (N_7039,N_6797,N_6788);
nor U7040 (N_7040,N_6925,N_7028);
or U7041 (N_7041,N_6885,N_6974);
nor U7042 (N_7042,N_7001,N_7035);
or U7043 (N_7043,N_6973,N_6921);
or U7044 (N_7044,N_6993,N_6918);
or U7045 (N_7045,N_6992,N_6898);
nor U7046 (N_7046,N_6887,N_6984);
nor U7047 (N_7047,N_6946,N_6922);
nor U7048 (N_7048,N_6965,N_6915);
xnor U7049 (N_7049,N_6935,N_6884);
and U7050 (N_7050,N_6897,N_6889);
nor U7051 (N_7051,N_6972,N_7003);
or U7052 (N_7052,N_6957,N_6987);
xor U7053 (N_7053,N_6999,N_6967);
nand U7054 (N_7054,N_6942,N_6986);
and U7055 (N_7055,N_6929,N_6933);
or U7056 (N_7056,N_7005,N_7026);
and U7057 (N_7057,N_6907,N_7002);
nor U7058 (N_7058,N_7023,N_6882);
and U7059 (N_7059,N_6940,N_7025);
nand U7060 (N_7060,N_7006,N_6880);
xnor U7061 (N_7061,N_6969,N_6980);
xnor U7062 (N_7062,N_6910,N_7018);
nor U7063 (N_7063,N_6961,N_7016);
xor U7064 (N_7064,N_6888,N_6890);
nor U7065 (N_7065,N_7022,N_7024);
and U7066 (N_7066,N_6923,N_7019);
nand U7067 (N_7067,N_6904,N_7036);
or U7068 (N_7068,N_6902,N_6892);
nand U7069 (N_7069,N_6894,N_7034);
or U7070 (N_7070,N_6954,N_6928);
nor U7071 (N_7071,N_6883,N_6951);
nor U7072 (N_7072,N_7038,N_6891);
and U7073 (N_7073,N_6909,N_6962);
or U7074 (N_7074,N_6955,N_7017);
and U7075 (N_7075,N_6994,N_6989);
xor U7076 (N_7076,N_6964,N_6938);
nand U7077 (N_7077,N_7030,N_6943);
xnor U7078 (N_7078,N_6930,N_6982);
xnor U7079 (N_7079,N_6977,N_6952);
or U7080 (N_7080,N_6949,N_6997);
xnor U7081 (N_7081,N_7033,N_7029);
xor U7082 (N_7082,N_7004,N_6975);
or U7083 (N_7083,N_6916,N_6966);
nor U7084 (N_7084,N_6926,N_6939);
or U7085 (N_7085,N_6908,N_6895);
xnor U7086 (N_7086,N_6995,N_7011);
nor U7087 (N_7087,N_6886,N_7031);
nor U7088 (N_7088,N_6920,N_6936);
xor U7089 (N_7089,N_6927,N_6953);
nor U7090 (N_7090,N_7009,N_6959);
xnor U7091 (N_7091,N_6978,N_6913);
nand U7092 (N_7092,N_6896,N_6996);
or U7093 (N_7093,N_6899,N_6998);
nor U7094 (N_7094,N_6917,N_7027);
xnor U7095 (N_7095,N_6893,N_7020);
nor U7096 (N_7096,N_7007,N_6937);
and U7097 (N_7097,N_7032,N_6970);
and U7098 (N_7098,N_6941,N_7000);
nor U7099 (N_7099,N_6911,N_6905);
or U7100 (N_7100,N_7039,N_6968);
and U7101 (N_7101,N_6932,N_6956);
or U7102 (N_7102,N_6919,N_6990);
xnor U7103 (N_7103,N_6924,N_6948);
nand U7104 (N_7104,N_6981,N_7021);
xor U7105 (N_7105,N_6963,N_6903);
xor U7106 (N_7106,N_6881,N_7037);
and U7107 (N_7107,N_6979,N_6914);
xor U7108 (N_7108,N_6985,N_7013);
and U7109 (N_7109,N_6988,N_6958);
and U7110 (N_7110,N_6945,N_6971);
or U7111 (N_7111,N_6960,N_7010);
or U7112 (N_7112,N_6912,N_6991);
nor U7113 (N_7113,N_6931,N_6976);
xor U7114 (N_7114,N_7012,N_6947);
or U7115 (N_7115,N_6950,N_6901);
and U7116 (N_7116,N_7014,N_6934);
or U7117 (N_7117,N_7008,N_6900);
nand U7118 (N_7118,N_6983,N_6944);
and U7119 (N_7119,N_6906,N_7015);
and U7120 (N_7120,N_6971,N_7021);
and U7121 (N_7121,N_6921,N_6892);
or U7122 (N_7122,N_6886,N_6899);
and U7123 (N_7123,N_6962,N_7033);
nor U7124 (N_7124,N_6924,N_6919);
xor U7125 (N_7125,N_7023,N_6908);
or U7126 (N_7126,N_6955,N_6941);
xnor U7127 (N_7127,N_6944,N_6954);
nor U7128 (N_7128,N_6909,N_7036);
nor U7129 (N_7129,N_6979,N_7039);
nand U7130 (N_7130,N_6897,N_6894);
xor U7131 (N_7131,N_6953,N_6971);
nand U7132 (N_7132,N_6886,N_6918);
nand U7133 (N_7133,N_6892,N_6981);
nor U7134 (N_7134,N_6940,N_6964);
nand U7135 (N_7135,N_6999,N_6894);
nand U7136 (N_7136,N_6976,N_7037);
xnor U7137 (N_7137,N_6973,N_6994);
nand U7138 (N_7138,N_6923,N_6919);
or U7139 (N_7139,N_6988,N_7020);
nand U7140 (N_7140,N_6896,N_6939);
xnor U7141 (N_7141,N_6880,N_6962);
nand U7142 (N_7142,N_6984,N_6965);
nor U7143 (N_7143,N_7020,N_6931);
or U7144 (N_7144,N_7026,N_6966);
and U7145 (N_7145,N_6885,N_6944);
nor U7146 (N_7146,N_6956,N_7019);
or U7147 (N_7147,N_7012,N_6948);
and U7148 (N_7148,N_7039,N_6933);
xnor U7149 (N_7149,N_7030,N_7039);
nor U7150 (N_7150,N_6900,N_6952);
nand U7151 (N_7151,N_6965,N_6922);
nor U7152 (N_7152,N_7037,N_7000);
or U7153 (N_7153,N_6890,N_6936);
xnor U7154 (N_7154,N_7030,N_6954);
xnor U7155 (N_7155,N_6931,N_7009);
or U7156 (N_7156,N_6901,N_6973);
nor U7157 (N_7157,N_6929,N_7030);
nand U7158 (N_7158,N_6880,N_6939);
xor U7159 (N_7159,N_7036,N_6992);
nand U7160 (N_7160,N_7020,N_6961);
and U7161 (N_7161,N_6931,N_6982);
nor U7162 (N_7162,N_6992,N_7017);
nor U7163 (N_7163,N_6983,N_6961);
and U7164 (N_7164,N_6965,N_6912);
nor U7165 (N_7165,N_6889,N_7019);
or U7166 (N_7166,N_7003,N_7016);
or U7167 (N_7167,N_6882,N_7021);
nor U7168 (N_7168,N_6914,N_7006);
nor U7169 (N_7169,N_6958,N_6881);
nor U7170 (N_7170,N_7009,N_6955);
or U7171 (N_7171,N_7008,N_7033);
or U7172 (N_7172,N_7024,N_6965);
and U7173 (N_7173,N_6958,N_6885);
or U7174 (N_7174,N_6883,N_6965);
and U7175 (N_7175,N_7033,N_7030);
nor U7176 (N_7176,N_6983,N_6895);
xnor U7177 (N_7177,N_6892,N_7026);
xor U7178 (N_7178,N_7006,N_6925);
or U7179 (N_7179,N_7014,N_6944);
nand U7180 (N_7180,N_6899,N_6936);
nor U7181 (N_7181,N_6969,N_6894);
xnor U7182 (N_7182,N_6967,N_7034);
xnor U7183 (N_7183,N_6913,N_6905);
nand U7184 (N_7184,N_7035,N_6943);
or U7185 (N_7185,N_6882,N_7003);
or U7186 (N_7186,N_7038,N_6905);
and U7187 (N_7187,N_6927,N_6980);
xnor U7188 (N_7188,N_6927,N_6933);
xor U7189 (N_7189,N_7007,N_6995);
xor U7190 (N_7190,N_6985,N_7021);
and U7191 (N_7191,N_6880,N_6908);
or U7192 (N_7192,N_6936,N_6952);
xor U7193 (N_7193,N_6884,N_7002);
nand U7194 (N_7194,N_6983,N_6984);
nand U7195 (N_7195,N_6955,N_7030);
nor U7196 (N_7196,N_7008,N_6893);
xor U7197 (N_7197,N_6979,N_7033);
nand U7198 (N_7198,N_6905,N_7004);
and U7199 (N_7199,N_6906,N_6949);
nor U7200 (N_7200,N_7194,N_7070);
nor U7201 (N_7201,N_7087,N_7051);
and U7202 (N_7202,N_7045,N_7074);
and U7203 (N_7203,N_7112,N_7047);
and U7204 (N_7204,N_7135,N_7115);
and U7205 (N_7205,N_7056,N_7170);
xnor U7206 (N_7206,N_7119,N_7108);
xor U7207 (N_7207,N_7175,N_7173);
nand U7208 (N_7208,N_7188,N_7198);
and U7209 (N_7209,N_7063,N_7163);
xnor U7210 (N_7210,N_7088,N_7094);
or U7211 (N_7211,N_7090,N_7145);
or U7212 (N_7212,N_7158,N_7162);
xnor U7213 (N_7213,N_7059,N_7103);
nand U7214 (N_7214,N_7072,N_7075);
or U7215 (N_7215,N_7091,N_7079);
nand U7216 (N_7216,N_7101,N_7160);
nand U7217 (N_7217,N_7132,N_7180);
xnor U7218 (N_7218,N_7073,N_7062);
nand U7219 (N_7219,N_7143,N_7078);
nand U7220 (N_7220,N_7191,N_7176);
and U7221 (N_7221,N_7076,N_7092);
and U7222 (N_7222,N_7152,N_7129);
xor U7223 (N_7223,N_7081,N_7064);
and U7224 (N_7224,N_7043,N_7124);
xnor U7225 (N_7225,N_7077,N_7041);
xor U7226 (N_7226,N_7100,N_7055);
or U7227 (N_7227,N_7057,N_7084);
xnor U7228 (N_7228,N_7172,N_7099);
nor U7229 (N_7229,N_7053,N_7161);
nand U7230 (N_7230,N_7187,N_7146);
and U7231 (N_7231,N_7111,N_7089);
nand U7232 (N_7232,N_7167,N_7104);
nand U7233 (N_7233,N_7121,N_7102);
nor U7234 (N_7234,N_7181,N_7114);
nor U7235 (N_7235,N_7110,N_7131);
and U7236 (N_7236,N_7117,N_7159);
nor U7237 (N_7237,N_7066,N_7154);
xnor U7238 (N_7238,N_7040,N_7182);
and U7239 (N_7239,N_7148,N_7106);
xnor U7240 (N_7240,N_7179,N_7085);
and U7241 (N_7241,N_7127,N_7177);
xnor U7242 (N_7242,N_7046,N_7137);
or U7243 (N_7243,N_7061,N_7150);
nor U7244 (N_7244,N_7171,N_7196);
and U7245 (N_7245,N_7098,N_7123);
and U7246 (N_7246,N_7133,N_7060);
nor U7247 (N_7247,N_7164,N_7178);
xnor U7248 (N_7248,N_7107,N_7149);
and U7249 (N_7249,N_7120,N_7130);
nand U7250 (N_7250,N_7096,N_7156);
xnor U7251 (N_7251,N_7097,N_7122);
nor U7252 (N_7252,N_7193,N_7069);
or U7253 (N_7253,N_7139,N_7184);
and U7254 (N_7254,N_7195,N_7197);
xnor U7255 (N_7255,N_7199,N_7168);
or U7256 (N_7256,N_7109,N_7189);
and U7257 (N_7257,N_7080,N_7153);
xnor U7258 (N_7258,N_7065,N_7050);
nand U7259 (N_7259,N_7042,N_7138);
xor U7260 (N_7260,N_7141,N_7067);
nor U7261 (N_7261,N_7174,N_7165);
nor U7262 (N_7262,N_7048,N_7113);
or U7263 (N_7263,N_7157,N_7058);
xnor U7264 (N_7264,N_7169,N_7068);
xnor U7265 (N_7265,N_7126,N_7142);
nand U7266 (N_7266,N_7155,N_7044);
nor U7267 (N_7267,N_7190,N_7093);
and U7268 (N_7268,N_7125,N_7049);
nand U7269 (N_7269,N_7186,N_7086);
and U7270 (N_7270,N_7083,N_7134);
or U7271 (N_7271,N_7147,N_7166);
xnor U7272 (N_7272,N_7136,N_7082);
or U7273 (N_7273,N_7151,N_7105);
and U7274 (N_7274,N_7140,N_7144);
nor U7275 (N_7275,N_7052,N_7185);
xor U7276 (N_7276,N_7071,N_7128);
nor U7277 (N_7277,N_7095,N_7116);
nand U7278 (N_7278,N_7118,N_7054);
and U7279 (N_7279,N_7192,N_7183);
or U7280 (N_7280,N_7140,N_7164);
xnor U7281 (N_7281,N_7168,N_7151);
and U7282 (N_7282,N_7167,N_7127);
nor U7283 (N_7283,N_7054,N_7148);
or U7284 (N_7284,N_7134,N_7056);
xnor U7285 (N_7285,N_7151,N_7121);
or U7286 (N_7286,N_7109,N_7173);
nor U7287 (N_7287,N_7146,N_7044);
or U7288 (N_7288,N_7157,N_7066);
nand U7289 (N_7289,N_7189,N_7141);
nor U7290 (N_7290,N_7143,N_7083);
nand U7291 (N_7291,N_7150,N_7081);
xnor U7292 (N_7292,N_7142,N_7136);
or U7293 (N_7293,N_7197,N_7040);
xnor U7294 (N_7294,N_7141,N_7160);
nand U7295 (N_7295,N_7056,N_7139);
nand U7296 (N_7296,N_7059,N_7121);
nor U7297 (N_7297,N_7080,N_7141);
nor U7298 (N_7298,N_7042,N_7161);
nand U7299 (N_7299,N_7094,N_7100);
xnor U7300 (N_7300,N_7196,N_7198);
nand U7301 (N_7301,N_7067,N_7119);
xnor U7302 (N_7302,N_7155,N_7189);
and U7303 (N_7303,N_7110,N_7087);
nor U7304 (N_7304,N_7090,N_7160);
nand U7305 (N_7305,N_7086,N_7176);
nand U7306 (N_7306,N_7111,N_7054);
nor U7307 (N_7307,N_7045,N_7093);
and U7308 (N_7308,N_7152,N_7112);
or U7309 (N_7309,N_7129,N_7148);
nor U7310 (N_7310,N_7068,N_7086);
or U7311 (N_7311,N_7157,N_7191);
and U7312 (N_7312,N_7140,N_7055);
or U7313 (N_7313,N_7120,N_7079);
or U7314 (N_7314,N_7103,N_7141);
or U7315 (N_7315,N_7042,N_7047);
xor U7316 (N_7316,N_7103,N_7107);
or U7317 (N_7317,N_7113,N_7049);
and U7318 (N_7318,N_7187,N_7049);
nand U7319 (N_7319,N_7199,N_7188);
and U7320 (N_7320,N_7057,N_7179);
or U7321 (N_7321,N_7113,N_7137);
and U7322 (N_7322,N_7078,N_7081);
nor U7323 (N_7323,N_7050,N_7145);
nor U7324 (N_7324,N_7107,N_7075);
nand U7325 (N_7325,N_7076,N_7150);
and U7326 (N_7326,N_7120,N_7085);
and U7327 (N_7327,N_7071,N_7182);
or U7328 (N_7328,N_7084,N_7076);
nor U7329 (N_7329,N_7137,N_7158);
and U7330 (N_7330,N_7146,N_7101);
nand U7331 (N_7331,N_7058,N_7178);
or U7332 (N_7332,N_7042,N_7085);
nand U7333 (N_7333,N_7156,N_7140);
and U7334 (N_7334,N_7082,N_7138);
nor U7335 (N_7335,N_7089,N_7099);
xnor U7336 (N_7336,N_7164,N_7059);
nand U7337 (N_7337,N_7157,N_7183);
or U7338 (N_7338,N_7099,N_7065);
nand U7339 (N_7339,N_7182,N_7085);
or U7340 (N_7340,N_7106,N_7054);
nor U7341 (N_7341,N_7198,N_7087);
and U7342 (N_7342,N_7154,N_7175);
nor U7343 (N_7343,N_7111,N_7112);
nor U7344 (N_7344,N_7187,N_7133);
xor U7345 (N_7345,N_7101,N_7132);
nand U7346 (N_7346,N_7176,N_7055);
xor U7347 (N_7347,N_7100,N_7191);
and U7348 (N_7348,N_7192,N_7113);
or U7349 (N_7349,N_7041,N_7097);
or U7350 (N_7350,N_7132,N_7077);
xnor U7351 (N_7351,N_7126,N_7104);
nor U7352 (N_7352,N_7061,N_7112);
and U7353 (N_7353,N_7107,N_7166);
nor U7354 (N_7354,N_7053,N_7082);
xnor U7355 (N_7355,N_7072,N_7194);
xor U7356 (N_7356,N_7097,N_7187);
nand U7357 (N_7357,N_7160,N_7180);
or U7358 (N_7358,N_7117,N_7157);
nand U7359 (N_7359,N_7085,N_7131);
or U7360 (N_7360,N_7203,N_7325);
xor U7361 (N_7361,N_7297,N_7222);
and U7362 (N_7362,N_7349,N_7265);
xor U7363 (N_7363,N_7315,N_7289);
nand U7364 (N_7364,N_7348,N_7359);
and U7365 (N_7365,N_7253,N_7319);
xnor U7366 (N_7366,N_7251,N_7217);
nand U7367 (N_7367,N_7329,N_7291);
and U7368 (N_7368,N_7332,N_7304);
xnor U7369 (N_7369,N_7275,N_7336);
nor U7370 (N_7370,N_7261,N_7308);
or U7371 (N_7371,N_7327,N_7307);
or U7372 (N_7372,N_7267,N_7284);
and U7373 (N_7373,N_7353,N_7320);
xor U7374 (N_7374,N_7252,N_7351);
or U7375 (N_7375,N_7312,N_7246);
or U7376 (N_7376,N_7343,N_7287);
xnor U7377 (N_7377,N_7305,N_7344);
nand U7378 (N_7378,N_7254,N_7273);
and U7379 (N_7379,N_7242,N_7316);
and U7380 (N_7380,N_7266,N_7262);
and U7381 (N_7381,N_7270,N_7328);
nor U7382 (N_7382,N_7260,N_7215);
nor U7383 (N_7383,N_7352,N_7220);
nor U7384 (N_7384,N_7229,N_7247);
and U7385 (N_7385,N_7339,N_7300);
and U7386 (N_7386,N_7214,N_7238);
nand U7387 (N_7387,N_7295,N_7347);
nor U7388 (N_7388,N_7245,N_7334);
nor U7389 (N_7389,N_7330,N_7216);
xor U7390 (N_7390,N_7241,N_7310);
and U7391 (N_7391,N_7299,N_7218);
nor U7392 (N_7392,N_7285,N_7322);
or U7393 (N_7393,N_7201,N_7358);
nand U7394 (N_7394,N_7306,N_7346);
and U7395 (N_7395,N_7282,N_7257);
or U7396 (N_7396,N_7314,N_7240);
xnor U7397 (N_7397,N_7255,N_7231);
and U7398 (N_7398,N_7233,N_7280);
xnor U7399 (N_7399,N_7237,N_7249);
or U7400 (N_7400,N_7200,N_7269);
or U7401 (N_7401,N_7236,N_7335);
xnor U7402 (N_7402,N_7235,N_7302);
nor U7403 (N_7403,N_7326,N_7298);
and U7404 (N_7404,N_7225,N_7259);
nand U7405 (N_7405,N_7293,N_7356);
nor U7406 (N_7406,N_7317,N_7228);
and U7407 (N_7407,N_7258,N_7234);
xnor U7408 (N_7408,N_7331,N_7221);
nor U7409 (N_7409,N_7207,N_7279);
or U7410 (N_7410,N_7283,N_7232);
or U7411 (N_7411,N_7323,N_7276);
nand U7412 (N_7412,N_7333,N_7294);
nor U7413 (N_7413,N_7213,N_7357);
nor U7414 (N_7414,N_7303,N_7281);
and U7415 (N_7415,N_7350,N_7209);
and U7416 (N_7416,N_7224,N_7341);
and U7417 (N_7417,N_7311,N_7272);
nand U7418 (N_7418,N_7206,N_7226);
xnor U7419 (N_7419,N_7274,N_7340);
or U7420 (N_7420,N_7248,N_7202);
nand U7421 (N_7421,N_7256,N_7243);
or U7422 (N_7422,N_7210,N_7219);
and U7423 (N_7423,N_7271,N_7208);
nand U7424 (N_7424,N_7321,N_7354);
nand U7425 (N_7425,N_7301,N_7268);
nor U7426 (N_7426,N_7342,N_7230);
xor U7427 (N_7427,N_7292,N_7355);
and U7428 (N_7428,N_7204,N_7278);
and U7429 (N_7429,N_7205,N_7223);
and U7430 (N_7430,N_7250,N_7211);
nor U7431 (N_7431,N_7264,N_7286);
nand U7432 (N_7432,N_7227,N_7309);
nor U7433 (N_7433,N_7324,N_7313);
or U7434 (N_7434,N_7288,N_7244);
xnor U7435 (N_7435,N_7263,N_7277);
nand U7436 (N_7436,N_7337,N_7345);
or U7437 (N_7437,N_7296,N_7338);
xnor U7438 (N_7438,N_7318,N_7239);
nand U7439 (N_7439,N_7212,N_7290);
nor U7440 (N_7440,N_7247,N_7283);
nand U7441 (N_7441,N_7225,N_7240);
and U7442 (N_7442,N_7248,N_7314);
xnor U7443 (N_7443,N_7297,N_7228);
nor U7444 (N_7444,N_7348,N_7291);
or U7445 (N_7445,N_7233,N_7246);
or U7446 (N_7446,N_7293,N_7313);
xnor U7447 (N_7447,N_7212,N_7323);
xor U7448 (N_7448,N_7346,N_7228);
xor U7449 (N_7449,N_7336,N_7358);
nand U7450 (N_7450,N_7216,N_7306);
and U7451 (N_7451,N_7321,N_7297);
xor U7452 (N_7452,N_7344,N_7313);
xnor U7453 (N_7453,N_7356,N_7334);
nand U7454 (N_7454,N_7325,N_7291);
nor U7455 (N_7455,N_7300,N_7222);
and U7456 (N_7456,N_7271,N_7341);
nor U7457 (N_7457,N_7275,N_7204);
or U7458 (N_7458,N_7325,N_7294);
and U7459 (N_7459,N_7216,N_7308);
nor U7460 (N_7460,N_7233,N_7271);
and U7461 (N_7461,N_7220,N_7327);
or U7462 (N_7462,N_7313,N_7229);
nor U7463 (N_7463,N_7285,N_7324);
nor U7464 (N_7464,N_7355,N_7273);
nand U7465 (N_7465,N_7246,N_7238);
nor U7466 (N_7466,N_7284,N_7229);
nor U7467 (N_7467,N_7338,N_7349);
and U7468 (N_7468,N_7345,N_7256);
nand U7469 (N_7469,N_7339,N_7297);
nand U7470 (N_7470,N_7259,N_7236);
nand U7471 (N_7471,N_7238,N_7221);
or U7472 (N_7472,N_7321,N_7272);
or U7473 (N_7473,N_7318,N_7344);
xnor U7474 (N_7474,N_7309,N_7202);
nand U7475 (N_7475,N_7350,N_7320);
nor U7476 (N_7476,N_7319,N_7333);
nor U7477 (N_7477,N_7342,N_7218);
and U7478 (N_7478,N_7286,N_7244);
nor U7479 (N_7479,N_7251,N_7343);
nand U7480 (N_7480,N_7288,N_7324);
or U7481 (N_7481,N_7226,N_7305);
nand U7482 (N_7482,N_7344,N_7270);
nand U7483 (N_7483,N_7357,N_7216);
xnor U7484 (N_7484,N_7239,N_7202);
nor U7485 (N_7485,N_7280,N_7345);
xnor U7486 (N_7486,N_7294,N_7332);
and U7487 (N_7487,N_7248,N_7220);
nor U7488 (N_7488,N_7204,N_7289);
and U7489 (N_7489,N_7302,N_7265);
nor U7490 (N_7490,N_7326,N_7222);
nor U7491 (N_7491,N_7212,N_7316);
or U7492 (N_7492,N_7225,N_7306);
and U7493 (N_7493,N_7353,N_7221);
and U7494 (N_7494,N_7245,N_7263);
nand U7495 (N_7495,N_7343,N_7256);
or U7496 (N_7496,N_7295,N_7225);
and U7497 (N_7497,N_7338,N_7278);
nor U7498 (N_7498,N_7337,N_7222);
nor U7499 (N_7499,N_7305,N_7349);
nor U7500 (N_7500,N_7291,N_7300);
xnor U7501 (N_7501,N_7312,N_7337);
xor U7502 (N_7502,N_7252,N_7350);
xor U7503 (N_7503,N_7211,N_7235);
and U7504 (N_7504,N_7292,N_7310);
xnor U7505 (N_7505,N_7324,N_7244);
nand U7506 (N_7506,N_7221,N_7250);
xor U7507 (N_7507,N_7320,N_7215);
xor U7508 (N_7508,N_7243,N_7205);
nand U7509 (N_7509,N_7298,N_7295);
xor U7510 (N_7510,N_7293,N_7211);
xnor U7511 (N_7511,N_7215,N_7219);
and U7512 (N_7512,N_7335,N_7202);
nor U7513 (N_7513,N_7203,N_7349);
or U7514 (N_7514,N_7340,N_7227);
nand U7515 (N_7515,N_7338,N_7217);
nand U7516 (N_7516,N_7201,N_7261);
xnor U7517 (N_7517,N_7335,N_7272);
nand U7518 (N_7518,N_7350,N_7216);
xor U7519 (N_7519,N_7343,N_7245);
and U7520 (N_7520,N_7458,N_7431);
nand U7521 (N_7521,N_7467,N_7429);
and U7522 (N_7522,N_7370,N_7447);
and U7523 (N_7523,N_7473,N_7362);
xnor U7524 (N_7524,N_7424,N_7364);
nor U7525 (N_7525,N_7387,N_7452);
and U7526 (N_7526,N_7404,N_7368);
xnor U7527 (N_7527,N_7517,N_7506);
nor U7528 (N_7528,N_7475,N_7392);
xnor U7529 (N_7529,N_7504,N_7425);
nand U7530 (N_7530,N_7405,N_7384);
xnor U7531 (N_7531,N_7441,N_7500);
and U7532 (N_7532,N_7513,N_7511);
nand U7533 (N_7533,N_7470,N_7514);
nor U7534 (N_7534,N_7481,N_7372);
nand U7535 (N_7535,N_7397,N_7519);
and U7536 (N_7536,N_7466,N_7510);
or U7537 (N_7537,N_7413,N_7406);
nor U7538 (N_7538,N_7361,N_7436);
nor U7539 (N_7539,N_7360,N_7508);
nand U7540 (N_7540,N_7480,N_7505);
and U7541 (N_7541,N_7408,N_7394);
nand U7542 (N_7542,N_7503,N_7399);
xor U7543 (N_7543,N_7459,N_7471);
xor U7544 (N_7544,N_7407,N_7414);
or U7545 (N_7545,N_7512,N_7415);
and U7546 (N_7546,N_7373,N_7400);
xnor U7547 (N_7547,N_7365,N_7501);
and U7548 (N_7548,N_7487,N_7396);
and U7549 (N_7549,N_7411,N_7455);
nor U7550 (N_7550,N_7419,N_7428);
nand U7551 (N_7551,N_7375,N_7507);
nor U7552 (N_7552,N_7378,N_7498);
or U7553 (N_7553,N_7494,N_7497);
xor U7554 (N_7554,N_7417,N_7516);
nor U7555 (N_7555,N_7418,N_7389);
or U7556 (N_7556,N_7383,N_7386);
nand U7557 (N_7557,N_7421,N_7430);
nor U7558 (N_7558,N_7435,N_7453);
nor U7559 (N_7559,N_7371,N_7433);
nor U7560 (N_7560,N_7492,N_7412);
nand U7561 (N_7561,N_7485,N_7496);
nand U7562 (N_7562,N_7488,N_7426);
xnor U7563 (N_7563,N_7381,N_7460);
or U7564 (N_7564,N_7420,N_7443);
nand U7565 (N_7565,N_7450,N_7422);
xor U7566 (N_7566,N_7366,N_7444);
xor U7567 (N_7567,N_7445,N_7403);
and U7568 (N_7568,N_7363,N_7456);
nor U7569 (N_7569,N_7463,N_7410);
xor U7570 (N_7570,N_7493,N_7442);
xor U7571 (N_7571,N_7476,N_7390);
nor U7572 (N_7572,N_7448,N_7367);
nor U7573 (N_7573,N_7423,N_7388);
nor U7574 (N_7574,N_7446,N_7495);
nand U7575 (N_7575,N_7468,N_7385);
or U7576 (N_7576,N_7464,N_7499);
and U7577 (N_7577,N_7509,N_7457);
or U7578 (N_7578,N_7369,N_7454);
and U7579 (N_7579,N_7462,N_7515);
or U7580 (N_7580,N_7379,N_7401);
or U7581 (N_7581,N_7393,N_7469);
or U7582 (N_7582,N_7491,N_7461);
and U7583 (N_7583,N_7440,N_7382);
or U7584 (N_7584,N_7479,N_7490);
nor U7585 (N_7585,N_7437,N_7377);
xor U7586 (N_7586,N_7451,N_7483);
nand U7587 (N_7587,N_7482,N_7438);
and U7588 (N_7588,N_7477,N_7484);
and U7589 (N_7589,N_7391,N_7376);
and U7590 (N_7590,N_7474,N_7465);
nor U7591 (N_7591,N_7472,N_7486);
or U7592 (N_7592,N_7409,N_7518);
xnor U7593 (N_7593,N_7432,N_7416);
nand U7594 (N_7594,N_7489,N_7478);
and U7595 (N_7595,N_7402,N_7380);
and U7596 (N_7596,N_7502,N_7398);
or U7597 (N_7597,N_7374,N_7434);
nor U7598 (N_7598,N_7427,N_7439);
and U7599 (N_7599,N_7449,N_7395);
nor U7600 (N_7600,N_7391,N_7450);
nand U7601 (N_7601,N_7452,N_7415);
nand U7602 (N_7602,N_7446,N_7368);
nor U7603 (N_7603,N_7400,N_7410);
and U7604 (N_7604,N_7516,N_7473);
nand U7605 (N_7605,N_7391,N_7447);
nand U7606 (N_7606,N_7411,N_7518);
nor U7607 (N_7607,N_7422,N_7391);
xnor U7608 (N_7608,N_7395,N_7478);
nor U7609 (N_7609,N_7465,N_7472);
or U7610 (N_7610,N_7409,N_7482);
xor U7611 (N_7611,N_7364,N_7482);
or U7612 (N_7612,N_7365,N_7480);
nor U7613 (N_7613,N_7444,N_7447);
nand U7614 (N_7614,N_7514,N_7512);
and U7615 (N_7615,N_7504,N_7376);
nand U7616 (N_7616,N_7481,N_7466);
xnor U7617 (N_7617,N_7502,N_7389);
or U7618 (N_7618,N_7464,N_7492);
nor U7619 (N_7619,N_7519,N_7483);
nand U7620 (N_7620,N_7488,N_7494);
nor U7621 (N_7621,N_7424,N_7503);
nand U7622 (N_7622,N_7496,N_7428);
and U7623 (N_7623,N_7401,N_7472);
or U7624 (N_7624,N_7516,N_7378);
nand U7625 (N_7625,N_7411,N_7464);
xnor U7626 (N_7626,N_7470,N_7364);
and U7627 (N_7627,N_7443,N_7361);
nor U7628 (N_7628,N_7405,N_7410);
or U7629 (N_7629,N_7427,N_7455);
nand U7630 (N_7630,N_7517,N_7432);
nor U7631 (N_7631,N_7478,N_7382);
or U7632 (N_7632,N_7413,N_7417);
nand U7633 (N_7633,N_7435,N_7398);
or U7634 (N_7634,N_7433,N_7385);
nand U7635 (N_7635,N_7460,N_7497);
nor U7636 (N_7636,N_7431,N_7487);
nor U7637 (N_7637,N_7372,N_7415);
nand U7638 (N_7638,N_7390,N_7516);
and U7639 (N_7639,N_7458,N_7519);
nor U7640 (N_7640,N_7367,N_7399);
xor U7641 (N_7641,N_7397,N_7462);
or U7642 (N_7642,N_7500,N_7516);
or U7643 (N_7643,N_7389,N_7497);
or U7644 (N_7644,N_7462,N_7385);
or U7645 (N_7645,N_7482,N_7435);
xnor U7646 (N_7646,N_7361,N_7368);
and U7647 (N_7647,N_7376,N_7450);
nor U7648 (N_7648,N_7408,N_7484);
xor U7649 (N_7649,N_7430,N_7376);
xnor U7650 (N_7650,N_7380,N_7444);
or U7651 (N_7651,N_7455,N_7483);
nor U7652 (N_7652,N_7429,N_7492);
xor U7653 (N_7653,N_7376,N_7433);
nor U7654 (N_7654,N_7468,N_7363);
nand U7655 (N_7655,N_7409,N_7415);
xor U7656 (N_7656,N_7427,N_7502);
nor U7657 (N_7657,N_7503,N_7393);
nand U7658 (N_7658,N_7448,N_7427);
or U7659 (N_7659,N_7428,N_7382);
and U7660 (N_7660,N_7400,N_7473);
and U7661 (N_7661,N_7500,N_7503);
xnor U7662 (N_7662,N_7383,N_7506);
and U7663 (N_7663,N_7401,N_7460);
nand U7664 (N_7664,N_7487,N_7388);
nor U7665 (N_7665,N_7452,N_7439);
nand U7666 (N_7666,N_7457,N_7479);
nor U7667 (N_7667,N_7424,N_7375);
and U7668 (N_7668,N_7475,N_7451);
or U7669 (N_7669,N_7476,N_7373);
or U7670 (N_7670,N_7499,N_7409);
or U7671 (N_7671,N_7507,N_7370);
nand U7672 (N_7672,N_7436,N_7490);
or U7673 (N_7673,N_7463,N_7417);
and U7674 (N_7674,N_7442,N_7440);
xnor U7675 (N_7675,N_7514,N_7389);
or U7676 (N_7676,N_7460,N_7452);
nand U7677 (N_7677,N_7443,N_7484);
or U7678 (N_7678,N_7361,N_7414);
nand U7679 (N_7679,N_7517,N_7474);
and U7680 (N_7680,N_7675,N_7596);
or U7681 (N_7681,N_7673,N_7581);
or U7682 (N_7682,N_7643,N_7627);
nand U7683 (N_7683,N_7559,N_7619);
and U7684 (N_7684,N_7557,N_7536);
xor U7685 (N_7685,N_7655,N_7629);
xor U7686 (N_7686,N_7616,N_7625);
or U7687 (N_7687,N_7669,N_7562);
and U7688 (N_7688,N_7661,N_7601);
and U7689 (N_7689,N_7637,N_7630);
or U7690 (N_7690,N_7543,N_7657);
nand U7691 (N_7691,N_7598,N_7544);
xor U7692 (N_7692,N_7615,N_7632);
nand U7693 (N_7693,N_7608,N_7610);
or U7694 (N_7694,N_7631,N_7587);
nand U7695 (N_7695,N_7532,N_7606);
nand U7696 (N_7696,N_7612,N_7531);
and U7697 (N_7697,N_7522,N_7555);
or U7698 (N_7698,N_7591,N_7564);
and U7699 (N_7699,N_7539,N_7617);
xnor U7700 (N_7700,N_7653,N_7524);
nand U7701 (N_7701,N_7609,N_7679);
or U7702 (N_7702,N_7548,N_7546);
and U7703 (N_7703,N_7640,N_7534);
and U7704 (N_7704,N_7649,N_7658);
nor U7705 (N_7705,N_7582,N_7584);
nor U7706 (N_7706,N_7571,N_7664);
nor U7707 (N_7707,N_7660,N_7662);
nand U7708 (N_7708,N_7590,N_7599);
nand U7709 (N_7709,N_7542,N_7639);
nor U7710 (N_7710,N_7621,N_7556);
xor U7711 (N_7711,N_7541,N_7538);
xnor U7712 (N_7712,N_7547,N_7520);
and U7713 (N_7713,N_7614,N_7523);
or U7714 (N_7714,N_7569,N_7654);
or U7715 (N_7715,N_7647,N_7549);
nand U7716 (N_7716,N_7650,N_7666);
and U7717 (N_7717,N_7565,N_7656);
nor U7718 (N_7718,N_7552,N_7580);
nor U7719 (N_7719,N_7579,N_7670);
nand U7720 (N_7720,N_7570,N_7628);
nor U7721 (N_7721,N_7636,N_7575);
nand U7722 (N_7722,N_7604,N_7545);
or U7723 (N_7723,N_7645,N_7525);
and U7724 (N_7724,N_7574,N_7588);
nand U7725 (N_7725,N_7641,N_7572);
or U7726 (N_7726,N_7633,N_7578);
nand U7727 (N_7727,N_7535,N_7529);
nand U7728 (N_7728,N_7568,N_7635);
or U7729 (N_7729,N_7560,N_7659);
or U7730 (N_7730,N_7642,N_7594);
nand U7731 (N_7731,N_7665,N_7597);
xor U7732 (N_7732,N_7623,N_7527);
nand U7733 (N_7733,N_7620,N_7678);
nor U7734 (N_7734,N_7602,N_7573);
nor U7735 (N_7735,N_7592,N_7576);
nand U7736 (N_7736,N_7607,N_7537);
nor U7737 (N_7737,N_7677,N_7583);
xnor U7738 (N_7738,N_7663,N_7554);
and U7739 (N_7739,N_7558,N_7644);
nor U7740 (N_7740,N_7553,N_7634);
and U7741 (N_7741,N_7530,N_7521);
and U7742 (N_7742,N_7563,N_7668);
or U7743 (N_7743,N_7613,N_7676);
or U7744 (N_7744,N_7667,N_7595);
nor U7745 (N_7745,N_7540,N_7646);
and U7746 (N_7746,N_7593,N_7533);
xor U7747 (N_7747,N_7586,N_7528);
nor U7748 (N_7748,N_7550,N_7671);
and U7749 (N_7749,N_7589,N_7561);
nor U7750 (N_7750,N_7652,N_7672);
and U7751 (N_7751,N_7566,N_7674);
nand U7752 (N_7752,N_7567,N_7638);
xor U7753 (N_7753,N_7551,N_7648);
or U7754 (N_7754,N_7577,N_7626);
and U7755 (N_7755,N_7526,N_7651);
or U7756 (N_7756,N_7605,N_7585);
or U7757 (N_7757,N_7611,N_7603);
nor U7758 (N_7758,N_7600,N_7624);
or U7759 (N_7759,N_7622,N_7618);
and U7760 (N_7760,N_7644,N_7653);
and U7761 (N_7761,N_7544,N_7675);
or U7762 (N_7762,N_7635,N_7675);
nand U7763 (N_7763,N_7528,N_7564);
or U7764 (N_7764,N_7653,N_7640);
and U7765 (N_7765,N_7667,N_7612);
nand U7766 (N_7766,N_7598,N_7566);
or U7767 (N_7767,N_7584,N_7649);
xnor U7768 (N_7768,N_7663,N_7550);
and U7769 (N_7769,N_7621,N_7669);
nor U7770 (N_7770,N_7576,N_7524);
nor U7771 (N_7771,N_7548,N_7592);
nand U7772 (N_7772,N_7546,N_7646);
xor U7773 (N_7773,N_7583,N_7631);
or U7774 (N_7774,N_7633,N_7554);
or U7775 (N_7775,N_7543,N_7589);
xor U7776 (N_7776,N_7589,N_7604);
and U7777 (N_7777,N_7526,N_7634);
nand U7778 (N_7778,N_7583,N_7649);
nor U7779 (N_7779,N_7638,N_7670);
and U7780 (N_7780,N_7658,N_7643);
or U7781 (N_7781,N_7592,N_7617);
and U7782 (N_7782,N_7651,N_7656);
nor U7783 (N_7783,N_7629,N_7667);
xor U7784 (N_7784,N_7528,N_7520);
nand U7785 (N_7785,N_7620,N_7578);
nor U7786 (N_7786,N_7660,N_7539);
or U7787 (N_7787,N_7676,N_7548);
nor U7788 (N_7788,N_7566,N_7633);
xnor U7789 (N_7789,N_7590,N_7562);
xnor U7790 (N_7790,N_7634,N_7568);
nand U7791 (N_7791,N_7585,N_7658);
or U7792 (N_7792,N_7598,N_7651);
nand U7793 (N_7793,N_7644,N_7641);
nor U7794 (N_7794,N_7665,N_7554);
nand U7795 (N_7795,N_7601,N_7537);
and U7796 (N_7796,N_7639,N_7569);
and U7797 (N_7797,N_7571,N_7618);
nand U7798 (N_7798,N_7620,N_7639);
nor U7799 (N_7799,N_7563,N_7636);
or U7800 (N_7800,N_7606,N_7675);
nor U7801 (N_7801,N_7553,N_7642);
nor U7802 (N_7802,N_7643,N_7586);
or U7803 (N_7803,N_7643,N_7544);
nand U7804 (N_7804,N_7672,N_7555);
or U7805 (N_7805,N_7521,N_7598);
xor U7806 (N_7806,N_7546,N_7559);
or U7807 (N_7807,N_7618,N_7612);
or U7808 (N_7808,N_7576,N_7583);
nor U7809 (N_7809,N_7662,N_7555);
xnor U7810 (N_7810,N_7550,N_7648);
nor U7811 (N_7811,N_7589,N_7660);
xor U7812 (N_7812,N_7604,N_7636);
xor U7813 (N_7813,N_7639,N_7675);
nor U7814 (N_7814,N_7581,N_7523);
nand U7815 (N_7815,N_7594,N_7538);
and U7816 (N_7816,N_7665,N_7662);
nand U7817 (N_7817,N_7595,N_7529);
and U7818 (N_7818,N_7520,N_7533);
nor U7819 (N_7819,N_7561,N_7563);
or U7820 (N_7820,N_7614,N_7546);
or U7821 (N_7821,N_7656,N_7540);
xnor U7822 (N_7822,N_7656,N_7673);
nor U7823 (N_7823,N_7551,N_7672);
or U7824 (N_7824,N_7573,N_7593);
nand U7825 (N_7825,N_7574,N_7546);
nand U7826 (N_7826,N_7600,N_7547);
and U7827 (N_7827,N_7640,N_7584);
xnor U7828 (N_7828,N_7553,N_7612);
nor U7829 (N_7829,N_7556,N_7661);
and U7830 (N_7830,N_7650,N_7587);
xor U7831 (N_7831,N_7632,N_7569);
and U7832 (N_7832,N_7596,N_7650);
and U7833 (N_7833,N_7675,N_7676);
nand U7834 (N_7834,N_7523,N_7655);
nand U7835 (N_7835,N_7657,N_7546);
xor U7836 (N_7836,N_7670,N_7540);
xor U7837 (N_7837,N_7535,N_7555);
and U7838 (N_7838,N_7652,N_7649);
nand U7839 (N_7839,N_7608,N_7618);
xnor U7840 (N_7840,N_7724,N_7699);
nand U7841 (N_7841,N_7700,N_7702);
or U7842 (N_7842,N_7693,N_7763);
xor U7843 (N_7843,N_7775,N_7765);
nand U7844 (N_7844,N_7833,N_7744);
nor U7845 (N_7845,N_7701,N_7760);
or U7846 (N_7846,N_7722,N_7687);
nand U7847 (N_7847,N_7821,N_7776);
nor U7848 (N_7848,N_7790,N_7816);
or U7849 (N_7849,N_7838,N_7809);
nor U7850 (N_7850,N_7718,N_7691);
nand U7851 (N_7851,N_7792,N_7717);
xnor U7852 (N_7852,N_7711,N_7825);
nor U7853 (N_7853,N_7777,N_7751);
nor U7854 (N_7854,N_7812,N_7743);
nand U7855 (N_7855,N_7817,N_7762);
nand U7856 (N_7856,N_7754,N_7803);
or U7857 (N_7857,N_7698,N_7682);
nor U7858 (N_7858,N_7719,N_7736);
or U7859 (N_7859,N_7692,N_7707);
xor U7860 (N_7860,N_7828,N_7795);
nor U7861 (N_7861,N_7735,N_7800);
xnor U7862 (N_7862,N_7780,N_7772);
xor U7863 (N_7863,N_7752,N_7696);
nor U7864 (N_7864,N_7808,N_7747);
nand U7865 (N_7865,N_7723,N_7690);
nor U7866 (N_7866,N_7713,N_7734);
and U7867 (N_7867,N_7708,N_7767);
or U7868 (N_7868,N_7826,N_7689);
nand U7869 (N_7869,N_7683,N_7807);
and U7870 (N_7870,N_7827,N_7784);
or U7871 (N_7871,N_7835,N_7771);
xnor U7872 (N_7872,N_7811,N_7716);
xor U7873 (N_7873,N_7834,N_7745);
nand U7874 (N_7874,N_7787,N_7755);
and U7875 (N_7875,N_7764,N_7750);
nand U7876 (N_7876,N_7789,N_7706);
or U7877 (N_7877,N_7732,N_7694);
nor U7878 (N_7878,N_7837,N_7820);
nor U7879 (N_7879,N_7810,N_7824);
or U7880 (N_7880,N_7756,N_7726);
or U7881 (N_7881,N_7788,N_7758);
and U7882 (N_7882,N_7778,N_7728);
xor U7883 (N_7883,N_7742,N_7799);
and U7884 (N_7884,N_7704,N_7684);
nor U7885 (N_7885,N_7783,N_7794);
and U7886 (N_7886,N_7814,N_7797);
and U7887 (N_7887,N_7705,N_7686);
or U7888 (N_7888,N_7685,N_7749);
or U7889 (N_7889,N_7798,N_7829);
and U7890 (N_7890,N_7753,N_7839);
nor U7891 (N_7891,N_7741,N_7695);
xor U7892 (N_7892,N_7738,N_7813);
nor U7893 (N_7893,N_7822,N_7731);
or U7894 (N_7894,N_7709,N_7681);
and U7895 (N_7895,N_7740,N_7781);
xnor U7896 (N_7896,N_7721,N_7805);
nand U7897 (N_7897,N_7737,N_7703);
nand U7898 (N_7898,N_7714,N_7801);
xor U7899 (N_7899,N_7791,N_7710);
or U7900 (N_7900,N_7773,N_7697);
nand U7901 (N_7901,N_7757,N_7761);
xor U7902 (N_7902,N_7715,N_7725);
nor U7903 (N_7903,N_7759,N_7831);
nand U7904 (N_7904,N_7748,N_7768);
xnor U7905 (N_7905,N_7730,N_7766);
nor U7906 (N_7906,N_7823,N_7746);
xor U7907 (N_7907,N_7836,N_7739);
xor U7908 (N_7908,N_7818,N_7769);
or U7909 (N_7909,N_7680,N_7712);
nor U7910 (N_7910,N_7727,N_7774);
nand U7911 (N_7911,N_7785,N_7819);
xnor U7912 (N_7912,N_7832,N_7688);
or U7913 (N_7913,N_7779,N_7796);
or U7914 (N_7914,N_7830,N_7729);
nand U7915 (N_7915,N_7720,N_7770);
nand U7916 (N_7916,N_7802,N_7782);
or U7917 (N_7917,N_7804,N_7733);
or U7918 (N_7918,N_7786,N_7806);
nand U7919 (N_7919,N_7793,N_7815);
or U7920 (N_7920,N_7774,N_7699);
nor U7921 (N_7921,N_7688,N_7759);
and U7922 (N_7922,N_7749,N_7839);
and U7923 (N_7923,N_7781,N_7815);
xnor U7924 (N_7924,N_7728,N_7809);
or U7925 (N_7925,N_7732,N_7838);
nand U7926 (N_7926,N_7839,N_7734);
nor U7927 (N_7927,N_7726,N_7781);
nand U7928 (N_7928,N_7829,N_7818);
nand U7929 (N_7929,N_7785,N_7801);
nor U7930 (N_7930,N_7794,N_7758);
xnor U7931 (N_7931,N_7709,N_7823);
and U7932 (N_7932,N_7720,N_7732);
and U7933 (N_7933,N_7779,N_7813);
nor U7934 (N_7934,N_7812,N_7738);
and U7935 (N_7935,N_7799,N_7837);
or U7936 (N_7936,N_7758,N_7753);
and U7937 (N_7937,N_7777,N_7805);
nand U7938 (N_7938,N_7719,N_7824);
xnor U7939 (N_7939,N_7785,N_7820);
nor U7940 (N_7940,N_7822,N_7776);
nand U7941 (N_7941,N_7760,N_7712);
xnor U7942 (N_7942,N_7793,N_7799);
or U7943 (N_7943,N_7808,N_7811);
nand U7944 (N_7944,N_7763,N_7692);
xor U7945 (N_7945,N_7814,N_7784);
nor U7946 (N_7946,N_7698,N_7700);
xnor U7947 (N_7947,N_7693,N_7681);
and U7948 (N_7948,N_7790,N_7806);
nand U7949 (N_7949,N_7808,N_7750);
xor U7950 (N_7950,N_7832,N_7754);
nor U7951 (N_7951,N_7730,N_7745);
or U7952 (N_7952,N_7817,N_7813);
nand U7953 (N_7953,N_7697,N_7809);
and U7954 (N_7954,N_7722,N_7795);
and U7955 (N_7955,N_7781,N_7690);
or U7956 (N_7956,N_7700,N_7680);
nand U7957 (N_7957,N_7743,N_7711);
and U7958 (N_7958,N_7784,N_7767);
nand U7959 (N_7959,N_7727,N_7810);
nand U7960 (N_7960,N_7741,N_7802);
or U7961 (N_7961,N_7757,N_7832);
xor U7962 (N_7962,N_7757,N_7825);
and U7963 (N_7963,N_7796,N_7697);
or U7964 (N_7964,N_7707,N_7782);
nand U7965 (N_7965,N_7771,N_7738);
and U7966 (N_7966,N_7702,N_7818);
or U7967 (N_7967,N_7837,N_7838);
nor U7968 (N_7968,N_7799,N_7790);
nor U7969 (N_7969,N_7731,N_7754);
nor U7970 (N_7970,N_7795,N_7752);
or U7971 (N_7971,N_7802,N_7813);
xnor U7972 (N_7972,N_7740,N_7695);
nor U7973 (N_7973,N_7737,N_7795);
xnor U7974 (N_7974,N_7743,N_7825);
nand U7975 (N_7975,N_7765,N_7836);
xor U7976 (N_7976,N_7769,N_7804);
xnor U7977 (N_7977,N_7706,N_7726);
or U7978 (N_7978,N_7741,N_7716);
nor U7979 (N_7979,N_7769,N_7765);
and U7980 (N_7980,N_7740,N_7732);
xor U7981 (N_7981,N_7752,N_7791);
xor U7982 (N_7982,N_7821,N_7836);
or U7983 (N_7983,N_7771,N_7789);
and U7984 (N_7984,N_7743,N_7827);
or U7985 (N_7985,N_7789,N_7779);
xnor U7986 (N_7986,N_7756,N_7759);
nor U7987 (N_7987,N_7727,N_7748);
nand U7988 (N_7988,N_7730,N_7819);
and U7989 (N_7989,N_7748,N_7818);
nand U7990 (N_7990,N_7824,N_7803);
nor U7991 (N_7991,N_7800,N_7749);
nand U7992 (N_7992,N_7707,N_7770);
xor U7993 (N_7993,N_7726,N_7753);
nor U7994 (N_7994,N_7745,N_7789);
nor U7995 (N_7995,N_7804,N_7744);
nor U7996 (N_7996,N_7799,N_7725);
nand U7997 (N_7997,N_7707,N_7813);
or U7998 (N_7998,N_7696,N_7812);
and U7999 (N_7999,N_7780,N_7759);
and U8000 (N_8000,N_7912,N_7962);
or U8001 (N_8001,N_7877,N_7949);
nand U8002 (N_8002,N_7847,N_7950);
and U8003 (N_8003,N_7959,N_7969);
xor U8004 (N_8004,N_7991,N_7935);
nor U8005 (N_8005,N_7924,N_7984);
and U8006 (N_8006,N_7998,N_7883);
or U8007 (N_8007,N_7996,N_7933);
nor U8008 (N_8008,N_7995,N_7856);
nand U8009 (N_8009,N_7964,N_7927);
nor U8010 (N_8010,N_7955,N_7852);
and U8011 (N_8011,N_7966,N_7869);
and U8012 (N_8012,N_7882,N_7893);
nor U8013 (N_8013,N_7853,N_7900);
nand U8014 (N_8014,N_7892,N_7859);
or U8015 (N_8015,N_7947,N_7979);
and U8016 (N_8016,N_7960,N_7889);
nand U8017 (N_8017,N_7946,N_7914);
or U8018 (N_8018,N_7910,N_7891);
and U8019 (N_8019,N_7937,N_7915);
nor U8020 (N_8020,N_7982,N_7978);
nor U8021 (N_8021,N_7862,N_7936);
and U8022 (N_8022,N_7952,N_7942);
and U8023 (N_8023,N_7993,N_7866);
xnor U8024 (N_8024,N_7896,N_7878);
nand U8025 (N_8025,N_7845,N_7986);
xor U8026 (N_8026,N_7855,N_7997);
nor U8027 (N_8027,N_7970,N_7972);
or U8028 (N_8028,N_7843,N_7928);
or U8029 (N_8029,N_7886,N_7961);
and U8030 (N_8030,N_7994,N_7911);
xnor U8031 (N_8031,N_7854,N_7873);
nand U8032 (N_8032,N_7887,N_7916);
or U8033 (N_8033,N_7963,N_7850);
nor U8034 (N_8034,N_7899,N_7930);
or U8035 (N_8035,N_7923,N_7934);
and U8036 (N_8036,N_7874,N_7973);
and U8037 (N_8037,N_7990,N_7988);
nor U8038 (N_8038,N_7871,N_7898);
or U8039 (N_8039,N_7926,N_7865);
nor U8040 (N_8040,N_7858,N_7909);
and U8041 (N_8041,N_7849,N_7872);
nor U8042 (N_8042,N_7840,N_7965);
xnor U8043 (N_8043,N_7976,N_7989);
or U8044 (N_8044,N_7857,N_7844);
nor U8045 (N_8045,N_7992,N_7999);
or U8046 (N_8046,N_7943,N_7931);
and U8047 (N_8047,N_7908,N_7903);
nand U8048 (N_8048,N_7980,N_7906);
nor U8049 (N_8049,N_7940,N_7864);
and U8050 (N_8050,N_7938,N_7948);
nand U8051 (N_8051,N_7968,N_7967);
nor U8052 (N_8052,N_7983,N_7870);
and U8053 (N_8053,N_7885,N_7902);
nor U8054 (N_8054,N_7879,N_7884);
xnor U8055 (N_8055,N_7880,N_7881);
and U8056 (N_8056,N_7941,N_7907);
and U8057 (N_8057,N_7974,N_7987);
nor U8058 (N_8058,N_7890,N_7842);
and U8059 (N_8059,N_7897,N_7913);
or U8060 (N_8060,N_7876,N_7975);
nor U8061 (N_8061,N_7868,N_7921);
xnor U8062 (N_8062,N_7977,N_7939);
nand U8063 (N_8063,N_7904,N_7848);
xor U8064 (N_8064,N_7958,N_7905);
nor U8065 (N_8065,N_7954,N_7919);
nand U8066 (N_8066,N_7851,N_7894);
nand U8067 (N_8067,N_7888,N_7981);
or U8068 (N_8068,N_7985,N_7956);
nor U8069 (N_8069,N_7846,N_7841);
xnor U8070 (N_8070,N_7875,N_7951);
nor U8071 (N_8071,N_7925,N_7867);
xor U8072 (N_8072,N_7901,N_7929);
or U8073 (N_8073,N_7920,N_7945);
xnor U8074 (N_8074,N_7953,N_7957);
and U8075 (N_8075,N_7971,N_7917);
xor U8076 (N_8076,N_7944,N_7860);
nand U8077 (N_8077,N_7863,N_7932);
and U8078 (N_8078,N_7895,N_7922);
and U8079 (N_8079,N_7918,N_7861);
nor U8080 (N_8080,N_7859,N_7891);
nor U8081 (N_8081,N_7922,N_7944);
and U8082 (N_8082,N_7931,N_7855);
nor U8083 (N_8083,N_7898,N_7885);
xor U8084 (N_8084,N_7934,N_7941);
and U8085 (N_8085,N_7996,N_7975);
nand U8086 (N_8086,N_7919,N_7855);
or U8087 (N_8087,N_7986,N_7929);
xor U8088 (N_8088,N_7935,N_7949);
nand U8089 (N_8089,N_7899,N_7880);
and U8090 (N_8090,N_7933,N_7915);
nand U8091 (N_8091,N_7936,N_7878);
and U8092 (N_8092,N_7916,N_7946);
xor U8093 (N_8093,N_7913,N_7888);
or U8094 (N_8094,N_7960,N_7940);
and U8095 (N_8095,N_7870,N_7912);
or U8096 (N_8096,N_7850,N_7974);
nor U8097 (N_8097,N_7999,N_7946);
xnor U8098 (N_8098,N_7990,N_7866);
nor U8099 (N_8099,N_7990,N_7915);
and U8100 (N_8100,N_7893,N_7972);
or U8101 (N_8101,N_7875,N_7913);
nand U8102 (N_8102,N_7926,N_7936);
xnor U8103 (N_8103,N_7937,N_7883);
or U8104 (N_8104,N_7995,N_7888);
xor U8105 (N_8105,N_7912,N_7893);
or U8106 (N_8106,N_7909,N_7974);
and U8107 (N_8107,N_7919,N_7894);
xor U8108 (N_8108,N_7948,N_7895);
xor U8109 (N_8109,N_7906,N_7870);
nand U8110 (N_8110,N_7904,N_7933);
nand U8111 (N_8111,N_7933,N_7995);
and U8112 (N_8112,N_7938,N_7927);
nand U8113 (N_8113,N_7945,N_7841);
nor U8114 (N_8114,N_7985,N_7841);
and U8115 (N_8115,N_7986,N_7940);
and U8116 (N_8116,N_7945,N_7888);
and U8117 (N_8117,N_7902,N_7927);
and U8118 (N_8118,N_7937,N_7884);
or U8119 (N_8119,N_7898,N_7988);
or U8120 (N_8120,N_7968,N_7876);
xor U8121 (N_8121,N_7959,N_7946);
nor U8122 (N_8122,N_7849,N_7871);
nor U8123 (N_8123,N_7915,N_7983);
xor U8124 (N_8124,N_7975,N_7880);
nor U8125 (N_8125,N_7968,N_7895);
xnor U8126 (N_8126,N_7926,N_7907);
nor U8127 (N_8127,N_7982,N_7915);
xnor U8128 (N_8128,N_7912,N_7906);
nand U8129 (N_8129,N_7842,N_7892);
and U8130 (N_8130,N_7878,N_7913);
xnor U8131 (N_8131,N_7959,N_7977);
or U8132 (N_8132,N_7881,N_7972);
xor U8133 (N_8133,N_7856,N_7976);
or U8134 (N_8134,N_7861,N_7916);
and U8135 (N_8135,N_7925,N_7996);
or U8136 (N_8136,N_7930,N_7910);
or U8137 (N_8137,N_7936,N_7937);
nand U8138 (N_8138,N_7899,N_7893);
or U8139 (N_8139,N_7890,N_7901);
nor U8140 (N_8140,N_7961,N_7984);
nor U8141 (N_8141,N_7983,N_7863);
nand U8142 (N_8142,N_7917,N_7983);
nor U8143 (N_8143,N_7984,N_7921);
nor U8144 (N_8144,N_7897,N_7960);
nor U8145 (N_8145,N_7873,N_7878);
xor U8146 (N_8146,N_7842,N_7961);
or U8147 (N_8147,N_7858,N_7872);
nand U8148 (N_8148,N_7913,N_7920);
xor U8149 (N_8149,N_7962,N_7841);
xnor U8150 (N_8150,N_7925,N_7885);
nor U8151 (N_8151,N_7958,N_7983);
nor U8152 (N_8152,N_7911,N_7848);
xor U8153 (N_8153,N_7929,N_7856);
or U8154 (N_8154,N_7904,N_7957);
or U8155 (N_8155,N_7853,N_7976);
nor U8156 (N_8156,N_7877,N_7856);
or U8157 (N_8157,N_7942,N_7885);
or U8158 (N_8158,N_7957,N_7931);
and U8159 (N_8159,N_7939,N_7979);
nor U8160 (N_8160,N_8045,N_8003);
and U8161 (N_8161,N_8017,N_8068);
and U8162 (N_8162,N_8152,N_8140);
nor U8163 (N_8163,N_8030,N_8020);
and U8164 (N_8164,N_8096,N_8047);
or U8165 (N_8165,N_8103,N_8148);
or U8166 (N_8166,N_8009,N_8104);
and U8167 (N_8167,N_8077,N_8046);
and U8168 (N_8168,N_8034,N_8101);
or U8169 (N_8169,N_8093,N_8133);
and U8170 (N_8170,N_8070,N_8087);
and U8171 (N_8171,N_8054,N_8125);
or U8172 (N_8172,N_8001,N_8135);
nand U8173 (N_8173,N_8022,N_8000);
xor U8174 (N_8174,N_8138,N_8010);
and U8175 (N_8175,N_8153,N_8074);
nor U8176 (N_8176,N_8050,N_8109);
nor U8177 (N_8177,N_8071,N_8043);
nor U8178 (N_8178,N_8076,N_8100);
nor U8179 (N_8179,N_8036,N_8112);
xnor U8180 (N_8180,N_8033,N_8118);
or U8181 (N_8181,N_8081,N_8062);
xnor U8182 (N_8182,N_8131,N_8052);
or U8183 (N_8183,N_8059,N_8005);
or U8184 (N_8184,N_8032,N_8019);
and U8185 (N_8185,N_8154,N_8099);
nor U8186 (N_8186,N_8027,N_8011);
or U8187 (N_8187,N_8060,N_8002);
nand U8188 (N_8188,N_8121,N_8040);
xnor U8189 (N_8189,N_8113,N_8091);
nor U8190 (N_8190,N_8129,N_8126);
and U8191 (N_8191,N_8024,N_8025);
or U8192 (N_8192,N_8145,N_8026);
and U8193 (N_8193,N_8119,N_8147);
and U8194 (N_8194,N_8114,N_8115);
nand U8195 (N_8195,N_8144,N_8137);
nor U8196 (N_8196,N_8108,N_8049);
or U8197 (N_8197,N_8098,N_8066);
nand U8198 (N_8198,N_8139,N_8082);
and U8199 (N_8199,N_8014,N_8128);
and U8200 (N_8200,N_8018,N_8088);
xor U8201 (N_8201,N_8072,N_8078);
nand U8202 (N_8202,N_8037,N_8086);
or U8203 (N_8203,N_8013,N_8141);
nand U8204 (N_8204,N_8061,N_8094);
nor U8205 (N_8205,N_8023,N_8048);
nor U8206 (N_8206,N_8067,N_8006);
or U8207 (N_8207,N_8041,N_8055);
and U8208 (N_8208,N_8085,N_8156);
nand U8209 (N_8209,N_8012,N_8042);
nand U8210 (N_8210,N_8079,N_8016);
xor U8211 (N_8211,N_8110,N_8080);
and U8212 (N_8212,N_8124,N_8083);
xor U8213 (N_8213,N_8031,N_8102);
and U8214 (N_8214,N_8107,N_8159);
or U8215 (N_8215,N_8004,N_8106);
xor U8216 (N_8216,N_8149,N_8065);
and U8217 (N_8217,N_8111,N_8151);
or U8218 (N_8218,N_8105,N_8015);
nand U8219 (N_8219,N_8063,N_8122);
nor U8220 (N_8220,N_8150,N_8120);
and U8221 (N_8221,N_8038,N_8090);
nand U8222 (N_8222,N_8069,N_8158);
and U8223 (N_8223,N_8084,N_8127);
or U8224 (N_8224,N_8117,N_8035);
nor U8225 (N_8225,N_8075,N_8092);
nor U8226 (N_8226,N_8134,N_8058);
and U8227 (N_8227,N_8028,N_8057);
nand U8228 (N_8228,N_8053,N_8064);
xnor U8229 (N_8229,N_8029,N_8095);
or U8230 (N_8230,N_8142,N_8143);
xor U8231 (N_8231,N_8089,N_8155);
or U8232 (N_8232,N_8146,N_8056);
or U8233 (N_8233,N_8116,N_8132);
nand U8234 (N_8234,N_8130,N_8051);
nor U8235 (N_8235,N_8044,N_8007);
nor U8236 (N_8236,N_8039,N_8157);
nand U8237 (N_8237,N_8008,N_8073);
and U8238 (N_8238,N_8021,N_8136);
xor U8239 (N_8239,N_8123,N_8097);
xor U8240 (N_8240,N_8105,N_8070);
nor U8241 (N_8241,N_8151,N_8037);
or U8242 (N_8242,N_8143,N_8119);
nand U8243 (N_8243,N_8044,N_8031);
nor U8244 (N_8244,N_8110,N_8159);
or U8245 (N_8245,N_8024,N_8144);
xnor U8246 (N_8246,N_8060,N_8059);
nand U8247 (N_8247,N_8117,N_8081);
xnor U8248 (N_8248,N_8145,N_8130);
nand U8249 (N_8249,N_8045,N_8156);
and U8250 (N_8250,N_8135,N_8065);
and U8251 (N_8251,N_8097,N_8144);
or U8252 (N_8252,N_8151,N_8080);
or U8253 (N_8253,N_8081,N_8005);
nand U8254 (N_8254,N_8038,N_8054);
xnor U8255 (N_8255,N_8122,N_8043);
nor U8256 (N_8256,N_8105,N_8067);
and U8257 (N_8257,N_8015,N_8067);
nand U8258 (N_8258,N_8073,N_8101);
nand U8259 (N_8259,N_8101,N_8077);
or U8260 (N_8260,N_8008,N_8101);
and U8261 (N_8261,N_8031,N_8148);
nand U8262 (N_8262,N_8034,N_8112);
nand U8263 (N_8263,N_8132,N_8135);
xnor U8264 (N_8264,N_8042,N_8129);
xnor U8265 (N_8265,N_8080,N_8061);
and U8266 (N_8266,N_8136,N_8051);
and U8267 (N_8267,N_8106,N_8026);
xnor U8268 (N_8268,N_8147,N_8045);
xor U8269 (N_8269,N_8044,N_8082);
or U8270 (N_8270,N_8055,N_8100);
or U8271 (N_8271,N_8054,N_8158);
xnor U8272 (N_8272,N_8081,N_8098);
and U8273 (N_8273,N_8037,N_8052);
nor U8274 (N_8274,N_8076,N_8125);
or U8275 (N_8275,N_8024,N_8066);
or U8276 (N_8276,N_8135,N_8046);
or U8277 (N_8277,N_8129,N_8105);
or U8278 (N_8278,N_8127,N_8068);
xor U8279 (N_8279,N_8110,N_8088);
nor U8280 (N_8280,N_8092,N_8036);
and U8281 (N_8281,N_8089,N_8131);
nand U8282 (N_8282,N_8133,N_8079);
or U8283 (N_8283,N_8151,N_8144);
xnor U8284 (N_8284,N_8138,N_8114);
or U8285 (N_8285,N_8082,N_8014);
and U8286 (N_8286,N_8146,N_8116);
and U8287 (N_8287,N_8121,N_8125);
xnor U8288 (N_8288,N_8054,N_8141);
and U8289 (N_8289,N_8122,N_8007);
nor U8290 (N_8290,N_8041,N_8053);
and U8291 (N_8291,N_8071,N_8039);
nand U8292 (N_8292,N_8147,N_8066);
nand U8293 (N_8293,N_8104,N_8061);
nand U8294 (N_8294,N_8079,N_8088);
or U8295 (N_8295,N_8047,N_8078);
or U8296 (N_8296,N_8041,N_8136);
xnor U8297 (N_8297,N_8121,N_8024);
nor U8298 (N_8298,N_8071,N_8021);
xnor U8299 (N_8299,N_8146,N_8016);
and U8300 (N_8300,N_8049,N_8116);
xor U8301 (N_8301,N_8086,N_8029);
nor U8302 (N_8302,N_8123,N_8048);
and U8303 (N_8303,N_8096,N_8122);
or U8304 (N_8304,N_8054,N_8085);
and U8305 (N_8305,N_8018,N_8033);
xnor U8306 (N_8306,N_8043,N_8031);
nand U8307 (N_8307,N_8152,N_8035);
and U8308 (N_8308,N_8087,N_8158);
xnor U8309 (N_8309,N_8144,N_8054);
or U8310 (N_8310,N_8005,N_8054);
nor U8311 (N_8311,N_8100,N_8130);
nor U8312 (N_8312,N_8022,N_8023);
and U8313 (N_8313,N_8002,N_8083);
nor U8314 (N_8314,N_8077,N_8151);
or U8315 (N_8315,N_8148,N_8030);
nand U8316 (N_8316,N_8051,N_8070);
nand U8317 (N_8317,N_8119,N_8094);
nor U8318 (N_8318,N_8047,N_8095);
nand U8319 (N_8319,N_8143,N_8100);
or U8320 (N_8320,N_8302,N_8239);
xor U8321 (N_8321,N_8202,N_8249);
xor U8322 (N_8322,N_8257,N_8297);
xnor U8323 (N_8323,N_8243,N_8295);
or U8324 (N_8324,N_8179,N_8253);
xor U8325 (N_8325,N_8244,N_8169);
nand U8326 (N_8326,N_8195,N_8219);
nor U8327 (N_8327,N_8285,N_8170);
nor U8328 (N_8328,N_8234,N_8296);
or U8329 (N_8329,N_8218,N_8181);
xor U8330 (N_8330,N_8176,N_8177);
or U8331 (N_8331,N_8270,N_8212);
xnor U8332 (N_8332,N_8204,N_8210);
and U8333 (N_8333,N_8268,N_8274);
and U8334 (N_8334,N_8319,N_8308);
nand U8335 (N_8335,N_8207,N_8260);
or U8336 (N_8336,N_8232,N_8272);
nand U8337 (N_8337,N_8199,N_8236);
or U8338 (N_8338,N_8192,N_8171);
xnor U8339 (N_8339,N_8304,N_8235);
nand U8340 (N_8340,N_8278,N_8190);
and U8341 (N_8341,N_8203,N_8281);
nand U8342 (N_8342,N_8317,N_8263);
xnor U8343 (N_8343,N_8208,N_8231);
and U8344 (N_8344,N_8241,N_8286);
or U8345 (N_8345,N_8289,N_8215);
nor U8346 (N_8346,N_8258,N_8227);
and U8347 (N_8347,N_8206,N_8303);
and U8348 (N_8348,N_8250,N_8167);
or U8349 (N_8349,N_8267,N_8284);
xnor U8350 (N_8350,N_8216,N_8201);
nand U8351 (N_8351,N_8174,N_8293);
nor U8352 (N_8352,N_8245,N_8275);
or U8353 (N_8353,N_8311,N_8254);
and U8354 (N_8354,N_8228,N_8175);
or U8355 (N_8355,N_8164,N_8173);
nor U8356 (N_8356,N_8279,N_8161);
or U8357 (N_8357,N_8280,N_8261);
xor U8358 (N_8358,N_8288,N_8220);
and U8359 (N_8359,N_8242,N_8310);
nor U8360 (N_8360,N_8265,N_8223);
and U8361 (N_8361,N_8309,N_8160);
and U8362 (N_8362,N_8191,N_8316);
or U8363 (N_8363,N_8271,N_8165);
xnor U8364 (N_8364,N_8184,N_8313);
xor U8365 (N_8365,N_8283,N_8307);
nor U8366 (N_8366,N_8198,N_8189);
nand U8367 (N_8367,N_8211,N_8266);
and U8368 (N_8368,N_8287,N_8209);
nand U8369 (N_8369,N_8226,N_8205);
nand U8370 (N_8370,N_8251,N_8214);
or U8371 (N_8371,N_8183,N_8168);
or U8372 (N_8372,N_8294,N_8256);
xor U8373 (N_8373,N_8224,N_8233);
nor U8374 (N_8374,N_8312,N_8282);
nor U8375 (N_8375,N_8182,N_8217);
nor U8376 (N_8376,N_8230,N_8318);
and U8377 (N_8377,N_8314,N_8298);
and U8378 (N_8378,N_8188,N_8229);
xor U8379 (N_8379,N_8200,N_8300);
xnor U8380 (N_8380,N_8255,N_8163);
or U8381 (N_8381,N_8222,N_8213);
nor U8382 (N_8382,N_8166,N_8259);
nor U8383 (N_8383,N_8315,N_8264);
nor U8384 (N_8384,N_8238,N_8305);
nand U8385 (N_8385,N_8291,N_8246);
and U8386 (N_8386,N_8299,N_8262);
or U8387 (N_8387,N_8292,N_8252);
xnor U8388 (N_8388,N_8240,N_8178);
and U8389 (N_8389,N_8277,N_8172);
nand U8390 (N_8390,N_8306,N_8193);
xor U8391 (N_8391,N_8194,N_8237);
and U8392 (N_8392,N_8269,N_8221);
nand U8393 (N_8393,N_8185,N_8197);
or U8394 (N_8394,N_8248,N_8273);
nand U8395 (N_8395,N_8290,N_8187);
nor U8396 (N_8396,N_8247,N_8186);
and U8397 (N_8397,N_8196,N_8301);
xor U8398 (N_8398,N_8162,N_8276);
nand U8399 (N_8399,N_8180,N_8225);
or U8400 (N_8400,N_8235,N_8293);
nand U8401 (N_8401,N_8193,N_8260);
or U8402 (N_8402,N_8188,N_8232);
or U8403 (N_8403,N_8268,N_8310);
xor U8404 (N_8404,N_8257,N_8304);
and U8405 (N_8405,N_8171,N_8308);
nand U8406 (N_8406,N_8291,N_8209);
and U8407 (N_8407,N_8297,N_8284);
xor U8408 (N_8408,N_8206,N_8256);
and U8409 (N_8409,N_8164,N_8162);
nor U8410 (N_8410,N_8231,N_8249);
nor U8411 (N_8411,N_8305,N_8181);
nor U8412 (N_8412,N_8198,N_8258);
and U8413 (N_8413,N_8284,N_8312);
or U8414 (N_8414,N_8230,N_8285);
and U8415 (N_8415,N_8317,N_8194);
nand U8416 (N_8416,N_8161,N_8216);
nand U8417 (N_8417,N_8278,N_8236);
nor U8418 (N_8418,N_8250,N_8271);
xnor U8419 (N_8419,N_8176,N_8288);
and U8420 (N_8420,N_8304,N_8316);
xor U8421 (N_8421,N_8180,N_8306);
nand U8422 (N_8422,N_8291,N_8199);
nand U8423 (N_8423,N_8193,N_8196);
and U8424 (N_8424,N_8208,N_8291);
nor U8425 (N_8425,N_8207,N_8306);
nor U8426 (N_8426,N_8181,N_8248);
or U8427 (N_8427,N_8227,N_8163);
or U8428 (N_8428,N_8252,N_8309);
nand U8429 (N_8429,N_8312,N_8224);
or U8430 (N_8430,N_8273,N_8197);
nor U8431 (N_8431,N_8230,N_8208);
nor U8432 (N_8432,N_8241,N_8229);
nand U8433 (N_8433,N_8206,N_8161);
and U8434 (N_8434,N_8188,N_8252);
xor U8435 (N_8435,N_8170,N_8289);
nor U8436 (N_8436,N_8221,N_8268);
nor U8437 (N_8437,N_8206,N_8232);
xnor U8438 (N_8438,N_8295,N_8180);
or U8439 (N_8439,N_8265,N_8201);
nor U8440 (N_8440,N_8273,N_8310);
xor U8441 (N_8441,N_8252,N_8294);
and U8442 (N_8442,N_8218,N_8277);
nand U8443 (N_8443,N_8207,N_8279);
nand U8444 (N_8444,N_8250,N_8303);
nor U8445 (N_8445,N_8236,N_8291);
nand U8446 (N_8446,N_8290,N_8315);
xor U8447 (N_8447,N_8250,N_8231);
nor U8448 (N_8448,N_8243,N_8302);
and U8449 (N_8449,N_8265,N_8192);
or U8450 (N_8450,N_8162,N_8174);
nor U8451 (N_8451,N_8201,N_8205);
xnor U8452 (N_8452,N_8258,N_8246);
or U8453 (N_8453,N_8199,N_8193);
or U8454 (N_8454,N_8205,N_8290);
and U8455 (N_8455,N_8186,N_8162);
and U8456 (N_8456,N_8302,N_8319);
xor U8457 (N_8457,N_8162,N_8210);
nand U8458 (N_8458,N_8198,N_8234);
nor U8459 (N_8459,N_8193,N_8282);
xor U8460 (N_8460,N_8252,N_8316);
xor U8461 (N_8461,N_8314,N_8242);
nand U8462 (N_8462,N_8289,N_8185);
or U8463 (N_8463,N_8316,N_8208);
and U8464 (N_8464,N_8309,N_8280);
nand U8465 (N_8465,N_8220,N_8208);
or U8466 (N_8466,N_8277,N_8222);
or U8467 (N_8467,N_8237,N_8275);
xor U8468 (N_8468,N_8171,N_8186);
xnor U8469 (N_8469,N_8185,N_8219);
xnor U8470 (N_8470,N_8279,N_8165);
nand U8471 (N_8471,N_8207,N_8297);
and U8472 (N_8472,N_8238,N_8277);
nor U8473 (N_8473,N_8193,N_8167);
and U8474 (N_8474,N_8309,N_8227);
nor U8475 (N_8475,N_8176,N_8255);
and U8476 (N_8476,N_8304,N_8287);
nand U8477 (N_8477,N_8282,N_8198);
nand U8478 (N_8478,N_8203,N_8314);
and U8479 (N_8479,N_8208,N_8286);
or U8480 (N_8480,N_8331,N_8321);
nand U8481 (N_8481,N_8441,N_8368);
or U8482 (N_8482,N_8468,N_8451);
nand U8483 (N_8483,N_8463,N_8475);
nor U8484 (N_8484,N_8428,N_8396);
and U8485 (N_8485,N_8389,N_8474);
and U8486 (N_8486,N_8372,N_8409);
or U8487 (N_8487,N_8477,N_8453);
xor U8488 (N_8488,N_8394,N_8433);
nand U8489 (N_8489,N_8388,N_8436);
or U8490 (N_8490,N_8338,N_8334);
nor U8491 (N_8491,N_8410,N_8379);
or U8492 (N_8492,N_8406,N_8356);
and U8493 (N_8493,N_8476,N_8454);
nand U8494 (N_8494,N_8429,N_8342);
xor U8495 (N_8495,N_8458,N_8450);
xnor U8496 (N_8496,N_8418,N_8430);
nand U8497 (N_8497,N_8395,N_8330);
and U8498 (N_8498,N_8327,N_8473);
xor U8499 (N_8499,N_8434,N_8391);
nor U8500 (N_8500,N_8399,N_8360);
nor U8501 (N_8501,N_8366,N_8402);
nand U8502 (N_8502,N_8457,N_8324);
nor U8503 (N_8503,N_8337,N_8355);
xor U8504 (N_8504,N_8320,N_8374);
or U8505 (N_8505,N_8416,N_8425);
and U8506 (N_8506,N_8415,N_8357);
xnor U8507 (N_8507,N_8365,N_8362);
xnor U8508 (N_8508,N_8341,N_8375);
or U8509 (N_8509,N_8478,N_8370);
or U8510 (N_8510,N_8479,N_8461);
or U8511 (N_8511,N_8412,N_8398);
nor U8512 (N_8512,N_8386,N_8384);
or U8513 (N_8513,N_8382,N_8335);
or U8514 (N_8514,N_8403,N_8380);
or U8515 (N_8515,N_8400,N_8371);
xor U8516 (N_8516,N_8329,N_8351);
or U8517 (N_8517,N_8359,N_8363);
or U8518 (N_8518,N_8340,N_8407);
nor U8519 (N_8519,N_8383,N_8377);
xnor U8520 (N_8520,N_8397,N_8413);
or U8521 (N_8521,N_8426,N_8420);
nor U8522 (N_8522,N_8354,N_8465);
nand U8523 (N_8523,N_8439,N_8449);
and U8524 (N_8524,N_8445,N_8456);
nor U8525 (N_8525,N_8447,N_8345);
xor U8526 (N_8526,N_8361,N_8385);
xor U8527 (N_8527,N_8381,N_8440);
nand U8528 (N_8528,N_8376,N_8422);
or U8529 (N_8529,N_8323,N_8364);
nor U8530 (N_8530,N_8401,N_8350);
nor U8531 (N_8531,N_8421,N_8333);
or U8532 (N_8532,N_8369,N_8392);
or U8533 (N_8533,N_8442,N_8431);
and U8534 (N_8534,N_8438,N_8470);
xnor U8535 (N_8535,N_8446,N_8435);
xor U8536 (N_8536,N_8336,N_8352);
or U8537 (N_8537,N_8326,N_8390);
or U8538 (N_8538,N_8404,N_8414);
or U8539 (N_8539,N_8373,N_8405);
and U8540 (N_8540,N_8459,N_8437);
nor U8541 (N_8541,N_8408,N_8393);
xor U8542 (N_8542,N_8332,N_8387);
nand U8543 (N_8543,N_8347,N_8339);
and U8544 (N_8544,N_8367,N_8466);
nand U8545 (N_8545,N_8448,N_8443);
xnor U8546 (N_8546,N_8343,N_8325);
nor U8547 (N_8547,N_8411,N_8349);
or U8548 (N_8548,N_8328,N_8460);
xor U8549 (N_8549,N_8344,N_8427);
or U8550 (N_8550,N_8353,N_8424);
nand U8551 (N_8551,N_8432,N_8322);
and U8552 (N_8552,N_8358,N_8346);
xor U8553 (N_8553,N_8467,N_8417);
or U8554 (N_8554,N_8472,N_8464);
or U8555 (N_8555,N_8378,N_8452);
nand U8556 (N_8556,N_8471,N_8469);
or U8557 (N_8557,N_8423,N_8419);
and U8558 (N_8558,N_8462,N_8455);
and U8559 (N_8559,N_8348,N_8444);
and U8560 (N_8560,N_8360,N_8430);
nor U8561 (N_8561,N_8435,N_8464);
and U8562 (N_8562,N_8378,N_8327);
nor U8563 (N_8563,N_8333,N_8426);
and U8564 (N_8564,N_8359,N_8461);
xor U8565 (N_8565,N_8449,N_8419);
and U8566 (N_8566,N_8422,N_8395);
nor U8567 (N_8567,N_8438,N_8353);
nand U8568 (N_8568,N_8442,N_8465);
or U8569 (N_8569,N_8325,N_8356);
and U8570 (N_8570,N_8375,N_8383);
nand U8571 (N_8571,N_8459,N_8441);
or U8572 (N_8572,N_8393,N_8322);
or U8573 (N_8573,N_8357,N_8395);
and U8574 (N_8574,N_8389,N_8433);
nor U8575 (N_8575,N_8425,N_8463);
and U8576 (N_8576,N_8360,N_8382);
nor U8577 (N_8577,N_8380,N_8462);
nor U8578 (N_8578,N_8474,N_8432);
nor U8579 (N_8579,N_8336,N_8335);
or U8580 (N_8580,N_8463,N_8441);
and U8581 (N_8581,N_8392,N_8454);
nor U8582 (N_8582,N_8441,N_8358);
nor U8583 (N_8583,N_8427,N_8386);
nand U8584 (N_8584,N_8328,N_8359);
xor U8585 (N_8585,N_8394,N_8351);
nand U8586 (N_8586,N_8479,N_8338);
or U8587 (N_8587,N_8384,N_8326);
or U8588 (N_8588,N_8350,N_8450);
nand U8589 (N_8589,N_8396,N_8407);
nand U8590 (N_8590,N_8421,N_8450);
and U8591 (N_8591,N_8420,N_8408);
and U8592 (N_8592,N_8459,N_8353);
nor U8593 (N_8593,N_8445,N_8442);
and U8594 (N_8594,N_8474,N_8385);
or U8595 (N_8595,N_8359,N_8479);
and U8596 (N_8596,N_8355,N_8321);
nand U8597 (N_8597,N_8416,N_8457);
xnor U8598 (N_8598,N_8400,N_8370);
and U8599 (N_8599,N_8440,N_8400);
and U8600 (N_8600,N_8454,N_8417);
and U8601 (N_8601,N_8342,N_8387);
or U8602 (N_8602,N_8383,N_8476);
xnor U8603 (N_8603,N_8321,N_8434);
or U8604 (N_8604,N_8398,N_8331);
or U8605 (N_8605,N_8381,N_8328);
nor U8606 (N_8606,N_8402,N_8425);
nand U8607 (N_8607,N_8324,N_8347);
nand U8608 (N_8608,N_8466,N_8399);
nor U8609 (N_8609,N_8348,N_8434);
and U8610 (N_8610,N_8322,N_8413);
nor U8611 (N_8611,N_8420,N_8446);
xnor U8612 (N_8612,N_8462,N_8354);
nor U8613 (N_8613,N_8406,N_8471);
xnor U8614 (N_8614,N_8441,N_8384);
nand U8615 (N_8615,N_8479,N_8372);
and U8616 (N_8616,N_8352,N_8391);
nor U8617 (N_8617,N_8385,N_8353);
nand U8618 (N_8618,N_8344,N_8374);
and U8619 (N_8619,N_8334,N_8349);
or U8620 (N_8620,N_8443,N_8440);
and U8621 (N_8621,N_8407,N_8397);
nor U8622 (N_8622,N_8464,N_8456);
nand U8623 (N_8623,N_8381,N_8420);
and U8624 (N_8624,N_8452,N_8439);
nand U8625 (N_8625,N_8389,N_8450);
or U8626 (N_8626,N_8478,N_8328);
and U8627 (N_8627,N_8386,N_8373);
and U8628 (N_8628,N_8473,N_8479);
and U8629 (N_8629,N_8380,N_8459);
nor U8630 (N_8630,N_8360,N_8449);
nor U8631 (N_8631,N_8437,N_8468);
xnor U8632 (N_8632,N_8432,N_8376);
nand U8633 (N_8633,N_8339,N_8449);
nand U8634 (N_8634,N_8383,N_8373);
nor U8635 (N_8635,N_8338,N_8320);
and U8636 (N_8636,N_8437,N_8355);
and U8637 (N_8637,N_8465,N_8365);
and U8638 (N_8638,N_8439,N_8432);
or U8639 (N_8639,N_8359,N_8411);
and U8640 (N_8640,N_8568,N_8603);
nor U8641 (N_8641,N_8512,N_8638);
nand U8642 (N_8642,N_8528,N_8495);
and U8643 (N_8643,N_8489,N_8578);
and U8644 (N_8644,N_8503,N_8569);
nor U8645 (N_8645,N_8635,N_8539);
or U8646 (N_8646,N_8585,N_8586);
and U8647 (N_8647,N_8560,N_8538);
nor U8648 (N_8648,N_8481,N_8570);
or U8649 (N_8649,N_8550,N_8488);
xor U8650 (N_8650,N_8541,N_8484);
and U8651 (N_8651,N_8629,N_8485);
and U8652 (N_8652,N_8624,N_8621);
nor U8653 (N_8653,N_8513,N_8532);
or U8654 (N_8654,N_8506,N_8514);
nor U8655 (N_8655,N_8627,N_8595);
nor U8656 (N_8656,N_8637,N_8483);
nor U8657 (N_8657,N_8566,N_8540);
or U8658 (N_8658,N_8599,N_8537);
nand U8659 (N_8659,N_8558,N_8553);
xor U8660 (N_8660,N_8497,N_8576);
or U8661 (N_8661,N_8623,N_8583);
nand U8662 (N_8662,N_8604,N_8554);
nor U8663 (N_8663,N_8557,N_8562);
nand U8664 (N_8664,N_8507,N_8622);
and U8665 (N_8665,N_8563,N_8504);
or U8666 (N_8666,N_8611,N_8609);
nor U8667 (N_8667,N_8620,N_8545);
nor U8668 (N_8668,N_8517,N_8527);
and U8669 (N_8669,N_8536,N_8574);
nor U8670 (N_8670,N_8582,N_8616);
nor U8671 (N_8671,N_8628,N_8602);
and U8672 (N_8672,N_8493,N_8480);
nor U8673 (N_8673,N_8523,N_8509);
nor U8674 (N_8674,N_8606,N_8525);
and U8675 (N_8675,N_8632,N_8533);
xnor U8676 (N_8676,N_8617,N_8519);
or U8677 (N_8677,N_8516,N_8605);
nor U8678 (N_8678,N_8494,N_8490);
xnor U8679 (N_8679,N_8577,N_8492);
nand U8680 (N_8680,N_8589,N_8598);
and U8681 (N_8681,N_8607,N_8587);
xnor U8682 (N_8682,N_8543,N_8564);
nand U8683 (N_8683,N_8592,N_8500);
and U8684 (N_8684,N_8594,N_8597);
nor U8685 (N_8685,N_8535,N_8588);
nor U8686 (N_8686,N_8548,N_8575);
nor U8687 (N_8687,N_8580,N_8612);
or U8688 (N_8688,N_8596,N_8501);
nor U8689 (N_8689,N_8498,N_8508);
nor U8690 (N_8690,N_8633,N_8505);
xnor U8691 (N_8691,N_8547,N_8534);
nand U8692 (N_8692,N_8613,N_8572);
nor U8693 (N_8693,N_8615,N_8549);
nand U8694 (N_8694,N_8515,N_8581);
and U8695 (N_8695,N_8551,N_8593);
or U8696 (N_8696,N_8531,N_8530);
and U8697 (N_8697,N_8482,N_8590);
nor U8698 (N_8698,N_8619,N_8639);
xor U8699 (N_8699,N_8510,N_8546);
or U8700 (N_8700,N_8556,N_8521);
or U8701 (N_8701,N_8511,N_8561);
nand U8702 (N_8702,N_8614,N_8610);
and U8703 (N_8703,N_8544,N_8567);
and U8704 (N_8704,N_8630,N_8542);
or U8705 (N_8705,N_8491,N_8486);
and U8706 (N_8706,N_8559,N_8573);
or U8707 (N_8707,N_8579,N_8502);
or U8708 (N_8708,N_8608,N_8600);
nand U8709 (N_8709,N_8526,N_8618);
nor U8710 (N_8710,N_8584,N_8522);
xor U8711 (N_8711,N_8626,N_8555);
nor U8712 (N_8712,N_8591,N_8631);
nand U8713 (N_8713,N_8524,N_8529);
nor U8714 (N_8714,N_8601,N_8634);
nor U8715 (N_8715,N_8496,N_8487);
nor U8716 (N_8716,N_8499,N_8636);
nor U8717 (N_8717,N_8571,N_8518);
and U8718 (N_8718,N_8565,N_8552);
nand U8719 (N_8719,N_8625,N_8520);
or U8720 (N_8720,N_8522,N_8511);
nor U8721 (N_8721,N_8591,N_8598);
and U8722 (N_8722,N_8610,N_8483);
nor U8723 (N_8723,N_8560,N_8624);
nor U8724 (N_8724,N_8633,N_8517);
or U8725 (N_8725,N_8488,N_8557);
nor U8726 (N_8726,N_8592,N_8590);
xnor U8727 (N_8727,N_8604,N_8553);
and U8728 (N_8728,N_8531,N_8485);
nor U8729 (N_8729,N_8498,N_8543);
and U8730 (N_8730,N_8569,N_8541);
or U8731 (N_8731,N_8489,N_8587);
nand U8732 (N_8732,N_8557,N_8495);
xor U8733 (N_8733,N_8579,N_8612);
and U8734 (N_8734,N_8496,N_8633);
nand U8735 (N_8735,N_8501,N_8575);
nand U8736 (N_8736,N_8513,N_8595);
xor U8737 (N_8737,N_8506,N_8573);
nor U8738 (N_8738,N_8583,N_8538);
nor U8739 (N_8739,N_8530,N_8635);
nor U8740 (N_8740,N_8599,N_8603);
nand U8741 (N_8741,N_8591,N_8639);
and U8742 (N_8742,N_8577,N_8490);
nor U8743 (N_8743,N_8588,N_8481);
and U8744 (N_8744,N_8513,N_8551);
nand U8745 (N_8745,N_8528,N_8497);
and U8746 (N_8746,N_8605,N_8549);
and U8747 (N_8747,N_8552,N_8595);
and U8748 (N_8748,N_8520,N_8493);
xor U8749 (N_8749,N_8490,N_8626);
nor U8750 (N_8750,N_8544,N_8556);
and U8751 (N_8751,N_8505,N_8504);
or U8752 (N_8752,N_8509,N_8585);
nor U8753 (N_8753,N_8496,N_8500);
or U8754 (N_8754,N_8595,N_8630);
or U8755 (N_8755,N_8590,N_8571);
or U8756 (N_8756,N_8491,N_8501);
and U8757 (N_8757,N_8606,N_8556);
nor U8758 (N_8758,N_8629,N_8559);
and U8759 (N_8759,N_8498,N_8535);
nand U8760 (N_8760,N_8505,N_8618);
or U8761 (N_8761,N_8569,N_8500);
and U8762 (N_8762,N_8612,N_8536);
nand U8763 (N_8763,N_8586,N_8592);
or U8764 (N_8764,N_8556,N_8500);
xor U8765 (N_8765,N_8524,N_8638);
or U8766 (N_8766,N_8630,N_8626);
nor U8767 (N_8767,N_8625,N_8541);
and U8768 (N_8768,N_8495,N_8608);
xnor U8769 (N_8769,N_8592,N_8622);
xor U8770 (N_8770,N_8556,N_8608);
and U8771 (N_8771,N_8599,N_8584);
or U8772 (N_8772,N_8515,N_8639);
and U8773 (N_8773,N_8534,N_8583);
xnor U8774 (N_8774,N_8499,N_8543);
xnor U8775 (N_8775,N_8517,N_8614);
or U8776 (N_8776,N_8619,N_8526);
nand U8777 (N_8777,N_8558,N_8581);
and U8778 (N_8778,N_8516,N_8530);
nand U8779 (N_8779,N_8482,N_8576);
and U8780 (N_8780,N_8499,N_8639);
nand U8781 (N_8781,N_8520,N_8539);
or U8782 (N_8782,N_8529,N_8559);
nor U8783 (N_8783,N_8635,N_8634);
nand U8784 (N_8784,N_8538,N_8629);
nand U8785 (N_8785,N_8516,N_8606);
and U8786 (N_8786,N_8498,N_8558);
and U8787 (N_8787,N_8588,N_8506);
xnor U8788 (N_8788,N_8489,N_8590);
nand U8789 (N_8789,N_8569,N_8630);
nor U8790 (N_8790,N_8497,N_8544);
and U8791 (N_8791,N_8606,N_8626);
nand U8792 (N_8792,N_8521,N_8611);
and U8793 (N_8793,N_8637,N_8523);
xor U8794 (N_8794,N_8638,N_8590);
nor U8795 (N_8795,N_8487,N_8489);
nand U8796 (N_8796,N_8589,N_8626);
or U8797 (N_8797,N_8639,N_8529);
nand U8798 (N_8798,N_8516,N_8531);
or U8799 (N_8799,N_8612,N_8550);
or U8800 (N_8800,N_8732,N_8698);
nand U8801 (N_8801,N_8670,N_8687);
nor U8802 (N_8802,N_8747,N_8699);
nor U8803 (N_8803,N_8682,N_8716);
xnor U8804 (N_8804,N_8713,N_8729);
nor U8805 (N_8805,N_8700,N_8757);
nor U8806 (N_8806,N_8706,N_8660);
and U8807 (N_8807,N_8701,N_8790);
and U8808 (N_8808,N_8694,N_8774);
nand U8809 (N_8809,N_8767,N_8691);
xnor U8810 (N_8810,N_8648,N_8715);
nor U8811 (N_8811,N_8754,N_8661);
nor U8812 (N_8812,N_8796,N_8748);
or U8813 (N_8813,N_8722,N_8772);
nand U8814 (N_8814,N_8656,N_8709);
xnor U8815 (N_8815,N_8725,N_8686);
xor U8816 (N_8816,N_8642,N_8766);
and U8817 (N_8817,N_8693,N_8647);
nand U8818 (N_8818,N_8668,N_8646);
nand U8819 (N_8819,N_8640,N_8741);
xor U8820 (N_8820,N_8692,N_8777);
nand U8821 (N_8821,N_8666,N_8650);
xor U8822 (N_8822,N_8655,N_8734);
or U8823 (N_8823,N_8778,N_8690);
nand U8824 (N_8824,N_8712,N_8679);
nand U8825 (N_8825,N_8753,N_8702);
nor U8826 (N_8826,N_8798,N_8781);
or U8827 (N_8827,N_8776,N_8685);
xor U8828 (N_8828,N_8703,N_8726);
nand U8829 (N_8829,N_8799,N_8784);
nor U8830 (N_8830,N_8676,N_8782);
xor U8831 (N_8831,N_8737,N_8762);
nor U8832 (N_8832,N_8675,N_8794);
and U8833 (N_8833,N_8704,N_8738);
and U8834 (N_8834,N_8736,N_8707);
nor U8835 (N_8835,N_8678,N_8688);
xnor U8836 (N_8836,N_8654,N_8758);
xnor U8837 (N_8837,N_8745,N_8728);
xor U8838 (N_8838,N_8651,N_8785);
nand U8839 (N_8839,N_8775,N_8789);
or U8840 (N_8840,N_8755,N_8756);
nand U8841 (N_8841,N_8730,N_8791);
or U8842 (N_8842,N_8669,N_8695);
or U8843 (N_8843,N_8718,N_8787);
or U8844 (N_8844,N_8770,N_8667);
nand U8845 (N_8845,N_8731,N_8733);
and U8846 (N_8846,N_8764,N_8793);
xnor U8847 (N_8847,N_8739,N_8657);
nor U8848 (N_8848,N_8743,N_8727);
or U8849 (N_8849,N_8689,N_8645);
and U8850 (N_8850,N_8721,N_8735);
or U8851 (N_8851,N_8644,N_8724);
or U8852 (N_8852,N_8740,N_8761);
nor U8853 (N_8853,N_8792,N_8786);
nand U8854 (N_8854,N_8677,N_8763);
nand U8855 (N_8855,N_8662,N_8674);
or U8856 (N_8856,N_8665,N_8795);
xnor U8857 (N_8857,N_8653,N_8765);
xnor U8858 (N_8858,N_8696,N_8769);
xor U8859 (N_8859,N_8750,N_8649);
and U8860 (N_8860,N_8671,N_8797);
xnor U8861 (N_8861,N_8759,N_8720);
and U8862 (N_8862,N_8672,N_8783);
nand U8863 (N_8863,N_8641,N_8719);
or U8864 (N_8864,N_8673,N_8683);
and U8865 (N_8865,N_8658,N_8717);
nand U8866 (N_8866,N_8681,N_8697);
nand U8867 (N_8867,N_8684,N_8652);
or U8868 (N_8868,N_8659,N_8788);
nor U8869 (N_8869,N_8708,N_8723);
nor U8870 (N_8870,N_8742,N_8680);
or U8871 (N_8871,N_8752,N_8643);
or U8872 (N_8872,N_8779,N_8746);
nor U8873 (N_8873,N_8780,N_8749);
and U8874 (N_8874,N_8710,N_8705);
or U8875 (N_8875,N_8664,N_8663);
or U8876 (N_8876,N_8744,N_8711);
nor U8877 (N_8877,N_8714,N_8768);
nor U8878 (N_8878,N_8760,N_8771);
or U8879 (N_8879,N_8773,N_8751);
nand U8880 (N_8880,N_8754,N_8640);
or U8881 (N_8881,N_8701,N_8776);
nor U8882 (N_8882,N_8791,N_8722);
xnor U8883 (N_8883,N_8644,N_8784);
nor U8884 (N_8884,N_8733,N_8643);
nand U8885 (N_8885,N_8674,N_8694);
xor U8886 (N_8886,N_8785,N_8775);
and U8887 (N_8887,N_8790,N_8786);
or U8888 (N_8888,N_8660,N_8790);
nand U8889 (N_8889,N_8657,N_8790);
xor U8890 (N_8890,N_8659,N_8662);
nand U8891 (N_8891,N_8771,N_8644);
nand U8892 (N_8892,N_8715,N_8650);
or U8893 (N_8893,N_8766,N_8755);
and U8894 (N_8894,N_8721,N_8755);
or U8895 (N_8895,N_8751,N_8744);
xnor U8896 (N_8896,N_8681,N_8727);
and U8897 (N_8897,N_8665,N_8755);
or U8898 (N_8898,N_8798,N_8711);
nand U8899 (N_8899,N_8682,N_8707);
xor U8900 (N_8900,N_8647,N_8682);
and U8901 (N_8901,N_8777,N_8789);
nor U8902 (N_8902,N_8682,N_8724);
nand U8903 (N_8903,N_8663,N_8681);
xor U8904 (N_8904,N_8774,N_8797);
or U8905 (N_8905,N_8688,N_8698);
xor U8906 (N_8906,N_8670,N_8756);
or U8907 (N_8907,N_8734,N_8771);
xnor U8908 (N_8908,N_8784,N_8695);
and U8909 (N_8909,N_8725,N_8713);
nor U8910 (N_8910,N_8772,N_8717);
nand U8911 (N_8911,N_8654,N_8762);
xnor U8912 (N_8912,N_8703,N_8679);
nor U8913 (N_8913,N_8659,N_8660);
xor U8914 (N_8914,N_8764,N_8651);
or U8915 (N_8915,N_8779,N_8705);
nand U8916 (N_8916,N_8732,N_8756);
and U8917 (N_8917,N_8760,N_8753);
xor U8918 (N_8918,N_8747,N_8652);
and U8919 (N_8919,N_8644,N_8681);
or U8920 (N_8920,N_8752,N_8653);
xor U8921 (N_8921,N_8791,N_8655);
nor U8922 (N_8922,N_8670,N_8713);
nand U8923 (N_8923,N_8788,N_8676);
or U8924 (N_8924,N_8723,N_8755);
xnor U8925 (N_8925,N_8716,N_8664);
or U8926 (N_8926,N_8734,N_8646);
nor U8927 (N_8927,N_8725,N_8735);
nor U8928 (N_8928,N_8757,N_8780);
and U8929 (N_8929,N_8645,N_8764);
xor U8930 (N_8930,N_8679,N_8716);
nor U8931 (N_8931,N_8667,N_8680);
nor U8932 (N_8932,N_8658,N_8684);
or U8933 (N_8933,N_8724,N_8749);
or U8934 (N_8934,N_8671,N_8756);
nor U8935 (N_8935,N_8654,N_8756);
nand U8936 (N_8936,N_8674,N_8726);
nand U8937 (N_8937,N_8670,N_8641);
and U8938 (N_8938,N_8748,N_8738);
and U8939 (N_8939,N_8792,N_8776);
or U8940 (N_8940,N_8794,N_8693);
and U8941 (N_8941,N_8745,N_8675);
xnor U8942 (N_8942,N_8766,N_8701);
nor U8943 (N_8943,N_8751,N_8668);
nor U8944 (N_8944,N_8650,N_8713);
and U8945 (N_8945,N_8768,N_8674);
and U8946 (N_8946,N_8760,N_8745);
or U8947 (N_8947,N_8773,N_8676);
or U8948 (N_8948,N_8768,N_8710);
and U8949 (N_8949,N_8689,N_8799);
or U8950 (N_8950,N_8698,N_8724);
nand U8951 (N_8951,N_8722,N_8787);
and U8952 (N_8952,N_8686,N_8720);
or U8953 (N_8953,N_8641,N_8659);
nand U8954 (N_8954,N_8692,N_8767);
or U8955 (N_8955,N_8788,N_8799);
nor U8956 (N_8956,N_8684,N_8755);
nand U8957 (N_8957,N_8792,N_8755);
nand U8958 (N_8958,N_8778,N_8779);
nand U8959 (N_8959,N_8754,N_8774);
nand U8960 (N_8960,N_8822,N_8810);
and U8961 (N_8961,N_8809,N_8949);
and U8962 (N_8962,N_8882,N_8944);
and U8963 (N_8963,N_8806,N_8837);
nor U8964 (N_8964,N_8878,N_8946);
and U8965 (N_8965,N_8803,N_8860);
nand U8966 (N_8966,N_8816,N_8853);
xnor U8967 (N_8967,N_8856,N_8802);
xor U8968 (N_8968,N_8814,N_8848);
or U8969 (N_8969,N_8825,N_8874);
nor U8970 (N_8970,N_8945,N_8903);
nand U8971 (N_8971,N_8935,N_8893);
nand U8972 (N_8972,N_8879,N_8915);
or U8973 (N_8973,N_8920,N_8885);
and U8974 (N_8974,N_8832,N_8890);
nor U8975 (N_8975,N_8954,N_8869);
nor U8976 (N_8976,N_8804,N_8900);
xnor U8977 (N_8977,N_8880,N_8896);
nand U8978 (N_8978,N_8957,N_8811);
nor U8979 (N_8979,N_8863,N_8948);
nor U8980 (N_8980,N_8892,N_8898);
or U8981 (N_8981,N_8934,N_8905);
nand U8982 (N_8982,N_8932,N_8858);
and U8983 (N_8983,N_8894,N_8844);
nand U8984 (N_8984,N_8836,N_8924);
xor U8985 (N_8985,N_8955,N_8897);
or U8986 (N_8986,N_8805,N_8818);
or U8987 (N_8987,N_8865,N_8851);
xor U8988 (N_8988,N_8927,N_8908);
and U8989 (N_8989,N_8956,N_8801);
nand U8990 (N_8990,N_8943,N_8936);
or U8991 (N_8991,N_8930,N_8847);
and U8992 (N_8992,N_8852,N_8928);
nor U8993 (N_8993,N_8872,N_8929);
and U8994 (N_8994,N_8933,N_8827);
nand U8995 (N_8995,N_8922,N_8888);
nand U8996 (N_8996,N_8800,N_8876);
xnor U8997 (N_8997,N_8891,N_8902);
xnor U8998 (N_8998,N_8895,N_8906);
nor U8999 (N_8999,N_8829,N_8864);
xor U9000 (N_9000,N_8862,N_8901);
and U9001 (N_9001,N_8839,N_8925);
nor U9002 (N_9002,N_8824,N_8889);
or U9003 (N_9003,N_8840,N_8833);
or U9004 (N_9004,N_8857,N_8884);
or U9005 (N_9005,N_8870,N_8831);
or U9006 (N_9006,N_8850,N_8821);
nor U9007 (N_9007,N_8812,N_8923);
or U9008 (N_9008,N_8849,N_8938);
and U9009 (N_9009,N_8947,N_8941);
xnor U9010 (N_9010,N_8913,N_8919);
and U9011 (N_9011,N_8859,N_8921);
or U9012 (N_9012,N_8912,N_8931);
or U9013 (N_9013,N_8939,N_8910);
nor U9014 (N_9014,N_8875,N_8917);
xor U9015 (N_9015,N_8907,N_8819);
and U9016 (N_9016,N_8820,N_8826);
nor U9017 (N_9017,N_8883,N_8861);
xor U9018 (N_9018,N_8873,N_8830);
xor U9019 (N_9019,N_8823,N_8942);
or U9020 (N_9020,N_8877,N_8911);
nor U9021 (N_9021,N_8855,N_8854);
and U9022 (N_9022,N_8886,N_8953);
and U9023 (N_9023,N_8807,N_8845);
nor U9024 (N_9024,N_8842,N_8959);
xor U9025 (N_9025,N_8843,N_8867);
and U9026 (N_9026,N_8828,N_8940);
nand U9027 (N_9027,N_8841,N_8916);
xor U9028 (N_9028,N_8899,N_8817);
nor U9029 (N_9029,N_8958,N_8926);
nand U9030 (N_9030,N_8918,N_8937);
xor U9031 (N_9031,N_8871,N_8951);
or U9032 (N_9032,N_8904,N_8881);
nor U9033 (N_9033,N_8813,N_8838);
xor U9034 (N_9034,N_8835,N_8909);
and U9035 (N_9035,N_8914,N_8834);
xnor U9036 (N_9036,N_8846,N_8887);
nand U9037 (N_9037,N_8808,N_8868);
nor U9038 (N_9038,N_8950,N_8866);
xor U9039 (N_9039,N_8952,N_8815);
or U9040 (N_9040,N_8890,N_8899);
or U9041 (N_9041,N_8819,N_8838);
or U9042 (N_9042,N_8800,N_8938);
and U9043 (N_9043,N_8815,N_8867);
nor U9044 (N_9044,N_8834,N_8836);
xnor U9045 (N_9045,N_8849,N_8817);
and U9046 (N_9046,N_8911,N_8958);
or U9047 (N_9047,N_8896,N_8939);
xnor U9048 (N_9048,N_8827,N_8925);
nand U9049 (N_9049,N_8845,N_8938);
xor U9050 (N_9050,N_8958,N_8852);
and U9051 (N_9051,N_8850,N_8829);
nand U9052 (N_9052,N_8837,N_8916);
xnor U9053 (N_9053,N_8891,N_8854);
nor U9054 (N_9054,N_8878,N_8875);
nand U9055 (N_9055,N_8865,N_8859);
xor U9056 (N_9056,N_8813,N_8802);
or U9057 (N_9057,N_8840,N_8900);
nor U9058 (N_9058,N_8917,N_8841);
nand U9059 (N_9059,N_8915,N_8876);
nand U9060 (N_9060,N_8861,N_8915);
and U9061 (N_9061,N_8828,N_8859);
nor U9062 (N_9062,N_8874,N_8951);
or U9063 (N_9063,N_8871,N_8859);
and U9064 (N_9064,N_8865,N_8950);
and U9065 (N_9065,N_8868,N_8800);
nand U9066 (N_9066,N_8952,N_8801);
and U9067 (N_9067,N_8896,N_8936);
and U9068 (N_9068,N_8921,N_8823);
and U9069 (N_9069,N_8940,N_8834);
and U9070 (N_9070,N_8896,N_8942);
nand U9071 (N_9071,N_8925,N_8895);
or U9072 (N_9072,N_8882,N_8902);
nand U9073 (N_9073,N_8873,N_8810);
xor U9074 (N_9074,N_8896,N_8841);
and U9075 (N_9075,N_8822,N_8953);
xnor U9076 (N_9076,N_8882,N_8814);
nor U9077 (N_9077,N_8924,N_8869);
xor U9078 (N_9078,N_8931,N_8891);
or U9079 (N_9079,N_8820,N_8920);
xor U9080 (N_9080,N_8914,N_8899);
xor U9081 (N_9081,N_8865,N_8829);
nand U9082 (N_9082,N_8940,N_8905);
nor U9083 (N_9083,N_8834,N_8821);
or U9084 (N_9084,N_8823,N_8886);
xor U9085 (N_9085,N_8947,N_8855);
nand U9086 (N_9086,N_8818,N_8885);
nor U9087 (N_9087,N_8882,N_8894);
and U9088 (N_9088,N_8861,N_8840);
xor U9089 (N_9089,N_8952,N_8842);
xor U9090 (N_9090,N_8859,N_8850);
or U9091 (N_9091,N_8875,N_8835);
or U9092 (N_9092,N_8943,N_8865);
nor U9093 (N_9093,N_8878,N_8948);
nor U9094 (N_9094,N_8804,N_8818);
xnor U9095 (N_9095,N_8942,N_8875);
nand U9096 (N_9096,N_8953,N_8925);
xnor U9097 (N_9097,N_8920,N_8875);
nor U9098 (N_9098,N_8865,N_8896);
nand U9099 (N_9099,N_8887,N_8804);
nand U9100 (N_9100,N_8947,N_8844);
xnor U9101 (N_9101,N_8890,N_8865);
nand U9102 (N_9102,N_8875,N_8934);
nand U9103 (N_9103,N_8829,N_8804);
nor U9104 (N_9104,N_8951,N_8904);
nor U9105 (N_9105,N_8955,N_8878);
or U9106 (N_9106,N_8930,N_8866);
xnor U9107 (N_9107,N_8856,N_8901);
xor U9108 (N_9108,N_8929,N_8898);
nand U9109 (N_9109,N_8922,N_8845);
and U9110 (N_9110,N_8884,N_8933);
and U9111 (N_9111,N_8909,N_8865);
nor U9112 (N_9112,N_8900,N_8929);
xor U9113 (N_9113,N_8941,N_8803);
and U9114 (N_9114,N_8949,N_8808);
nand U9115 (N_9115,N_8900,N_8823);
or U9116 (N_9116,N_8940,N_8835);
and U9117 (N_9117,N_8809,N_8893);
nand U9118 (N_9118,N_8943,N_8873);
nand U9119 (N_9119,N_8919,N_8902);
xnor U9120 (N_9120,N_9017,N_8990);
nor U9121 (N_9121,N_9119,N_8962);
nand U9122 (N_9122,N_9022,N_9108);
or U9123 (N_9123,N_9019,N_9035);
nor U9124 (N_9124,N_9070,N_8961);
nor U9125 (N_9125,N_9029,N_9015);
nand U9126 (N_9126,N_9067,N_9002);
or U9127 (N_9127,N_9095,N_9089);
xor U9128 (N_9128,N_9050,N_9071);
nand U9129 (N_9129,N_9012,N_9052);
and U9130 (N_9130,N_9093,N_9109);
nand U9131 (N_9131,N_9030,N_9091);
nor U9132 (N_9132,N_9110,N_9044);
nand U9133 (N_9133,N_9032,N_8984);
nand U9134 (N_9134,N_8987,N_9046);
and U9135 (N_9135,N_9008,N_9049);
and U9136 (N_9136,N_9018,N_9006);
nor U9137 (N_9137,N_9073,N_8971);
and U9138 (N_9138,N_9026,N_9083);
and U9139 (N_9139,N_9085,N_9025);
xnor U9140 (N_9140,N_8993,N_8965);
nand U9141 (N_9141,N_8996,N_9078);
nand U9142 (N_9142,N_9102,N_8985);
or U9143 (N_9143,N_9097,N_8999);
nor U9144 (N_9144,N_9003,N_9082);
and U9145 (N_9145,N_9031,N_9023);
or U9146 (N_9146,N_9028,N_8963);
or U9147 (N_9147,N_8982,N_8981);
and U9148 (N_9148,N_9105,N_9053);
and U9149 (N_9149,N_9090,N_9024);
nand U9150 (N_9150,N_9036,N_9034);
or U9151 (N_9151,N_9103,N_8973);
xnor U9152 (N_9152,N_9021,N_9057);
or U9153 (N_9153,N_9088,N_9084);
and U9154 (N_9154,N_8977,N_9069);
or U9155 (N_9155,N_8967,N_9045);
and U9156 (N_9156,N_8966,N_9016);
nand U9157 (N_9157,N_9059,N_9062);
nor U9158 (N_9158,N_9096,N_9063);
and U9159 (N_9159,N_9117,N_9099);
nor U9160 (N_9160,N_9094,N_9043);
xnor U9161 (N_9161,N_8989,N_8986);
or U9162 (N_9162,N_9011,N_9007);
and U9163 (N_9163,N_9041,N_9054);
or U9164 (N_9164,N_8969,N_8994);
nor U9165 (N_9165,N_9040,N_9081);
nor U9166 (N_9166,N_9009,N_9113);
and U9167 (N_9167,N_8960,N_9056);
nand U9168 (N_9168,N_9000,N_9051);
xnor U9169 (N_9169,N_9020,N_8978);
xor U9170 (N_9170,N_8972,N_9039);
and U9171 (N_9171,N_8964,N_9013);
or U9172 (N_9172,N_9076,N_9004);
or U9173 (N_9173,N_8983,N_9107);
xor U9174 (N_9174,N_9037,N_8988);
or U9175 (N_9175,N_8992,N_9106);
or U9176 (N_9176,N_9058,N_9101);
or U9177 (N_9177,N_9112,N_8980);
xor U9178 (N_9178,N_9072,N_9048);
nand U9179 (N_9179,N_8968,N_8976);
nor U9180 (N_9180,N_8974,N_9060);
and U9181 (N_9181,N_9042,N_9114);
and U9182 (N_9182,N_8995,N_9116);
and U9183 (N_9183,N_8991,N_9092);
nor U9184 (N_9184,N_9001,N_9080);
nor U9185 (N_9185,N_9074,N_9055);
xnor U9186 (N_9186,N_9047,N_9033);
and U9187 (N_9187,N_9077,N_9061);
or U9188 (N_9188,N_9005,N_9027);
or U9189 (N_9189,N_9118,N_9010);
and U9190 (N_9190,N_9066,N_9111);
nor U9191 (N_9191,N_9075,N_9065);
nor U9192 (N_9192,N_9079,N_9064);
or U9193 (N_9193,N_9098,N_8979);
nand U9194 (N_9194,N_9038,N_9115);
and U9195 (N_9195,N_9087,N_9086);
or U9196 (N_9196,N_9014,N_9100);
nand U9197 (N_9197,N_9104,N_8998);
nor U9198 (N_9198,N_9068,N_8970);
and U9199 (N_9199,N_8997,N_8975);
nor U9200 (N_9200,N_8984,N_9085);
nor U9201 (N_9201,N_9048,N_9074);
or U9202 (N_9202,N_9056,N_9108);
nand U9203 (N_9203,N_8992,N_8988);
nand U9204 (N_9204,N_8975,N_9108);
and U9205 (N_9205,N_8989,N_9090);
nand U9206 (N_9206,N_9102,N_9023);
or U9207 (N_9207,N_9039,N_9103);
nand U9208 (N_9208,N_8992,N_9027);
xnor U9209 (N_9209,N_8998,N_9096);
or U9210 (N_9210,N_9119,N_8996);
xnor U9211 (N_9211,N_9066,N_9034);
nor U9212 (N_9212,N_9109,N_9085);
nand U9213 (N_9213,N_9014,N_9086);
or U9214 (N_9214,N_9024,N_9021);
or U9215 (N_9215,N_9033,N_9116);
xor U9216 (N_9216,N_9095,N_9010);
nor U9217 (N_9217,N_9051,N_9061);
xnor U9218 (N_9218,N_9079,N_9018);
xor U9219 (N_9219,N_9112,N_8992);
nand U9220 (N_9220,N_9095,N_9066);
and U9221 (N_9221,N_8964,N_9034);
nor U9222 (N_9222,N_9111,N_9057);
xor U9223 (N_9223,N_9031,N_9115);
and U9224 (N_9224,N_9101,N_9030);
and U9225 (N_9225,N_9041,N_8972);
nand U9226 (N_9226,N_9083,N_9119);
nor U9227 (N_9227,N_9093,N_9070);
and U9228 (N_9228,N_8964,N_9041);
nand U9229 (N_9229,N_9082,N_9006);
nand U9230 (N_9230,N_9067,N_9081);
nand U9231 (N_9231,N_9075,N_9099);
nand U9232 (N_9232,N_9112,N_9102);
xnor U9233 (N_9233,N_9069,N_9088);
nand U9234 (N_9234,N_9024,N_9105);
xor U9235 (N_9235,N_9093,N_9086);
nand U9236 (N_9236,N_8974,N_9117);
and U9237 (N_9237,N_9090,N_8986);
and U9238 (N_9238,N_9072,N_9035);
nor U9239 (N_9239,N_9052,N_9092);
or U9240 (N_9240,N_9021,N_8972);
nand U9241 (N_9241,N_9000,N_9068);
or U9242 (N_9242,N_8994,N_9098);
xnor U9243 (N_9243,N_9119,N_9047);
and U9244 (N_9244,N_9069,N_9100);
and U9245 (N_9245,N_8989,N_9032);
nor U9246 (N_9246,N_9118,N_9054);
nor U9247 (N_9247,N_9058,N_8980);
nand U9248 (N_9248,N_9105,N_8997);
nor U9249 (N_9249,N_8965,N_9034);
xnor U9250 (N_9250,N_9018,N_8995);
nand U9251 (N_9251,N_8967,N_9099);
xnor U9252 (N_9252,N_8987,N_9068);
nor U9253 (N_9253,N_9019,N_9016);
xor U9254 (N_9254,N_9119,N_8984);
nand U9255 (N_9255,N_9008,N_9093);
and U9256 (N_9256,N_8960,N_8975);
nand U9257 (N_9257,N_8980,N_8978);
nand U9258 (N_9258,N_9027,N_8994);
and U9259 (N_9259,N_9008,N_8982);
and U9260 (N_9260,N_9102,N_9012);
nand U9261 (N_9261,N_9021,N_9012);
and U9262 (N_9262,N_9076,N_9037);
nand U9263 (N_9263,N_9113,N_9109);
or U9264 (N_9264,N_9043,N_8971);
nand U9265 (N_9265,N_9024,N_9083);
xnor U9266 (N_9266,N_9111,N_9034);
nor U9267 (N_9267,N_8995,N_8990);
nor U9268 (N_9268,N_8997,N_8993);
nand U9269 (N_9269,N_8965,N_8975);
nand U9270 (N_9270,N_9076,N_9024);
nor U9271 (N_9271,N_9116,N_8992);
nor U9272 (N_9272,N_9117,N_8999);
nor U9273 (N_9273,N_9086,N_9066);
nand U9274 (N_9274,N_9047,N_8960);
nand U9275 (N_9275,N_8994,N_9065);
and U9276 (N_9276,N_8985,N_9103);
nor U9277 (N_9277,N_9099,N_9028);
and U9278 (N_9278,N_9085,N_9081);
and U9279 (N_9279,N_9096,N_9019);
nand U9280 (N_9280,N_9124,N_9260);
xnor U9281 (N_9281,N_9166,N_9185);
or U9282 (N_9282,N_9203,N_9188);
or U9283 (N_9283,N_9164,N_9227);
nand U9284 (N_9284,N_9231,N_9120);
nor U9285 (N_9285,N_9208,N_9222);
nor U9286 (N_9286,N_9234,N_9244);
or U9287 (N_9287,N_9235,N_9254);
or U9288 (N_9288,N_9159,N_9137);
xnor U9289 (N_9289,N_9195,N_9276);
nand U9290 (N_9290,N_9155,N_9136);
nand U9291 (N_9291,N_9247,N_9245);
and U9292 (N_9292,N_9153,N_9125);
and U9293 (N_9293,N_9233,N_9157);
or U9294 (N_9294,N_9211,N_9161);
or U9295 (N_9295,N_9266,N_9206);
xor U9296 (N_9296,N_9148,N_9241);
nand U9297 (N_9297,N_9184,N_9144);
or U9298 (N_9298,N_9189,N_9232);
nor U9299 (N_9299,N_9223,N_9123);
nand U9300 (N_9300,N_9174,N_9221);
nor U9301 (N_9301,N_9212,N_9228);
and U9302 (N_9302,N_9261,N_9275);
and U9303 (N_9303,N_9214,N_9200);
nand U9304 (N_9304,N_9230,N_9171);
nor U9305 (N_9305,N_9135,N_9187);
and U9306 (N_9306,N_9173,N_9249);
and U9307 (N_9307,N_9240,N_9140);
xor U9308 (N_9308,N_9237,N_9149);
xor U9309 (N_9309,N_9224,N_9186);
nor U9310 (N_9310,N_9251,N_9156);
nand U9311 (N_9311,N_9197,N_9277);
xor U9312 (N_9312,N_9278,N_9257);
nand U9313 (N_9313,N_9150,N_9246);
xor U9314 (N_9314,N_9128,N_9215);
xor U9315 (N_9315,N_9194,N_9141);
and U9316 (N_9316,N_9170,N_9252);
nand U9317 (N_9317,N_9178,N_9248);
nand U9318 (N_9318,N_9134,N_9145);
nor U9319 (N_9319,N_9272,N_9122);
nor U9320 (N_9320,N_9167,N_9250);
nor U9321 (N_9321,N_9218,N_9265);
nand U9322 (N_9322,N_9151,N_9169);
nor U9323 (N_9323,N_9210,N_9191);
xnor U9324 (N_9324,N_9269,N_9179);
xnor U9325 (N_9325,N_9152,N_9274);
nor U9326 (N_9326,N_9273,N_9130);
xnor U9327 (N_9327,N_9243,N_9142);
nand U9328 (N_9328,N_9263,N_9193);
and U9329 (N_9329,N_9176,N_9138);
xnor U9330 (N_9330,N_9143,N_9132);
nand U9331 (N_9331,N_9204,N_9201);
nor U9332 (N_9332,N_9239,N_9207);
xor U9333 (N_9333,N_9262,N_9205);
or U9334 (N_9334,N_9270,N_9147);
or U9335 (N_9335,N_9220,N_9202);
xnor U9336 (N_9336,N_9271,N_9238);
or U9337 (N_9337,N_9253,N_9180);
nand U9338 (N_9338,N_9177,N_9217);
nand U9339 (N_9339,N_9264,N_9259);
or U9340 (N_9340,N_9213,N_9139);
xor U9341 (N_9341,N_9216,N_9183);
and U9342 (N_9342,N_9255,N_9160);
xnor U9343 (N_9343,N_9225,N_9163);
and U9344 (N_9344,N_9154,N_9229);
nand U9345 (N_9345,N_9198,N_9181);
or U9346 (N_9346,N_9162,N_9258);
nor U9347 (N_9347,N_9256,N_9127);
and U9348 (N_9348,N_9190,N_9192);
and U9349 (N_9349,N_9267,N_9209);
and U9350 (N_9350,N_9121,N_9182);
xor U9351 (N_9351,N_9196,N_9165);
and U9352 (N_9352,N_9268,N_9129);
xnor U9353 (N_9353,N_9199,N_9279);
nor U9354 (N_9354,N_9219,N_9126);
nor U9355 (N_9355,N_9226,N_9133);
nand U9356 (N_9356,N_9131,N_9175);
and U9357 (N_9357,N_9158,N_9172);
xnor U9358 (N_9358,N_9146,N_9242);
nor U9359 (N_9359,N_9236,N_9168);
nor U9360 (N_9360,N_9130,N_9194);
nand U9361 (N_9361,N_9158,N_9131);
xor U9362 (N_9362,N_9133,N_9275);
nor U9363 (N_9363,N_9261,N_9203);
nor U9364 (N_9364,N_9211,N_9160);
and U9365 (N_9365,N_9167,N_9232);
nor U9366 (N_9366,N_9265,N_9262);
or U9367 (N_9367,N_9201,N_9236);
nor U9368 (N_9368,N_9263,N_9258);
nand U9369 (N_9369,N_9243,N_9205);
nand U9370 (N_9370,N_9226,N_9236);
xnor U9371 (N_9371,N_9202,N_9144);
and U9372 (N_9372,N_9195,N_9147);
and U9373 (N_9373,N_9127,N_9162);
nand U9374 (N_9374,N_9225,N_9248);
nor U9375 (N_9375,N_9165,N_9240);
xnor U9376 (N_9376,N_9186,N_9278);
and U9377 (N_9377,N_9266,N_9234);
xor U9378 (N_9378,N_9138,N_9203);
and U9379 (N_9379,N_9196,N_9150);
and U9380 (N_9380,N_9257,N_9262);
nand U9381 (N_9381,N_9252,N_9164);
and U9382 (N_9382,N_9228,N_9224);
and U9383 (N_9383,N_9229,N_9139);
xor U9384 (N_9384,N_9250,N_9247);
and U9385 (N_9385,N_9148,N_9204);
xnor U9386 (N_9386,N_9186,N_9195);
and U9387 (N_9387,N_9124,N_9152);
and U9388 (N_9388,N_9155,N_9185);
nor U9389 (N_9389,N_9251,N_9220);
nor U9390 (N_9390,N_9258,N_9239);
or U9391 (N_9391,N_9154,N_9185);
or U9392 (N_9392,N_9154,N_9263);
or U9393 (N_9393,N_9240,N_9147);
xnor U9394 (N_9394,N_9214,N_9244);
or U9395 (N_9395,N_9169,N_9172);
nand U9396 (N_9396,N_9257,N_9279);
and U9397 (N_9397,N_9214,N_9151);
nor U9398 (N_9398,N_9181,N_9209);
xnor U9399 (N_9399,N_9271,N_9182);
xnor U9400 (N_9400,N_9147,N_9170);
or U9401 (N_9401,N_9124,N_9217);
nor U9402 (N_9402,N_9211,N_9183);
nor U9403 (N_9403,N_9127,N_9179);
nand U9404 (N_9404,N_9228,N_9155);
nand U9405 (N_9405,N_9211,N_9247);
nand U9406 (N_9406,N_9148,N_9213);
or U9407 (N_9407,N_9175,N_9123);
or U9408 (N_9408,N_9214,N_9155);
xor U9409 (N_9409,N_9127,N_9128);
nand U9410 (N_9410,N_9256,N_9160);
xor U9411 (N_9411,N_9219,N_9153);
nand U9412 (N_9412,N_9279,N_9222);
nand U9413 (N_9413,N_9234,N_9224);
xor U9414 (N_9414,N_9177,N_9147);
and U9415 (N_9415,N_9153,N_9191);
or U9416 (N_9416,N_9186,N_9215);
xnor U9417 (N_9417,N_9250,N_9193);
nand U9418 (N_9418,N_9212,N_9153);
xor U9419 (N_9419,N_9171,N_9196);
nand U9420 (N_9420,N_9140,N_9270);
and U9421 (N_9421,N_9211,N_9257);
xor U9422 (N_9422,N_9134,N_9146);
nor U9423 (N_9423,N_9147,N_9135);
xor U9424 (N_9424,N_9268,N_9192);
and U9425 (N_9425,N_9204,N_9260);
nor U9426 (N_9426,N_9187,N_9132);
and U9427 (N_9427,N_9261,N_9186);
and U9428 (N_9428,N_9165,N_9215);
and U9429 (N_9429,N_9261,N_9258);
nor U9430 (N_9430,N_9150,N_9248);
and U9431 (N_9431,N_9199,N_9246);
nor U9432 (N_9432,N_9228,N_9136);
nor U9433 (N_9433,N_9163,N_9232);
and U9434 (N_9434,N_9261,N_9125);
nor U9435 (N_9435,N_9249,N_9143);
xor U9436 (N_9436,N_9183,N_9195);
or U9437 (N_9437,N_9120,N_9223);
xnor U9438 (N_9438,N_9132,N_9235);
and U9439 (N_9439,N_9159,N_9192);
nor U9440 (N_9440,N_9365,N_9317);
nand U9441 (N_9441,N_9327,N_9383);
nor U9442 (N_9442,N_9298,N_9427);
nor U9443 (N_9443,N_9303,N_9407);
nand U9444 (N_9444,N_9429,N_9409);
xnor U9445 (N_9445,N_9307,N_9325);
nand U9446 (N_9446,N_9357,N_9356);
nor U9447 (N_9447,N_9311,N_9399);
nand U9448 (N_9448,N_9377,N_9355);
xnor U9449 (N_9449,N_9374,N_9305);
and U9450 (N_9450,N_9284,N_9351);
nor U9451 (N_9451,N_9406,N_9397);
or U9452 (N_9452,N_9359,N_9439);
nor U9453 (N_9453,N_9358,N_9432);
nor U9454 (N_9454,N_9371,N_9372);
nor U9455 (N_9455,N_9316,N_9391);
nand U9456 (N_9456,N_9425,N_9438);
and U9457 (N_9457,N_9286,N_9283);
xnor U9458 (N_9458,N_9296,N_9402);
and U9459 (N_9459,N_9349,N_9414);
nor U9460 (N_9460,N_9424,N_9426);
xnor U9461 (N_9461,N_9434,N_9423);
xnor U9462 (N_9462,N_9321,N_9376);
and U9463 (N_9463,N_9300,N_9430);
or U9464 (N_9464,N_9369,N_9341);
nor U9465 (N_9465,N_9422,N_9361);
and U9466 (N_9466,N_9313,N_9353);
nand U9467 (N_9467,N_9431,N_9331);
nor U9468 (N_9468,N_9398,N_9363);
xnor U9469 (N_9469,N_9337,N_9392);
nor U9470 (N_9470,N_9435,N_9345);
xnor U9471 (N_9471,N_9322,N_9396);
xnor U9472 (N_9472,N_9304,N_9410);
nand U9473 (N_9473,N_9384,N_9417);
nand U9474 (N_9474,N_9285,N_9437);
nor U9475 (N_9475,N_9360,N_9312);
nor U9476 (N_9476,N_9385,N_9290);
nand U9477 (N_9477,N_9389,N_9299);
xnor U9478 (N_9478,N_9289,N_9366);
nand U9479 (N_9479,N_9338,N_9315);
nor U9480 (N_9480,N_9401,N_9343);
nand U9481 (N_9481,N_9352,N_9308);
nand U9482 (N_9482,N_9326,N_9293);
and U9483 (N_9483,N_9387,N_9280);
xnor U9484 (N_9484,N_9403,N_9421);
nor U9485 (N_9485,N_9428,N_9332);
nand U9486 (N_9486,N_9301,N_9368);
or U9487 (N_9487,N_9405,N_9388);
and U9488 (N_9488,N_9318,N_9418);
xor U9489 (N_9489,N_9333,N_9281);
xnor U9490 (N_9490,N_9306,N_9297);
nor U9491 (N_9491,N_9314,N_9292);
nor U9492 (N_9492,N_9394,N_9320);
nand U9493 (N_9493,N_9287,N_9393);
xor U9494 (N_9494,N_9404,N_9294);
or U9495 (N_9495,N_9324,N_9302);
and U9496 (N_9496,N_9346,N_9330);
and U9497 (N_9497,N_9334,N_9339);
or U9498 (N_9498,N_9408,N_9362);
nand U9499 (N_9499,N_9347,N_9319);
xnor U9500 (N_9500,N_9386,N_9354);
or U9501 (N_9501,N_9413,N_9411);
and U9502 (N_9502,N_9379,N_9323);
and U9503 (N_9503,N_9415,N_9350);
and U9504 (N_9504,N_9364,N_9310);
nor U9505 (N_9505,N_9309,N_9335);
and U9506 (N_9506,N_9381,N_9390);
and U9507 (N_9507,N_9342,N_9433);
or U9508 (N_9508,N_9419,N_9378);
xor U9509 (N_9509,N_9367,N_9382);
or U9510 (N_9510,N_9288,N_9412);
or U9511 (N_9511,N_9373,N_9329);
nand U9512 (N_9512,N_9380,N_9375);
nor U9513 (N_9513,N_9291,N_9370);
or U9514 (N_9514,N_9416,N_9340);
nor U9515 (N_9515,N_9282,N_9336);
nor U9516 (N_9516,N_9328,N_9400);
nand U9517 (N_9517,N_9344,N_9348);
and U9518 (N_9518,N_9420,N_9295);
and U9519 (N_9519,N_9436,N_9395);
nand U9520 (N_9520,N_9403,N_9288);
xnor U9521 (N_9521,N_9394,N_9289);
xor U9522 (N_9522,N_9436,N_9388);
nor U9523 (N_9523,N_9325,N_9341);
nor U9524 (N_9524,N_9289,N_9409);
nor U9525 (N_9525,N_9339,N_9358);
xor U9526 (N_9526,N_9293,N_9350);
and U9527 (N_9527,N_9415,N_9339);
or U9528 (N_9528,N_9338,N_9331);
nand U9529 (N_9529,N_9379,N_9410);
xnor U9530 (N_9530,N_9412,N_9420);
nand U9531 (N_9531,N_9365,N_9325);
xor U9532 (N_9532,N_9309,N_9340);
or U9533 (N_9533,N_9405,N_9386);
nand U9534 (N_9534,N_9371,N_9406);
and U9535 (N_9535,N_9333,N_9350);
and U9536 (N_9536,N_9287,N_9347);
and U9537 (N_9537,N_9397,N_9387);
nor U9538 (N_9538,N_9378,N_9303);
or U9539 (N_9539,N_9403,N_9293);
or U9540 (N_9540,N_9385,N_9313);
and U9541 (N_9541,N_9436,N_9349);
nor U9542 (N_9542,N_9358,N_9294);
nor U9543 (N_9543,N_9346,N_9305);
nor U9544 (N_9544,N_9392,N_9287);
nor U9545 (N_9545,N_9287,N_9326);
nand U9546 (N_9546,N_9394,N_9294);
nand U9547 (N_9547,N_9382,N_9419);
nand U9548 (N_9548,N_9326,N_9354);
xor U9549 (N_9549,N_9283,N_9315);
and U9550 (N_9550,N_9349,N_9409);
nand U9551 (N_9551,N_9365,N_9345);
nor U9552 (N_9552,N_9399,N_9397);
or U9553 (N_9553,N_9384,N_9370);
xor U9554 (N_9554,N_9422,N_9328);
and U9555 (N_9555,N_9387,N_9316);
and U9556 (N_9556,N_9421,N_9299);
nand U9557 (N_9557,N_9330,N_9300);
nand U9558 (N_9558,N_9342,N_9402);
or U9559 (N_9559,N_9294,N_9335);
nor U9560 (N_9560,N_9427,N_9343);
or U9561 (N_9561,N_9395,N_9331);
nand U9562 (N_9562,N_9376,N_9297);
nand U9563 (N_9563,N_9380,N_9364);
nand U9564 (N_9564,N_9309,N_9372);
nand U9565 (N_9565,N_9289,N_9379);
and U9566 (N_9566,N_9411,N_9326);
nor U9567 (N_9567,N_9400,N_9394);
xor U9568 (N_9568,N_9285,N_9431);
nand U9569 (N_9569,N_9401,N_9285);
and U9570 (N_9570,N_9396,N_9382);
xnor U9571 (N_9571,N_9394,N_9406);
nor U9572 (N_9572,N_9418,N_9349);
and U9573 (N_9573,N_9283,N_9428);
xor U9574 (N_9574,N_9298,N_9347);
nor U9575 (N_9575,N_9377,N_9289);
nand U9576 (N_9576,N_9283,N_9423);
and U9577 (N_9577,N_9344,N_9407);
xnor U9578 (N_9578,N_9377,N_9317);
xnor U9579 (N_9579,N_9318,N_9424);
and U9580 (N_9580,N_9357,N_9312);
and U9581 (N_9581,N_9323,N_9313);
xnor U9582 (N_9582,N_9396,N_9392);
and U9583 (N_9583,N_9357,N_9406);
and U9584 (N_9584,N_9427,N_9303);
nor U9585 (N_9585,N_9299,N_9373);
and U9586 (N_9586,N_9331,N_9293);
nor U9587 (N_9587,N_9331,N_9354);
and U9588 (N_9588,N_9421,N_9286);
nand U9589 (N_9589,N_9345,N_9406);
and U9590 (N_9590,N_9366,N_9420);
nand U9591 (N_9591,N_9299,N_9360);
and U9592 (N_9592,N_9401,N_9319);
and U9593 (N_9593,N_9385,N_9364);
xnor U9594 (N_9594,N_9347,N_9330);
and U9595 (N_9595,N_9372,N_9423);
nand U9596 (N_9596,N_9292,N_9394);
nor U9597 (N_9597,N_9319,N_9304);
xor U9598 (N_9598,N_9399,N_9305);
or U9599 (N_9599,N_9375,N_9333);
nand U9600 (N_9600,N_9501,N_9553);
nand U9601 (N_9601,N_9567,N_9493);
nor U9602 (N_9602,N_9488,N_9500);
nor U9603 (N_9603,N_9471,N_9504);
nand U9604 (N_9604,N_9562,N_9495);
and U9605 (N_9605,N_9584,N_9579);
nor U9606 (N_9606,N_9558,N_9590);
or U9607 (N_9607,N_9552,N_9492);
nand U9608 (N_9608,N_9587,N_9597);
nor U9609 (N_9609,N_9469,N_9539);
nor U9610 (N_9610,N_9536,N_9525);
or U9611 (N_9611,N_9476,N_9441);
xor U9612 (N_9612,N_9545,N_9447);
nand U9613 (N_9613,N_9559,N_9454);
and U9614 (N_9614,N_9581,N_9522);
nand U9615 (N_9615,N_9474,N_9575);
and U9616 (N_9616,N_9440,N_9513);
or U9617 (N_9617,N_9464,N_9445);
xor U9618 (N_9618,N_9534,N_9556);
nand U9619 (N_9619,N_9551,N_9446);
nor U9620 (N_9620,N_9570,N_9475);
xnor U9621 (N_9621,N_9451,N_9453);
or U9622 (N_9622,N_9598,N_9472);
nand U9623 (N_9623,N_9569,N_9494);
nand U9624 (N_9624,N_9489,N_9596);
nand U9625 (N_9625,N_9457,N_9482);
and U9626 (N_9626,N_9555,N_9554);
nand U9627 (N_9627,N_9468,N_9563);
nand U9628 (N_9628,N_9467,N_9508);
xnor U9629 (N_9629,N_9546,N_9487);
and U9630 (N_9630,N_9455,N_9531);
and U9631 (N_9631,N_9444,N_9568);
xnor U9632 (N_9632,N_9524,N_9519);
nor U9633 (N_9633,N_9532,N_9517);
nand U9634 (N_9634,N_9586,N_9547);
xnor U9635 (N_9635,N_9459,N_9561);
or U9636 (N_9636,N_9502,N_9450);
nand U9637 (N_9637,N_9583,N_9460);
nand U9638 (N_9638,N_9473,N_9564);
nor U9639 (N_9639,N_9542,N_9548);
and U9640 (N_9640,N_9511,N_9509);
nand U9641 (N_9641,N_9479,N_9588);
nand U9642 (N_9642,N_9518,N_9505);
nand U9643 (N_9643,N_9520,N_9490);
and U9644 (N_9644,N_9507,N_9449);
or U9645 (N_9645,N_9480,N_9484);
and U9646 (N_9646,N_9594,N_9571);
nor U9647 (N_9647,N_9595,N_9550);
nand U9648 (N_9648,N_9442,N_9544);
xnor U9649 (N_9649,N_9529,N_9582);
xor U9650 (N_9650,N_9535,N_9443);
and U9651 (N_9651,N_9463,N_9491);
or U9652 (N_9652,N_9541,N_9452);
nor U9653 (N_9653,N_9486,N_9528);
and U9654 (N_9654,N_9576,N_9593);
or U9655 (N_9655,N_9573,N_9506);
nor U9656 (N_9656,N_9572,N_9512);
nand U9657 (N_9657,N_9585,N_9574);
and U9658 (N_9658,N_9448,N_9516);
xor U9659 (N_9659,N_9527,N_9523);
or U9660 (N_9660,N_9560,N_9514);
or U9661 (N_9661,N_9483,N_9510);
and U9662 (N_9662,N_9578,N_9466);
nor U9663 (N_9663,N_9496,N_9521);
and U9664 (N_9664,N_9470,N_9589);
xor U9665 (N_9665,N_9537,N_9456);
xor U9666 (N_9666,N_9498,N_9577);
or U9667 (N_9667,N_9538,N_9461);
or U9668 (N_9668,N_9526,N_9515);
nand U9669 (N_9669,N_9462,N_9580);
and U9670 (N_9670,N_9543,N_9477);
nor U9671 (N_9671,N_9478,N_9549);
xnor U9672 (N_9672,N_9565,N_9503);
xnor U9673 (N_9673,N_9497,N_9458);
or U9674 (N_9674,N_9481,N_9499);
xnor U9675 (N_9675,N_9591,N_9592);
nand U9676 (N_9676,N_9540,N_9465);
nor U9677 (N_9677,N_9557,N_9485);
nor U9678 (N_9678,N_9530,N_9533);
xnor U9679 (N_9679,N_9599,N_9566);
nor U9680 (N_9680,N_9446,N_9482);
xnor U9681 (N_9681,N_9511,N_9462);
xor U9682 (N_9682,N_9535,N_9451);
or U9683 (N_9683,N_9468,N_9519);
xnor U9684 (N_9684,N_9542,N_9572);
xor U9685 (N_9685,N_9460,N_9463);
nand U9686 (N_9686,N_9568,N_9466);
and U9687 (N_9687,N_9479,N_9481);
nor U9688 (N_9688,N_9479,N_9502);
or U9689 (N_9689,N_9487,N_9483);
nor U9690 (N_9690,N_9556,N_9537);
nand U9691 (N_9691,N_9489,N_9471);
nor U9692 (N_9692,N_9568,N_9478);
or U9693 (N_9693,N_9465,N_9591);
or U9694 (N_9694,N_9453,N_9537);
nor U9695 (N_9695,N_9539,N_9491);
and U9696 (N_9696,N_9502,N_9572);
nand U9697 (N_9697,N_9596,N_9459);
nor U9698 (N_9698,N_9588,N_9540);
or U9699 (N_9699,N_9598,N_9559);
nor U9700 (N_9700,N_9479,N_9549);
nor U9701 (N_9701,N_9524,N_9532);
or U9702 (N_9702,N_9440,N_9586);
nand U9703 (N_9703,N_9588,N_9463);
xnor U9704 (N_9704,N_9519,N_9457);
or U9705 (N_9705,N_9599,N_9519);
nor U9706 (N_9706,N_9567,N_9464);
xnor U9707 (N_9707,N_9529,N_9533);
xnor U9708 (N_9708,N_9443,N_9562);
and U9709 (N_9709,N_9482,N_9460);
xnor U9710 (N_9710,N_9471,N_9544);
or U9711 (N_9711,N_9564,N_9525);
xor U9712 (N_9712,N_9581,N_9540);
nand U9713 (N_9713,N_9493,N_9499);
nand U9714 (N_9714,N_9470,N_9510);
and U9715 (N_9715,N_9532,N_9472);
or U9716 (N_9716,N_9475,N_9531);
nor U9717 (N_9717,N_9496,N_9582);
xnor U9718 (N_9718,N_9466,N_9443);
nor U9719 (N_9719,N_9577,N_9562);
and U9720 (N_9720,N_9598,N_9550);
nor U9721 (N_9721,N_9556,N_9514);
nand U9722 (N_9722,N_9564,N_9508);
and U9723 (N_9723,N_9472,N_9490);
nand U9724 (N_9724,N_9582,N_9544);
nor U9725 (N_9725,N_9508,N_9553);
or U9726 (N_9726,N_9540,N_9534);
xnor U9727 (N_9727,N_9576,N_9506);
and U9728 (N_9728,N_9490,N_9446);
nor U9729 (N_9729,N_9505,N_9493);
nand U9730 (N_9730,N_9529,N_9544);
nor U9731 (N_9731,N_9508,N_9456);
nor U9732 (N_9732,N_9581,N_9523);
or U9733 (N_9733,N_9466,N_9505);
xor U9734 (N_9734,N_9485,N_9596);
nand U9735 (N_9735,N_9462,N_9573);
nor U9736 (N_9736,N_9534,N_9558);
xor U9737 (N_9737,N_9490,N_9535);
or U9738 (N_9738,N_9591,N_9453);
nor U9739 (N_9739,N_9515,N_9582);
and U9740 (N_9740,N_9550,N_9450);
nor U9741 (N_9741,N_9584,N_9568);
nand U9742 (N_9742,N_9548,N_9519);
xor U9743 (N_9743,N_9470,N_9463);
and U9744 (N_9744,N_9503,N_9542);
nand U9745 (N_9745,N_9494,N_9559);
or U9746 (N_9746,N_9540,N_9500);
or U9747 (N_9747,N_9502,N_9512);
and U9748 (N_9748,N_9522,N_9583);
nor U9749 (N_9749,N_9479,N_9517);
and U9750 (N_9750,N_9503,N_9576);
nand U9751 (N_9751,N_9596,N_9478);
or U9752 (N_9752,N_9471,N_9538);
or U9753 (N_9753,N_9595,N_9503);
xnor U9754 (N_9754,N_9497,N_9448);
nand U9755 (N_9755,N_9518,N_9508);
nor U9756 (N_9756,N_9443,N_9459);
nand U9757 (N_9757,N_9569,N_9518);
nand U9758 (N_9758,N_9460,N_9445);
nor U9759 (N_9759,N_9488,N_9459);
xnor U9760 (N_9760,N_9662,N_9674);
nor U9761 (N_9761,N_9634,N_9679);
nand U9762 (N_9762,N_9652,N_9712);
xnor U9763 (N_9763,N_9715,N_9628);
nand U9764 (N_9764,N_9687,N_9707);
or U9765 (N_9765,N_9758,N_9617);
nand U9766 (N_9766,N_9602,N_9744);
and U9767 (N_9767,N_9632,N_9751);
nor U9768 (N_9768,N_9667,N_9635);
xor U9769 (N_9769,N_9742,N_9629);
nand U9770 (N_9770,N_9727,N_9619);
xnor U9771 (N_9771,N_9620,N_9701);
nand U9772 (N_9772,N_9604,N_9731);
nand U9773 (N_9773,N_9650,N_9735);
and U9774 (N_9774,N_9605,N_9697);
or U9775 (N_9775,N_9637,N_9677);
nor U9776 (N_9776,N_9738,N_9753);
nor U9777 (N_9777,N_9626,N_9621);
or U9778 (N_9778,N_9639,N_9622);
or U9779 (N_9779,N_9666,N_9683);
nand U9780 (N_9780,N_9725,N_9651);
xnor U9781 (N_9781,N_9729,N_9644);
nor U9782 (N_9782,N_9714,N_9733);
xor U9783 (N_9783,N_9685,N_9702);
nand U9784 (N_9784,N_9695,N_9710);
and U9785 (N_9785,N_9638,N_9670);
and U9786 (N_9786,N_9706,N_9700);
nor U9787 (N_9787,N_9759,N_9606);
xnor U9788 (N_9788,N_9703,N_9681);
and U9789 (N_9789,N_9609,N_9636);
nand U9790 (N_9790,N_9719,N_9658);
nor U9791 (N_9791,N_9705,N_9752);
nand U9792 (N_9792,N_9743,N_9640);
nand U9793 (N_9793,N_9699,N_9633);
xor U9794 (N_9794,N_9680,N_9717);
nor U9795 (N_9795,N_9721,N_9641);
nor U9796 (N_9796,N_9646,N_9716);
nand U9797 (N_9797,N_9686,N_9739);
xor U9798 (N_9798,N_9655,N_9740);
or U9799 (N_9799,N_9718,N_9600);
xnor U9800 (N_9800,N_9745,N_9724);
nor U9801 (N_9801,N_9648,N_9664);
or U9802 (N_9802,N_9656,N_9671);
xor U9803 (N_9803,N_9746,N_9696);
nand U9804 (N_9804,N_9660,N_9693);
nand U9805 (N_9805,N_9627,N_9623);
xnor U9806 (N_9806,N_9665,N_9625);
xnor U9807 (N_9807,N_9726,N_9708);
or U9808 (N_9808,N_9613,N_9737);
and U9809 (N_9809,N_9704,N_9654);
nand U9810 (N_9810,N_9691,N_9631);
xor U9811 (N_9811,N_9747,N_9614);
xnor U9812 (N_9812,N_9748,N_9754);
or U9813 (N_9813,N_9657,N_9736);
and U9814 (N_9814,N_9607,N_9653);
or U9815 (N_9815,N_9675,N_9615);
nor U9816 (N_9816,N_9612,N_9678);
or U9817 (N_9817,N_9692,N_9611);
xnor U9818 (N_9818,N_9741,N_9730);
xnor U9819 (N_9819,N_9661,N_9723);
xor U9820 (N_9820,N_9734,N_9676);
or U9821 (N_9821,N_9659,N_9682);
and U9822 (N_9822,N_9601,N_9690);
xor U9823 (N_9823,N_9728,N_9663);
xnor U9824 (N_9824,N_9750,N_9669);
or U9825 (N_9825,N_9668,N_9732);
nor U9826 (N_9826,N_9608,N_9757);
or U9827 (N_9827,N_9603,N_9722);
nor U9828 (N_9828,N_9711,N_9610);
xor U9829 (N_9829,N_9616,N_9755);
nor U9830 (N_9830,N_9645,N_9688);
or U9831 (N_9831,N_9720,N_9749);
xnor U9832 (N_9832,N_9698,N_9684);
or U9833 (N_9833,N_9673,N_9647);
xnor U9834 (N_9834,N_9624,N_9672);
nand U9835 (N_9835,N_9713,N_9756);
and U9836 (N_9836,N_9618,N_9642);
xnor U9837 (N_9837,N_9709,N_9630);
or U9838 (N_9838,N_9649,N_9643);
nor U9839 (N_9839,N_9689,N_9694);
nor U9840 (N_9840,N_9745,N_9719);
or U9841 (N_9841,N_9710,N_9664);
nand U9842 (N_9842,N_9701,N_9673);
or U9843 (N_9843,N_9608,N_9633);
nor U9844 (N_9844,N_9684,N_9625);
or U9845 (N_9845,N_9721,N_9620);
nand U9846 (N_9846,N_9652,N_9666);
or U9847 (N_9847,N_9686,N_9624);
and U9848 (N_9848,N_9759,N_9664);
or U9849 (N_9849,N_9737,N_9726);
xnor U9850 (N_9850,N_9659,N_9697);
and U9851 (N_9851,N_9714,N_9611);
nor U9852 (N_9852,N_9667,N_9738);
xor U9853 (N_9853,N_9640,N_9688);
xnor U9854 (N_9854,N_9602,N_9696);
nor U9855 (N_9855,N_9726,N_9740);
nand U9856 (N_9856,N_9713,N_9635);
or U9857 (N_9857,N_9695,N_9650);
or U9858 (N_9858,N_9729,N_9751);
nor U9859 (N_9859,N_9743,N_9632);
or U9860 (N_9860,N_9729,N_9652);
and U9861 (N_9861,N_9616,N_9673);
and U9862 (N_9862,N_9714,N_9740);
nor U9863 (N_9863,N_9709,N_9670);
or U9864 (N_9864,N_9608,N_9696);
or U9865 (N_9865,N_9609,N_9742);
nand U9866 (N_9866,N_9643,N_9624);
nor U9867 (N_9867,N_9601,N_9712);
nand U9868 (N_9868,N_9612,N_9727);
nand U9869 (N_9869,N_9691,N_9715);
and U9870 (N_9870,N_9619,N_9649);
or U9871 (N_9871,N_9695,N_9609);
xnor U9872 (N_9872,N_9743,N_9665);
nor U9873 (N_9873,N_9650,N_9655);
xor U9874 (N_9874,N_9691,N_9644);
and U9875 (N_9875,N_9647,N_9630);
or U9876 (N_9876,N_9619,N_9758);
or U9877 (N_9877,N_9643,N_9687);
and U9878 (N_9878,N_9718,N_9728);
nand U9879 (N_9879,N_9725,N_9627);
or U9880 (N_9880,N_9672,N_9731);
and U9881 (N_9881,N_9601,N_9745);
xor U9882 (N_9882,N_9702,N_9747);
nor U9883 (N_9883,N_9652,N_9637);
nor U9884 (N_9884,N_9738,N_9602);
nor U9885 (N_9885,N_9609,N_9669);
nor U9886 (N_9886,N_9667,N_9606);
or U9887 (N_9887,N_9674,N_9727);
nor U9888 (N_9888,N_9755,N_9725);
nand U9889 (N_9889,N_9755,N_9735);
and U9890 (N_9890,N_9672,N_9630);
nand U9891 (N_9891,N_9617,N_9612);
or U9892 (N_9892,N_9738,N_9682);
xor U9893 (N_9893,N_9714,N_9607);
nor U9894 (N_9894,N_9653,N_9712);
nor U9895 (N_9895,N_9735,N_9646);
or U9896 (N_9896,N_9630,N_9733);
xnor U9897 (N_9897,N_9638,N_9652);
and U9898 (N_9898,N_9681,N_9673);
and U9899 (N_9899,N_9752,N_9681);
or U9900 (N_9900,N_9648,N_9627);
xnor U9901 (N_9901,N_9672,N_9724);
xnor U9902 (N_9902,N_9602,N_9673);
nand U9903 (N_9903,N_9738,N_9606);
and U9904 (N_9904,N_9725,N_9692);
nor U9905 (N_9905,N_9723,N_9755);
nand U9906 (N_9906,N_9715,N_9637);
nand U9907 (N_9907,N_9754,N_9709);
and U9908 (N_9908,N_9744,N_9662);
nor U9909 (N_9909,N_9652,N_9631);
or U9910 (N_9910,N_9694,N_9700);
or U9911 (N_9911,N_9708,N_9673);
and U9912 (N_9912,N_9752,N_9755);
xor U9913 (N_9913,N_9611,N_9691);
or U9914 (N_9914,N_9652,N_9726);
nand U9915 (N_9915,N_9709,N_9753);
or U9916 (N_9916,N_9723,N_9676);
nor U9917 (N_9917,N_9730,N_9664);
xor U9918 (N_9918,N_9609,N_9727);
or U9919 (N_9919,N_9705,N_9732);
xnor U9920 (N_9920,N_9918,N_9816);
nor U9921 (N_9921,N_9872,N_9912);
and U9922 (N_9922,N_9890,N_9800);
or U9923 (N_9923,N_9852,N_9915);
xnor U9924 (N_9924,N_9914,N_9897);
or U9925 (N_9925,N_9821,N_9831);
and U9926 (N_9926,N_9889,N_9873);
nor U9927 (N_9927,N_9868,N_9902);
nand U9928 (N_9928,N_9845,N_9882);
and U9929 (N_9929,N_9847,N_9789);
nand U9930 (N_9930,N_9824,N_9878);
nor U9931 (N_9931,N_9913,N_9894);
nor U9932 (N_9932,N_9783,N_9883);
or U9933 (N_9933,N_9782,N_9766);
and U9934 (N_9934,N_9811,N_9874);
or U9935 (N_9935,N_9919,N_9858);
xnor U9936 (N_9936,N_9765,N_9813);
or U9937 (N_9937,N_9784,N_9860);
or U9938 (N_9938,N_9832,N_9899);
nor U9939 (N_9939,N_9837,N_9909);
and U9940 (N_9940,N_9888,N_9817);
nor U9941 (N_9941,N_9795,N_9844);
and U9942 (N_9942,N_9903,N_9807);
xnor U9943 (N_9943,N_9814,N_9778);
or U9944 (N_9944,N_9825,N_9773);
xor U9945 (N_9945,N_9900,N_9810);
or U9946 (N_9946,N_9850,N_9863);
xor U9947 (N_9947,N_9822,N_9891);
nor U9948 (N_9948,N_9791,N_9818);
or U9949 (N_9949,N_9774,N_9801);
and U9950 (N_9950,N_9771,N_9796);
xnor U9951 (N_9951,N_9809,N_9916);
nand U9952 (N_9952,N_9797,N_9854);
or U9953 (N_9953,N_9827,N_9780);
nand U9954 (N_9954,N_9790,N_9805);
nor U9955 (N_9955,N_9871,N_9779);
and U9956 (N_9956,N_9861,N_9768);
xor U9957 (N_9957,N_9866,N_9901);
nor U9958 (N_9958,N_9880,N_9804);
xor U9959 (N_9959,N_9893,N_9851);
and U9960 (N_9960,N_9876,N_9906);
nor U9961 (N_9961,N_9911,N_9806);
xor U9962 (N_9962,N_9907,N_9846);
and U9963 (N_9963,N_9828,N_9910);
nand U9964 (N_9964,N_9764,N_9877);
and U9965 (N_9965,N_9802,N_9879);
and U9966 (N_9966,N_9829,N_9830);
xor U9967 (N_9967,N_9867,N_9781);
and U9968 (N_9968,N_9862,N_9785);
xnor U9969 (N_9969,N_9770,N_9808);
or U9970 (N_9970,N_9763,N_9823);
or U9971 (N_9971,N_9792,N_9870);
or U9972 (N_9972,N_9865,N_9857);
or U9973 (N_9973,N_9885,N_9776);
xor U9974 (N_9974,N_9761,N_9836);
xnor U9975 (N_9975,N_9833,N_9820);
xnor U9976 (N_9976,N_9856,N_9905);
nor U9977 (N_9977,N_9769,N_9819);
nand U9978 (N_9978,N_9840,N_9812);
or U9979 (N_9979,N_9841,N_9762);
xnor U9980 (N_9980,N_9815,N_9760);
nor U9981 (N_9981,N_9859,N_9896);
and U9982 (N_9982,N_9777,N_9849);
and U9983 (N_9983,N_9798,N_9898);
xor U9984 (N_9984,N_9842,N_9881);
and U9985 (N_9985,N_9786,N_9917);
nand U9986 (N_9986,N_9835,N_9875);
xor U9987 (N_9987,N_9794,N_9767);
and U9988 (N_9988,N_9853,N_9788);
xor U9989 (N_9989,N_9826,N_9787);
or U9990 (N_9990,N_9838,N_9904);
nand U9991 (N_9991,N_9887,N_9799);
nand U9992 (N_9992,N_9869,N_9834);
or U9993 (N_9993,N_9772,N_9895);
xor U9994 (N_9994,N_9839,N_9864);
nor U9995 (N_9995,N_9848,N_9843);
nor U9996 (N_9996,N_9793,N_9884);
nand U9997 (N_9997,N_9886,N_9855);
and U9998 (N_9998,N_9908,N_9803);
xor U9999 (N_9999,N_9892,N_9775);
and U10000 (N_10000,N_9831,N_9863);
xor U10001 (N_10001,N_9847,N_9783);
and U10002 (N_10002,N_9806,N_9764);
nand U10003 (N_10003,N_9906,N_9854);
and U10004 (N_10004,N_9814,N_9827);
or U10005 (N_10005,N_9849,N_9800);
and U10006 (N_10006,N_9773,N_9847);
nor U10007 (N_10007,N_9768,N_9785);
xnor U10008 (N_10008,N_9886,N_9919);
nand U10009 (N_10009,N_9904,N_9889);
and U10010 (N_10010,N_9900,N_9771);
nor U10011 (N_10011,N_9915,N_9878);
and U10012 (N_10012,N_9844,N_9787);
and U10013 (N_10013,N_9805,N_9836);
or U10014 (N_10014,N_9760,N_9809);
nor U10015 (N_10015,N_9854,N_9919);
or U10016 (N_10016,N_9880,N_9908);
nor U10017 (N_10017,N_9775,N_9868);
and U10018 (N_10018,N_9879,N_9866);
and U10019 (N_10019,N_9867,N_9875);
and U10020 (N_10020,N_9827,N_9826);
nand U10021 (N_10021,N_9787,N_9859);
xnor U10022 (N_10022,N_9782,N_9878);
or U10023 (N_10023,N_9855,N_9763);
nand U10024 (N_10024,N_9815,N_9884);
nand U10025 (N_10025,N_9803,N_9880);
nand U10026 (N_10026,N_9827,N_9864);
nor U10027 (N_10027,N_9871,N_9864);
nor U10028 (N_10028,N_9897,N_9764);
xnor U10029 (N_10029,N_9786,N_9902);
nor U10030 (N_10030,N_9903,N_9910);
nand U10031 (N_10031,N_9787,N_9815);
nor U10032 (N_10032,N_9852,N_9864);
xor U10033 (N_10033,N_9785,N_9830);
or U10034 (N_10034,N_9905,N_9891);
xor U10035 (N_10035,N_9888,N_9768);
nand U10036 (N_10036,N_9815,N_9842);
nand U10037 (N_10037,N_9877,N_9844);
and U10038 (N_10038,N_9845,N_9771);
and U10039 (N_10039,N_9796,N_9852);
and U10040 (N_10040,N_9883,N_9797);
xor U10041 (N_10041,N_9767,N_9865);
or U10042 (N_10042,N_9862,N_9834);
nor U10043 (N_10043,N_9914,N_9873);
and U10044 (N_10044,N_9897,N_9900);
nand U10045 (N_10045,N_9822,N_9771);
xnor U10046 (N_10046,N_9796,N_9817);
or U10047 (N_10047,N_9899,N_9790);
or U10048 (N_10048,N_9864,N_9906);
nor U10049 (N_10049,N_9877,N_9880);
nand U10050 (N_10050,N_9800,N_9766);
or U10051 (N_10051,N_9861,N_9801);
or U10052 (N_10052,N_9814,N_9831);
nor U10053 (N_10053,N_9807,N_9855);
or U10054 (N_10054,N_9890,N_9831);
nand U10055 (N_10055,N_9823,N_9888);
and U10056 (N_10056,N_9766,N_9778);
or U10057 (N_10057,N_9845,N_9875);
nand U10058 (N_10058,N_9811,N_9895);
nor U10059 (N_10059,N_9912,N_9881);
xnor U10060 (N_10060,N_9899,N_9866);
or U10061 (N_10061,N_9911,N_9769);
nor U10062 (N_10062,N_9882,N_9838);
xnor U10063 (N_10063,N_9845,N_9910);
or U10064 (N_10064,N_9763,N_9905);
nand U10065 (N_10065,N_9824,N_9779);
and U10066 (N_10066,N_9787,N_9909);
nor U10067 (N_10067,N_9765,N_9781);
xor U10068 (N_10068,N_9793,N_9876);
nand U10069 (N_10069,N_9762,N_9866);
nand U10070 (N_10070,N_9857,N_9779);
xor U10071 (N_10071,N_9780,N_9906);
nor U10072 (N_10072,N_9764,N_9771);
nand U10073 (N_10073,N_9860,N_9839);
and U10074 (N_10074,N_9826,N_9813);
nand U10075 (N_10075,N_9760,N_9841);
nor U10076 (N_10076,N_9841,N_9812);
nor U10077 (N_10077,N_9855,N_9799);
xnor U10078 (N_10078,N_9864,N_9819);
xnor U10079 (N_10079,N_9797,N_9861);
and U10080 (N_10080,N_9931,N_9987);
xor U10081 (N_10081,N_9975,N_10030);
and U10082 (N_10082,N_10040,N_10064);
xor U10083 (N_10083,N_9980,N_9958);
xnor U10084 (N_10084,N_10016,N_9969);
xor U10085 (N_10085,N_9936,N_10068);
nor U10086 (N_10086,N_10004,N_10054);
xnor U10087 (N_10087,N_9935,N_10023);
or U10088 (N_10088,N_9997,N_10017);
xnor U10089 (N_10089,N_10007,N_10024);
nor U10090 (N_10090,N_9930,N_9921);
nand U10091 (N_10091,N_10034,N_9998);
nand U10092 (N_10092,N_9920,N_9965);
and U10093 (N_10093,N_9991,N_10069);
xnor U10094 (N_10094,N_9960,N_9947);
or U10095 (N_10095,N_9977,N_9957);
nand U10096 (N_10096,N_9962,N_10013);
nor U10097 (N_10097,N_10078,N_9959);
nor U10098 (N_10098,N_9927,N_10020);
nor U10099 (N_10099,N_10047,N_10031);
nor U10100 (N_10100,N_9984,N_10070);
nor U10101 (N_10101,N_9976,N_10073);
or U10102 (N_10102,N_10035,N_9968);
and U10103 (N_10103,N_10027,N_9923);
xor U10104 (N_10104,N_9966,N_9963);
nand U10105 (N_10105,N_9941,N_10014);
nand U10106 (N_10106,N_9988,N_9986);
or U10107 (N_10107,N_9961,N_9993);
xnor U10108 (N_10108,N_10067,N_10041);
nand U10109 (N_10109,N_10057,N_9952);
xnor U10110 (N_10110,N_10029,N_9933);
nand U10111 (N_10111,N_9937,N_10075);
nor U10112 (N_10112,N_10011,N_9999);
nor U10113 (N_10113,N_10008,N_9970);
nor U10114 (N_10114,N_9979,N_9955);
nor U10115 (N_10115,N_10046,N_10037);
xnor U10116 (N_10116,N_9942,N_9978);
xnor U10117 (N_10117,N_10026,N_10071);
and U10118 (N_10118,N_9950,N_9925);
or U10119 (N_10119,N_10056,N_10038);
nand U10120 (N_10120,N_9985,N_10025);
xor U10121 (N_10121,N_9945,N_10021);
nand U10122 (N_10122,N_9992,N_10033);
nor U10123 (N_10123,N_10063,N_10055);
and U10124 (N_10124,N_9949,N_9926);
or U10125 (N_10125,N_9971,N_10012);
xnor U10126 (N_10126,N_9964,N_10042);
and U10127 (N_10127,N_10060,N_9948);
nor U10128 (N_10128,N_9994,N_10077);
or U10129 (N_10129,N_10002,N_10052);
nor U10130 (N_10130,N_9946,N_10050);
nor U10131 (N_10131,N_10009,N_9944);
nand U10132 (N_10132,N_9938,N_10058);
xor U10133 (N_10133,N_10018,N_9953);
nand U10134 (N_10134,N_10015,N_10022);
and U10135 (N_10135,N_9932,N_9996);
or U10136 (N_10136,N_10053,N_9990);
nor U10137 (N_10137,N_10001,N_10049);
nand U10138 (N_10138,N_10076,N_9989);
nor U10139 (N_10139,N_10061,N_10074);
xor U10140 (N_10140,N_9940,N_9981);
and U10141 (N_10141,N_10079,N_9934);
nor U10142 (N_10142,N_10072,N_9995);
and U10143 (N_10143,N_10066,N_10032);
nor U10144 (N_10144,N_9939,N_9982);
xnor U10145 (N_10145,N_10044,N_9974);
nand U10146 (N_10146,N_10006,N_10051);
nor U10147 (N_10147,N_10045,N_9972);
xor U10148 (N_10148,N_10003,N_9983);
xnor U10149 (N_10149,N_9954,N_10000);
and U10150 (N_10150,N_9967,N_10019);
nand U10151 (N_10151,N_9922,N_9951);
nand U10152 (N_10152,N_10062,N_10010);
nand U10153 (N_10153,N_10036,N_10059);
nand U10154 (N_10154,N_10043,N_10065);
and U10155 (N_10155,N_9929,N_9928);
or U10156 (N_10156,N_9973,N_9943);
nand U10157 (N_10157,N_9924,N_9956);
xnor U10158 (N_10158,N_10005,N_10039);
nor U10159 (N_10159,N_10028,N_10048);
xor U10160 (N_10160,N_10021,N_9927);
nor U10161 (N_10161,N_10017,N_10040);
and U10162 (N_10162,N_9976,N_10072);
xor U10163 (N_10163,N_10052,N_9954);
nand U10164 (N_10164,N_9983,N_10042);
nor U10165 (N_10165,N_10062,N_9983);
xnor U10166 (N_10166,N_10065,N_9961);
or U10167 (N_10167,N_9935,N_9969);
or U10168 (N_10168,N_9925,N_9972);
xor U10169 (N_10169,N_10060,N_10020);
nand U10170 (N_10170,N_10015,N_9921);
nor U10171 (N_10171,N_10044,N_10002);
and U10172 (N_10172,N_9992,N_10030);
nand U10173 (N_10173,N_9953,N_10076);
xor U10174 (N_10174,N_10055,N_10072);
and U10175 (N_10175,N_9970,N_9980);
or U10176 (N_10176,N_9953,N_9990);
xnor U10177 (N_10177,N_10035,N_9976);
nand U10178 (N_10178,N_9998,N_10066);
xor U10179 (N_10179,N_9923,N_10002);
and U10180 (N_10180,N_10017,N_9980);
xnor U10181 (N_10181,N_9964,N_9990);
or U10182 (N_10182,N_9925,N_10001);
nor U10183 (N_10183,N_9927,N_9935);
or U10184 (N_10184,N_10059,N_10050);
or U10185 (N_10185,N_9943,N_9989);
nor U10186 (N_10186,N_9972,N_10052);
and U10187 (N_10187,N_9926,N_10042);
nand U10188 (N_10188,N_9992,N_10032);
or U10189 (N_10189,N_10030,N_10057);
xnor U10190 (N_10190,N_10077,N_10062);
xnor U10191 (N_10191,N_10054,N_10079);
or U10192 (N_10192,N_10006,N_10033);
nor U10193 (N_10193,N_10028,N_10029);
and U10194 (N_10194,N_9922,N_9947);
and U10195 (N_10195,N_10007,N_10071);
or U10196 (N_10196,N_10044,N_9960);
or U10197 (N_10197,N_9995,N_10009);
xnor U10198 (N_10198,N_9966,N_9978);
nand U10199 (N_10199,N_9930,N_10039);
nand U10200 (N_10200,N_9953,N_10000);
nand U10201 (N_10201,N_9946,N_10012);
nor U10202 (N_10202,N_10012,N_9943);
xnor U10203 (N_10203,N_9939,N_10043);
or U10204 (N_10204,N_10071,N_9996);
and U10205 (N_10205,N_9940,N_10013);
and U10206 (N_10206,N_10077,N_9939);
and U10207 (N_10207,N_9925,N_9952);
or U10208 (N_10208,N_9936,N_9966);
nor U10209 (N_10209,N_9941,N_9983);
or U10210 (N_10210,N_9986,N_9991);
nor U10211 (N_10211,N_9942,N_10027);
or U10212 (N_10212,N_9941,N_9988);
xor U10213 (N_10213,N_9985,N_9937);
or U10214 (N_10214,N_9935,N_10049);
and U10215 (N_10215,N_10017,N_9928);
nor U10216 (N_10216,N_10000,N_9998);
nor U10217 (N_10217,N_9950,N_9951);
and U10218 (N_10218,N_10049,N_10075);
or U10219 (N_10219,N_10012,N_10064);
or U10220 (N_10220,N_9972,N_9980);
xnor U10221 (N_10221,N_10009,N_10022);
or U10222 (N_10222,N_9943,N_10067);
xor U10223 (N_10223,N_9993,N_9996);
nand U10224 (N_10224,N_9941,N_10072);
and U10225 (N_10225,N_10008,N_9980);
xnor U10226 (N_10226,N_10000,N_9920);
xnor U10227 (N_10227,N_9967,N_10068);
or U10228 (N_10228,N_10006,N_10053);
xor U10229 (N_10229,N_9979,N_10050);
or U10230 (N_10230,N_10062,N_10015);
or U10231 (N_10231,N_9925,N_10057);
nor U10232 (N_10232,N_9975,N_10028);
nand U10233 (N_10233,N_9941,N_10051);
xor U10234 (N_10234,N_9964,N_9948);
nand U10235 (N_10235,N_9948,N_10034);
xnor U10236 (N_10236,N_10075,N_9945);
nand U10237 (N_10237,N_9982,N_9943);
nand U10238 (N_10238,N_9950,N_10017);
nand U10239 (N_10239,N_10000,N_10033);
nor U10240 (N_10240,N_10171,N_10198);
nand U10241 (N_10241,N_10157,N_10153);
nor U10242 (N_10242,N_10233,N_10098);
and U10243 (N_10243,N_10146,N_10179);
and U10244 (N_10244,N_10236,N_10197);
nand U10245 (N_10245,N_10137,N_10087);
or U10246 (N_10246,N_10194,N_10191);
nand U10247 (N_10247,N_10130,N_10166);
nor U10248 (N_10248,N_10117,N_10207);
and U10249 (N_10249,N_10232,N_10185);
or U10250 (N_10250,N_10169,N_10100);
nand U10251 (N_10251,N_10135,N_10108);
nor U10252 (N_10252,N_10097,N_10156);
nor U10253 (N_10253,N_10205,N_10192);
and U10254 (N_10254,N_10145,N_10189);
xnor U10255 (N_10255,N_10096,N_10129);
xor U10256 (N_10256,N_10162,N_10213);
nand U10257 (N_10257,N_10190,N_10159);
and U10258 (N_10258,N_10126,N_10172);
xor U10259 (N_10259,N_10167,N_10085);
xor U10260 (N_10260,N_10106,N_10237);
or U10261 (N_10261,N_10092,N_10200);
nand U10262 (N_10262,N_10149,N_10143);
or U10263 (N_10263,N_10221,N_10230);
or U10264 (N_10264,N_10125,N_10140);
nor U10265 (N_10265,N_10134,N_10142);
nor U10266 (N_10266,N_10082,N_10229);
and U10267 (N_10267,N_10083,N_10219);
nor U10268 (N_10268,N_10091,N_10128);
and U10269 (N_10269,N_10196,N_10113);
nor U10270 (N_10270,N_10136,N_10155);
nor U10271 (N_10271,N_10115,N_10138);
nand U10272 (N_10272,N_10170,N_10188);
and U10273 (N_10273,N_10132,N_10195);
and U10274 (N_10274,N_10088,N_10084);
nor U10275 (N_10275,N_10187,N_10223);
or U10276 (N_10276,N_10206,N_10180);
nor U10277 (N_10277,N_10182,N_10114);
nor U10278 (N_10278,N_10220,N_10093);
xnor U10279 (N_10279,N_10154,N_10127);
nor U10280 (N_10280,N_10199,N_10238);
or U10281 (N_10281,N_10105,N_10204);
and U10282 (N_10282,N_10120,N_10203);
nand U10283 (N_10283,N_10109,N_10217);
and U10284 (N_10284,N_10133,N_10112);
xnor U10285 (N_10285,N_10175,N_10147);
nor U10286 (N_10286,N_10186,N_10151);
and U10287 (N_10287,N_10165,N_10222);
xnor U10288 (N_10288,N_10224,N_10193);
nor U10289 (N_10289,N_10144,N_10161);
xor U10290 (N_10290,N_10123,N_10176);
nand U10291 (N_10291,N_10212,N_10168);
or U10292 (N_10292,N_10226,N_10103);
xor U10293 (N_10293,N_10227,N_10184);
or U10294 (N_10294,N_10225,N_10231);
nor U10295 (N_10295,N_10181,N_10210);
nand U10296 (N_10296,N_10080,N_10102);
nand U10297 (N_10297,N_10090,N_10148);
nor U10298 (N_10298,N_10095,N_10104);
nand U10299 (N_10299,N_10174,N_10086);
xnor U10300 (N_10300,N_10234,N_10164);
xor U10301 (N_10301,N_10239,N_10183);
xnor U10302 (N_10302,N_10139,N_10089);
or U10303 (N_10303,N_10094,N_10216);
nor U10304 (N_10304,N_10118,N_10235);
xnor U10305 (N_10305,N_10150,N_10173);
nand U10306 (N_10306,N_10111,N_10228);
and U10307 (N_10307,N_10124,N_10131);
and U10308 (N_10308,N_10201,N_10208);
xor U10309 (N_10309,N_10152,N_10099);
nand U10310 (N_10310,N_10178,N_10214);
nor U10311 (N_10311,N_10119,N_10116);
and U10312 (N_10312,N_10121,N_10101);
and U10313 (N_10313,N_10218,N_10141);
xnor U10314 (N_10314,N_10211,N_10215);
or U10315 (N_10315,N_10177,N_10163);
and U10316 (N_10316,N_10107,N_10158);
nor U10317 (N_10317,N_10081,N_10110);
nand U10318 (N_10318,N_10209,N_10122);
nand U10319 (N_10319,N_10160,N_10202);
xnor U10320 (N_10320,N_10097,N_10212);
nand U10321 (N_10321,N_10158,N_10100);
or U10322 (N_10322,N_10108,N_10211);
xnor U10323 (N_10323,N_10145,N_10155);
and U10324 (N_10324,N_10167,N_10106);
xnor U10325 (N_10325,N_10182,N_10189);
xor U10326 (N_10326,N_10104,N_10172);
nand U10327 (N_10327,N_10220,N_10226);
and U10328 (N_10328,N_10182,N_10126);
xnor U10329 (N_10329,N_10097,N_10178);
xor U10330 (N_10330,N_10220,N_10230);
nand U10331 (N_10331,N_10136,N_10134);
nand U10332 (N_10332,N_10212,N_10230);
or U10333 (N_10333,N_10097,N_10191);
nand U10334 (N_10334,N_10111,N_10233);
or U10335 (N_10335,N_10159,N_10165);
xor U10336 (N_10336,N_10188,N_10202);
or U10337 (N_10337,N_10149,N_10165);
xnor U10338 (N_10338,N_10124,N_10227);
and U10339 (N_10339,N_10200,N_10191);
nor U10340 (N_10340,N_10142,N_10151);
xnor U10341 (N_10341,N_10098,N_10089);
xor U10342 (N_10342,N_10211,N_10146);
xnor U10343 (N_10343,N_10216,N_10233);
and U10344 (N_10344,N_10228,N_10139);
nand U10345 (N_10345,N_10134,N_10150);
nand U10346 (N_10346,N_10167,N_10226);
or U10347 (N_10347,N_10215,N_10178);
xnor U10348 (N_10348,N_10088,N_10217);
or U10349 (N_10349,N_10217,N_10126);
nand U10350 (N_10350,N_10130,N_10171);
xor U10351 (N_10351,N_10203,N_10183);
xnor U10352 (N_10352,N_10191,N_10107);
and U10353 (N_10353,N_10106,N_10152);
nand U10354 (N_10354,N_10122,N_10235);
xnor U10355 (N_10355,N_10099,N_10137);
and U10356 (N_10356,N_10151,N_10115);
nand U10357 (N_10357,N_10176,N_10100);
and U10358 (N_10358,N_10212,N_10174);
nor U10359 (N_10359,N_10130,N_10081);
nand U10360 (N_10360,N_10081,N_10224);
and U10361 (N_10361,N_10228,N_10211);
nand U10362 (N_10362,N_10213,N_10159);
nand U10363 (N_10363,N_10102,N_10163);
and U10364 (N_10364,N_10129,N_10127);
nand U10365 (N_10365,N_10178,N_10143);
or U10366 (N_10366,N_10104,N_10102);
nand U10367 (N_10367,N_10097,N_10190);
nor U10368 (N_10368,N_10109,N_10199);
nor U10369 (N_10369,N_10147,N_10206);
or U10370 (N_10370,N_10099,N_10138);
xnor U10371 (N_10371,N_10085,N_10207);
nand U10372 (N_10372,N_10128,N_10162);
nand U10373 (N_10373,N_10109,N_10135);
xnor U10374 (N_10374,N_10115,N_10125);
and U10375 (N_10375,N_10190,N_10226);
and U10376 (N_10376,N_10211,N_10142);
xnor U10377 (N_10377,N_10183,N_10090);
nand U10378 (N_10378,N_10139,N_10081);
xnor U10379 (N_10379,N_10118,N_10081);
nor U10380 (N_10380,N_10150,N_10101);
or U10381 (N_10381,N_10210,N_10140);
and U10382 (N_10382,N_10216,N_10138);
xor U10383 (N_10383,N_10104,N_10122);
and U10384 (N_10384,N_10174,N_10081);
or U10385 (N_10385,N_10142,N_10221);
or U10386 (N_10386,N_10135,N_10156);
xor U10387 (N_10387,N_10089,N_10135);
nor U10388 (N_10388,N_10112,N_10104);
nor U10389 (N_10389,N_10196,N_10101);
and U10390 (N_10390,N_10207,N_10210);
or U10391 (N_10391,N_10138,N_10112);
and U10392 (N_10392,N_10163,N_10186);
nand U10393 (N_10393,N_10217,N_10229);
and U10394 (N_10394,N_10090,N_10160);
and U10395 (N_10395,N_10128,N_10179);
xnor U10396 (N_10396,N_10230,N_10129);
or U10397 (N_10397,N_10166,N_10098);
nand U10398 (N_10398,N_10239,N_10199);
xnor U10399 (N_10399,N_10202,N_10093);
nand U10400 (N_10400,N_10385,N_10386);
and U10401 (N_10401,N_10318,N_10274);
nand U10402 (N_10402,N_10317,N_10316);
or U10403 (N_10403,N_10387,N_10283);
and U10404 (N_10404,N_10359,N_10258);
xor U10405 (N_10405,N_10332,N_10330);
nand U10406 (N_10406,N_10375,N_10260);
and U10407 (N_10407,N_10348,N_10281);
and U10408 (N_10408,N_10379,N_10391);
nor U10409 (N_10409,N_10290,N_10371);
nor U10410 (N_10410,N_10355,N_10397);
and U10411 (N_10411,N_10304,N_10322);
nor U10412 (N_10412,N_10395,N_10356);
nor U10413 (N_10413,N_10370,N_10364);
nor U10414 (N_10414,N_10392,N_10377);
nand U10415 (N_10415,N_10287,N_10279);
and U10416 (N_10416,N_10381,N_10362);
nand U10417 (N_10417,N_10338,N_10272);
nor U10418 (N_10418,N_10372,N_10259);
nor U10419 (N_10419,N_10329,N_10250);
xor U10420 (N_10420,N_10343,N_10366);
or U10421 (N_10421,N_10264,N_10323);
xor U10422 (N_10422,N_10378,N_10340);
or U10423 (N_10423,N_10383,N_10321);
or U10424 (N_10424,N_10257,N_10285);
nand U10425 (N_10425,N_10396,N_10265);
xor U10426 (N_10426,N_10350,N_10301);
nand U10427 (N_10427,N_10277,N_10252);
xnor U10428 (N_10428,N_10365,N_10312);
nor U10429 (N_10429,N_10334,N_10254);
xor U10430 (N_10430,N_10246,N_10289);
nand U10431 (N_10431,N_10314,N_10345);
or U10432 (N_10432,N_10311,N_10303);
nand U10433 (N_10433,N_10354,N_10327);
and U10434 (N_10434,N_10337,N_10399);
or U10435 (N_10435,N_10335,N_10315);
and U10436 (N_10436,N_10336,N_10331);
and U10437 (N_10437,N_10253,N_10302);
or U10438 (N_10438,N_10309,N_10273);
and U10439 (N_10439,N_10267,N_10294);
or U10440 (N_10440,N_10282,N_10384);
or U10441 (N_10441,N_10296,N_10393);
nor U10442 (N_10442,N_10278,N_10339);
nor U10443 (N_10443,N_10280,N_10240);
xnor U10444 (N_10444,N_10245,N_10389);
xnor U10445 (N_10445,N_10319,N_10374);
nor U10446 (N_10446,N_10244,N_10368);
nor U10447 (N_10447,N_10373,N_10341);
nor U10448 (N_10448,N_10293,N_10353);
and U10449 (N_10449,N_10310,N_10398);
xnor U10450 (N_10450,N_10358,N_10276);
xor U10451 (N_10451,N_10360,N_10266);
nor U10452 (N_10452,N_10307,N_10263);
or U10453 (N_10453,N_10363,N_10320);
nand U10454 (N_10454,N_10388,N_10361);
nand U10455 (N_10455,N_10268,N_10347);
xnor U10456 (N_10456,N_10313,N_10300);
nor U10457 (N_10457,N_10284,N_10270);
or U10458 (N_10458,N_10326,N_10308);
and U10459 (N_10459,N_10394,N_10261);
nand U10460 (N_10460,N_10346,N_10251);
xnor U10461 (N_10461,N_10298,N_10306);
and U10462 (N_10462,N_10269,N_10349);
xor U10463 (N_10463,N_10248,N_10380);
and U10464 (N_10464,N_10367,N_10369);
nor U10465 (N_10465,N_10292,N_10288);
nand U10466 (N_10466,N_10243,N_10275);
and U10467 (N_10467,N_10249,N_10262);
nor U10468 (N_10468,N_10351,N_10291);
or U10469 (N_10469,N_10342,N_10357);
xor U10470 (N_10470,N_10333,N_10241);
nor U10471 (N_10471,N_10295,N_10305);
and U10472 (N_10472,N_10376,N_10247);
and U10473 (N_10473,N_10328,N_10242);
nand U10474 (N_10474,N_10344,N_10324);
or U10475 (N_10475,N_10286,N_10299);
or U10476 (N_10476,N_10255,N_10390);
nand U10477 (N_10477,N_10382,N_10325);
nor U10478 (N_10478,N_10297,N_10256);
nand U10479 (N_10479,N_10271,N_10352);
or U10480 (N_10480,N_10393,N_10258);
nand U10481 (N_10481,N_10379,N_10271);
xnor U10482 (N_10482,N_10391,N_10253);
and U10483 (N_10483,N_10241,N_10321);
and U10484 (N_10484,N_10354,N_10250);
nand U10485 (N_10485,N_10322,N_10293);
nor U10486 (N_10486,N_10351,N_10283);
nand U10487 (N_10487,N_10251,N_10288);
nor U10488 (N_10488,N_10377,N_10261);
and U10489 (N_10489,N_10318,N_10383);
nand U10490 (N_10490,N_10366,N_10313);
and U10491 (N_10491,N_10392,N_10311);
nand U10492 (N_10492,N_10325,N_10288);
and U10493 (N_10493,N_10279,N_10362);
and U10494 (N_10494,N_10348,N_10296);
and U10495 (N_10495,N_10378,N_10360);
nor U10496 (N_10496,N_10368,N_10333);
nor U10497 (N_10497,N_10279,N_10316);
nor U10498 (N_10498,N_10268,N_10343);
nor U10499 (N_10499,N_10258,N_10363);
nor U10500 (N_10500,N_10394,N_10373);
xor U10501 (N_10501,N_10262,N_10361);
or U10502 (N_10502,N_10287,N_10241);
nand U10503 (N_10503,N_10267,N_10365);
nor U10504 (N_10504,N_10245,N_10352);
nand U10505 (N_10505,N_10351,N_10381);
or U10506 (N_10506,N_10313,N_10356);
and U10507 (N_10507,N_10395,N_10289);
and U10508 (N_10508,N_10344,N_10271);
xor U10509 (N_10509,N_10331,N_10342);
and U10510 (N_10510,N_10283,N_10240);
nand U10511 (N_10511,N_10316,N_10332);
nand U10512 (N_10512,N_10249,N_10339);
or U10513 (N_10513,N_10399,N_10240);
or U10514 (N_10514,N_10274,N_10388);
or U10515 (N_10515,N_10374,N_10389);
nor U10516 (N_10516,N_10372,N_10293);
xnor U10517 (N_10517,N_10332,N_10348);
and U10518 (N_10518,N_10321,N_10284);
xor U10519 (N_10519,N_10323,N_10337);
nor U10520 (N_10520,N_10262,N_10310);
nand U10521 (N_10521,N_10268,N_10379);
nor U10522 (N_10522,N_10344,N_10325);
or U10523 (N_10523,N_10329,N_10338);
nor U10524 (N_10524,N_10272,N_10381);
xnor U10525 (N_10525,N_10255,N_10359);
and U10526 (N_10526,N_10356,N_10287);
nand U10527 (N_10527,N_10349,N_10362);
nor U10528 (N_10528,N_10262,N_10392);
nand U10529 (N_10529,N_10304,N_10389);
nor U10530 (N_10530,N_10279,N_10246);
xnor U10531 (N_10531,N_10383,N_10300);
and U10532 (N_10532,N_10299,N_10329);
and U10533 (N_10533,N_10263,N_10332);
xnor U10534 (N_10534,N_10243,N_10297);
nand U10535 (N_10535,N_10280,N_10247);
and U10536 (N_10536,N_10330,N_10373);
nand U10537 (N_10537,N_10383,N_10361);
nand U10538 (N_10538,N_10363,N_10297);
and U10539 (N_10539,N_10326,N_10383);
and U10540 (N_10540,N_10244,N_10256);
nand U10541 (N_10541,N_10305,N_10314);
or U10542 (N_10542,N_10250,N_10240);
xor U10543 (N_10543,N_10349,N_10280);
nand U10544 (N_10544,N_10352,N_10242);
nor U10545 (N_10545,N_10261,N_10352);
or U10546 (N_10546,N_10394,N_10360);
nand U10547 (N_10547,N_10392,N_10382);
and U10548 (N_10548,N_10351,N_10378);
nor U10549 (N_10549,N_10274,N_10399);
or U10550 (N_10550,N_10395,N_10323);
nor U10551 (N_10551,N_10345,N_10258);
nand U10552 (N_10552,N_10324,N_10323);
and U10553 (N_10553,N_10341,N_10392);
xnor U10554 (N_10554,N_10289,N_10269);
xor U10555 (N_10555,N_10332,N_10318);
and U10556 (N_10556,N_10383,N_10376);
nand U10557 (N_10557,N_10303,N_10278);
nand U10558 (N_10558,N_10322,N_10362);
and U10559 (N_10559,N_10290,N_10291);
xnor U10560 (N_10560,N_10547,N_10507);
nor U10561 (N_10561,N_10541,N_10419);
and U10562 (N_10562,N_10484,N_10546);
and U10563 (N_10563,N_10526,N_10498);
nor U10564 (N_10564,N_10400,N_10515);
nor U10565 (N_10565,N_10417,N_10533);
nor U10566 (N_10566,N_10513,N_10475);
xor U10567 (N_10567,N_10540,N_10415);
and U10568 (N_10568,N_10481,N_10503);
or U10569 (N_10569,N_10413,N_10539);
nand U10570 (N_10570,N_10459,N_10402);
or U10571 (N_10571,N_10416,N_10428);
nor U10572 (N_10572,N_10509,N_10504);
or U10573 (N_10573,N_10544,N_10512);
or U10574 (N_10574,N_10514,N_10441);
xnor U10575 (N_10575,N_10496,N_10545);
and U10576 (N_10576,N_10494,N_10437);
or U10577 (N_10577,N_10427,N_10470);
and U10578 (N_10578,N_10421,N_10550);
nand U10579 (N_10579,N_10471,N_10432);
nand U10580 (N_10580,N_10534,N_10491);
and U10581 (N_10581,N_10442,N_10527);
xnor U10582 (N_10582,N_10450,N_10429);
or U10583 (N_10583,N_10476,N_10552);
and U10584 (N_10584,N_10436,N_10487);
nor U10585 (N_10585,N_10488,N_10521);
and U10586 (N_10586,N_10493,N_10492);
nand U10587 (N_10587,N_10465,N_10499);
and U10588 (N_10588,N_10501,N_10406);
xnor U10589 (N_10589,N_10511,N_10422);
xor U10590 (N_10590,N_10469,N_10449);
nor U10591 (N_10591,N_10500,N_10425);
and U10592 (N_10592,N_10472,N_10532);
and U10593 (N_10593,N_10559,N_10439);
and U10594 (N_10594,N_10423,N_10447);
and U10595 (N_10595,N_10489,N_10490);
xnor U10596 (N_10596,N_10495,N_10457);
nand U10597 (N_10597,N_10531,N_10418);
nand U10598 (N_10598,N_10536,N_10505);
nand U10599 (N_10599,N_10460,N_10463);
nand U10600 (N_10600,N_10497,N_10519);
or U10601 (N_10601,N_10410,N_10404);
and U10602 (N_10602,N_10440,N_10420);
and U10603 (N_10603,N_10530,N_10522);
and U10604 (N_10604,N_10480,N_10549);
nor U10605 (N_10605,N_10453,N_10434);
xnor U10606 (N_10606,N_10518,N_10537);
nand U10607 (N_10607,N_10485,N_10454);
nand U10608 (N_10608,N_10523,N_10548);
or U10609 (N_10609,N_10542,N_10478);
nor U10610 (N_10610,N_10426,N_10464);
xor U10611 (N_10611,N_10444,N_10466);
xnor U10612 (N_10612,N_10482,N_10448);
nand U10613 (N_10613,N_10520,N_10435);
nor U10614 (N_10614,N_10458,N_10555);
and U10615 (N_10615,N_10462,N_10433);
nor U10616 (N_10616,N_10477,N_10455);
or U10617 (N_10617,N_10405,N_10502);
nor U10618 (N_10618,N_10517,N_10486);
or U10619 (N_10619,N_10543,N_10557);
and U10620 (N_10620,N_10473,N_10529);
xor U10621 (N_10621,N_10452,N_10414);
nand U10622 (N_10622,N_10411,N_10467);
or U10623 (N_10623,N_10468,N_10409);
nand U10624 (N_10624,N_10424,N_10431);
xor U10625 (N_10625,N_10412,N_10524);
and U10626 (N_10626,N_10483,N_10528);
and U10627 (N_10627,N_10407,N_10451);
nand U10628 (N_10628,N_10551,N_10445);
and U10629 (N_10629,N_10558,N_10456);
nand U10630 (N_10630,N_10525,N_10446);
nand U10631 (N_10631,N_10408,N_10506);
nor U10632 (N_10632,N_10479,N_10516);
xor U10633 (N_10633,N_10556,N_10430);
and U10634 (N_10634,N_10538,N_10554);
xor U10635 (N_10635,N_10508,N_10438);
nand U10636 (N_10636,N_10553,N_10474);
nor U10637 (N_10637,N_10510,N_10443);
nor U10638 (N_10638,N_10403,N_10401);
and U10639 (N_10639,N_10535,N_10461);
and U10640 (N_10640,N_10473,N_10445);
nor U10641 (N_10641,N_10543,N_10485);
and U10642 (N_10642,N_10451,N_10458);
or U10643 (N_10643,N_10453,N_10506);
nor U10644 (N_10644,N_10499,N_10456);
nand U10645 (N_10645,N_10557,N_10418);
and U10646 (N_10646,N_10428,N_10478);
xnor U10647 (N_10647,N_10481,N_10505);
and U10648 (N_10648,N_10474,N_10410);
or U10649 (N_10649,N_10494,N_10515);
or U10650 (N_10650,N_10509,N_10532);
nor U10651 (N_10651,N_10555,N_10516);
xnor U10652 (N_10652,N_10542,N_10471);
xor U10653 (N_10653,N_10532,N_10518);
nor U10654 (N_10654,N_10409,N_10519);
and U10655 (N_10655,N_10502,N_10535);
nor U10656 (N_10656,N_10462,N_10477);
xnor U10657 (N_10657,N_10435,N_10423);
xnor U10658 (N_10658,N_10448,N_10507);
nand U10659 (N_10659,N_10482,N_10497);
nand U10660 (N_10660,N_10522,N_10487);
nand U10661 (N_10661,N_10467,N_10553);
nor U10662 (N_10662,N_10523,N_10471);
nor U10663 (N_10663,N_10528,N_10489);
or U10664 (N_10664,N_10410,N_10532);
or U10665 (N_10665,N_10484,N_10459);
xor U10666 (N_10666,N_10478,N_10489);
or U10667 (N_10667,N_10456,N_10543);
or U10668 (N_10668,N_10400,N_10441);
nor U10669 (N_10669,N_10448,N_10514);
xnor U10670 (N_10670,N_10410,N_10483);
and U10671 (N_10671,N_10498,N_10470);
nor U10672 (N_10672,N_10485,N_10476);
nor U10673 (N_10673,N_10493,N_10547);
xnor U10674 (N_10674,N_10490,N_10504);
or U10675 (N_10675,N_10451,N_10504);
or U10676 (N_10676,N_10546,N_10532);
nor U10677 (N_10677,N_10489,N_10458);
or U10678 (N_10678,N_10536,N_10533);
and U10679 (N_10679,N_10424,N_10553);
or U10680 (N_10680,N_10437,N_10405);
or U10681 (N_10681,N_10475,N_10477);
nand U10682 (N_10682,N_10557,N_10470);
and U10683 (N_10683,N_10450,N_10405);
nand U10684 (N_10684,N_10425,N_10518);
or U10685 (N_10685,N_10470,N_10512);
xor U10686 (N_10686,N_10503,N_10479);
nand U10687 (N_10687,N_10545,N_10405);
and U10688 (N_10688,N_10496,N_10429);
nand U10689 (N_10689,N_10501,N_10405);
xor U10690 (N_10690,N_10403,N_10523);
nand U10691 (N_10691,N_10510,N_10460);
nand U10692 (N_10692,N_10550,N_10437);
nor U10693 (N_10693,N_10437,N_10412);
nand U10694 (N_10694,N_10469,N_10444);
xor U10695 (N_10695,N_10432,N_10445);
and U10696 (N_10696,N_10541,N_10511);
nor U10697 (N_10697,N_10526,N_10479);
or U10698 (N_10698,N_10537,N_10425);
nor U10699 (N_10699,N_10509,N_10458);
nor U10700 (N_10700,N_10469,N_10430);
or U10701 (N_10701,N_10432,N_10542);
xor U10702 (N_10702,N_10417,N_10497);
nand U10703 (N_10703,N_10528,N_10411);
nor U10704 (N_10704,N_10438,N_10518);
nand U10705 (N_10705,N_10491,N_10436);
or U10706 (N_10706,N_10458,N_10449);
nand U10707 (N_10707,N_10444,N_10415);
nor U10708 (N_10708,N_10544,N_10437);
nand U10709 (N_10709,N_10448,N_10528);
xnor U10710 (N_10710,N_10522,N_10420);
nand U10711 (N_10711,N_10411,N_10412);
xnor U10712 (N_10712,N_10557,N_10486);
nor U10713 (N_10713,N_10511,N_10433);
xnor U10714 (N_10714,N_10426,N_10471);
or U10715 (N_10715,N_10535,N_10442);
nor U10716 (N_10716,N_10544,N_10449);
nand U10717 (N_10717,N_10457,N_10436);
and U10718 (N_10718,N_10487,N_10559);
and U10719 (N_10719,N_10411,N_10549);
and U10720 (N_10720,N_10718,N_10596);
and U10721 (N_10721,N_10594,N_10710);
nand U10722 (N_10722,N_10579,N_10578);
nand U10723 (N_10723,N_10619,N_10623);
and U10724 (N_10724,N_10646,N_10700);
or U10725 (N_10725,N_10681,N_10632);
or U10726 (N_10726,N_10657,N_10649);
or U10727 (N_10727,N_10691,N_10670);
and U10728 (N_10728,N_10690,N_10680);
nand U10729 (N_10729,N_10610,N_10659);
nor U10730 (N_10730,N_10641,N_10609);
and U10731 (N_10731,N_10573,N_10585);
xor U10732 (N_10732,N_10638,N_10713);
nand U10733 (N_10733,N_10591,N_10622);
xor U10734 (N_10734,N_10574,N_10589);
xor U10735 (N_10735,N_10561,N_10607);
xnor U10736 (N_10736,N_10715,N_10648);
or U10737 (N_10737,N_10592,N_10689);
and U10738 (N_10738,N_10667,N_10697);
and U10739 (N_10739,N_10582,N_10616);
or U10740 (N_10740,N_10629,N_10673);
and U10741 (N_10741,N_10562,N_10686);
or U10742 (N_10742,N_10640,N_10627);
nand U10743 (N_10743,N_10664,N_10630);
nor U10744 (N_10744,N_10599,N_10620);
nor U10745 (N_10745,N_10633,N_10661);
xor U10746 (N_10746,N_10569,N_10605);
nor U10747 (N_10747,N_10636,N_10564);
nand U10748 (N_10748,N_10590,N_10675);
nand U10749 (N_10749,N_10625,N_10666);
or U10750 (N_10750,N_10601,N_10575);
nand U10751 (N_10751,N_10603,N_10653);
and U10752 (N_10752,N_10598,N_10708);
and U10753 (N_10753,N_10679,N_10634);
nor U10754 (N_10754,N_10665,N_10705);
nor U10755 (N_10755,N_10674,N_10647);
nand U10756 (N_10756,N_10606,N_10572);
xnor U10757 (N_10757,N_10677,N_10684);
or U10758 (N_10758,N_10597,N_10614);
xnor U10759 (N_10759,N_10602,N_10699);
or U10760 (N_10760,N_10683,N_10698);
xnor U10761 (N_10761,N_10624,N_10621);
nor U10762 (N_10762,N_10707,N_10586);
xnor U10763 (N_10763,N_10650,N_10608);
nor U10764 (N_10764,N_10701,N_10628);
xor U10765 (N_10765,N_10583,N_10612);
or U10766 (N_10766,N_10672,N_10711);
nand U10767 (N_10767,N_10671,N_10717);
xor U10768 (N_10768,N_10694,N_10617);
nor U10769 (N_10769,N_10678,N_10600);
nand U10770 (N_10770,N_10669,N_10662);
xor U10771 (N_10771,N_10639,N_10702);
nand U10772 (N_10772,N_10695,N_10709);
nand U10773 (N_10773,N_10626,N_10567);
or U10774 (N_10774,N_10563,N_10696);
and U10775 (N_10775,N_10618,N_10645);
and U10776 (N_10776,N_10581,N_10584);
xor U10777 (N_10777,N_10663,N_10642);
nor U10778 (N_10778,N_10637,N_10651);
or U10779 (N_10779,N_10688,N_10676);
and U10780 (N_10780,N_10685,N_10643);
or U10781 (N_10781,N_10613,N_10615);
nor U10782 (N_10782,N_10692,N_10658);
or U10783 (N_10783,N_10588,N_10654);
xor U10784 (N_10784,N_10712,N_10682);
nand U10785 (N_10785,N_10580,N_10577);
nand U10786 (N_10786,N_10706,N_10593);
xnor U10787 (N_10787,N_10660,N_10604);
xnor U10788 (N_10788,N_10595,N_10652);
nand U10789 (N_10789,N_10668,N_10656);
and U10790 (N_10790,N_10576,N_10644);
or U10791 (N_10791,N_10566,N_10704);
nor U10792 (N_10792,N_10687,N_10714);
xor U10793 (N_10793,N_10571,N_10703);
nand U10794 (N_10794,N_10716,N_10560);
xnor U10795 (N_10795,N_10719,N_10635);
xnor U10796 (N_10796,N_10568,N_10565);
xor U10797 (N_10797,N_10693,N_10570);
nor U10798 (N_10798,N_10587,N_10655);
nor U10799 (N_10799,N_10611,N_10631);
nand U10800 (N_10800,N_10682,N_10688);
xnor U10801 (N_10801,N_10617,N_10560);
or U10802 (N_10802,N_10713,N_10602);
xor U10803 (N_10803,N_10676,N_10707);
nor U10804 (N_10804,N_10609,N_10578);
xor U10805 (N_10805,N_10660,N_10705);
and U10806 (N_10806,N_10652,N_10670);
nor U10807 (N_10807,N_10583,N_10685);
nor U10808 (N_10808,N_10675,N_10684);
nand U10809 (N_10809,N_10693,N_10628);
nand U10810 (N_10810,N_10710,N_10711);
xnor U10811 (N_10811,N_10565,N_10605);
nand U10812 (N_10812,N_10654,N_10644);
or U10813 (N_10813,N_10597,N_10609);
and U10814 (N_10814,N_10615,N_10623);
or U10815 (N_10815,N_10606,N_10688);
or U10816 (N_10816,N_10620,N_10665);
xnor U10817 (N_10817,N_10683,N_10707);
nand U10818 (N_10818,N_10590,N_10706);
and U10819 (N_10819,N_10584,N_10696);
or U10820 (N_10820,N_10620,N_10581);
or U10821 (N_10821,N_10637,N_10712);
nor U10822 (N_10822,N_10640,N_10641);
nor U10823 (N_10823,N_10595,N_10605);
nand U10824 (N_10824,N_10581,N_10611);
nand U10825 (N_10825,N_10590,N_10687);
and U10826 (N_10826,N_10600,N_10693);
xor U10827 (N_10827,N_10581,N_10621);
xnor U10828 (N_10828,N_10627,N_10620);
xnor U10829 (N_10829,N_10586,N_10597);
or U10830 (N_10830,N_10698,N_10661);
xnor U10831 (N_10831,N_10596,N_10641);
nand U10832 (N_10832,N_10696,N_10673);
xor U10833 (N_10833,N_10683,N_10597);
xor U10834 (N_10834,N_10602,N_10645);
nor U10835 (N_10835,N_10603,N_10621);
nand U10836 (N_10836,N_10630,N_10684);
and U10837 (N_10837,N_10636,N_10662);
or U10838 (N_10838,N_10713,N_10631);
nor U10839 (N_10839,N_10684,N_10646);
or U10840 (N_10840,N_10575,N_10591);
and U10841 (N_10841,N_10599,N_10566);
nand U10842 (N_10842,N_10601,N_10600);
xor U10843 (N_10843,N_10672,N_10675);
nor U10844 (N_10844,N_10701,N_10684);
xor U10845 (N_10845,N_10673,N_10643);
and U10846 (N_10846,N_10605,N_10696);
nor U10847 (N_10847,N_10670,N_10635);
nor U10848 (N_10848,N_10573,N_10656);
nand U10849 (N_10849,N_10565,N_10564);
or U10850 (N_10850,N_10679,N_10578);
nor U10851 (N_10851,N_10671,N_10706);
and U10852 (N_10852,N_10657,N_10630);
xor U10853 (N_10853,N_10696,N_10679);
nand U10854 (N_10854,N_10642,N_10602);
nor U10855 (N_10855,N_10690,N_10709);
nor U10856 (N_10856,N_10712,N_10718);
or U10857 (N_10857,N_10599,N_10657);
nor U10858 (N_10858,N_10632,N_10566);
nand U10859 (N_10859,N_10614,N_10667);
nor U10860 (N_10860,N_10677,N_10714);
xnor U10861 (N_10861,N_10602,N_10576);
nand U10862 (N_10862,N_10712,N_10635);
or U10863 (N_10863,N_10626,N_10579);
or U10864 (N_10864,N_10685,N_10639);
xnor U10865 (N_10865,N_10633,N_10708);
and U10866 (N_10866,N_10620,N_10562);
or U10867 (N_10867,N_10584,N_10661);
or U10868 (N_10868,N_10681,N_10674);
and U10869 (N_10869,N_10667,N_10715);
and U10870 (N_10870,N_10684,N_10597);
nor U10871 (N_10871,N_10652,N_10711);
xnor U10872 (N_10872,N_10629,N_10661);
or U10873 (N_10873,N_10667,N_10634);
nand U10874 (N_10874,N_10660,N_10627);
and U10875 (N_10875,N_10621,N_10571);
nand U10876 (N_10876,N_10620,N_10719);
nand U10877 (N_10877,N_10579,N_10600);
or U10878 (N_10878,N_10601,N_10590);
xnor U10879 (N_10879,N_10561,N_10678);
or U10880 (N_10880,N_10793,N_10784);
or U10881 (N_10881,N_10877,N_10720);
and U10882 (N_10882,N_10808,N_10835);
nand U10883 (N_10883,N_10876,N_10726);
nand U10884 (N_10884,N_10841,N_10815);
and U10885 (N_10885,N_10727,N_10852);
and U10886 (N_10886,N_10828,N_10741);
xnor U10887 (N_10887,N_10811,N_10824);
xnor U10888 (N_10888,N_10774,N_10779);
xnor U10889 (N_10889,N_10776,N_10758);
and U10890 (N_10890,N_10754,N_10753);
nor U10891 (N_10891,N_10782,N_10761);
nor U10892 (N_10892,N_10867,N_10866);
xnor U10893 (N_10893,N_10833,N_10851);
xnor U10894 (N_10894,N_10735,N_10829);
nand U10895 (N_10895,N_10752,N_10757);
nor U10896 (N_10896,N_10874,N_10818);
nand U10897 (N_10897,N_10799,N_10781);
nor U10898 (N_10898,N_10763,N_10842);
or U10899 (N_10899,N_10821,N_10791);
or U10900 (N_10900,N_10839,N_10856);
and U10901 (N_10901,N_10834,N_10858);
nand U10902 (N_10902,N_10816,N_10859);
or U10903 (N_10903,N_10838,N_10790);
nand U10904 (N_10904,N_10743,N_10728);
nand U10905 (N_10905,N_10783,N_10853);
nand U10906 (N_10906,N_10854,N_10809);
xnor U10907 (N_10907,N_10827,N_10813);
and U10908 (N_10908,N_10855,N_10810);
nand U10909 (N_10909,N_10857,N_10734);
nand U10910 (N_10910,N_10739,N_10806);
nand U10911 (N_10911,N_10765,N_10875);
or U10912 (N_10912,N_10729,N_10733);
nor U10913 (N_10913,N_10770,N_10848);
xor U10914 (N_10914,N_10803,N_10814);
xor U10915 (N_10915,N_10836,N_10830);
xnor U10916 (N_10916,N_10766,N_10863);
and U10917 (N_10917,N_10843,N_10879);
xnor U10918 (N_10918,N_10736,N_10747);
nand U10919 (N_10919,N_10749,N_10724);
nand U10920 (N_10920,N_10723,N_10725);
or U10921 (N_10921,N_10801,N_10837);
or U10922 (N_10922,N_10764,N_10796);
and U10923 (N_10923,N_10844,N_10798);
nand U10924 (N_10924,N_10750,N_10751);
or U10925 (N_10925,N_10772,N_10759);
nand U10926 (N_10926,N_10831,N_10804);
and U10927 (N_10927,N_10742,N_10785);
nor U10928 (N_10928,N_10744,N_10862);
nand U10929 (N_10929,N_10777,N_10840);
nand U10930 (N_10930,N_10786,N_10760);
nor U10931 (N_10931,N_10871,N_10771);
nor U10932 (N_10932,N_10878,N_10778);
or U10933 (N_10933,N_10792,N_10850);
nor U10934 (N_10934,N_10773,N_10870);
xor U10935 (N_10935,N_10794,N_10769);
or U10936 (N_10936,N_10789,N_10787);
nand U10937 (N_10937,N_10748,N_10788);
nor U10938 (N_10938,N_10802,N_10817);
or U10939 (N_10939,N_10807,N_10846);
nand U10940 (N_10940,N_10861,N_10860);
and U10941 (N_10941,N_10780,N_10865);
and U10942 (N_10942,N_10812,N_10746);
nor U10943 (N_10943,N_10868,N_10832);
nor U10944 (N_10944,N_10737,N_10849);
and U10945 (N_10945,N_10762,N_10847);
xor U10946 (N_10946,N_10797,N_10823);
xnor U10947 (N_10947,N_10819,N_10775);
xor U10948 (N_10948,N_10805,N_10732);
nor U10949 (N_10949,N_10722,N_10795);
xnor U10950 (N_10950,N_10731,N_10820);
and U10951 (N_10951,N_10738,N_10756);
xor U10952 (N_10952,N_10869,N_10864);
nand U10953 (N_10953,N_10755,N_10730);
nand U10954 (N_10954,N_10845,N_10721);
and U10955 (N_10955,N_10872,N_10822);
and U10956 (N_10956,N_10825,N_10826);
and U10957 (N_10957,N_10745,N_10767);
xor U10958 (N_10958,N_10800,N_10768);
and U10959 (N_10959,N_10873,N_10740);
and U10960 (N_10960,N_10800,N_10727);
nor U10961 (N_10961,N_10871,N_10740);
xnor U10962 (N_10962,N_10735,N_10744);
or U10963 (N_10963,N_10771,N_10753);
nor U10964 (N_10964,N_10862,N_10726);
or U10965 (N_10965,N_10808,N_10738);
xnor U10966 (N_10966,N_10847,N_10808);
or U10967 (N_10967,N_10818,N_10737);
or U10968 (N_10968,N_10812,N_10841);
xor U10969 (N_10969,N_10779,N_10724);
or U10970 (N_10970,N_10726,N_10756);
and U10971 (N_10971,N_10742,N_10853);
and U10972 (N_10972,N_10737,N_10721);
xnor U10973 (N_10973,N_10798,N_10726);
and U10974 (N_10974,N_10721,N_10729);
and U10975 (N_10975,N_10796,N_10768);
and U10976 (N_10976,N_10774,N_10860);
xor U10977 (N_10977,N_10742,N_10795);
xnor U10978 (N_10978,N_10807,N_10767);
nand U10979 (N_10979,N_10826,N_10764);
nor U10980 (N_10980,N_10797,N_10766);
nand U10981 (N_10981,N_10800,N_10824);
nor U10982 (N_10982,N_10748,N_10868);
nor U10983 (N_10983,N_10817,N_10733);
nor U10984 (N_10984,N_10846,N_10879);
and U10985 (N_10985,N_10751,N_10757);
or U10986 (N_10986,N_10773,N_10770);
nor U10987 (N_10987,N_10850,N_10741);
and U10988 (N_10988,N_10867,N_10808);
xor U10989 (N_10989,N_10819,N_10874);
nor U10990 (N_10990,N_10854,N_10790);
and U10991 (N_10991,N_10725,N_10779);
nand U10992 (N_10992,N_10774,N_10780);
nor U10993 (N_10993,N_10815,N_10750);
and U10994 (N_10994,N_10801,N_10740);
or U10995 (N_10995,N_10776,N_10836);
or U10996 (N_10996,N_10777,N_10758);
and U10997 (N_10997,N_10862,N_10783);
nor U10998 (N_10998,N_10764,N_10799);
nand U10999 (N_10999,N_10800,N_10736);
and U11000 (N_11000,N_10740,N_10744);
or U11001 (N_11001,N_10797,N_10722);
or U11002 (N_11002,N_10833,N_10786);
nor U11003 (N_11003,N_10804,N_10806);
nand U11004 (N_11004,N_10806,N_10770);
or U11005 (N_11005,N_10720,N_10845);
nor U11006 (N_11006,N_10827,N_10792);
xor U11007 (N_11007,N_10760,N_10858);
xor U11008 (N_11008,N_10793,N_10785);
nor U11009 (N_11009,N_10811,N_10821);
nand U11010 (N_11010,N_10866,N_10756);
nand U11011 (N_11011,N_10722,N_10746);
xor U11012 (N_11012,N_10783,N_10824);
and U11013 (N_11013,N_10863,N_10839);
nand U11014 (N_11014,N_10775,N_10846);
nor U11015 (N_11015,N_10771,N_10866);
and U11016 (N_11016,N_10722,N_10863);
and U11017 (N_11017,N_10829,N_10849);
or U11018 (N_11018,N_10737,N_10724);
or U11019 (N_11019,N_10763,N_10766);
nand U11020 (N_11020,N_10825,N_10843);
nor U11021 (N_11021,N_10794,N_10788);
xor U11022 (N_11022,N_10801,N_10862);
nand U11023 (N_11023,N_10855,N_10793);
or U11024 (N_11024,N_10747,N_10763);
nand U11025 (N_11025,N_10765,N_10785);
or U11026 (N_11026,N_10730,N_10823);
and U11027 (N_11027,N_10731,N_10848);
and U11028 (N_11028,N_10848,N_10773);
and U11029 (N_11029,N_10849,N_10818);
or U11030 (N_11030,N_10809,N_10838);
nand U11031 (N_11031,N_10828,N_10754);
nor U11032 (N_11032,N_10826,N_10809);
nand U11033 (N_11033,N_10815,N_10864);
or U11034 (N_11034,N_10867,N_10811);
nand U11035 (N_11035,N_10799,N_10867);
nand U11036 (N_11036,N_10831,N_10773);
and U11037 (N_11037,N_10866,N_10742);
nand U11038 (N_11038,N_10847,N_10835);
or U11039 (N_11039,N_10803,N_10873);
nand U11040 (N_11040,N_10935,N_10965);
and U11041 (N_11041,N_10948,N_10962);
and U11042 (N_11042,N_10911,N_10886);
or U11043 (N_11043,N_10989,N_10956);
nand U11044 (N_11044,N_10926,N_11031);
nand U11045 (N_11045,N_10949,N_10998);
xor U11046 (N_11046,N_10982,N_10999);
xor U11047 (N_11047,N_10921,N_10990);
nand U11048 (N_11048,N_11017,N_10928);
nor U11049 (N_11049,N_10986,N_10975);
xnor U11050 (N_11050,N_10993,N_10942);
nor U11051 (N_11051,N_11009,N_10915);
or U11052 (N_11052,N_10970,N_10918);
and U11053 (N_11053,N_10973,N_11038);
and U11054 (N_11054,N_10932,N_10909);
xnor U11055 (N_11055,N_10937,N_11004);
xnor U11056 (N_11056,N_11013,N_10945);
xnor U11057 (N_11057,N_10951,N_11008);
nand U11058 (N_11058,N_10997,N_10946);
or U11059 (N_11059,N_11016,N_10978);
xnor U11060 (N_11060,N_11039,N_10923);
nor U11061 (N_11061,N_10938,N_11032);
and U11062 (N_11062,N_11026,N_10972);
xnor U11063 (N_11063,N_10985,N_10930);
xor U11064 (N_11064,N_10910,N_10924);
xnor U11065 (N_11065,N_10885,N_10908);
and U11066 (N_11066,N_11023,N_11018);
or U11067 (N_11067,N_11007,N_11027);
nor U11068 (N_11068,N_11014,N_10901);
or U11069 (N_11069,N_11021,N_10905);
nor U11070 (N_11070,N_10936,N_10967);
and U11071 (N_11071,N_10958,N_11000);
nand U11072 (N_11072,N_10934,N_11001);
nor U11073 (N_11073,N_11024,N_11020);
and U11074 (N_11074,N_10880,N_10960);
nand U11075 (N_11075,N_10996,N_11036);
and U11076 (N_11076,N_10898,N_10953);
and U11077 (N_11077,N_10884,N_10976);
or U11078 (N_11078,N_11010,N_10919);
xor U11079 (N_11079,N_11002,N_10897);
nor U11080 (N_11080,N_10920,N_10927);
nand U11081 (N_11081,N_10912,N_10891);
xnor U11082 (N_11082,N_10979,N_10964);
xnor U11083 (N_11083,N_10994,N_10944);
or U11084 (N_11084,N_10933,N_10947);
nor U11085 (N_11085,N_10955,N_10968);
and U11086 (N_11086,N_11029,N_11033);
and U11087 (N_11087,N_10974,N_10903);
and U11088 (N_11088,N_10889,N_10957);
or U11089 (N_11089,N_10896,N_10882);
nand U11090 (N_11090,N_10992,N_11015);
or U11091 (N_11091,N_10907,N_10987);
and U11092 (N_11092,N_10939,N_10913);
nand U11093 (N_11093,N_10980,N_10925);
xor U11094 (N_11094,N_11034,N_10916);
xor U11095 (N_11095,N_10963,N_10900);
nor U11096 (N_11096,N_10940,N_10902);
nor U11097 (N_11097,N_10892,N_11003);
xnor U11098 (N_11098,N_10991,N_10883);
xor U11099 (N_11099,N_10931,N_11028);
xnor U11100 (N_11100,N_10922,N_10961);
nand U11101 (N_11101,N_11035,N_10929);
or U11102 (N_11102,N_10943,N_10971);
nand U11103 (N_11103,N_11019,N_10966);
xor U11104 (N_11104,N_11022,N_10969);
or U11105 (N_11105,N_10887,N_10952);
nand U11106 (N_11106,N_11012,N_11005);
or U11107 (N_11107,N_11037,N_10983);
and U11108 (N_11108,N_10890,N_10950);
nor U11109 (N_11109,N_10984,N_10893);
xnor U11110 (N_11110,N_10899,N_10904);
xor U11111 (N_11111,N_10977,N_10895);
nor U11112 (N_11112,N_10906,N_10917);
nor U11113 (N_11113,N_10894,N_10914);
and U11114 (N_11114,N_11011,N_10959);
xor U11115 (N_11115,N_10981,N_11030);
nand U11116 (N_11116,N_10888,N_10941);
or U11117 (N_11117,N_11025,N_11006);
nand U11118 (N_11118,N_10881,N_10995);
and U11119 (N_11119,N_10954,N_10988);
xnor U11120 (N_11120,N_10929,N_11011);
nor U11121 (N_11121,N_10899,N_11036);
xor U11122 (N_11122,N_10966,N_10942);
nand U11123 (N_11123,N_10967,N_10977);
nor U11124 (N_11124,N_10930,N_10894);
xnor U11125 (N_11125,N_10906,N_10909);
or U11126 (N_11126,N_11025,N_11020);
xnor U11127 (N_11127,N_10882,N_11013);
xnor U11128 (N_11128,N_10991,N_11038);
nor U11129 (N_11129,N_10998,N_10942);
xnor U11130 (N_11130,N_11008,N_10922);
nand U11131 (N_11131,N_10946,N_10984);
and U11132 (N_11132,N_11003,N_10887);
xor U11133 (N_11133,N_10936,N_10992);
nor U11134 (N_11134,N_10927,N_10990);
nor U11135 (N_11135,N_10935,N_11017);
xnor U11136 (N_11136,N_10943,N_11008);
or U11137 (N_11137,N_11033,N_11038);
nor U11138 (N_11138,N_10956,N_10915);
nand U11139 (N_11139,N_10957,N_10934);
nand U11140 (N_11140,N_10907,N_11021);
xnor U11141 (N_11141,N_10908,N_10946);
nand U11142 (N_11142,N_11012,N_10977);
nor U11143 (N_11143,N_11008,N_11038);
nand U11144 (N_11144,N_10977,N_11020);
or U11145 (N_11145,N_10934,N_11005);
and U11146 (N_11146,N_10919,N_10971);
and U11147 (N_11147,N_11023,N_10927);
nand U11148 (N_11148,N_10889,N_10986);
or U11149 (N_11149,N_11026,N_11003);
and U11150 (N_11150,N_10956,N_10897);
or U11151 (N_11151,N_10901,N_11039);
nor U11152 (N_11152,N_10980,N_10931);
and U11153 (N_11153,N_10946,N_10974);
or U11154 (N_11154,N_10909,N_10882);
and U11155 (N_11155,N_11004,N_10917);
and U11156 (N_11156,N_10965,N_11001);
xor U11157 (N_11157,N_10978,N_10959);
or U11158 (N_11158,N_10983,N_11035);
and U11159 (N_11159,N_10915,N_10913);
and U11160 (N_11160,N_11022,N_10999);
or U11161 (N_11161,N_11038,N_10900);
and U11162 (N_11162,N_11012,N_10943);
xnor U11163 (N_11163,N_10889,N_10942);
xor U11164 (N_11164,N_10926,N_10891);
or U11165 (N_11165,N_10964,N_11031);
or U11166 (N_11166,N_10959,N_11020);
nor U11167 (N_11167,N_10951,N_10994);
nor U11168 (N_11168,N_10948,N_10944);
nand U11169 (N_11169,N_10959,N_11034);
and U11170 (N_11170,N_10957,N_10907);
xnor U11171 (N_11171,N_11022,N_10931);
nor U11172 (N_11172,N_11032,N_10936);
or U11173 (N_11173,N_10943,N_11017);
xor U11174 (N_11174,N_11011,N_10888);
nand U11175 (N_11175,N_10908,N_10979);
and U11176 (N_11176,N_11018,N_10898);
nand U11177 (N_11177,N_10930,N_10914);
xnor U11178 (N_11178,N_11016,N_11019);
xnor U11179 (N_11179,N_11001,N_10999);
nand U11180 (N_11180,N_10900,N_10971);
nand U11181 (N_11181,N_10900,N_10975);
nor U11182 (N_11182,N_10920,N_11024);
and U11183 (N_11183,N_10980,N_10986);
and U11184 (N_11184,N_10950,N_10960);
and U11185 (N_11185,N_10899,N_11024);
xnor U11186 (N_11186,N_10888,N_10988);
nor U11187 (N_11187,N_10951,N_10979);
or U11188 (N_11188,N_10911,N_11021);
nand U11189 (N_11189,N_11026,N_11031);
nor U11190 (N_11190,N_10913,N_11012);
nor U11191 (N_11191,N_10919,N_10956);
nand U11192 (N_11192,N_10952,N_10969);
xor U11193 (N_11193,N_10902,N_10891);
and U11194 (N_11194,N_10999,N_10913);
and U11195 (N_11195,N_10941,N_10957);
and U11196 (N_11196,N_10952,N_10987);
xnor U11197 (N_11197,N_10990,N_10951);
and U11198 (N_11198,N_10881,N_11010);
or U11199 (N_11199,N_10980,N_10910);
nor U11200 (N_11200,N_11168,N_11195);
xnor U11201 (N_11201,N_11192,N_11092);
xnor U11202 (N_11202,N_11095,N_11115);
or U11203 (N_11203,N_11136,N_11066);
or U11204 (N_11204,N_11041,N_11125);
and U11205 (N_11205,N_11098,N_11104);
nand U11206 (N_11206,N_11132,N_11176);
xnor U11207 (N_11207,N_11061,N_11078);
nand U11208 (N_11208,N_11122,N_11193);
xnor U11209 (N_11209,N_11081,N_11045);
or U11210 (N_11210,N_11067,N_11179);
nand U11211 (N_11211,N_11171,N_11180);
nand U11212 (N_11212,N_11099,N_11172);
nand U11213 (N_11213,N_11077,N_11083);
nor U11214 (N_11214,N_11184,N_11135);
or U11215 (N_11215,N_11189,N_11147);
nor U11216 (N_11216,N_11134,N_11120);
xnor U11217 (N_11217,N_11127,N_11182);
xor U11218 (N_11218,N_11177,N_11074);
nand U11219 (N_11219,N_11137,N_11054);
and U11220 (N_11220,N_11194,N_11052);
nor U11221 (N_11221,N_11173,N_11086);
or U11222 (N_11222,N_11129,N_11149);
and U11223 (N_11223,N_11040,N_11152);
or U11224 (N_11224,N_11091,N_11139);
and U11225 (N_11225,N_11146,N_11148);
nor U11226 (N_11226,N_11117,N_11118);
nand U11227 (N_11227,N_11153,N_11069);
xor U11228 (N_11228,N_11053,N_11130);
nor U11229 (N_11229,N_11043,N_11113);
or U11230 (N_11230,N_11063,N_11112);
nand U11231 (N_11231,N_11105,N_11072);
and U11232 (N_11232,N_11065,N_11056);
and U11233 (N_11233,N_11191,N_11109);
and U11234 (N_11234,N_11094,N_11181);
nor U11235 (N_11235,N_11140,N_11158);
nand U11236 (N_11236,N_11150,N_11143);
nor U11237 (N_11237,N_11196,N_11082);
or U11238 (N_11238,N_11154,N_11107);
nand U11239 (N_11239,N_11062,N_11163);
nor U11240 (N_11240,N_11089,N_11198);
xor U11241 (N_11241,N_11073,N_11049);
nand U11242 (N_11242,N_11151,N_11197);
nor U11243 (N_11243,N_11123,N_11126);
xor U11244 (N_11244,N_11157,N_11183);
and U11245 (N_11245,N_11097,N_11080);
nor U11246 (N_11246,N_11048,N_11188);
nand U11247 (N_11247,N_11050,N_11046);
nand U11248 (N_11248,N_11145,N_11161);
xnor U11249 (N_11249,N_11075,N_11068);
nor U11250 (N_11250,N_11190,N_11199);
nor U11251 (N_11251,N_11090,N_11055);
and U11252 (N_11252,N_11131,N_11141);
or U11253 (N_11253,N_11174,N_11100);
xnor U11254 (N_11254,N_11165,N_11114);
and U11255 (N_11255,N_11169,N_11044);
nand U11256 (N_11256,N_11133,N_11087);
or U11257 (N_11257,N_11144,N_11166);
and U11258 (N_11258,N_11138,N_11101);
nand U11259 (N_11259,N_11121,N_11128);
and U11260 (N_11260,N_11108,N_11096);
xor U11261 (N_11261,N_11186,N_11103);
nand U11262 (N_11262,N_11059,N_11106);
and U11263 (N_11263,N_11124,N_11110);
xor U11264 (N_11264,N_11058,N_11116);
xor U11265 (N_11265,N_11111,N_11071);
nor U11266 (N_11266,N_11076,N_11060);
and U11267 (N_11267,N_11162,N_11156);
nor U11268 (N_11268,N_11160,N_11187);
or U11269 (N_11269,N_11093,N_11057);
nor U11270 (N_11270,N_11119,N_11088);
nand U11271 (N_11271,N_11185,N_11178);
nor U11272 (N_11272,N_11102,N_11042);
nor U11273 (N_11273,N_11051,N_11047);
nand U11274 (N_11274,N_11142,N_11085);
nor U11275 (N_11275,N_11164,N_11070);
and U11276 (N_11276,N_11167,N_11064);
nor U11277 (N_11277,N_11170,N_11079);
xor U11278 (N_11278,N_11155,N_11175);
or U11279 (N_11279,N_11159,N_11084);
or U11280 (N_11280,N_11148,N_11069);
nand U11281 (N_11281,N_11094,N_11115);
nor U11282 (N_11282,N_11140,N_11199);
nor U11283 (N_11283,N_11075,N_11056);
nand U11284 (N_11284,N_11197,N_11142);
and U11285 (N_11285,N_11083,N_11113);
nor U11286 (N_11286,N_11095,N_11192);
and U11287 (N_11287,N_11055,N_11070);
or U11288 (N_11288,N_11049,N_11191);
nor U11289 (N_11289,N_11106,N_11056);
or U11290 (N_11290,N_11160,N_11199);
nand U11291 (N_11291,N_11164,N_11123);
nor U11292 (N_11292,N_11126,N_11098);
nand U11293 (N_11293,N_11081,N_11107);
xor U11294 (N_11294,N_11193,N_11127);
xor U11295 (N_11295,N_11166,N_11087);
or U11296 (N_11296,N_11154,N_11116);
and U11297 (N_11297,N_11137,N_11181);
xnor U11298 (N_11298,N_11048,N_11082);
and U11299 (N_11299,N_11115,N_11167);
nand U11300 (N_11300,N_11041,N_11068);
xor U11301 (N_11301,N_11056,N_11197);
or U11302 (N_11302,N_11137,N_11079);
xnor U11303 (N_11303,N_11061,N_11161);
nand U11304 (N_11304,N_11084,N_11109);
xor U11305 (N_11305,N_11176,N_11043);
xnor U11306 (N_11306,N_11145,N_11088);
or U11307 (N_11307,N_11087,N_11165);
xnor U11308 (N_11308,N_11113,N_11048);
nor U11309 (N_11309,N_11151,N_11068);
and U11310 (N_11310,N_11185,N_11116);
xnor U11311 (N_11311,N_11189,N_11196);
xnor U11312 (N_11312,N_11082,N_11194);
xor U11313 (N_11313,N_11155,N_11107);
xnor U11314 (N_11314,N_11129,N_11103);
nor U11315 (N_11315,N_11155,N_11103);
xor U11316 (N_11316,N_11083,N_11163);
or U11317 (N_11317,N_11178,N_11120);
nand U11318 (N_11318,N_11114,N_11048);
nand U11319 (N_11319,N_11148,N_11054);
or U11320 (N_11320,N_11183,N_11070);
and U11321 (N_11321,N_11098,N_11101);
and U11322 (N_11322,N_11083,N_11056);
xnor U11323 (N_11323,N_11080,N_11194);
nand U11324 (N_11324,N_11068,N_11161);
or U11325 (N_11325,N_11057,N_11144);
nor U11326 (N_11326,N_11157,N_11143);
nand U11327 (N_11327,N_11144,N_11126);
or U11328 (N_11328,N_11158,N_11053);
nand U11329 (N_11329,N_11169,N_11067);
and U11330 (N_11330,N_11044,N_11111);
nand U11331 (N_11331,N_11069,N_11175);
or U11332 (N_11332,N_11185,N_11127);
nor U11333 (N_11333,N_11135,N_11198);
or U11334 (N_11334,N_11171,N_11052);
or U11335 (N_11335,N_11048,N_11198);
nor U11336 (N_11336,N_11117,N_11086);
xnor U11337 (N_11337,N_11081,N_11147);
nor U11338 (N_11338,N_11046,N_11043);
nor U11339 (N_11339,N_11064,N_11084);
nor U11340 (N_11340,N_11172,N_11169);
nor U11341 (N_11341,N_11199,N_11197);
nor U11342 (N_11342,N_11084,N_11040);
and U11343 (N_11343,N_11135,N_11104);
xnor U11344 (N_11344,N_11070,N_11082);
or U11345 (N_11345,N_11056,N_11199);
and U11346 (N_11346,N_11190,N_11167);
xnor U11347 (N_11347,N_11162,N_11051);
or U11348 (N_11348,N_11125,N_11103);
nand U11349 (N_11349,N_11104,N_11193);
or U11350 (N_11350,N_11076,N_11091);
or U11351 (N_11351,N_11180,N_11168);
and U11352 (N_11352,N_11117,N_11148);
nand U11353 (N_11353,N_11177,N_11084);
and U11354 (N_11354,N_11188,N_11167);
xnor U11355 (N_11355,N_11080,N_11089);
nor U11356 (N_11356,N_11092,N_11149);
or U11357 (N_11357,N_11194,N_11042);
xor U11358 (N_11358,N_11162,N_11059);
xor U11359 (N_11359,N_11126,N_11198);
and U11360 (N_11360,N_11270,N_11257);
nor U11361 (N_11361,N_11242,N_11286);
nand U11362 (N_11362,N_11230,N_11273);
nor U11363 (N_11363,N_11333,N_11272);
and U11364 (N_11364,N_11305,N_11251);
nor U11365 (N_11365,N_11347,N_11319);
or U11366 (N_11366,N_11239,N_11307);
nor U11367 (N_11367,N_11342,N_11244);
nand U11368 (N_11368,N_11229,N_11262);
xnor U11369 (N_11369,N_11339,N_11241);
nor U11370 (N_11370,N_11250,N_11329);
nor U11371 (N_11371,N_11265,N_11285);
xor U11372 (N_11372,N_11247,N_11224);
and U11373 (N_11373,N_11222,N_11240);
nor U11374 (N_11374,N_11353,N_11304);
or U11375 (N_11375,N_11284,N_11253);
and U11376 (N_11376,N_11358,N_11261);
xor U11377 (N_11377,N_11323,N_11238);
nor U11378 (N_11378,N_11302,N_11288);
and U11379 (N_11379,N_11298,N_11200);
nand U11380 (N_11380,N_11279,N_11255);
and U11381 (N_11381,N_11225,N_11281);
and U11382 (N_11382,N_11337,N_11275);
and U11383 (N_11383,N_11325,N_11228);
or U11384 (N_11384,N_11259,N_11231);
xnor U11385 (N_11385,N_11248,N_11219);
xor U11386 (N_11386,N_11343,N_11268);
and U11387 (N_11387,N_11296,N_11233);
xor U11388 (N_11388,N_11292,N_11301);
xor U11389 (N_11389,N_11269,N_11293);
nor U11390 (N_11390,N_11313,N_11356);
and U11391 (N_11391,N_11349,N_11338);
and U11392 (N_11392,N_11266,N_11320);
nor U11393 (N_11393,N_11274,N_11202);
xor U11394 (N_11394,N_11314,N_11263);
nor U11395 (N_11395,N_11352,N_11326);
xnor U11396 (N_11396,N_11341,N_11345);
nor U11397 (N_11397,N_11316,N_11237);
or U11398 (N_11398,N_11297,N_11318);
or U11399 (N_11399,N_11346,N_11232);
and U11400 (N_11400,N_11243,N_11271);
xnor U11401 (N_11401,N_11290,N_11215);
nor U11402 (N_11402,N_11209,N_11223);
and U11403 (N_11403,N_11221,N_11249);
nand U11404 (N_11404,N_11203,N_11310);
nor U11405 (N_11405,N_11324,N_11294);
nor U11406 (N_11406,N_11227,N_11252);
and U11407 (N_11407,N_11201,N_11254);
and U11408 (N_11408,N_11303,N_11214);
nor U11409 (N_11409,N_11277,N_11213);
nand U11410 (N_11410,N_11295,N_11308);
xnor U11411 (N_11411,N_11210,N_11246);
xor U11412 (N_11412,N_11334,N_11354);
and U11413 (N_11413,N_11258,N_11217);
nand U11414 (N_11414,N_11315,N_11260);
nand U11415 (N_11415,N_11218,N_11317);
xor U11416 (N_11416,N_11321,N_11283);
nor U11417 (N_11417,N_11336,N_11299);
nand U11418 (N_11418,N_11267,N_11206);
or U11419 (N_11419,N_11351,N_11300);
and U11420 (N_11420,N_11208,N_11234);
nand U11421 (N_11421,N_11235,N_11291);
nand U11422 (N_11422,N_11245,N_11306);
and U11423 (N_11423,N_11327,N_11212);
or U11424 (N_11424,N_11348,N_11340);
and U11425 (N_11425,N_11328,N_11236);
and U11426 (N_11426,N_11204,N_11331);
or U11427 (N_11427,N_11220,N_11322);
and U11428 (N_11428,N_11216,N_11205);
nand U11429 (N_11429,N_11289,N_11330);
nand U11430 (N_11430,N_11359,N_11287);
xnor U11431 (N_11431,N_11282,N_11357);
xnor U11432 (N_11432,N_11278,N_11344);
nor U11433 (N_11433,N_11355,N_11207);
or U11434 (N_11434,N_11264,N_11280);
nor U11435 (N_11435,N_11276,N_11332);
or U11436 (N_11436,N_11312,N_11350);
xor U11437 (N_11437,N_11309,N_11256);
xnor U11438 (N_11438,N_11311,N_11226);
xor U11439 (N_11439,N_11211,N_11335);
or U11440 (N_11440,N_11315,N_11287);
or U11441 (N_11441,N_11343,N_11351);
or U11442 (N_11442,N_11235,N_11351);
and U11443 (N_11443,N_11258,N_11201);
nand U11444 (N_11444,N_11244,N_11332);
xor U11445 (N_11445,N_11211,N_11219);
nor U11446 (N_11446,N_11221,N_11287);
and U11447 (N_11447,N_11211,N_11304);
nor U11448 (N_11448,N_11207,N_11255);
nor U11449 (N_11449,N_11254,N_11307);
xnor U11450 (N_11450,N_11231,N_11309);
nand U11451 (N_11451,N_11342,N_11287);
xnor U11452 (N_11452,N_11248,N_11216);
nand U11453 (N_11453,N_11338,N_11259);
nor U11454 (N_11454,N_11241,N_11352);
or U11455 (N_11455,N_11209,N_11240);
xnor U11456 (N_11456,N_11306,N_11250);
and U11457 (N_11457,N_11232,N_11267);
nor U11458 (N_11458,N_11238,N_11306);
nand U11459 (N_11459,N_11222,N_11314);
nand U11460 (N_11460,N_11359,N_11211);
and U11461 (N_11461,N_11314,N_11233);
nor U11462 (N_11462,N_11275,N_11209);
or U11463 (N_11463,N_11309,N_11338);
xnor U11464 (N_11464,N_11224,N_11357);
or U11465 (N_11465,N_11217,N_11298);
or U11466 (N_11466,N_11356,N_11309);
nor U11467 (N_11467,N_11275,N_11314);
and U11468 (N_11468,N_11239,N_11352);
nand U11469 (N_11469,N_11213,N_11212);
nor U11470 (N_11470,N_11259,N_11319);
or U11471 (N_11471,N_11205,N_11238);
or U11472 (N_11472,N_11292,N_11333);
or U11473 (N_11473,N_11333,N_11227);
and U11474 (N_11474,N_11209,N_11307);
nand U11475 (N_11475,N_11270,N_11278);
and U11476 (N_11476,N_11251,N_11269);
nand U11477 (N_11477,N_11221,N_11218);
nor U11478 (N_11478,N_11278,N_11323);
and U11479 (N_11479,N_11246,N_11209);
xor U11480 (N_11480,N_11232,N_11256);
or U11481 (N_11481,N_11270,N_11295);
nand U11482 (N_11482,N_11298,N_11288);
or U11483 (N_11483,N_11303,N_11299);
nand U11484 (N_11484,N_11338,N_11262);
and U11485 (N_11485,N_11355,N_11206);
nor U11486 (N_11486,N_11204,N_11332);
nand U11487 (N_11487,N_11231,N_11248);
or U11488 (N_11488,N_11321,N_11293);
nor U11489 (N_11489,N_11261,N_11272);
or U11490 (N_11490,N_11305,N_11283);
nand U11491 (N_11491,N_11213,N_11294);
nor U11492 (N_11492,N_11307,N_11233);
xor U11493 (N_11493,N_11323,N_11235);
nor U11494 (N_11494,N_11231,N_11303);
nand U11495 (N_11495,N_11283,N_11350);
and U11496 (N_11496,N_11266,N_11206);
nand U11497 (N_11497,N_11215,N_11237);
and U11498 (N_11498,N_11338,N_11257);
and U11499 (N_11499,N_11232,N_11235);
nor U11500 (N_11500,N_11293,N_11206);
or U11501 (N_11501,N_11357,N_11305);
or U11502 (N_11502,N_11278,N_11274);
xnor U11503 (N_11503,N_11319,N_11314);
nor U11504 (N_11504,N_11256,N_11217);
nand U11505 (N_11505,N_11266,N_11286);
xnor U11506 (N_11506,N_11257,N_11269);
xor U11507 (N_11507,N_11227,N_11292);
or U11508 (N_11508,N_11300,N_11249);
or U11509 (N_11509,N_11233,N_11204);
or U11510 (N_11510,N_11255,N_11256);
nand U11511 (N_11511,N_11215,N_11301);
nor U11512 (N_11512,N_11303,N_11223);
or U11513 (N_11513,N_11213,N_11233);
nand U11514 (N_11514,N_11294,N_11329);
xnor U11515 (N_11515,N_11265,N_11292);
or U11516 (N_11516,N_11203,N_11290);
nand U11517 (N_11517,N_11211,N_11273);
nor U11518 (N_11518,N_11277,N_11306);
nor U11519 (N_11519,N_11327,N_11309);
or U11520 (N_11520,N_11406,N_11444);
nor U11521 (N_11521,N_11364,N_11397);
xor U11522 (N_11522,N_11401,N_11494);
and U11523 (N_11523,N_11509,N_11470);
and U11524 (N_11524,N_11395,N_11402);
xor U11525 (N_11525,N_11475,N_11400);
nor U11526 (N_11526,N_11491,N_11483);
nand U11527 (N_11527,N_11378,N_11504);
or U11528 (N_11528,N_11394,N_11512);
nand U11529 (N_11529,N_11452,N_11375);
xnor U11530 (N_11530,N_11510,N_11431);
nor U11531 (N_11531,N_11481,N_11453);
nand U11532 (N_11532,N_11461,N_11390);
xor U11533 (N_11533,N_11518,N_11478);
and U11534 (N_11534,N_11437,N_11460);
or U11535 (N_11535,N_11404,N_11422);
nor U11536 (N_11536,N_11489,N_11362);
xnor U11537 (N_11537,N_11389,N_11467);
or U11538 (N_11538,N_11502,N_11411);
nand U11539 (N_11539,N_11474,N_11454);
nor U11540 (N_11540,N_11449,N_11407);
and U11541 (N_11541,N_11487,N_11516);
and U11542 (N_11542,N_11365,N_11499);
or U11543 (N_11543,N_11371,N_11488);
nor U11544 (N_11544,N_11519,N_11408);
nand U11545 (N_11545,N_11485,N_11438);
or U11546 (N_11546,N_11514,N_11373);
xnor U11547 (N_11547,N_11459,N_11505);
nor U11548 (N_11548,N_11420,N_11445);
nand U11549 (N_11549,N_11496,N_11451);
xnor U11550 (N_11550,N_11419,N_11398);
and U11551 (N_11551,N_11434,N_11477);
nand U11552 (N_11552,N_11476,N_11486);
nand U11553 (N_11553,N_11480,N_11428);
nand U11554 (N_11554,N_11412,N_11429);
nor U11555 (N_11555,N_11513,N_11403);
xor U11556 (N_11556,N_11497,N_11376);
or U11557 (N_11557,N_11457,N_11501);
nor U11558 (N_11558,N_11368,N_11415);
nand U11559 (N_11559,N_11442,N_11500);
nor U11560 (N_11560,N_11440,N_11462);
and U11561 (N_11561,N_11482,N_11456);
xnor U11562 (N_11562,N_11433,N_11507);
or U11563 (N_11563,N_11423,N_11447);
nor U11564 (N_11564,N_11387,N_11466);
or U11565 (N_11565,N_11490,N_11413);
nand U11566 (N_11566,N_11381,N_11464);
nand U11567 (N_11567,N_11409,N_11424);
nand U11568 (N_11568,N_11430,N_11472);
nor U11569 (N_11569,N_11410,N_11463);
xnor U11570 (N_11570,N_11511,N_11498);
and U11571 (N_11571,N_11372,N_11436);
nand U11572 (N_11572,N_11388,N_11484);
and U11573 (N_11573,N_11468,N_11448);
nor U11574 (N_11574,N_11515,N_11503);
xor U11575 (N_11575,N_11446,N_11435);
xor U11576 (N_11576,N_11379,N_11366);
nor U11577 (N_11577,N_11361,N_11382);
or U11578 (N_11578,N_11506,N_11405);
or U11579 (N_11579,N_11416,N_11426);
nor U11580 (N_11580,N_11414,N_11465);
xor U11581 (N_11581,N_11374,N_11369);
or U11582 (N_11582,N_11418,N_11384);
xnor U11583 (N_11583,N_11396,N_11425);
nand U11584 (N_11584,N_11508,N_11471);
and U11585 (N_11585,N_11517,N_11360);
and U11586 (N_11586,N_11385,N_11455);
or U11587 (N_11587,N_11443,N_11439);
nand U11588 (N_11588,N_11383,N_11367);
and U11589 (N_11589,N_11391,N_11386);
nand U11590 (N_11590,N_11393,N_11377);
and U11591 (N_11591,N_11417,N_11370);
nor U11592 (N_11592,N_11473,N_11392);
nand U11593 (N_11593,N_11479,N_11492);
and U11594 (N_11594,N_11469,N_11493);
nor U11595 (N_11595,N_11495,N_11399);
or U11596 (N_11596,N_11450,N_11458);
xor U11597 (N_11597,N_11380,N_11421);
nand U11598 (N_11598,N_11427,N_11441);
or U11599 (N_11599,N_11363,N_11432);
and U11600 (N_11600,N_11476,N_11516);
or U11601 (N_11601,N_11387,N_11452);
and U11602 (N_11602,N_11448,N_11447);
nor U11603 (N_11603,N_11372,N_11490);
or U11604 (N_11604,N_11424,N_11492);
and U11605 (N_11605,N_11497,N_11364);
or U11606 (N_11606,N_11448,N_11411);
nand U11607 (N_11607,N_11431,N_11497);
nor U11608 (N_11608,N_11406,N_11370);
and U11609 (N_11609,N_11458,N_11510);
nor U11610 (N_11610,N_11506,N_11416);
xor U11611 (N_11611,N_11475,N_11412);
nand U11612 (N_11612,N_11439,N_11469);
nor U11613 (N_11613,N_11514,N_11461);
nor U11614 (N_11614,N_11373,N_11428);
or U11615 (N_11615,N_11443,N_11382);
nand U11616 (N_11616,N_11412,N_11507);
nor U11617 (N_11617,N_11517,N_11507);
and U11618 (N_11618,N_11500,N_11456);
nand U11619 (N_11619,N_11472,N_11481);
or U11620 (N_11620,N_11463,N_11381);
and U11621 (N_11621,N_11456,N_11519);
nor U11622 (N_11622,N_11389,N_11413);
and U11623 (N_11623,N_11502,N_11480);
xnor U11624 (N_11624,N_11466,N_11496);
or U11625 (N_11625,N_11469,N_11387);
xnor U11626 (N_11626,N_11519,N_11480);
nor U11627 (N_11627,N_11510,N_11460);
or U11628 (N_11628,N_11381,N_11412);
nand U11629 (N_11629,N_11493,N_11430);
nand U11630 (N_11630,N_11372,N_11371);
nor U11631 (N_11631,N_11471,N_11387);
xor U11632 (N_11632,N_11456,N_11462);
or U11633 (N_11633,N_11391,N_11417);
nor U11634 (N_11634,N_11486,N_11470);
or U11635 (N_11635,N_11421,N_11509);
nor U11636 (N_11636,N_11465,N_11499);
nor U11637 (N_11637,N_11499,N_11395);
and U11638 (N_11638,N_11446,N_11449);
or U11639 (N_11639,N_11477,N_11461);
or U11640 (N_11640,N_11370,N_11493);
nor U11641 (N_11641,N_11485,N_11361);
nand U11642 (N_11642,N_11502,N_11505);
nor U11643 (N_11643,N_11466,N_11512);
and U11644 (N_11644,N_11428,N_11482);
and U11645 (N_11645,N_11431,N_11480);
nor U11646 (N_11646,N_11380,N_11448);
xor U11647 (N_11647,N_11398,N_11476);
xnor U11648 (N_11648,N_11482,N_11361);
nor U11649 (N_11649,N_11366,N_11411);
nand U11650 (N_11650,N_11446,N_11367);
and U11651 (N_11651,N_11518,N_11369);
nand U11652 (N_11652,N_11474,N_11451);
nor U11653 (N_11653,N_11511,N_11500);
nand U11654 (N_11654,N_11400,N_11437);
nand U11655 (N_11655,N_11514,N_11386);
xor U11656 (N_11656,N_11381,N_11513);
and U11657 (N_11657,N_11516,N_11390);
xnor U11658 (N_11658,N_11367,N_11518);
nand U11659 (N_11659,N_11501,N_11438);
and U11660 (N_11660,N_11363,N_11439);
and U11661 (N_11661,N_11473,N_11418);
nor U11662 (N_11662,N_11388,N_11514);
nand U11663 (N_11663,N_11517,N_11433);
and U11664 (N_11664,N_11395,N_11480);
nor U11665 (N_11665,N_11488,N_11437);
and U11666 (N_11666,N_11499,N_11472);
or U11667 (N_11667,N_11434,N_11363);
nor U11668 (N_11668,N_11495,N_11510);
xnor U11669 (N_11669,N_11433,N_11482);
or U11670 (N_11670,N_11386,N_11431);
nand U11671 (N_11671,N_11462,N_11482);
nand U11672 (N_11672,N_11414,N_11413);
nor U11673 (N_11673,N_11387,N_11394);
nand U11674 (N_11674,N_11517,N_11465);
xor U11675 (N_11675,N_11496,N_11500);
and U11676 (N_11676,N_11414,N_11399);
xnor U11677 (N_11677,N_11511,N_11460);
nand U11678 (N_11678,N_11496,N_11369);
nand U11679 (N_11679,N_11519,N_11455);
nor U11680 (N_11680,N_11548,N_11648);
nor U11681 (N_11681,N_11566,N_11625);
nand U11682 (N_11682,N_11677,N_11656);
xor U11683 (N_11683,N_11575,N_11543);
and U11684 (N_11684,N_11520,N_11572);
and U11685 (N_11685,N_11624,N_11598);
nor U11686 (N_11686,N_11580,N_11675);
nand U11687 (N_11687,N_11650,N_11556);
nand U11688 (N_11688,N_11521,N_11576);
nor U11689 (N_11689,N_11557,N_11615);
and U11690 (N_11690,N_11593,N_11545);
nor U11691 (N_11691,N_11619,N_11551);
and U11692 (N_11692,N_11607,N_11562);
or U11693 (N_11693,N_11589,N_11643);
nor U11694 (N_11694,N_11555,N_11629);
nor U11695 (N_11695,N_11622,N_11561);
xnor U11696 (N_11696,N_11670,N_11582);
and U11697 (N_11697,N_11570,N_11620);
xnor U11698 (N_11698,N_11617,N_11621);
xor U11699 (N_11699,N_11639,N_11553);
xnor U11700 (N_11700,N_11671,N_11541);
or U11701 (N_11701,N_11649,N_11550);
nor U11702 (N_11702,N_11601,N_11596);
nor U11703 (N_11703,N_11638,N_11569);
xor U11704 (N_11704,N_11532,N_11535);
and U11705 (N_11705,N_11546,N_11667);
nor U11706 (N_11706,N_11531,N_11544);
nor U11707 (N_11707,N_11653,N_11529);
and U11708 (N_11708,N_11537,N_11586);
xnor U11709 (N_11709,N_11608,N_11633);
and U11710 (N_11710,N_11573,N_11577);
nor U11711 (N_11711,N_11669,N_11567);
nor U11712 (N_11712,N_11602,N_11534);
nand U11713 (N_11713,N_11554,N_11604);
and U11714 (N_11714,N_11610,N_11642);
and U11715 (N_11715,N_11590,N_11563);
xnor U11716 (N_11716,N_11655,N_11628);
xor U11717 (N_11717,N_11581,N_11672);
xnor U11718 (N_11718,N_11522,N_11578);
nor U11719 (N_11719,N_11536,N_11658);
nand U11720 (N_11720,N_11528,N_11665);
and U11721 (N_11721,N_11565,N_11525);
xnor U11722 (N_11722,N_11645,N_11636);
nor U11723 (N_11723,N_11647,N_11540);
nor U11724 (N_11724,N_11652,N_11668);
xor U11725 (N_11725,N_11614,N_11646);
nor U11726 (N_11726,N_11660,N_11592);
nand U11727 (N_11727,N_11552,N_11631);
xnor U11728 (N_11728,N_11626,N_11523);
xor U11729 (N_11729,N_11630,N_11588);
or U11730 (N_11730,N_11587,N_11605);
and U11731 (N_11731,N_11659,N_11591);
nor U11732 (N_11732,N_11676,N_11603);
or U11733 (N_11733,N_11526,N_11651);
or U11734 (N_11734,N_11595,N_11558);
or U11735 (N_11735,N_11564,N_11634);
nand U11736 (N_11736,N_11549,N_11606);
nand U11737 (N_11737,N_11533,N_11635);
nand U11738 (N_11738,N_11663,N_11585);
nand U11739 (N_11739,N_11679,N_11644);
or U11740 (N_11740,N_11661,N_11616);
nand U11741 (N_11741,N_11538,N_11597);
xnor U11742 (N_11742,N_11571,N_11641);
or U11743 (N_11743,N_11611,N_11613);
nand U11744 (N_11744,N_11527,N_11662);
and U11745 (N_11745,N_11574,N_11568);
nor U11746 (N_11746,N_11637,N_11654);
xnor U11747 (N_11747,N_11657,N_11664);
xnor U11748 (N_11748,N_11560,N_11579);
xor U11749 (N_11749,N_11559,N_11612);
or U11750 (N_11750,N_11609,N_11594);
nor U11751 (N_11751,N_11539,N_11542);
xor U11752 (N_11752,N_11627,N_11584);
nor U11753 (N_11753,N_11618,N_11600);
xnor U11754 (N_11754,N_11547,N_11583);
nand U11755 (N_11755,N_11674,N_11623);
and U11756 (N_11756,N_11640,N_11678);
nor U11757 (N_11757,N_11666,N_11524);
or U11758 (N_11758,N_11632,N_11673);
nor U11759 (N_11759,N_11599,N_11530);
xor U11760 (N_11760,N_11632,N_11660);
nor U11761 (N_11761,N_11585,N_11527);
or U11762 (N_11762,N_11565,N_11621);
xor U11763 (N_11763,N_11679,N_11664);
or U11764 (N_11764,N_11554,N_11642);
nor U11765 (N_11765,N_11625,N_11592);
nand U11766 (N_11766,N_11666,N_11548);
nor U11767 (N_11767,N_11674,N_11678);
and U11768 (N_11768,N_11651,N_11595);
nand U11769 (N_11769,N_11545,N_11575);
or U11770 (N_11770,N_11590,N_11565);
or U11771 (N_11771,N_11561,N_11630);
or U11772 (N_11772,N_11576,N_11668);
and U11773 (N_11773,N_11607,N_11663);
xnor U11774 (N_11774,N_11637,N_11609);
nor U11775 (N_11775,N_11586,N_11675);
and U11776 (N_11776,N_11678,N_11626);
nor U11777 (N_11777,N_11648,N_11606);
or U11778 (N_11778,N_11538,N_11574);
nand U11779 (N_11779,N_11574,N_11605);
and U11780 (N_11780,N_11664,N_11640);
xor U11781 (N_11781,N_11563,N_11648);
nor U11782 (N_11782,N_11577,N_11642);
or U11783 (N_11783,N_11597,N_11593);
nand U11784 (N_11784,N_11531,N_11620);
or U11785 (N_11785,N_11626,N_11527);
nand U11786 (N_11786,N_11585,N_11644);
and U11787 (N_11787,N_11645,N_11618);
nand U11788 (N_11788,N_11654,N_11520);
and U11789 (N_11789,N_11556,N_11543);
nor U11790 (N_11790,N_11677,N_11520);
xnor U11791 (N_11791,N_11595,N_11652);
or U11792 (N_11792,N_11679,N_11620);
nor U11793 (N_11793,N_11563,N_11646);
and U11794 (N_11794,N_11607,N_11621);
or U11795 (N_11795,N_11630,N_11653);
or U11796 (N_11796,N_11554,N_11530);
xor U11797 (N_11797,N_11603,N_11641);
nand U11798 (N_11798,N_11593,N_11530);
or U11799 (N_11799,N_11585,N_11639);
or U11800 (N_11800,N_11620,N_11555);
xnor U11801 (N_11801,N_11629,N_11668);
and U11802 (N_11802,N_11636,N_11622);
nor U11803 (N_11803,N_11520,N_11594);
nand U11804 (N_11804,N_11529,N_11569);
nand U11805 (N_11805,N_11636,N_11534);
and U11806 (N_11806,N_11670,N_11660);
nor U11807 (N_11807,N_11589,N_11641);
xor U11808 (N_11808,N_11650,N_11577);
and U11809 (N_11809,N_11655,N_11531);
or U11810 (N_11810,N_11545,N_11537);
nor U11811 (N_11811,N_11620,N_11602);
or U11812 (N_11812,N_11587,N_11663);
nor U11813 (N_11813,N_11569,N_11623);
xnor U11814 (N_11814,N_11610,N_11646);
and U11815 (N_11815,N_11669,N_11613);
nor U11816 (N_11816,N_11522,N_11616);
or U11817 (N_11817,N_11589,N_11546);
nor U11818 (N_11818,N_11547,N_11539);
or U11819 (N_11819,N_11536,N_11652);
and U11820 (N_11820,N_11527,N_11584);
xnor U11821 (N_11821,N_11664,N_11627);
xnor U11822 (N_11822,N_11651,N_11553);
nand U11823 (N_11823,N_11676,N_11678);
nand U11824 (N_11824,N_11540,N_11602);
xnor U11825 (N_11825,N_11661,N_11627);
xnor U11826 (N_11826,N_11544,N_11675);
xnor U11827 (N_11827,N_11520,N_11562);
xnor U11828 (N_11828,N_11642,N_11674);
and U11829 (N_11829,N_11632,N_11527);
xnor U11830 (N_11830,N_11627,N_11570);
nand U11831 (N_11831,N_11563,N_11628);
or U11832 (N_11832,N_11643,N_11671);
and U11833 (N_11833,N_11620,N_11658);
xor U11834 (N_11834,N_11582,N_11615);
and U11835 (N_11835,N_11645,N_11646);
and U11836 (N_11836,N_11600,N_11552);
nand U11837 (N_11837,N_11640,N_11576);
and U11838 (N_11838,N_11634,N_11638);
or U11839 (N_11839,N_11586,N_11526);
nand U11840 (N_11840,N_11766,N_11830);
xnor U11841 (N_11841,N_11726,N_11781);
or U11842 (N_11842,N_11764,N_11790);
or U11843 (N_11843,N_11829,N_11804);
nor U11844 (N_11844,N_11687,N_11736);
xor U11845 (N_11845,N_11729,N_11775);
nor U11846 (N_11846,N_11691,N_11753);
and U11847 (N_11847,N_11724,N_11796);
and U11848 (N_11848,N_11718,N_11803);
or U11849 (N_11849,N_11744,N_11686);
and U11850 (N_11850,N_11778,N_11794);
nand U11851 (N_11851,N_11770,N_11811);
or U11852 (N_11852,N_11838,N_11784);
and U11853 (N_11853,N_11730,N_11831);
and U11854 (N_11854,N_11695,N_11828);
nand U11855 (N_11855,N_11700,N_11772);
or U11856 (N_11856,N_11745,N_11692);
or U11857 (N_11857,N_11740,N_11735);
or U11858 (N_11858,N_11743,N_11754);
or U11859 (N_11859,N_11833,N_11777);
nor U11860 (N_11860,N_11731,N_11683);
nor U11861 (N_11861,N_11819,N_11806);
or U11862 (N_11862,N_11779,N_11768);
and U11863 (N_11863,N_11818,N_11782);
nand U11864 (N_11864,N_11705,N_11802);
xnor U11865 (N_11865,N_11693,N_11721);
or U11866 (N_11866,N_11680,N_11732);
nor U11867 (N_11867,N_11799,N_11719);
or U11868 (N_11868,N_11767,N_11760);
nand U11869 (N_11869,N_11747,N_11688);
nand U11870 (N_11870,N_11698,N_11707);
or U11871 (N_11871,N_11708,N_11765);
and U11872 (N_11872,N_11715,N_11762);
or U11873 (N_11873,N_11773,N_11706);
nand U11874 (N_11874,N_11684,N_11734);
xor U11875 (N_11875,N_11751,N_11815);
xor U11876 (N_11876,N_11822,N_11834);
or U11877 (N_11877,N_11791,N_11723);
xnor U11878 (N_11878,N_11826,N_11788);
or U11879 (N_11879,N_11716,N_11701);
and U11880 (N_11880,N_11789,N_11824);
xor U11881 (N_11881,N_11816,N_11758);
xnor U11882 (N_11882,N_11714,N_11807);
and U11883 (N_11883,N_11738,N_11769);
nand U11884 (N_11884,N_11713,N_11711);
or U11885 (N_11885,N_11812,N_11703);
xnor U11886 (N_11886,N_11800,N_11783);
nor U11887 (N_11887,N_11685,N_11746);
xnor U11888 (N_11888,N_11820,N_11697);
nand U11889 (N_11889,N_11709,N_11725);
or U11890 (N_11890,N_11710,N_11756);
nor U11891 (N_11891,N_11681,N_11763);
xor U11892 (N_11892,N_11798,N_11809);
xnor U11893 (N_11893,N_11810,N_11696);
nor U11894 (N_11894,N_11827,N_11817);
xnor U11895 (N_11895,N_11771,N_11717);
nor U11896 (N_11896,N_11759,N_11823);
xor U11897 (N_11897,N_11702,N_11786);
nor U11898 (N_11898,N_11792,N_11814);
or U11899 (N_11899,N_11720,N_11739);
nor U11900 (N_11900,N_11780,N_11813);
xnor U11901 (N_11901,N_11748,N_11749);
xor U11902 (N_11902,N_11808,N_11839);
xor U11903 (N_11903,N_11837,N_11712);
xor U11904 (N_11904,N_11699,N_11755);
xnor U11905 (N_11905,N_11832,N_11776);
nand U11906 (N_11906,N_11821,N_11689);
and U11907 (N_11907,N_11757,N_11805);
or U11908 (N_11908,N_11787,N_11752);
xor U11909 (N_11909,N_11797,N_11737);
or U11910 (N_11910,N_11750,N_11704);
nor U11911 (N_11911,N_11727,N_11785);
nand U11912 (N_11912,N_11694,N_11795);
xnor U11913 (N_11913,N_11722,N_11774);
nand U11914 (N_11914,N_11836,N_11793);
xor U11915 (N_11915,N_11741,N_11761);
and U11916 (N_11916,N_11742,N_11835);
and U11917 (N_11917,N_11682,N_11690);
or U11918 (N_11918,N_11728,N_11825);
and U11919 (N_11919,N_11733,N_11801);
xnor U11920 (N_11920,N_11800,N_11714);
nand U11921 (N_11921,N_11705,N_11838);
and U11922 (N_11922,N_11737,N_11752);
and U11923 (N_11923,N_11796,N_11744);
nor U11924 (N_11924,N_11706,N_11681);
xor U11925 (N_11925,N_11717,N_11786);
and U11926 (N_11926,N_11826,N_11719);
or U11927 (N_11927,N_11775,N_11753);
nor U11928 (N_11928,N_11705,N_11829);
nand U11929 (N_11929,N_11747,N_11812);
and U11930 (N_11930,N_11799,N_11715);
or U11931 (N_11931,N_11685,N_11836);
xor U11932 (N_11932,N_11680,N_11742);
xor U11933 (N_11933,N_11700,N_11833);
nand U11934 (N_11934,N_11827,N_11784);
nand U11935 (N_11935,N_11748,N_11762);
xnor U11936 (N_11936,N_11839,N_11832);
and U11937 (N_11937,N_11788,N_11798);
nand U11938 (N_11938,N_11835,N_11815);
nor U11939 (N_11939,N_11760,N_11783);
and U11940 (N_11940,N_11733,N_11732);
or U11941 (N_11941,N_11737,N_11817);
nand U11942 (N_11942,N_11703,N_11808);
xnor U11943 (N_11943,N_11756,N_11735);
nand U11944 (N_11944,N_11715,N_11809);
nand U11945 (N_11945,N_11786,N_11804);
nand U11946 (N_11946,N_11749,N_11743);
nand U11947 (N_11947,N_11759,N_11812);
nand U11948 (N_11948,N_11821,N_11802);
nor U11949 (N_11949,N_11826,N_11713);
nand U11950 (N_11950,N_11824,N_11750);
and U11951 (N_11951,N_11689,N_11771);
nand U11952 (N_11952,N_11785,N_11830);
xor U11953 (N_11953,N_11828,N_11811);
nand U11954 (N_11954,N_11693,N_11724);
or U11955 (N_11955,N_11694,N_11757);
nand U11956 (N_11956,N_11796,N_11701);
nor U11957 (N_11957,N_11770,N_11690);
nand U11958 (N_11958,N_11712,N_11813);
nand U11959 (N_11959,N_11686,N_11748);
nor U11960 (N_11960,N_11788,N_11685);
xnor U11961 (N_11961,N_11836,N_11771);
and U11962 (N_11962,N_11706,N_11754);
nor U11963 (N_11963,N_11686,N_11826);
nor U11964 (N_11964,N_11741,N_11748);
and U11965 (N_11965,N_11723,N_11747);
nand U11966 (N_11966,N_11806,N_11699);
or U11967 (N_11967,N_11781,N_11825);
nand U11968 (N_11968,N_11704,N_11733);
and U11969 (N_11969,N_11784,N_11743);
xor U11970 (N_11970,N_11786,N_11809);
or U11971 (N_11971,N_11741,N_11809);
or U11972 (N_11972,N_11765,N_11802);
nor U11973 (N_11973,N_11764,N_11716);
and U11974 (N_11974,N_11750,N_11733);
or U11975 (N_11975,N_11688,N_11798);
nand U11976 (N_11976,N_11695,N_11747);
xnor U11977 (N_11977,N_11760,N_11825);
nand U11978 (N_11978,N_11694,N_11693);
nand U11979 (N_11979,N_11836,N_11816);
nand U11980 (N_11980,N_11689,N_11686);
nand U11981 (N_11981,N_11766,N_11685);
or U11982 (N_11982,N_11819,N_11740);
nand U11983 (N_11983,N_11826,N_11684);
or U11984 (N_11984,N_11767,N_11740);
nor U11985 (N_11985,N_11794,N_11777);
nor U11986 (N_11986,N_11812,N_11776);
nor U11987 (N_11987,N_11754,N_11685);
or U11988 (N_11988,N_11750,N_11818);
xor U11989 (N_11989,N_11702,N_11728);
and U11990 (N_11990,N_11753,N_11836);
or U11991 (N_11991,N_11714,N_11827);
xor U11992 (N_11992,N_11749,N_11721);
nor U11993 (N_11993,N_11744,N_11780);
xnor U11994 (N_11994,N_11763,N_11794);
and U11995 (N_11995,N_11757,N_11766);
xor U11996 (N_11996,N_11755,N_11698);
and U11997 (N_11997,N_11705,N_11805);
or U11998 (N_11998,N_11825,N_11818);
xnor U11999 (N_11999,N_11830,N_11836);
xnor U12000 (N_12000,N_11855,N_11984);
nand U12001 (N_12001,N_11926,N_11890);
or U12002 (N_12002,N_11887,N_11970);
xor U12003 (N_12003,N_11871,N_11892);
or U12004 (N_12004,N_11967,N_11917);
and U12005 (N_12005,N_11928,N_11941);
and U12006 (N_12006,N_11988,N_11929);
nor U12007 (N_12007,N_11897,N_11888);
nand U12008 (N_12008,N_11850,N_11921);
and U12009 (N_12009,N_11977,N_11965);
nand U12010 (N_12010,N_11969,N_11859);
nor U12011 (N_12011,N_11955,N_11920);
or U12012 (N_12012,N_11936,N_11865);
or U12013 (N_12013,N_11885,N_11842);
nor U12014 (N_12014,N_11944,N_11933);
nand U12015 (N_12015,N_11915,N_11895);
and U12016 (N_12016,N_11978,N_11957);
and U12017 (N_12017,N_11996,N_11923);
nor U12018 (N_12018,N_11878,N_11953);
nand U12019 (N_12019,N_11930,N_11992);
or U12020 (N_12020,N_11877,N_11873);
nor U12021 (N_12021,N_11975,N_11924);
and U12022 (N_12022,N_11863,N_11862);
and U12023 (N_12023,N_11946,N_11896);
xor U12024 (N_12024,N_11952,N_11971);
and U12025 (N_12025,N_11904,N_11854);
nand U12026 (N_12026,N_11851,N_11905);
xor U12027 (N_12027,N_11907,N_11991);
nor U12028 (N_12028,N_11961,N_11937);
nand U12029 (N_12029,N_11932,N_11857);
nand U12030 (N_12030,N_11900,N_11940);
nand U12031 (N_12031,N_11943,N_11879);
xor U12032 (N_12032,N_11945,N_11880);
and U12033 (N_12033,N_11852,N_11968);
xor U12034 (N_12034,N_11976,N_11962);
xnor U12035 (N_12035,N_11919,N_11973);
nand U12036 (N_12036,N_11882,N_11910);
and U12037 (N_12037,N_11939,N_11986);
and U12038 (N_12038,N_11860,N_11899);
nand U12039 (N_12039,N_11954,N_11960);
and U12040 (N_12040,N_11869,N_11989);
and U12041 (N_12041,N_11909,N_11918);
xor U12042 (N_12042,N_11934,N_11901);
xor U12043 (N_12043,N_11980,N_11902);
xnor U12044 (N_12044,N_11868,N_11974);
or U12045 (N_12045,N_11886,N_11853);
xnor U12046 (N_12046,N_11981,N_11874);
nand U12047 (N_12047,N_11883,N_11999);
nor U12048 (N_12048,N_11964,N_11891);
nand U12049 (N_12049,N_11903,N_11949);
xor U12050 (N_12050,N_11956,N_11914);
or U12051 (N_12051,N_11950,N_11972);
or U12052 (N_12052,N_11844,N_11959);
and U12053 (N_12053,N_11938,N_11947);
or U12054 (N_12054,N_11958,N_11846);
or U12055 (N_12055,N_11864,N_11983);
and U12056 (N_12056,N_11935,N_11963);
or U12057 (N_12057,N_11870,N_11966);
nor U12058 (N_12058,N_11998,N_11893);
xor U12059 (N_12059,N_11876,N_11995);
or U12060 (N_12060,N_11861,N_11990);
or U12061 (N_12061,N_11927,N_11913);
xnor U12062 (N_12062,N_11898,N_11866);
nand U12063 (N_12063,N_11849,N_11858);
xor U12064 (N_12064,N_11906,N_11997);
xor U12065 (N_12065,N_11845,N_11911);
xor U12066 (N_12066,N_11922,N_11908);
nand U12067 (N_12067,N_11925,N_11894);
nand U12068 (N_12068,N_11951,N_11942);
nor U12069 (N_12069,N_11948,N_11889);
xor U12070 (N_12070,N_11993,N_11982);
xor U12071 (N_12071,N_11987,N_11848);
xnor U12072 (N_12072,N_11840,N_11843);
and U12073 (N_12073,N_11881,N_11979);
xor U12074 (N_12074,N_11867,N_11985);
nand U12075 (N_12075,N_11912,N_11841);
nor U12076 (N_12076,N_11916,N_11872);
nand U12077 (N_12077,N_11856,N_11994);
xnor U12078 (N_12078,N_11931,N_11875);
nor U12079 (N_12079,N_11847,N_11884);
or U12080 (N_12080,N_11918,N_11934);
xnor U12081 (N_12081,N_11970,N_11856);
nor U12082 (N_12082,N_11920,N_11900);
and U12083 (N_12083,N_11892,N_11894);
or U12084 (N_12084,N_11916,N_11873);
xnor U12085 (N_12085,N_11954,N_11929);
nand U12086 (N_12086,N_11994,N_11913);
nor U12087 (N_12087,N_11903,N_11971);
and U12088 (N_12088,N_11994,N_11916);
nand U12089 (N_12089,N_11953,N_11924);
xnor U12090 (N_12090,N_11980,N_11895);
and U12091 (N_12091,N_11886,N_11977);
or U12092 (N_12092,N_11968,N_11932);
and U12093 (N_12093,N_11992,N_11867);
nor U12094 (N_12094,N_11951,N_11950);
nand U12095 (N_12095,N_11991,N_11849);
nand U12096 (N_12096,N_11929,N_11940);
nor U12097 (N_12097,N_11998,N_11864);
xor U12098 (N_12098,N_11922,N_11971);
nor U12099 (N_12099,N_11924,N_11997);
or U12100 (N_12100,N_11887,N_11968);
nand U12101 (N_12101,N_11941,N_11890);
xor U12102 (N_12102,N_11967,N_11892);
nand U12103 (N_12103,N_11914,N_11911);
nand U12104 (N_12104,N_11972,N_11899);
or U12105 (N_12105,N_11933,N_11941);
xor U12106 (N_12106,N_11968,N_11940);
and U12107 (N_12107,N_11924,N_11923);
nand U12108 (N_12108,N_11939,N_11858);
nand U12109 (N_12109,N_11917,N_11961);
xor U12110 (N_12110,N_11968,N_11862);
nand U12111 (N_12111,N_11890,N_11956);
nor U12112 (N_12112,N_11975,N_11845);
nand U12113 (N_12113,N_11857,N_11956);
nand U12114 (N_12114,N_11986,N_11845);
nand U12115 (N_12115,N_11991,N_11968);
nor U12116 (N_12116,N_11918,N_11911);
xor U12117 (N_12117,N_11931,N_11877);
and U12118 (N_12118,N_11954,N_11970);
nand U12119 (N_12119,N_11856,N_11857);
xnor U12120 (N_12120,N_11953,N_11974);
nand U12121 (N_12121,N_11888,N_11866);
nand U12122 (N_12122,N_11903,N_11841);
and U12123 (N_12123,N_11861,N_11867);
nor U12124 (N_12124,N_11996,N_11932);
xor U12125 (N_12125,N_11921,N_11941);
and U12126 (N_12126,N_11933,N_11900);
or U12127 (N_12127,N_11841,N_11860);
xnor U12128 (N_12128,N_11844,N_11943);
and U12129 (N_12129,N_11921,N_11938);
xor U12130 (N_12130,N_11886,N_11984);
and U12131 (N_12131,N_11990,N_11953);
nand U12132 (N_12132,N_11879,N_11885);
or U12133 (N_12133,N_11920,N_11865);
or U12134 (N_12134,N_11840,N_11981);
xor U12135 (N_12135,N_11997,N_11934);
and U12136 (N_12136,N_11926,N_11861);
or U12137 (N_12137,N_11991,N_11853);
or U12138 (N_12138,N_11996,N_11868);
nor U12139 (N_12139,N_11988,N_11927);
and U12140 (N_12140,N_11892,N_11901);
xnor U12141 (N_12141,N_11879,N_11905);
or U12142 (N_12142,N_11908,N_11976);
or U12143 (N_12143,N_11842,N_11934);
and U12144 (N_12144,N_11947,N_11942);
or U12145 (N_12145,N_11875,N_11962);
or U12146 (N_12146,N_11963,N_11956);
and U12147 (N_12147,N_11897,N_11915);
or U12148 (N_12148,N_11981,N_11887);
nor U12149 (N_12149,N_11978,N_11845);
xnor U12150 (N_12150,N_11872,N_11852);
nor U12151 (N_12151,N_11940,N_11939);
nor U12152 (N_12152,N_11994,N_11966);
or U12153 (N_12153,N_11996,N_11952);
nand U12154 (N_12154,N_11907,N_11904);
and U12155 (N_12155,N_11947,N_11954);
nand U12156 (N_12156,N_11896,N_11848);
nor U12157 (N_12157,N_11879,N_11861);
nor U12158 (N_12158,N_11878,N_11881);
nand U12159 (N_12159,N_11863,N_11939);
nand U12160 (N_12160,N_12042,N_12151);
and U12161 (N_12161,N_12146,N_12069);
nand U12162 (N_12162,N_12095,N_12027);
and U12163 (N_12163,N_12031,N_12093);
and U12164 (N_12164,N_12136,N_12020);
nor U12165 (N_12165,N_12054,N_12132);
xor U12166 (N_12166,N_12137,N_12080);
or U12167 (N_12167,N_12120,N_12060);
and U12168 (N_12168,N_12158,N_12133);
and U12169 (N_12169,N_12083,N_12111);
and U12170 (N_12170,N_12105,N_12110);
nor U12171 (N_12171,N_12068,N_12026);
and U12172 (N_12172,N_12021,N_12157);
or U12173 (N_12173,N_12088,N_12032);
or U12174 (N_12174,N_12097,N_12098);
xor U12175 (N_12175,N_12102,N_12138);
nand U12176 (N_12176,N_12152,N_12127);
xor U12177 (N_12177,N_12091,N_12147);
and U12178 (N_12178,N_12126,N_12086);
xor U12179 (N_12179,N_12008,N_12063);
nand U12180 (N_12180,N_12092,N_12051);
nor U12181 (N_12181,N_12022,N_12104);
and U12182 (N_12182,N_12028,N_12061);
nand U12183 (N_12183,N_12155,N_12002);
and U12184 (N_12184,N_12124,N_12082);
or U12185 (N_12185,N_12016,N_12119);
or U12186 (N_12186,N_12106,N_12050);
nor U12187 (N_12187,N_12077,N_12039);
and U12188 (N_12188,N_12135,N_12040);
nor U12189 (N_12189,N_12000,N_12023);
and U12190 (N_12190,N_12056,N_12018);
or U12191 (N_12191,N_12103,N_12059);
and U12192 (N_12192,N_12084,N_12094);
nand U12193 (N_12193,N_12129,N_12153);
nand U12194 (N_12194,N_12145,N_12079);
nor U12195 (N_12195,N_12113,N_12148);
and U12196 (N_12196,N_12053,N_12101);
or U12197 (N_12197,N_12035,N_12122);
and U12198 (N_12198,N_12078,N_12072);
nand U12199 (N_12199,N_12066,N_12012);
xnor U12200 (N_12200,N_12114,N_12123);
nor U12201 (N_12201,N_12150,N_12055);
or U12202 (N_12202,N_12115,N_12048);
or U12203 (N_12203,N_12070,N_12067);
xnor U12204 (N_12204,N_12041,N_12149);
or U12205 (N_12205,N_12052,N_12045);
xor U12206 (N_12206,N_12089,N_12030);
or U12207 (N_12207,N_12007,N_12112);
nand U12208 (N_12208,N_12001,N_12081);
or U12209 (N_12209,N_12076,N_12009);
and U12210 (N_12210,N_12128,N_12038);
nand U12211 (N_12211,N_12043,N_12010);
xor U12212 (N_12212,N_12116,N_12090);
xor U12213 (N_12213,N_12017,N_12003);
nand U12214 (N_12214,N_12049,N_12005);
or U12215 (N_12215,N_12019,N_12134);
xnor U12216 (N_12216,N_12074,N_12014);
nand U12217 (N_12217,N_12046,N_12071);
nor U12218 (N_12218,N_12065,N_12006);
nor U12219 (N_12219,N_12141,N_12064);
or U12220 (N_12220,N_12131,N_12159);
xnor U12221 (N_12221,N_12109,N_12142);
xnor U12222 (N_12222,N_12117,N_12034);
or U12223 (N_12223,N_12024,N_12058);
xor U12224 (N_12224,N_12015,N_12062);
nor U12225 (N_12225,N_12139,N_12004);
or U12226 (N_12226,N_12108,N_12044);
nor U12227 (N_12227,N_12057,N_12154);
nor U12228 (N_12228,N_12036,N_12140);
and U12229 (N_12229,N_12118,N_12073);
xor U12230 (N_12230,N_12130,N_12144);
nor U12231 (N_12231,N_12037,N_12100);
nand U12232 (N_12232,N_12156,N_12125);
nor U12233 (N_12233,N_12033,N_12075);
nor U12234 (N_12234,N_12029,N_12096);
nand U12235 (N_12235,N_12121,N_12143);
nor U12236 (N_12236,N_12099,N_12085);
or U12237 (N_12237,N_12047,N_12011);
nand U12238 (N_12238,N_12087,N_12013);
or U12239 (N_12239,N_12025,N_12107);
nor U12240 (N_12240,N_12080,N_12078);
nor U12241 (N_12241,N_12031,N_12052);
nand U12242 (N_12242,N_12122,N_12093);
and U12243 (N_12243,N_12142,N_12127);
xor U12244 (N_12244,N_12027,N_12034);
xor U12245 (N_12245,N_12073,N_12101);
or U12246 (N_12246,N_12005,N_12078);
xor U12247 (N_12247,N_12011,N_12145);
and U12248 (N_12248,N_12059,N_12106);
nand U12249 (N_12249,N_12064,N_12070);
nand U12250 (N_12250,N_12158,N_12157);
nand U12251 (N_12251,N_12042,N_12019);
and U12252 (N_12252,N_12024,N_12013);
and U12253 (N_12253,N_12067,N_12096);
or U12254 (N_12254,N_12058,N_12033);
or U12255 (N_12255,N_12122,N_12009);
and U12256 (N_12256,N_12146,N_12156);
or U12257 (N_12257,N_12132,N_12004);
nor U12258 (N_12258,N_12076,N_12124);
or U12259 (N_12259,N_12067,N_12057);
xor U12260 (N_12260,N_12060,N_12088);
and U12261 (N_12261,N_12127,N_12141);
and U12262 (N_12262,N_12066,N_12119);
nand U12263 (N_12263,N_12106,N_12142);
and U12264 (N_12264,N_12123,N_12038);
and U12265 (N_12265,N_12032,N_12151);
xnor U12266 (N_12266,N_12085,N_12113);
or U12267 (N_12267,N_12016,N_12153);
nor U12268 (N_12268,N_12129,N_12105);
and U12269 (N_12269,N_12123,N_12044);
or U12270 (N_12270,N_12001,N_12057);
and U12271 (N_12271,N_12092,N_12060);
xnor U12272 (N_12272,N_12154,N_12121);
nor U12273 (N_12273,N_12031,N_12101);
and U12274 (N_12274,N_12025,N_12106);
nand U12275 (N_12275,N_12111,N_12089);
xor U12276 (N_12276,N_12130,N_12069);
and U12277 (N_12277,N_12088,N_12105);
nand U12278 (N_12278,N_12076,N_12136);
and U12279 (N_12279,N_12145,N_12151);
and U12280 (N_12280,N_12137,N_12109);
or U12281 (N_12281,N_12154,N_12133);
and U12282 (N_12282,N_12107,N_12014);
and U12283 (N_12283,N_12085,N_12106);
nand U12284 (N_12284,N_12025,N_12102);
or U12285 (N_12285,N_12134,N_12025);
nor U12286 (N_12286,N_12039,N_12024);
nand U12287 (N_12287,N_12060,N_12053);
nor U12288 (N_12288,N_12062,N_12044);
and U12289 (N_12289,N_12050,N_12008);
nor U12290 (N_12290,N_12122,N_12049);
xnor U12291 (N_12291,N_12019,N_12056);
xnor U12292 (N_12292,N_12010,N_12147);
or U12293 (N_12293,N_12146,N_12002);
xor U12294 (N_12294,N_12137,N_12154);
nand U12295 (N_12295,N_12052,N_12131);
nor U12296 (N_12296,N_12145,N_12142);
nor U12297 (N_12297,N_12023,N_12106);
nor U12298 (N_12298,N_12040,N_12108);
nand U12299 (N_12299,N_12008,N_12035);
and U12300 (N_12300,N_12061,N_12020);
nand U12301 (N_12301,N_12089,N_12109);
and U12302 (N_12302,N_12079,N_12013);
nor U12303 (N_12303,N_12061,N_12098);
and U12304 (N_12304,N_12031,N_12131);
nand U12305 (N_12305,N_12123,N_12141);
nor U12306 (N_12306,N_12087,N_12023);
or U12307 (N_12307,N_12092,N_12133);
and U12308 (N_12308,N_12106,N_12054);
nor U12309 (N_12309,N_12087,N_12120);
nor U12310 (N_12310,N_12008,N_12101);
and U12311 (N_12311,N_12083,N_12032);
nand U12312 (N_12312,N_12075,N_12135);
nor U12313 (N_12313,N_12146,N_12025);
nand U12314 (N_12314,N_12032,N_12055);
xnor U12315 (N_12315,N_12020,N_12102);
nor U12316 (N_12316,N_12152,N_12047);
xor U12317 (N_12317,N_12080,N_12065);
nor U12318 (N_12318,N_12026,N_12146);
or U12319 (N_12319,N_12012,N_12097);
nor U12320 (N_12320,N_12265,N_12197);
nand U12321 (N_12321,N_12235,N_12192);
nor U12322 (N_12322,N_12285,N_12240);
nand U12323 (N_12323,N_12239,N_12252);
xor U12324 (N_12324,N_12180,N_12243);
xor U12325 (N_12325,N_12165,N_12225);
or U12326 (N_12326,N_12250,N_12266);
nand U12327 (N_12327,N_12164,N_12276);
or U12328 (N_12328,N_12217,N_12284);
nand U12329 (N_12329,N_12302,N_12220);
xnor U12330 (N_12330,N_12222,N_12189);
xor U12331 (N_12331,N_12274,N_12298);
xor U12332 (N_12332,N_12245,N_12186);
and U12333 (N_12333,N_12288,N_12241);
nor U12334 (N_12334,N_12292,N_12272);
nor U12335 (N_12335,N_12271,N_12261);
and U12336 (N_12336,N_12208,N_12234);
or U12337 (N_12337,N_12258,N_12167);
nor U12338 (N_12338,N_12256,N_12215);
or U12339 (N_12339,N_12269,N_12175);
xor U12340 (N_12340,N_12221,N_12238);
nor U12341 (N_12341,N_12228,N_12275);
nand U12342 (N_12342,N_12190,N_12198);
nor U12343 (N_12343,N_12178,N_12244);
or U12344 (N_12344,N_12211,N_12248);
or U12345 (N_12345,N_12204,N_12295);
xnor U12346 (N_12346,N_12308,N_12251);
xor U12347 (N_12347,N_12278,N_12316);
or U12348 (N_12348,N_12314,N_12277);
nand U12349 (N_12349,N_12296,N_12309);
nand U12350 (N_12350,N_12168,N_12199);
and U12351 (N_12351,N_12206,N_12160);
and U12352 (N_12352,N_12305,N_12306);
or U12353 (N_12353,N_12249,N_12286);
and U12354 (N_12354,N_12259,N_12182);
xor U12355 (N_12355,N_12268,N_12254);
nor U12356 (N_12356,N_12267,N_12231);
nand U12357 (N_12357,N_12227,N_12280);
and U12358 (N_12358,N_12303,N_12166);
or U12359 (N_12359,N_12290,N_12184);
nor U12360 (N_12360,N_12201,N_12287);
and U12361 (N_12361,N_12297,N_12226);
nand U12362 (N_12362,N_12171,N_12289);
and U12363 (N_12363,N_12179,N_12230);
and U12364 (N_12364,N_12181,N_12293);
and U12365 (N_12365,N_12279,N_12253);
nor U12366 (N_12366,N_12209,N_12205);
xnor U12367 (N_12367,N_12236,N_12216);
or U12368 (N_12368,N_12172,N_12237);
xor U12369 (N_12369,N_12273,N_12169);
xor U12370 (N_12370,N_12185,N_12299);
nand U12371 (N_12371,N_12247,N_12301);
or U12372 (N_12372,N_12317,N_12176);
nand U12373 (N_12373,N_12183,N_12213);
and U12374 (N_12374,N_12260,N_12257);
xnor U12375 (N_12375,N_12224,N_12218);
nor U12376 (N_12376,N_12310,N_12177);
xor U12377 (N_12377,N_12187,N_12307);
nand U12378 (N_12378,N_12262,N_12174);
nand U12379 (N_12379,N_12161,N_12202);
nor U12380 (N_12380,N_12313,N_12233);
xnor U12381 (N_12381,N_12200,N_12229);
and U12382 (N_12382,N_12194,N_12319);
and U12383 (N_12383,N_12173,N_12255);
nor U12384 (N_12384,N_12223,N_12212);
and U12385 (N_12385,N_12210,N_12219);
xor U12386 (N_12386,N_12191,N_12246);
and U12387 (N_12387,N_12315,N_12193);
xnor U12388 (N_12388,N_12300,N_12282);
nor U12389 (N_12389,N_12304,N_12195);
xnor U12390 (N_12390,N_12188,N_12170);
or U12391 (N_12391,N_12311,N_12291);
xor U12392 (N_12392,N_12163,N_12312);
nor U12393 (N_12393,N_12214,N_12263);
and U12394 (N_12394,N_12232,N_12270);
xnor U12395 (N_12395,N_12264,N_12203);
xor U12396 (N_12396,N_12207,N_12196);
and U12397 (N_12397,N_12242,N_12281);
nor U12398 (N_12398,N_12162,N_12283);
xor U12399 (N_12399,N_12318,N_12294);
xnor U12400 (N_12400,N_12236,N_12299);
xnor U12401 (N_12401,N_12166,N_12317);
xor U12402 (N_12402,N_12249,N_12167);
and U12403 (N_12403,N_12163,N_12194);
nor U12404 (N_12404,N_12297,N_12206);
and U12405 (N_12405,N_12214,N_12209);
and U12406 (N_12406,N_12228,N_12198);
nand U12407 (N_12407,N_12222,N_12297);
nor U12408 (N_12408,N_12247,N_12168);
xor U12409 (N_12409,N_12246,N_12170);
nor U12410 (N_12410,N_12257,N_12212);
nand U12411 (N_12411,N_12301,N_12180);
nor U12412 (N_12412,N_12221,N_12310);
or U12413 (N_12413,N_12220,N_12282);
nand U12414 (N_12414,N_12299,N_12295);
nand U12415 (N_12415,N_12291,N_12302);
nand U12416 (N_12416,N_12306,N_12250);
and U12417 (N_12417,N_12241,N_12194);
nor U12418 (N_12418,N_12185,N_12295);
nand U12419 (N_12419,N_12311,N_12304);
nor U12420 (N_12420,N_12239,N_12187);
or U12421 (N_12421,N_12308,N_12310);
and U12422 (N_12422,N_12167,N_12259);
or U12423 (N_12423,N_12214,N_12294);
nor U12424 (N_12424,N_12173,N_12183);
and U12425 (N_12425,N_12223,N_12259);
nor U12426 (N_12426,N_12228,N_12214);
nor U12427 (N_12427,N_12227,N_12303);
or U12428 (N_12428,N_12276,N_12242);
nand U12429 (N_12429,N_12195,N_12205);
xor U12430 (N_12430,N_12308,N_12276);
nor U12431 (N_12431,N_12316,N_12314);
or U12432 (N_12432,N_12311,N_12246);
or U12433 (N_12433,N_12266,N_12299);
nand U12434 (N_12434,N_12285,N_12207);
and U12435 (N_12435,N_12235,N_12225);
or U12436 (N_12436,N_12197,N_12168);
or U12437 (N_12437,N_12228,N_12309);
nand U12438 (N_12438,N_12174,N_12240);
or U12439 (N_12439,N_12204,N_12287);
or U12440 (N_12440,N_12168,N_12257);
or U12441 (N_12441,N_12283,N_12169);
nand U12442 (N_12442,N_12305,N_12273);
or U12443 (N_12443,N_12246,N_12212);
xnor U12444 (N_12444,N_12205,N_12161);
nand U12445 (N_12445,N_12222,N_12188);
or U12446 (N_12446,N_12272,N_12201);
nand U12447 (N_12447,N_12292,N_12246);
or U12448 (N_12448,N_12293,N_12206);
or U12449 (N_12449,N_12199,N_12273);
nor U12450 (N_12450,N_12255,N_12292);
nor U12451 (N_12451,N_12275,N_12196);
or U12452 (N_12452,N_12166,N_12275);
and U12453 (N_12453,N_12260,N_12211);
nand U12454 (N_12454,N_12180,N_12303);
nor U12455 (N_12455,N_12283,N_12263);
xnor U12456 (N_12456,N_12238,N_12318);
or U12457 (N_12457,N_12164,N_12214);
and U12458 (N_12458,N_12243,N_12236);
xnor U12459 (N_12459,N_12293,N_12310);
and U12460 (N_12460,N_12304,N_12193);
and U12461 (N_12461,N_12312,N_12280);
or U12462 (N_12462,N_12195,N_12295);
nor U12463 (N_12463,N_12241,N_12189);
or U12464 (N_12464,N_12308,N_12183);
and U12465 (N_12465,N_12272,N_12224);
and U12466 (N_12466,N_12217,N_12303);
xnor U12467 (N_12467,N_12272,N_12182);
nor U12468 (N_12468,N_12304,N_12222);
and U12469 (N_12469,N_12198,N_12187);
nand U12470 (N_12470,N_12233,N_12268);
nand U12471 (N_12471,N_12276,N_12292);
xor U12472 (N_12472,N_12283,N_12238);
xnor U12473 (N_12473,N_12216,N_12279);
and U12474 (N_12474,N_12258,N_12279);
nor U12475 (N_12475,N_12300,N_12268);
nor U12476 (N_12476,N_12225,N_12214);
nor U12477 (N_12477,N_12206,N_12214);
nor U12478 (N_12478,N_12314,N_12199);
xnor U12479 (N_12479,N_12213,N_12185);
and U12480 (N_12480,N_12351,N_12446);
and U12481 (N_12481,N_12366,N_12372);
xor U12482 (N_12482,N_12382,N_12399);
nand U12483 (N_12483,N_12473,N_12355);
nand U12484 (N_12484,N_12439,N_12468);
and U12485 (N_12485,N_12371,N_12367);
nor U12486 (N_12486,N_12411,N_12357);
nor U12487 (N_12487,N_12471,N_12341);
xor U12488 (N_12488,N_12417,N_12349);
or U12489 (N_12489,N_12356,N_12416);
or U12490 (N_12490,N_12458,N_12373);
xnor U12491 (N_12491,N_12470,N_12405);
xnor U12492 (N_12492,N_12377,N_12456);
nor U12493 (N_12493,N_12343,N_12453);
xor U12494 (N_12494,N_12395,N_12328);
and U12495 (N_12495,N_12323,N_12360);
xor U12496 (N_12496,N_12326,N_12332);
nor U12497 (N_12497,N_12379,N_12454);
nand U12498 (N_12498,N_12350,N_12472);
and U12499 (N_12499,N_12347,N_12440);
or U12500 (N_12500,N_12327,N_12346);
xnor U12501 (N_12501,N_12414,N_12422);
nor U12502 (N_12502,N_12428,N_12429);
nand U12503 (N_12503,N_12469,N_12370);
nor U12504 (N_12504,N_12400,N_12401);
and U12505 (N_12505,N_12434,N_12419);
and U12506 (N_12506,N_12352,N_12359);
xnor U12507 (N_12507,N_12410,N_12361);
or U12508 (N_12508,N_12435,N_12385);
xor U12509 (N_12509,N_12418,N_12375);
and U12510 (N_12510,N_12397,N_12477);
xor U12511 (N_12511,N_12386,N_12336);
xor U12512 (N_12512,N_12475,N_12461);
nor U12513 (N_12513,N_12450,N_12431);
or U12514 (N_12514,N_12369,N_12465);
xor U12515 (N_12515,N_12345,N_12476);
nor U12516 (N_12516,N_12427,N_12335);
and U12517 (N_12517,N_12398,N_12329);
or U12518 (N_12518,N_12449,N_12358);
and U12519 (N_12519,N_12415,N_12474);
xor U12520 (N_12520,N_12374,N_12325);
nand U12521 (N_12521,N_12437,N_12442);
nor U12522 (N_12522,N_12388,N_12333);
and U12523 (N_12523,N_12432,N_12334);
xor U12524 (N_12524,N_12365,N_12424);
or U12525 (N_12525,N_12354,N_12402);
nand U12526 (N_12526,N_12436,N_12479);
and U12527 (N_12527,N_12466,N_12451);
nor U12528 (N_12528,N_12324,N_12464);
xnor U12529 (N_12529,N_12421,N_12392);
nand U12530 (N_12530,N_12463,N_12452);
or U12531 (N_12531,N_12348,N_12447);
and U12532 (N_12532,N_12403,N_12404);
and U12533 (N_12533,N_12460,N_12390);
and U12534 (N_12534,N_12462,N_12467);
nor U12535 (N_12535,N_12406,N_12363);
nand U12536 (N_12536,N_12445,N_12455);
nor U12537 (N_12537,N_12407,N_12337);
and U12538 (N_12538,N_12430,N_12444);
nand U12539 (N_12539,N_12457,N_12433);
nor U12540 (N_12540,N_12443,N_12459);
nand U12541 (N_12541,N_12321,N_12441);
xor U12542 (N_12542,N_12340,N_12393);
nor U12543 (N_12543,N_12391,N_12420);
or U12544 (N_12544,N_12381,N_12426);
nand U12545 (N_12545,N_12322,N_12383);
nand U12546 (N_12546,N_12425,N_12364);
nor U12547 (N_12547,N_12413,N_12423);
and U12548 (N_12548,N_12378,N_12380);
nand U12549 (N_12549,N_12320,N_12389);
nand U12550 (N_12550,N_12330,N_12478);
nand U12551 (N_12551,N_12394,N_12331);
or U12552 (N_12552,N_12409,N_12338);
xnor U12553 (N_12553,N_12412,N_12344);
and U12554 (N_12554,N_12387,N_12342);
or U12555 (N_12555,N_12368,N_12438);
and U12556 (N_12556,N_12339,N_12376);
xor U12557 (N_12557,N_12408,N_12384);
nand U12558 (N_12558,N_12396,N_12448);
xor U12559 (N_12559,N_12362,N_12353);
xor U12560 (N_12560,N_12468,N_12436);
and U12561 (N_12561,N_12370,N_12372);
nor U12562 (N_12562,N_12390,N_12388);
or U12563 (N_12563,N_12409,N_12479);
xnor U12564 (N_12564,N_12474,N_12344);
nand U12565 (N_12565,N_12384,N_12357);
xnor U12566 (N_12566,N_12429,N_12385);
nand U12567 (N_12567,N_12339,N_12379);
xnor U12568 (N_12568,N_12424,N_12417);
or U12569 (N_12569,N_12399,N_12355);
nand U12570 (N_12570,N_12381,N_12460);
nor U12571 (N_12571,N_12380,N_12365);
nand U12572 (N_12572,N_12348,N_12339);
nor U12573 (N_12573,N_12402,N_12364);
and U12574 (N_12574,N_12395,N_12475);
or U12575 (N_12575,N_12445,N_12419);
and U12576 (N_12576,N_12383,N_12375);
xnor U12577 (N_12577,N_12352,N_12431);
xor U12578 (N_12578,N_12403,N_12418);
nor U12579 (N_12579,N_12378,N_12385);
nand U12580 (N_12580,N_12467,N_12457);
nand U12581 (N_12581,N_12438,N_12379);
nor U12582 (N_12582,N_12410,N_12429);
nor U12583 (N_12583,N_12446,N_12321);
nor U12584 (N_12584,N_12479,N_12355);
xor U12585 (N_12585,N_12465,N_12459);
nor U12586 (N_12586,N_12456,N_12330);
xor U12587 (N_12587,N_12473,N_12366);
nor U12588 (N_12588,N_12412,N_12336);
and U12589 (N_12589,N_12470,N_12379);
and U12590 (N_12590,N_12477,N_12471);
nand U12591 (N_12591,N_12396,N_12380);
and U12592 (N_12592,N_12385,N_12361);
nor U12593 (N_12593,N_12470,N_12466);
and U12594 (N_12594,N_12374,N_12415);
nand U12595 (N_12595,N_12433,N_12337);
nor U12596 (N_12596,N_12408,N_12415);
nand U12597 (N_12597,N_12412,N_12463);
xnor U12598 (N_12598,N_12381,N_12422);
and U12599 (N_12599,N_12457,N_12431);
nor U12600 (N_12600,N_12383,N_12417);
nand U12601 (N_12601,N_12424,N_12372);
xnor U12602 (N_12602,N_12332,N_12327);
nor U12603 (N_12603,N_12430,N_12321);
nor U12604 (N_12604,N_12343,N_12424);
nor U12605 (N_12605,N_12385,N_12390);
and U12606 (N_12606,N_12468,N_12336);
xnor U12607 (N_12607,N_12326,N_12380);
and U12608 (N_12608,N_12337,N_12392);
or U12609 (N_12609,N_12370,N_12418);
nor U12610 (N_12610,N_12393,N_12362);
and U12611 (N_12611,N_12397,N_12385);
and U12612 (N_12612,N_12373,N_12438);
nor U12613 (N_12613,N_12431,N_12356);
nor U12614 (N_12614,N_12437,N_12335);
and U12615 (N_12615,N_12334,N_12426);
xnor U12616 (N_12616,N_12327,N_12347);
nand U12617 (N_12617,N_12418,N_12451);
nand U12618 (N_12618,N_12466,N_12322);
nor U12619 (N_12619,N_12326,N_12446);
xor U12620 (N_12620,N_12462,N_12322);
nor U12621 (N_12621,N_12323,N_12445);
nand U12622 (N_12622,N_12432,N_12346);
xor U12623 (N_12623,N_12474,N_12328);
or U12624 (N_12624,N_12366,N_12347);
nor U12625 (N_12625,N_12392,N_12474);
or U12626 (N_12626,N_12394,N_12440);
nand U12627 (N_12627,N_12349,N_12422);
and U12628 (N_12628,N_12373,N_12380);
xnor U12629 (N_12629,N_12348,N_12382);
xor U12630 (N_12630,N_12455,N_12324);
and U12631 (N_12631,N_12354,N_12406);
xnor U12632 (N_12632,N_12411,N_12344);
nor U12633 (N_12633,N_12382,N_12448);
or U12634 (N_12634,N_12402,N_12347);
nor U12635 (N_12635,N_12368,N_12349);
nor U12636 (N_12636,N_12359,N_12338);
nand U12637 (N_12637,N_12384,N_12468);
xnor U12638 (N_12638,N_12469,N_12452);
or U12639 (N_12639,N_12395,N_12321);
nor U12640 (N_12640,N_12571,N_12581);
and U12641 (N_12641,N_12619,N_12558);
nor U12642 (N_12642,N_12491,N_12639);
nand U12643 (N_12643,N_12624,N_12503);
nor U12644 (N_12644,N_12511,N_12485);
and U12645 (N_12645,N_12500,N_12528);
or U12646 (N_12646,N_12609,N_12494);
nor U12647 (N_12647,N_12541,N_12549);
nor U12648 (N_12648,N_12622,N_12554);
nor U12649 (N_12649,N_12506,N_12516);
nor U12650 (N_12650,N_12623,N_12557);
or U12651 (N_12651,N_12522,N_12498);
nand U12652 (N_12652,N_12590,N_12493);
xnor U12653 (N_12653,N_12533,N_12607);
nand U12654 (N_12654,N_12556,N_12602);
nand U12655 (N_12655,N_12605,N_12582);
or U12656 (N_12656,N_12538,N_12489);
and U12657 (N_12657,N_12534,N_12548);
nand U12658 (N_12658,N_12614,N_12637);
and U12659 (N_12659,N_12560,N_12501);
or U12660 (N_12660,N_12536,N_12518);
nand U12661 (N_12661,N_12540,N_12564);
and U12662 (N_12662,N_12603,N_12630);
nand U12663 (N_12663,N_12600,N_12562);
and U12664 (N_12664,N_12569,N_12632);
nor U12665 (N_12665,N_12591,N_12559);
nand U12666 (N_12666,N_12525,N_12589);
or U12667 (N_12667,N_12596,N_12505);
xnor U12668 (N_12668,N_12545,N_12551);
or U12669 (N_12669,N_12620,N_12484);
xnor U12670 (N_12670,N_12553,N_12612);
and U12671 (N_12671,N_12574,N_12509);
nor U12672 (N_12672,N_12585,N_12629);
xnor U12673 (N_12673,N_12520,N_12628);
or U12674 (N_12674,N_12544,N_12586);
nand U12675 (N_12675,N_12576,N_12572);
and U12676 (N_12676,N_12508,N_12567);
xor U12677 (N_12677,N_12561,N_12626);
xnor U12678 (N_12678,N_12621,N_12584);
and U12679 (N_12679,N_12552,N_12601);
or U12680 (N_12680,N_12532,N_12555);
nand U12681 (N_12681,N_12578,N_12638);
nor U12682 (N_12682,N_12517,N_12502);
nor U12683 (N_12683,N_12481,N_12593);
and U12684 (N_12684,N_12592,N_12529);
or U12685 (N_12685,N_12595,N_12631);
and U12686 (N_12686,N_12539,N_12570);
nor U12687 (N_12687,N_12610,N_12537);
nor U12688 (N_12688,N_12566,N_12483);
nor U12689 (N_12689,N_12627,N_12636);
or U12690 (N_12690,N_12594,N_12634);
and U12691 (N_12691,N_12521,N_12512);
nor U12692 (N_12692,N_12615,N_12526);
or U12693 (N_12693,N_12496,N_12568);
xor U12694 (N_12694,N_12499,N_12515);
nand U12695 (N_12695,N_12507,N_12514);
nor U12696 (N_12696,N_12523,N_12598);
or U12697 (N_12697,N_12606,N_12575);
nand U12698 (N_12698,N_12563,N_12577);
nor U12699 (N_12699,N_12611,N_12482);
xnor U12700 (N_12700,N_12490,N_12604);
nor U12701 (N_12701,N_12542,N_12492);
and U12702 (N_12702,N_12488,N_12599);
xnor U12703 (N_12703,N_12519,N_12486);
nand U12704 (N_12704,N_12613,N_12547);
xnor U12705 (N_12705,N_12580,N_12497);
and U12706 (N_12706,N_12487,N_12583);
nor U12707 (N_12707,N_12617,N_12531);
or U12708 (N_12708,N_12510,N_12480);
and U12709 (N_12709,N_12530,N_12543);
or U12710 (N_12710,N_12625,N_12546);
and U12711 (N_12711,N_12579,N_12527);
nand U12712 (N_12712,N_12573,N_12616);
or U12713 (N_12713,N_12504,N_12495);
nand U12714 (N_12714,N_12635,N_12618);
and U12715 (N_12715,N_12550,N_12524);
nor U12716 (N_12716,N_12608,N_12597);
and U12717 (N_12717,N_12633,N_12535);
and U12718 (N_12718,N_12588,N_12513);
or U12719 (N_12719,N_12587,N_12565);
nand U12720 (N_12720,N_12565,N_12624);
nor U12721 (N_12721,N_12517,N_12599);
xnor U12722 (N_12722,N_12562,N_12561);
and U12723 (N_12723,N_12593,N_12615);
and U12724 (N_12724,N_12550,N_12492);
nor U12725 (N_12725,N_12482,N_12486);
nand U12726 (N_12726,N_12516,N_12480);
nor U12727 (N_12727,N_12530,N_12604);
nand U12728 (N_12728,N_12557,N_12523);
xnor U12729 (N_12729,N_12503,N_12616);
or U12730 (N_12730,N_12525,N_12562);
nand U12731 (N_12731,N_12570,N_12536);
or U12732 (N_12732,N_12590,N_12631);
nand U12733 (N_12733,N_12505,N_12528);
xor U12734 (N_12734,N_12625,N_12560);
nor U12735 (N_12735,N_12564,N_12620);
or U12736 (N_12736,N_12499,N_12557);
and U12737 (N_12737,N_12538,N_12555);
or U12738 (N_12738,N_12606,N_12528);
or U12739 (N_12739,N_12521,N_12622);
nand U12740 (N_12740,N_12595,N_12523);
nor U12741 (N_12741,N_12481,N_12516);
or U12742 (N_12742,N_12539,N_12523);
and U12743 (N_12743,N_12639,N_12603);
nor U12744 (N_12744,N_12577,N_12592);
and U12745 (N_12745,N_12587,N_12581);
and U12746 (N_12746,N_12624,N_12481);
or U12747 (N_12747,N_12530,N_12524);
xnor U12748 (N_12748,N_12512,N_12562);
and U12749 (N_12749,N_12623,N_12510);
nor U12750 (N_12750,N_12485,N_12482);
xnor U12751 (N_12751,N_12636,N_12492);
or U12752 (N_12752,N_12613,N_12605);
nand U12753 (N_12753,N_12580,N_12583);
nand U12754 (N_12754,N_12546,N_12529);
or U12755 (N_12755,N_12619,N_12499);
xnor U12756 (N_12756,N_12527,N_12542);
xor U12757 (N_12757,N_12631,N_12573);
nand U12758 (N_12758,N_12621,N_12556);
nor U12759 (N_12759,N_12550,N_12521);
or U12760 (N_12760,N_12594,N_12480);
nand U12761 (N_12761,N_12483,N_12527);
nor U12762 (N_12762,N_12559,N_12602);
xnor U12763 (N_12763,N_12543,N_12519);
xnor U12764 (N_12764,N_12619,N_12497);
xor U12765 (N_12765,N_12533,N_12518);
nand U12766 (N_12766,N_12546,N_12632);
or U12767 (N_12767,N_12609,N_12525);
nand U12768 (N_12768,N_12490,N_12538);
and U12769 (N_12769,N_12489,N_12602);
nor U12770 (N_12770,N_12569,N_12611);
and U12771 (N_12771,N_12560,N_12549);
xor U12772 (N_12772,N_12638,N_12569);
xnor U12773 (N_12773,N_12506,N_12482);
nand U12774 (N_12774,N_12616,N_12635);
nand U12775 (N_12775,N_12561,N_12525);
xnor U12776 (N_12776,N_12522,N_12512);
or U12777 (N_12777,N_12624,N_12492);
nand U12778 (N_12778,N_12611,N_12605);
nand U12779 (N_12779,N_12537,N_12523);
nor U12780 (N_12780,N_12619,N_12549);
or U12781 (N_12781,N_12515,N_12529);
and U12782 (N_12782,N_12583,N_12557);
and U12783 (N_12783,N_12607,N_12593);
nor U12784 (N_12784,N_12631,N_12568);
or U12785 (N_12785,N_12578,N_12532);
and U12786 (N_12786,N_12619,N_12548);
nand U12787 (N_12787,N_12577,N_12508);
xnor U12788 (N_12788,N_12516,N_12555);
nand U12789 (N_12789,N_12585,N_12567);
nand U12790 (N_12790,N_12586,N_12569);
or U12791 (N_12791,N_12489,N_12617);
nand U12792 (N_12792,N_12564,N_12627);
xor U12793 (N_12793,N_12525,N_12513);
nand U12794 (N_12794,N_12486,N_12621);
xor U12795 (N_12795,N_12582,N_12560);
xor U12796 (N_12796,N_12558,N_12523);
or U12797 (N_12797,N_12622,N_12624);
or U12798 (N_12798,N_12496,N_12561);
and U12799 (N_12799,N_12606,N_12577);
nor U12800 (N_12800,N_12683,N_12763);
nand U12801 (N_12801,N_12708,N_12647);
xor U12802 (N_12802,N_12688,N_12640);
nor U12803 (N_12803,N_12723,N_12744);
xnor U12804 (N_12804,N_12690,N_12650);
or U12805 (N_12805,N_12715,N_12768);
or U12806 (N_12806,N_12746,N_12652);
nor U12807 (N_12807,N_12783,N_12782);
or U12808 (N_12808,N_12656,N_12777);
and U12809 (N_12809,N_12753,N_12681);
nor U12810 (N_12810,N_12734,N_12790);
or U12811 (N_12811,N_12685,N_12674);
or U12812 (N_12812,N_12743,N_12761);
nor U12813 (N_12813,N_12731,N_12717);
nor U12814 (N_12814,N_12646,N_12781);
nand U12815 (N_12815,N_12742,N_12795);
or U12816 (N_12816,N_12691,N_12778);
xnor U12817 (N_12817,N_12721,N_12735);
and U12818 (N_12818,N_12658,N_12798);
nand U12819 (N_12819,N_12724,N_12752);
xor U12820 (N_12820,N_12707,N_12668);
nand U12821 (N_12821,N_12712,N_12667);
or U12822 (N_12822,N_12722,N_12703);
nand U12823 (N_12823,N_12706,N_12695);
nor U12824 (N_12824,N_12792,N_12678);
or U12825 (N_12825,N_12769,N_12787);
xor U12826 (N_12826,N_12726,N_12755);
or U12827 (N_12827,N_12740,N_12728);
and U12828 (N_12828,N_12758,N_12682);
and U12829 (N_12829,N_12770,N_12757);
and U12830 (N_12830,N_12654,N_12732);
xor U12831 (N_12831,N_12775,N_12672);
nor U12832 (N_12832,N_12747,N_12750);
nand U12833 (N_12833,N_12791,N_12694);
xor U12834 (N_12834,N_12796,N_12642);
and U12835 (N_12835,N_12680,N_12754);
or U12836 (N_12836,N_12705,N_12733);
xor U12837 (N_12837,N_12710,N_12711);
nor U12838 (N_12838,N_12773,N_12725);
or U12839 (N_12839,N_12786,N_12692);
nand U12840 (N_12840,N_12739,N_12756);
xor U12841 (N_12841,N_12762,N_12797);
nor U12842 (N_12842,N_12716,N_12669);
or U12843 (N_12843,N_12749,N_12702);
nand U12844 (N_12844,N_12727,N_12697);
and U12845 (N_12845,N_12675,N_12799);
nor U12846 (N_12846,N_12663,N_12779);
and U12847 (N_12847,N_12774,N_12693);
xor U12848 (N_12848,N_12655,N_12671);
and U12849 (N_12849,N_12748,N_12643);
xnor U12850 (N_12850,N_12745,N_12696);
or U12851 (N_12851,N_12771,N_12653);
nand U12852 (N_12852,N_12730,N_12673);
or U12853 (N_12853,N_12662,N_12718);
or U12854 (N_12854,N_12659,N_12741);
and U12855 (N_12855,N_12641,N_12666);
nor U12856 (N_12856,N_12785,N_12736);
nand U12857 (N_12857,N_12737,N_12660);
and U12858 (N_12858,N_12767,N_12676);
xnor U12859 (N_12859,N_12719,N_12665);
and U12860 (N_12860,N_12714,N_12686);
xnor U12861 (N_12861,N_12729,N_12764);
and U12862 (N_12862,N_12765,N_12793);
and U12863 (N_12863,N_12794,N_12709);
xnor U12864 (N_12864,N_12766,N_12684);
nor U12865 (N_12865,N_12772,N_12699);
or U12866 (N_12866,N_12644,N_12645);
nor U12867 (N_12867,N_12784,N_12657);
and U12868 (N_12868,N_12738,N_12664);
nor U12869 (N_12869,N_12651,N_12780);
and U12870 (N_12870,N_12649,N_12698);
or U12871 (N_12871,N_12700,N_12670);
nand U12872 (N_12872,N_12713,N_12677);
nand U12873 (N_12873,N_12661,N_12759);
nor U12874 (N_12874,N_12704,N_12776);
or U12875 (N_12875,N_12760,N_12687);
nand U12876 (N_12876,N_12751,N_12788);
nor U12877 (N_12877,N_12720,N_12648);
and U12878 (N_12878,N_12701,N_12679);
nor U12879 (N_12879,N_12689,N_12789);
nor U12880 (N_12880,N_12734,N_12700);
or U12881 (N_12881,N_12679,N_12771);
nor U12882 (N_12882,N_12641,N_12722);
nor U12883 (N_12883,N_12771,N_12680);
nand U12884 (N_12884,N_12793,N_12680);
or U12885 (N_12885,N_12641,N_12646);
or U12886 (N_12886,N_12718,N_12680);
nand U12887 (N_12887,N_12750,N_12684);
or U12888 (N_12888,N_12765,N_12743);
nand U12889 (N_12889,N_12794,N_12697);
or U12890 (N_12890,N_12687,N_12771);
and U12891 (N_12891,N_12706,N_12736);
nor U12892 (N_12892,N_12799,N_12658);
nand U12893 (N_12893,N_12762,N_12720);
xor U12894 (N_12894,N_12717,N_12775);
or U12895 (N_12895,N_12762,N_12651);
or U12896 (N_12896,N_12689,N_12703);
or U12897 (N_12897,N_12650,N_12642);
nand U12898 (N_12898,N_12653,N_12795);
and U12899 (N_12899,N_12669,N_12762);
and U12900 (N_12900,N_12725,N_12684);
nand U12901 (N_12901,N_12684,N_12694);
nand U12902 (N_12902,N_12797,N_12793);
and U12903 (N_12903,N_12789,N_12702);
xnor U12904 (N_12904,N_12656,N_12696);
nor U12905 (N_12905,N_12650,N_12781);
nor U12906 (N_12906,N_12767,N_12752);
or U12907 (N_12907,N_12650,N_12732);
nor U12908 (N_12908,N_12762,N_12649);
xor U12909 (N_12909,N_12765,N_12795);
xnor U12910 (N_12910,N_12760,N_12654);
and U12911 (N_12911,N_12741,N_12692);
xnor U12912 (N_12912,N_12693,N_12650);
xor U12913 (N_12913,N_12669,N_12706);
and U12914 (N_12914,N_12767,N_12757);
xor U12915 (N_12915,N_12754,N_12649);
and U12916 (N_12916,N_12701,N_12654);
and U12917 (N_12917,N_12709,N_12745);
and U12918 (N_12918,N_12734,N_12786);
or U12919 (N_12919,N_12678,N_12743);
nor U12920 (N_12920,N_12642,N_12719);
nor U12921 (N_12921,N_12686,N_12789);
or U12922 (N_12922,N_12679,N_12732);
nand U12923 (N_12923,N_12782,N_12701);
xnor U12924 (N_12924,N_12790,N_12791);
and U12925 (N_12925,N_12761,N_12784);
nand U12926 (N_12926,N_12799,N_12651);
xnor U12927 (N_12927,N_12684,N_12772);
or U12928 (N_12928,N_12782,N_12697);
nand U12929 (N_12929,N_12701,N_12675);
and U12930 (N_12930,N_12732,N_12757);
xnor U12931 (N_12931,N_12650,N_12771);
or U12932 (N_12932,N_12681,N_12790);
and U12933 (N_12933,N_12668,N_12792);
or U12934 (N_12934,N_12728,N_12763);
or U12935 (N_12935,N_12659,N_12701);
or U12936 (N_12936,N_12738,N_12742);
or U12937 (N_12937,N_12672,N_12793);
or U12938 (N_12938,N_12681,N_12654);
or U12939 (N_12939,N_12684,N_12668);
nand U12940 (N_12940,N_12777,N_12688);
nand U12941 (N_12941,N_12654,N_12796);
nor U12942 (N_12942,N_12691,N_12768);
nand U12943 (N_12943,N_12642,N_12739);
nor U12944 (N_12944,N_12662,N_12755);
nor U12945 (N_12945,N_12710,N_12796);
xnor U12946 (N_12946,N_12764,N_12728);
nor U12947 (N_12947,N_12776,N_12700);
or U12948 (N_12948,N_12692,N_12769);
and U12949 (N_12949,N_12671,N_12776);
nor U12950 (N_12950,N_12699,N_12659);
and U12951 (N_12951,N_12696,N_12731);
xnor U12952 (N_12952,N_12658,N_12711);
or U12953 (N_12953,N_12723,N_12677);
nor U12954 (N_12954,N_12756,N_12762);
nand U12955 (N_12955,N_12691,N_12645);
and U12956 (N_12956,N_12686,N_12706);
xnor U12957 (N_12957,N_12763,N_12748);
and U12958 (N_12958,N_12650,N_12687);
or U12959 (N_12959,N_12777,N_12660);
nand U12960 (N_12960,N_12834,N_12850);
and U12961 (N_12961,N_12915,N_12955);
nand U12962 (N_12962,N_12932,N_12909);
xnor U12963 (N_12963,N_12865,N_12847);
nand U12964 (N_12964,N_12935,N_12947);
or U12965 (N_12965,N_12950,N_12958);
nand U12966 (N_12966,N_12824,N_12877);
xnor U12967 (N_12967,N_12867,N_12807);
or U12968 (N_12968,N_12891,N_12871);
or U12969 (N_12969,N_12884,N_12885);
and U12970 (N_12970,N_12904,N_12878);
and U12971 (N_12971,N_12908,N_12822);
or U12972 (N_12972,N_12920,N_12945);
nand U12973 (N_12973,N_12811,N_12954);
and U12974 (N_12974,N_12952,N_12846);
nand U12975 (N_12975,N_12889,N_12874);
xnor U12976 (N_12976,N_12845,N_12859);
xor U12977 (N_12977,N_12911,N_12857);
and U12978 (N_12978,N_12815,N_12886);
and U12979 (N_12979,N_12821,N_12808);
and U12980 (N_12980,N_12882,N_12870);
nand U12981 (N_12981,N_12829,N_12812);
xnor U12982 (N_12982,N_12910,N_12906);
or U12983 (N_12983,N_12901,N_12931);
nand U12984 (N_12984,N_12861,N_12890);
nand U12985 (N_12985,N_12835,N_12925);
and U12986 (N_12986,N_12875,N_12905);
and U12987 (N_12987,N_12802,N_12848);
nor U12988 (N_12988,N_12862,N_12953);
and U12989 (N_12989,N_12959,N_12948);
and U12990 (N_12990,N_12839,N_12881);
and U12991 (N_12991,N_12926,N_12898);
nand U12992 (N_12992,N_12918,N_12844);
or U12993 (N_12993,N_12903,N_12944);
xor U12994 (N_12994,N_12856,N_12826);
nand U12995 (N_12995,N_12924,N_12809);
xor U12996 (N_12996,N_12817,N_12912);
nor U12997 (N_12997,N_12827,N_12917);
and U12998 (N_12998,N_12810,N_12853);
nor U12999 (N_12999,N_12818,N_12836);
nand U13000 (N_13000,N_12900,N_12921);
nand U13001 (N_13001,N_12940,N_12951);
nor U13002 (N_13002,N_12893,N_12914);
or U13003 (N_13003,N_12831,N_12928);
xor U13004 (N_13004,N_12828,N_12896);
xnor U13005 (N_13005,N_12942,N_12816);
and U13006 (N_13006,N_12841,N_12883);
xnor U13007 (N_13007,N_12800,N_12840);
xor U13008 (N_13008,N_12838,N_12919);
xnor U13009 (N_13009,N_12860,N_12927);
xnor U13010 (N_13010,N_12814,N_12879);
xor U13011 (N_13011,N_12922,N_12813);
nand U13012 (N_13012,N_12923,N_12902);
nor U13013 (N_13013,N_12897,N_12820);
or U13014 (N_13014,N_12849,N_12837);
and U13015 (N_13015,N_12843,N_12933);
and U13016 (N_13016,N_12852,N_12936);
nand U13017 (N_13017,N_12916,N_12866);
or U13018 (N_13018,N_12823,N_12899);
or U13019 (N_13019,N_12880,N_12876);
and U13020 (N_13020,N_12949,N_12832);
nor U13021 (N_13021,N_12842,N_12872);
and U13022 (N_13022,N_12851,N_12819);
xor U13023 (N_13023,N_12907,N_12863);
xor U13024 (N_13024,N_12854,N_12869);
nand U13025 (N_13025,N_12892,N_12868);
and U13026 (N_13026,N_12946,N_12833);
nor U13027 (N_13027,N_12894,N_12806);
or U13028 (N_13028,N_12930,N_12858);
or U13029 (N_13029,N_12803,N_12938);
and U13030 (N_13030,N_12830,N_12804);
or U13031 (N_13031,N_12873,N_12929);
xnor U13032 (N_13032,N_12855,N_12887);
xor U13033 (N_13033,N_12913,N_12939);
nor U13034 (N_13034,N_12805,N_12801);
nor U13035 (N_13035,N_12957,N_12895);
nor U13036 (N_13036,N_12888,N_12956);
nor U13037 (N_13037,N_12943,N_12934);
nor U13038 (N_13038,N_12864,N_12825);
and U13039 (N_13039,N_12937,N_12941);
or U13040 (N_13040,N_12930,N_12879);
or U13041 (N_13041,N_12901,N_12922);
or U13042 (N_13042,N_12934,N_12833);
and U13043 (N_13043,N_12884,N_12939);
or U13044 (N_13044,N_12901,N_12804);
and U13045 (N_13045,N_12891,N_12845);
nand U13046 (N_13046,N_12810,N_12873);
nor U13047 (N_13047,N_12835,N_12933);
or U13048 (N_13048,N_12888,N_12903);
xnor U13049 (N_13049,N_12807,N_12873);
nand U13050 (N_13050,N_12922,N_12893);
nor U13051 (N_13051,N_12848,N_12860);
nor U13052 (N_13052,N_12836,N_12865);
and U13053 (N_13053,N_12913,N_12883);
xor U13054 (N_13054,N_12909,N_12921);
nor U13055 (N_13055,N_12879,N_12822);
and U13056 (N_13056,N_12811,N_12846);
nand U13057 (N_13057,N_12800,N_12929);
and U13058 (N_13058,N_12837,N_12935);
nand U13059 (N_13059,N_12942,N_12862);
nor U13060 (N_13060,N_12800,N_12889);
xor U13061 (N_13061,N_12940,N_12922);
nor U13062 (N_13062,N_12860,N_12856);
nor U13063 (N_13063,N_12900,N_12865);
nand U13064 (N_13064,N_12931,N_12842);
xor U13065 (N_13065,N_12955,N_12834);
xnor U13066 (N_13066,N_12878,N_12836);
xor U13067 (N_13067,N_12908,N_12947);
or U13068 (N_13068,N_12895,N_12942);
nor U13069 (N_13069,N_12947,N_12813);
nor U13070 (N_13070,N_12844,N_12932);
nor U13071 (N_13071,N_12837,N_12865);
and U13072 (N_13072,N_12836,N_12869);
nand U13073 (N_13073,N_12955,N_12950);
nand U13074 (N_13074,N_12906,N_12823);
or U13075 (N_13075,N_12897,N_12836);
or U13076 (N_13076,N_12953,N_12801);
xnor U13077 (N_13077,N_12827,N_12825);
or U13078 (N_13078,N_12939,N_12908);
nor U13079 (N_13079,N_12956,N_12926);
or U13080 (N_13080,N_12873,N_12865);
nor U13081 (N_13081,N_12810,N_12901);
nand U13082 (N_13082,N_12830,N_12821);
nor U13083 (N_13083,N_12844,N_12955);
or U13084 (N_13084,N_12820,N_12873);
nand U13085 (N_13085,N_12894,N_12924);
and U13086 (N_13086,N_12889,N_12896);
nand U13087 (N_13087,N_12859,N_12906);
nand U13088 (N_13088,N_12916,N_12873);
nand U13089 (N_13089,N_12845,N_12912);
or U13090 (N_13090,N_12854,N_12846);
xnor U13091 (N_13091,N_12848,N_12862);
nand U13092 (N_13092,N_12877,N_12815);
or U13093 (N_13093,N_12865,N_12933);
nor U13094 (N_13094,N_12954,N_12912);
nand U13095 (N_13095,N_12826,N_12847);
nand U13096 (N_13096,N_12956,N_12892);
nor U13097 (N_13097,N_12870,N_12957);
nand U13098 (N_13098,N_12907,N_12866);
nand U13099 (N_13099,N_12945,N_12805);
xnor U13100 (N_13100,N_12929,N_12801);
nor U13101 (N_13101,N_12878,N_12807);
nor U13102 (N_13102,N_12881,N_12944);
or U13103 (N_13103,N_12933,N_12847);
xor U13104 (N_13104,N_12857,N_12950);
and U13105 (N_13105,N_12903,N_12851);
or U13106 (N_13106,N_12919,N_12934);
nor U13107 (N_13107,N_12914,N_12857);
nand U13108 (N_13108,N_12903,N_12905);
nor U13109 (N_13109,N_12852,N_12801);
nor U13110 (N_13110,N_12871,N_12920);
xor U13111 (N_13111,N_12935,N_12930);
nor U13112 (N_13112,N_12832,N_12815);
xnor U13113 (N_13113,N_12893,N_12821);
nor U13114 (N_13114,N_12827,N_12847);
xor U13115 (N_13115,N_12900,N_12878);
or U13116 (N_13116,N_12921,N_12870);
or U13117 (N_13117,N_12954,N_12808);
nor U13118 (N_13118,N_12843,N_12899);
or U13119 (N_13119,N_12927,N_12895);
or U13120 (N_13120,N_13056,N_13030);
or U13121 (N_13121,N_13067,N_13042);
or U13122 (N_13122,N_13084,N_13105);
or U13123 (N_13123,N_12980,N_12976);
or U13124 (N_13124,N_13029,N_13046);
xor U13125 (N_13125,N_13111,N_13022);
nand U13126 (N_13126,N_13043,N_13002);
and U13127 (N_13127,N_13109,N_13061);
nor U13128 (N_13128,N_13076,N_13013);
and U13129 (N_13129,N_13009,N_13048);
xor U13130 (N_13130,N_13008,N_13086);
nand U13131 (N_13131,N_13017,N_13071);
and U13132 (N_13132,N_13080,N_13090);
nor U13133 (N_13133,N_13110,N_12983);
nand U13134 (N_13134,N_13024,N_13023);
or U13135 (N_13135,N_13005,N_13102);
and U13136 (N_13136,N_12993,N_13052);
or U13137 (N_13137,N_13100,N_13053);
xnor U13138 (N_13138,N_13000,N_13117);
or U13139 (N_13139,N_13108,N_12988);
nor U13140 (N_13140,N_12984,N_13055);
xor U13141 (N_13141,N_13088,N_12973);
nor U13142 (N_13142,N_12977,N_13116);
nand U13143 (N_13143,N_12979,N_13031);
nor U13144 (N_13144,N_12974,N_13113);
and U13145 (N_13145,N_13097,N_13092);
xor U13146 (N_13146,N_13025,N_13119);
nor U13147 (N_13147,N_13021,N_13035);
and U13148 (N_13148,N_13107,N_13037);
xor U13149 (N_13149,N_13099,N_13003);
nor U13150 (N_13150,N_13041,N_13065);
nand U13151 (N_13151,N_12961,N_13094);
nand U13152 (N_13152,N_13103,N_13077);
and U13153 (N_13153,N_13089,N_13069);
and U13154 (N_13154,N_12964,N_12998);
xor U13155 (N_13155,N_12978,N_12986);
nand U13156 (N_13156,N_13034,N_12997);
and U13157 (N_13157,N_13057,N_13016);
nand U13158 (N_13158,N_12991,N_12989);
and U13159 (N_13159,N_13106,N_13033);
and U13160 (N_13160,N_13078,N_13020);
nand U13161 (N_13161,N_13040,N_13087);
and U13162 (N_13162,N_13091,N_13051);
nor U13163 (N_13163,N_13012,N_13060);
or U13164 (N_13164,N_13032,N_13028);
or U13165 (N_13165,N_13112,N_12970);
nand U13166 (N_13166,N_13081,N_13049);
or U13167 (N_13167,N_13050,N_13072);
nand U13168 (N_13168,N_13019,N_13014);
or U13169 (N_13169,N_12963,N_13114);
nor U13170 (N_13170,N_12967,N_13026);
xnor U13171 (N_13171,N_12965,N_13007);
xor U13172 (N_13172,N_12982,N_13073);
nor U13173 (N_13173,N_13018,N_13079);
xnor U13174 (N_13174,N_13068,N_13064);
nand U13175 (N_13175,N_13095,N_13085);
nand U13176 (N_13176,N_13010,N_12972);
nand U13177 (N_13177,N_12996,N_13006);
or U13178 (N_13178,N_12960,N_13038);
and U13179 (N_13179,N_13066,N_13044);
and U13180 (N_13180,N_13054,N_12971);
nand U13181 (N_13181,N_13075,N_13083);
nand U13182 (N_13182,N_12985,N_12990);
xnor U13183 (N_13183,N_12992,N_13045);
xnor U13184 (N_13184,N_12975,N_13039);
or U13185 (N_13185,N_12994,N_13101);
xnor U13186 (N_13186,N_12968,N_13063);
or U13187 (N_13187,N_12966,N_13001);
nor U13188 (N_13188,N_12962,N_12981);
or U13189 (N_13189,N_12987,N_13062);
and U13190 (N_13190,N_13098,N_13082);
or U13191 (N_13191,N_13011,N_13115);
or U13192 (N_13192,N_13074,N_13104);
and U13193 (N_13193,N_13036,N_13027);
nand U13194 (N_13194,N_12969,N_13015);
and U13195 (N_13195,N_13070,N_13059);
and U13196 (N_13196,N_12999,N_13047);
nor U13197 (N_13197,N_12995,N_13096);
and U13198 (N_13198,N_13093,N_13004);
and U13199 (N_13199,N_13058,N_13118);
and U13200 (N_13200,N_13024,N_13114);
nand U13201 (N_13201,N_13061,N_13009);
or U13202 (N_13202,N_13079,N_12971);
or U13203 (N_13203,N_13006,N_13095);
nor U13204 (N_13204,N_13014,N_13034);
and U13205 (N_13205,N_13043,N_13073);
and U13206 (N_13206,N_13047,N_12967);
xor U13207 (N_13207,N_13077,N_13020);
xnor U13208 (N_13208,N_13092,N_13028);
xor U13209 (N_13209,N_13076,N_13073);
xor U13210 (N_13210,N_13054,N_13037);
xnor U13211 (N_13211,N_13113,N_12968);
or U13212 (N_13212,N_13099,N_13040);
and U13213 (N_13213,N_13060,N_13092);
xnor U13214 (N_13214,N_13093,N_13062);
nand U13215 (N_13215,N_13050,N_12962);
nand U13216 (N_13216,N_13055,N_13087);
xnor U13217 (N_13217,N_13096,N_12965);
xor U13218 (N_13218,N_13067,N_13089);
or U13219 (N_13219,N_13014,N_12981);
nand U13220 (N_13220,N_12964,N_13086);
and U13221 (N_13221,N_13069,N_13014);
nand U13222 (N_13222,N_13021,N_13076);
xnor U13223 (N_13223,N_13051,N_13035);
or U13224 (N_13224,N_12986,N_13100);
nand U13225 (N_13225,N_13022,N_13103);
and U13226 (N_13226,N_13043,N_13013);
nor U13227 (N_13227,N_13027,N_12975);
or U13228 (N_13228,N_12978,N_13097);
nand U13229 (N_13229,N_13031,N_13116);
and U13230 (N_13230,N_13041,N_13056);
xor U13231 (N_13231,N_13052,N_13040);
nor U13232 (N_13232,N_13035,N_13113);
xnor U13233 (N_13233,N_13093,N_13085);
xnor U13234 (N_13234,N_13024,N_13069);
or U13235 (N_13235,N_13034,N_13077);
or U13236 (N_13236,N_13055,N_13012);
and U13237 (N_13237,N_13029,N_12984);
nor U13238 (N_13238,N_13084,N_13069);
or U13239 (N_13239,N_13075,N_12978);
and U13240 (N_13240,N_13107,N_12996);
or U13241 (N_13241,N_13027,N_13063);
nand U13242 (N_13242,N_13006,N_12989);
nand U13243 (N_13243,N_13088,N_13007);
and U13244 (N_13244,N_13006,N_12990);
and U13245 (N_13245,N_13015,N_13095);
xor U13246 (N_13246,N_13000,N_12979);
nor U13247 (N_13247,N_13077,N_13012);
and U13248 (N_13248,N_13038,N_13115);
nor U13249 (N_13249,N_13041,N_13010);
nor U13250 (N_13250,N_13006,N_13057);
or U13251 (N_13251,N_12996,N_13028);
and U13252 (N_13252,N_13000,N_13070);
or U13253 (N_13253,N_12999,N_12964);
and U13254 (N_13254,N_13098,N_13075);
nor U13255 (N_13255,N_13072,N_13107);
xor U13256 (N_13256,N_12980,N_12967);
or U13257 (N_13257,N_13059,N_12973);
nor U13258 (N_13258,N_13095,N_13011);
or U13259 (N_13259,N_12985,N_13086);
xnor U13260 (N_13260,N_12976,N_12992);
xnor U13261 (N_13261,N_13048,N_13060);
nand U13262 (N_13262,N_13063,N_13074);
and U13263 (N_13263,N_13077,N_13090);
and U13264 (N_13264,N_13038,N_13023);
xnor U13265 (N_13265,N_12962,N_13103);
xnor U13266 (N_13266,N_13109,N_12964);
xor U13267 (N_13267,N_12981,N_13046);
xor U13268 (N_13268,N_13089,N_13033);
or U13269 (N_13269,N_12961,N_13055);
and U13270 (N_13270,N_13102,N_12976);
and U13271 (N_13271,N_12976,N_13046);
and U13272 (N_13272,N_13049,N_12964);
nand U13273 (N_13273,N_12995,N_13015);
nor U13274 (N_13274,N_13042,N_13104);
nor U13275 (N_13275,N_12976,N_12974);
nor U13276 (N_13276,N_12980,N_13100);
or U13277 (N_13277,N_12981,N_13017);
nor U13278 (N_13278,N_13049,N_13103);
nand U13279 (N_13279,N_12962,N_13112);
nand U13280 (N_13280,N_13189,N_13223);
nand U13281 (N_13281,N_13234,N_13265);
and U13282 (N_13282,N_13174,N_13196);
nor U13283 (N_13283,N_13181,N_13248);
nand U13284 (N_13284,N_13128,N_13216);
nor U13285 (N_13285,N_13209,N_13177);
and U13286 (N_13286,N_13271,N_13121);
xor U13287 (N_13287,N_13122,N_13137);
nand U13288 (N_13288,N_13127,N_13144);
nor U13289 (N_13289,N_13160,N_13131);
and U13290 (N_13290,N_13191,N_13171);
nand U13291 (N_13291,N_13237,N_13240);
nor U13292 (N_13292,N_13123,N_13238);
xnor U13293 (N_13293,N_13233,N_13200);
nor U13294 (N_13294,N_13151,N_13262);
xor U13295 (N_13295,N_13199,N_13190);
or U13296 (N_13296,N_13264,N_13168);
nor U13297 (N_13297,N_13273,N_13165);
or U13298 (N_13298,N_13229,N_13249);
xor U13299 (N_13299,N_13244,N_13232);
nand U13300 (N_13300,N_13134,N_13213);
nor U13301 (N_13301,N_13226,N_13178);
nor U13302 (N_13302,N_13241,N_13173);
and U13303 (N_13303,N_13263,N_13203);
xnor U13304 (N_13304,N_13217,N_13207);
xor U13305 (N_13305,N_13225,N_13138);
and U13306 (N_13306,N_13182,N_13198);
and U13307 (N_13307,N_13239,N_13253);
and U13308 (N_13308,N_13242,N_13246);
nor U13309 (N_13309,N_13201,N_13268);
and U13310 (N_13310,N_13183,N_13208);
nand U13311 (N_13311,N_13205,N_13252);
or U13312 (N_13312,N_13243,N_13277);
and U13313 (N_13313,N_13143,N_13156);
and U13314 (N_13314,N_13167,N_13154);
and U13315 (N_13315,N_13188,N_13194);
nand U13316 (N_13316,N_13254,N_13222);
or U13317 (N_13317,N_13135,N_13140);
nor U13318 (N_13318,N_13125,N_13228);
nand U13319 (N_13319,N_13129,N_13270);
and U13320 (N_13320,N_13120,N_13235);
or U13321 (N_13321,N_13192,N_13231);
xor U13322 (N_13322,N_13250,N_13149);
nor U13323 (N_13323,N_13275,N_13152);
nand U13324 (N_13324,N_13202,N_13220);
xnor U13325 (N_13325,N_13276,N_13153);
nor U13326 (N_13326,N_13150,N_13141);
nand U13327 (N_13327,N_13204,N_13179);
nor U13328 (N_13328,N_13219,N_13175);
or U13329 (N_13329,N_13158,N_13251);
nor U13330 (N_13330,N_13146,N_13256);
and U13331 (N_13331,N_13130,N_13162);
nand U13332 (N_13332,N_13230,N_13187);
or U13333 (N_13333,N_13260,N_13170);
nand U13334 (N_13334,N_13159,N_13157);
nor U13335 (N_13335,N_13163,N_13269);
and U13336 (N_13336,N_13267,N_13147);
and U13337 (N_13337,N_13180,N_13139);
nor U13338 (N_13338,N_13161,N_13197);
nand U13339 (N_13339,N_13278,N_13221);
xnor U13340 (N_13340,N_13266,N_13210);
and U13341 (N_13341,N_13124,N_13245);
xnor U13342 (N_13342,N_13176,N_13195);
or U13343 (N_13343,N_13184,N_13172);
xnor U13344 (N_13344,N_13224,N_13148);
xor U13345 (N_13345,N_13133,N_13132);
and U13346 (N_13346,N_13236,N_13261);
or U13347 (N_13347,N_13274,N_13255);
nand U13348 (N_13348,N_13169,N_13136);
nand U13349 (N_13349,N_13142,N_13257);
xor U13350 (N_13350,N_13272,N_13164);
nand U13351 (N_13351,N_13155,N_13214);
and U13352 (N_13352,N_13259,N_13227);
and U13353 (N_13353,N_13166,N_13145);
and U13354 (N_13354,N_13212,N_13218);
and U13355 (N_13355,N_13258,N_13193);
and U13356 (N_13356,N_13211,N_13206);
xnor U13357 (N_13357,N_13215,N_13186);
nor U13358 (N_13358,N_13247,N_13279);
or U13359 (N_13359,N_13126,N_13185);
nor U13360 (N_13360,N_13229,N_13209);
or U13361 (N_13361,N_13179,N_13180);
or U13362 (N_13362,N_13245,N_13269);
xnor U13363 (N_13363,N_13194,N_13277);
nor U13364 (N_13364,N_13274,N_13145);
and U13365 (N_13365,N_13200,N_13191);
nand U13366 (N_13366,N_13161,N_13131);
nor U13367 (N_13367,N_13274,N_13188);
or U13368 (N_13368,N_13184,N_13226);
and U13369 (N_13369,N_13205,N_13209);
nand U13370 (N_13370,N_13222,N_13148);
nor U13371 (N_13371,N_13204,N_13196);
nor U13372 (N_13372,N_13273,N_13162);
nand U13373 (N_13373,N_13230,N_13232);
or U13374 (N_13374,N_13158,N_13157);
nand U13375 (N_13375,N_13279,N_13272);
nand U13376 (N_13376,N_13208,N_13126);
or U13377 (N_13377,N_13259,N_13264);
xnor U13378 (N_13378,N_13236,N_13134);
xor U13379 (N_13379,N_13184,N_13211);
or U13380 (N_13380,N_13271,N_13135);
nand U13381 (N_13381,N_13262,N_13273);
xnor U13382 (N_13382,N_13225,N_13245);
or U13383 (N_13383,N_13180,N_13208);
or U13384 (N_13384,N_13139,N_13263);
xnor U13385 (N_13385,N_13169,N_13242);
nor U13386 (N_13386,N_13187,N_13259);
or U13387 (N_13387,N_13249,N_13258);
xnor U13388 (N_13388,N_13132,N_13143);
xnor U13389 (N_13389,N_13194,N_13206);
xor U13390 (N_13390,N_13167,N_13232);
or U13391 (N_13391,N_13144,N_13132);
nand U13392 (N_13392,N_13127,N_13211);
xor U13393 (N_13393,N_13158,N_13138);
xnor U13394 (N_13394,N_13158,N_13204);
nor U13395 (N_13395,N_13217,N_13232);
xor U13396 (N_13396,N_13220,N_13203);
or U13397 (N_13397,N_13159,N_13232);
nor U13398 (N_13398,N_13209,N_13122);
and U13399 (N_13399,N_13237,N_13189);
nand U13400 (N_13400,N_13121,N_13218);
or U13401 (N_13401,N_13229,N_13176);
xor U13402 (N_13402,N_13162,N_13196);
xnor U13403 (N_13403,N_13220,N_13248);
nand U13404 (N_13404,N_13273,N_13133);
nor U13405 (N_13405,N_13143,N_13123);
nand U13406 (N_13406,N_13152,N_13155);
or U13407 (N_13407,N_13133,N_13162);
and U13408 (N_13408,N_13133,N_13230);
and U13409 (N_13409,N_13229,N_13179);
nand U13410 (N_13410,N_13148,N_13144);
nor U13411 (N_13411,N_13182,N_13258);
nand U13412 (N_13412,N_13207,N_13147);
nand U13413 (N_13413,N_13232,N_13210);
xor U13414 (N_13414,N_13150,N_13199);
and U13415 (N_13415,N_13195,N_13206);
or U13416 (N_13416,N_13264,N_13183);
nand U13417 (N_13417,N_13212,N_13188);
xnor U13418 (N_13418,N_13273,N_13150);
nor U13419 (N_13419,N_13151,N_13186);
xor U13420 (N_13420,N_13137,N_13252);
nand U13421 (N_13421,N_13263,N_13130);
nand U13422 (N_13422,N_13233,N_13142);
nand U13423 (N_13423,N_13239,N_13273);
or U13424 (N_13424,N_13121,N_13198);
or U13425 (N_13425,N_13120,N_13258);
and U13426 (N_13426,N_13148,N_13152);
or U13427 (N_13427,N_13125,N_13183);
and U13428 (N_13428,N_13187,N_13174);
and U13429 (N_13429,N_13277,N_13222);
nand U13430 (N_13430,N_13201,N_13246);
xor U13431 (N_13431,N_13235,N_13154);
xor U13432 (N_13432,N_13224,N_13160);
xnor U13433 (N_13433,N_13276,N_13128);
or U13434 (N_13434,N_13197,N_13270);
or U13435 (N_13435,N_13173,N_13127);
xnor U13436 (N_13436,N_13212,N_13201);
xor U13437 (N_13437,N_13121,N_13235);
xor U13438 (N_13438,N_13177,N_13197);
nor U13439 (N_13439,N_13213,N_13194);
or U13440 (N_13440,N_13394,N_13332);
and U13441 (N_13441,N_13367,N_13283);
nand U13442 (N_13442,N_13307,N_13333);
xor U13443 (N_13443,N_13434,N_13430);
xnor U13444 (N_13444,N_13408,N_13431);
and U13445 (N_13445,N_13422,N_13366);
nor U13446 (N_13446,N_13315,N_13403);
nor U13447 (N_13447,N_13288,N_13340);
and U13448 (N_13448,N_13327,N_13380);
nand U13449 (N_13449,N_13316,N_13391);
xor U13450 (N_13450,N_13382,N_13309);
or U13451 (N_13451,N_13397,N_13323);
xnor U13452 (N_13452,N_13420,N_13411);
and U13453 (N_13453,N_13427,N_13405);
xor U13454 (N_13454,N_13344,N_13436);
nor U13455 (N_13455,N_13348,N_13387);
and U13456 (N_13456,N_13304,N_13302);
or U13457 (N_13457,N_13365,N_13414);
nor U13458 (N_13458,N_13418,N_13284);
and U13459 (N_13459,N_13341,N_13299);
and U13460 (N_13460,N_13329,N_13407);
nor U13461 (N_13461,N_13416,N_13346);
xor U13462 (N_13462,N_13437,N_13317);
or U13463 (N_13463,N_13339,N_13303);
or U13464 (N_13464,N_13372,N_13334);
nor U13465 (N_13465,N_13395,N_13301);
or U13466 (N_13466,N_13285,N_13392);
nand U13467 (N_13467,N_13331,N_13406);
xor U13468 (N_13468,N_13359,N_13324);
xnor U13469 (N_13469,N_13353,N_13362);
nor U13470 (N_13470,N_13377,N_13381);
xor U13471 (N_13471,N_13393,N_13345);
nand U13472 (N_13472,N_13413,N_13310);
and U13473 (N_13473,N_13401,N_13298);
nor U13474 (N_13474,N_13371,N_13281);
or U13475 (N_13475,N_13426,N_13398);
nor U13476 (N_13476,N_13305,N_13336);
nor U13477 (N_13477,N_13425,N_13386);
xor U13478 (N_13478,N_13389,N_13357);
and U13479 (N_13479,N_13330,N_13421);
xnor U13480 (N_13480,N_13338,N_13297);
nand U13481 (N_13481,N_13356,N_13360);
or U13482 (N_13482,N_13294,N_13280);
nor U13483 (N_13483,N_13321,N_13385);
or U13484 (N_13484,N_13312,N_13311);
xor U13485 (N_13485,N_13373,N_13319);
nand U13486 (N_13486,N_13396,N_13383);
nor U13487 (N_13487,N_13290,N_13355);
nor U13488 (N_13488,N_13388,N_13342);
nand U13489 (N_13489,N_13409,N_13337);
or U13490 (N_13490,N_13378,N_13322);
or U13491 (N_13491,N_13350,N_13368);
xnor U13492 (N_13492,N_13291,N_13410);
and U13493 (N_13493,N_13415,N_13320);
or U13494 (N_13494,N_13314,N_13379);
and U13495 (N_13495,N_13374,N_13428);
nor U13496 (N_13496,N_13352,N_13423);
and U13497 (N_13497,N_13361,N_13335);
and U13498 (N_13498,N_13400,N_13432);
xnor U13499 (N_13499,N_13296,N_13325);
nor U13500 (N_13500,N_13363,N_13424);
nor U13501 (N_13501,N_13282,N_13364);
xnor U13502 (N_13502,N_13369,N_13349);
and U13503 (N_13503,N_13328,N_13318);
and U13504 (N_13504,N_13351,N_13343);
xor U13505 (N_13505,N_13439,N_13376);
nor U13506 (N_13506,N_13295,N_13313);
nor U13507 (N_13507,N_13402,N_13289);
or U13508 (N_13508,N_13390,N_13293);
nand U13509 (N_13509,N_13399,N_13433);
xnor U13510 (N_13510,N_13429,N_13435);
and U13511 (N_13511,N_13358,N_13412);
or U13512 (N_13512,N_13287,N_13300);
or U13513 (N_13513,N_13306,N_13354);
or U13514 (N_13514,N_13404,N_13292);
xnor U13515 (N_13515,N_13370,N_13308);
and U13516 (N_13516,N_13419,N_13384);
xor U13517 (N_13517,N_13326,N_13375);
xnor U13518 (N_13518,N_13417,N_13438);
nor U13519 (N_13519,N_13347,N_13286);
or U13520 (N_13520,N_13367,N_13394);
nor U13521 (N_13521,N_13433,N_13354);
and U13522 (N_13522,N_13282,N_13366);
and U13523 (N_13523,N_13439,N_13432);
nand U13524 (N_13524,N_13398,N_13286);
or U13525 (N_13525,N_13411,N_13363);
nand U13526 (N_13526,N_13306,N_13414);
or U13527 (N_13527,N_13433,N_13411);
and U13528 (N_13528,N_13384,N_13289);
or U13529 (N_13529,N_13427,N_13390);
xor U13530 (N_13530,N_13325,N_13372);
xnor U13531 (N_13531,N_13414,N_13331);
and U13532 (N_13532,N_13424,N_13314);
or U13533 (N_13533,N_13348,N_13361);
nor U13534 (N_13534,N_13330,N_13409);
nand U13535 (N_13535,N_13364,N_13423);
nand U13536 (N_13536,N_13365,N_13367);
or U13537 (N_13537,N_13390,N_13343);
xor U13538 (N_13538,N_13321,N_13307);
nor U13539 (N_13539,N_13428,N_13346);
nor U13540 (N_13540,N_13345,N_13332);
and U13541 (N_13541,N_13313,N_13375);
and U13542 (N_13542,N_13395,N_13422);
nor U13543 (N_13543,N_13319,N_13416);
xnor U13544 (N_13544,N_13385,N_13344);
nor U13545 (N_13545,N_13305,N_13281);
and U13546 (N_13546,N_13296,N_13401);
and U13547 (N_13547,N_13293,N_13420);
or U13548 (N_13548,N_13355,N_13364);
nand U13549 (N_13549,N_13304,N_13379);
nand U13550 (N_13550,N_13338,N_13350);
or U13551 (N_13551,N_13412,N_13284);
or U13552 (N_13552,N_13368,N_13355);
or U13553 (N_13553,N_13319,N_13382);
or U13554 (N_13554,N_13346,N_13356);
or U13555 (N_13555,N_13324,N_13418);
nand U13556 (N_13556,N_13357,N_13400);
nor U13557 (N_13557,N_13376,N_13282);
nand U13558 (N_13558,N_13429,N_13424);
and U13559 (N_13559,N_13296,N_13317);
or U13560 (N_13560,N_13428,N_13402);
xnor U13561 (N_13561,N_13392,N_13412);
xor U13562 (N_13562,N_13316,N_13299);
and U13563 (N_13563,N_13413,N_13352);
nor U13564 (N_13564,N_13368,N_13411);
or U13565 (N_13565,N_13401,N_13283);
and U13566 (N_13566,N_13393,N_13285);
and U13567 (N_13567,N_13349,N_13353);
xnor U13568 (N_13568,N_13434,N_13349);
and U13569 (N_13569,N_13415,N_13339);
nor U13570 (N_13570,N_13424,N_13328);
and U13571 (N_13571,N_13351,N_13294);
nand U13572 (N_13572,N_13432,N_13434);
xnor U13573 (N_13573,N_13431,N_13318);
nand U13574 (N_13574,N_13414,N_13371);
xnor U13575 (N_13575,N_13295,N_13430);
or U13576 (N_13576,N_13358,N_13310);
xor U13577 (N_13577,N_13432,N_13415);
nor U13578 (N_13578,N_13344,N_13387);
xor U13579 (N_13579,N_13420,N_13282);
or U13580 (N_13580,N_13351,N_13435);
and U13581 (N_13581,N_13397,N_13334);
and U13582 (N_13582,N_13317,N_13347);
or U13583 (N_13583,N_13352,N_13309);
xor U13584 (N_13584,N_13411,N_13364);
nand U13585 (N_13585,N_13413,N_13366);
xnor U13586 (N_13586,N_13394,N_13348);
and U13587 (N_13587,N_13314,N_13341);
nor U13588 (N_13588,N_13368,N_13289);
xnor U13589 (N_13589,N_13323,N_13385);
xor U13590 (N_13590,N_13327,N_13421);
xnor U13591 (N_13591,N_13437,N_13436);
or U13592 (N_13592,N_13404,N_13312);
nand U13593 (N_13593,N_13326,N_13358);
nand U13594 (N_13594,N_13345,N_13366);
nor U13595 (N_13595,N_13319,N_13333);
xnor U13596 (N_13596,N_13353,N_13314);
or U13597 (N_13597,N_13411,N_13412);
or U13598 (N_13598,N_13291,N_13296);
nor U13599 (N_13599,N_13400,N_13294);
nor U13600 (N_13600,N_13564,N_13463);
xor U13601 (N_13601,N_13502,N_13448);
or U13602 (N_13602,N_13500,N_13582);
or U13603 (N_13603,N_13568,N_13520);
nor U13604 (N_13604,N_13498,N_13598);
and U13605 (N_13605,N_13515,N_13566);
and U13606 (N_13606,N_13473,N_13548);
and U13607 (N_13607,N_13487,N_13546);
and U13608 (N_13608,N_13586,N_13489);
nand U13609 (N_13609,N_13554,N_13486);
nand U13610 (N_13610,N_13467,N_13596);
and U13611 (N_13611,N_13465,N_13480);
xnor U13612 (N_13612,N_13589,N_13492);
and U13613 (N_13613,N_13481,N_13584);
nand U13614 (N_13614,N_13495,N_13545);
nor U13615 (N_13615,N_13585,N_13471);
xnor U13616 (N_13616,N_13539,N_13510);
or U13617 (N_13617,N_13529,N_13578);
nor U13618 (N_13618,N_13597,N_13535);
nand U13619 (N_13619,N_13577,N_13587);
nor U13620 (N_13620,N_13457,N_13511);
nor U13621 (N_13621,N_13464,N_13475);
xnor U13622 (N_13622,N_13454,N_13549);
or U13623 (N_13623,N_13460,N_13483);
or U13624 (N_13624,N_13455,N_13506);
nand U13625 (N_13625,N_13469,N_13521);
nand U13626 (N_13626,N_13494,N_13524);
xor U13627 (N_13627,N_13499,N_13580);
nand U13628 (N_13628,N_13474,N_13461);
nand U13629 (N_13629,N_13588,N_13556);
or U13630 (N_13630,N_13547,N_13449);
or U13631 (N_13631,N_13594,N_13555);
xnor U13632 (N_13632,N_13579,N_13592);
nand U13633 (N_13633,N_13537,N_13488);
nor U13634 (N_13634,N_13522,N_13512);
or U13635 (N_13635,N_13450,N_13516);
and U13636 (N_13636,N_13575,N_13466);
nor U13637 (N_13637,N_13538,N_13552);
nor U13638 (N_13638,N_13479,N_13451);
xor U13639 (N_13639,N_13542,N_13497);
xnor U13640 (N_13640,N_13528,N_13572);
or U13641 (N_13641,N_13441,N_13543);
and U13642 (N_13642,N_13496,N_13553);
xor U13643 (N_13643,N_13443,N_13567);
nand U13644 (N_13644,N_13562,N_13517);
or U13645 (N_13645,N_13501,N_13541);
xor U13646 (N_13646,N_13459,N_13490);
and U13647 (N_13647,N_13595,N_13550);
nor U13648 (N_13648,N_13442,N_13563);
nand U13649 (N_13649,N_13445,N_13583);
xnor U13650 (N_13650,N_13505,N_13485);
nor U13651 (N_13651,N_13525,N_13581);
xnor U13652 (N_13652,N_13453,N_13532);
nor U13653 (N_13653,N_13508,N_13558);
or U13654 (N_13654,N_13569,N_13468);
and U13655 (N_13655,N_13540,N_13447);
nand U13656 (N_13656,N_13576,N_13530);
or U13657 (N_13657,N_13570,N_13536);
nor U13658 (N_13658,N_13476,N_13590);
and U13659 (N_13659,N_13557,N_13561);
nand U13660 (N_13660,N_13551,N_13593);
or U13661 (N_13661,N_13472,N_13573);
or U13662 (N_13662,N_13456,N_13503);
nand U13663 (N_13663,N_13531,N_13560);
nor U13664 (N_13664,N_13574,N_13565);
and U13665 (N_13665,N_13446,N_13452);
nand U13666 (N_13666,N_13526,N_13504);
nor U13667 (N_13667,N_13571,N_13513);
nand U13668 (N_13668,N_13534,N_13478);
and U13669 (N_13669,N_13507,N_13591);
or U13670 (N_13670,N_13440,N_13527);
nor U13671 (N_13671,N_13514,N_13599);
nand U13672 (N_13672,N_13519,N_13559);
and U13673 (N_13673,N_13470,N_13509);
or U13674 (N_13674,N_13462,N_13523);
nor U13675 (N_13675,N_13518,N_13484);
xnor U13676 (N_13676,N_13491,N_13477);
and U13677 (N_13677,N_13533,N_13482);
nor U13678 (N_13678,N_13544,N_13493);
xnor U13679 (N_13679,N_13458,N_13444);
nand U13680 (N_13680,N_13459,N_13543);
nand U13681 (N_13681,N_13542,N_13566);
and U13682 (N_13682,N_13492,N_13567);
nor U13683 (N_13683,N_13517,N_13474);
and U13684 (N_13684,N_13473,N_13507);
or U13685 (N_13685,N_13597,N_13583);
nor U13686 (N_13686,N_13444,N_13459);
and U13687 (N_13687,N_13469,N_13503);
xnor U13688 (N_13688,N_13551,N_13486);
nand U13689 (N_13689,N_13483,N_13440);
nand U13690 (N_13690,N_13449,N_13528);
and U13691 (N_13691,N_13500,N_13492);
nand U13692 (N_13692,N_13484,N_13463);
and U13693 (N_13693,N_13562,N_13493);
nor U13694 (N_13694,N_13558,N_13451);
xnor U13695 (N_13695,N_13488,N_13463);
xor U13696 (N_13696,N_13486,N_13561);
nor U13697 (N_13697,N_13555,N_13596);
xor U13698 (N_13698,N_13512,N_13441);
xnor U13699 (N_13699,N_13473,N_13518);
xnor U13700 (N_13700,N_13501,N_13554);
nand U13701 (N_13701,N_13596,N_13445);
xor U13702 (N_13702,N_13455,N_13495);
xnor U13703 (N_13703,N_13582,N_13464);
nor U13704 (N_13704,N_13521,N_13563);
or U13705 (N_13705,N_13498,N_13550);
nor U13706 (N_13706,N_13472,N_13583);
or U13707 (N_13707,N_13545,N_13565);
and U13708 (N_13708,N_13527,N_13520);
nor U13709 (N_13709,N_13472,N_13474);
or U13710 (N_13710,N_13580,N_13465);
or U13711 (N_13711,N_13565,N_13483);
xor U13712 (N_13712,N_13579,N_13440);
nand U13713 (N_13713,N_13520,N_13557);
nor U13714 (N_13714,N_13524,N_13457);
and U13715 (N_13715,N_13571,N_13581);
xor U13716 (N_13716,N_13514,N_13508);
or U13717 (N_13717,N_13502,N_13531);
or U13718 (N_13718,N_13506,N_13501);
xnor U13719 (N_13719,N_13530,N_13490);
nand U13720 (N_13720,N_13584,N_13463);
and U13721 (N_13721,N_13568,N_13573);
xnor U13722 (N_13722,N_13571,N_13470);
and U13723 (N_13723,N_13549,N_13479);
nor U13724 (N_13724,N_13582,N_13517);
nand U13725 (N_13725,N_13512,N_13529);
nor U13726 (N_13726,N_13562,N_13568);
xor U13727 (N_13727,N_13441,N_13515);
or U13728 (N_13728,N_13486,N_13540);
nor U13729 (N_13729,N_13440,N_13572);
and U13730 (N_13730,N_13570,N_13555);
or U13731 (N_13731,N_13556,N_13448);
nor U13732 (N_13732,N_13443,N_13563);
xor U13733 (N_13733,N_13533,N_13578);
xor U13734 (N_13734,N_13539,N_13503);
and U13735 (N_13735,N_13448,N_13533);
nand U13736 (N_13736,N_13540,N_13563);
nor U13737 (N_13737,N_13477,N_13488);
and U13738 (N_13738,N_13470,N_13478);
nor U13739 (N_13739,N_13481,N_13488);
nand U13740 (N_13740,N_13572,N_13533);
nor U13741 (N_13741,N_13466,N_13561);
and U13742 (N_13742,N_13553,N_13594);
and U13743 (N_13743,N_13577,N_13462);
nor U13744 (N_13744,N_13552,N_13458);
nor U13745 (N_13745,N_13525,N_13443);
nand U13746 (N_13746,N_13525,N_13451);
xor U13747 (N_13747,N_13530,N_13533);
nand U13748 (N_13748,N_13515,N_13541);
and U13749 (N_13749,N_13597,N_13449);
or U13750 (N_13750,N_13565,N_13584);
xnor U13751 (N_13751,N_13583,N_13507);
nor U13752 (N_13752,N_13474,N_13529);
nand U13753 (N_13753,N_13521,N_13501);
xor U13754 (N_13754,N_13468,N_13547);
nand U13755 (N_13755,N_13593,N_13508);
xnor U13756 (N_13756,N_13548,N_13583);
and U13757 (N_13757,N_13452,N_13468);
or U13758 (N_13758,N_13455,N_13459);
nor U13759 (N_13759,N_13518,N_13502);
and U13760 (N_13760,N_13732,N_13733);
nor U13761 (N_13761,N_13662,N_13656);
or U13762 (N_13762,N_13632,N_13611);
nand U13763 (N_13763,N_13758,N_13711);
and U13764 (N_13764,N_13637,N_13643);
or U13765 (N_13765,N_13685,N_13699);
xor U13766 (N_13766,N_13649,N_13694);
nand U13767 (N_13767,N_13686,N_13625);
or U13768 (N_13768,N_13620,N_13674);
or U13769 (N_13769,N_13600,N_13728);
nor U13770 (N_13770,N_13705,N_13629);
nor U13771 (N_13771,N_13659,N_13669);
or U13772 (N_13772,N_13742,N_13676);
xnor U13773 (N_13773,N_13755,N_13745);
or U13774 (N_13774,N_13603,N_13719);
nor U13775 (N_13775,N_13683,N_13718);
and U13776 (N_13776,N_13636,N_13697);
and U13777 (N_13777,N_13757,N_13663);
nand U13778 (N_13778,N_13743,N_13695);
and U13779 (N_13779,N_13731,N_13654);
and U13780 (N_13780,N_13621,N_13640);
xnor U13781 (N_13781,N_13619,N_13673);
xor U13782 (N_13782,N_13668,N_13675);
nand U13783 (N_13783,N_13751,N_13730);
or U13784 (N_13784,N_13723,N_13689);
or U13785 (N_13785,N_13759,N_13642);
and U13786 (N_13786,N_13672,N_13688);
nand U13787 (N_13787,N_13752,N_13708);
and U13788 (N_13788,N_13749,N_13613);
nor U13789 (N_13789,N_13739,N_13646);
nor U13790 (N_13790,N_13703,N_13616);
nor U13791 (N_13791,N_13720,N_13658);
xor U13792 (N_13792,N_13707,N_13618);
nor U13793 (N_13793,N_13712,N_13753);
nand U13794 (N_13794,N_13671,N_13687);
xnor U13795 (N_13795,N_13638,N_13666);
nor U13796 (N_13796,N_13641,N_13680);
and U13797 (N_13797,N_13679,N_13748);
xor U13798 (N_13798,N_13655,N_13609);
or U13799 (N_13799,N_13608,N_13704);
or U13800 (N_13800,N_13710,N_13665);
nor U13801 (N_13801,N_13681,N_13729);
or U13802 (N_13802,N_13756,N_13651);
nand U13803 (N_13803,N_13635,N_13606);
and U13804 (N_13804,N_13701,N_13738);
nor U13805 (N_13805,N_13648,N_13660);
nor U13806 (N_13806,N_13670,N_13627);
xnor U13807 (N_13807,N_13664,N_13639);
nand U13808 (N_13808,N_13661,N_13750);
nor U13809 (N_13809,N_13717,N_13630);
nand U13810 (N_13810,N_13678,N_13667);
nor U13811 (N_13811,N_13754,N_13612);
nor U13812 (N_13812,N_13604,N_13605);
nor U13813 (N_13813,N_13722,N_13607);
and U13814 (N_13814,N_13677,N_13716);
and U13815 (N_13815,N_13650,N_13631);
or U13816 (N_13816,N_13696,N_13724);
xnor U13817 (N_13817,N_13734,N_13715);
and U13818 (N_13818,N_13706,N_13698);
nor U13819 (N_13819,N_13614,N_13709);
and U13820 (N_13820,N_13744,N_13601);
or U13821 (N_13821,N_13726,N_13740);
and U13822 (N_13822,N_13692,N_13746);
nor U13823 (N_13823,N_13747,N_13737);
and U13824 (N_13824,N_13626,N_13645);
nor U13825 (N_13825,N_13634,N_13684);
nor U13826 (N_13826,N_13713,N_13727);
or U13827 (N_13827,N_13647,N_13610);
xor U13828 (N_13828,N_13615,N_13682);
and U13829 (N_13829,N_13736,N_13700);
xnor U13830 (N_13830,N_13624,N_13628);
xnor U13831 (N_13831,N_13617,N_13702);
and U13832 (N_13832,N_13652,N_13602);
nand U13833 (N_13833,N_13721,N_13741);
xnor U13834 (N_13834,N_13622,N_13623);
xnor U13835 (N_13835,N_13691,N_13714);
xor U13836 (N_13836,N_13725,N_13690);
nand U13837 (N_13837,N_13693,N_13653);
xnor U13838 (N_13838,N_13657,N_13633);
and U13839 (N_13839,N_13644,N_13735);
and U13840 (N_13840,N_13688,N_13650);
nand U13841 (N_13841,N_13639,N_13603);
xnor U13842 (N_13842,N_13606,N_13682);
xor U13843 (N_13843,N_13679,N_13636);
nand U13844 (N_13844,N_13610,N_13664);
xor U13845 (N_13845,N_13737,N_13603);
xor U13846 (N_13846,N_13685,N_13656);
and U13847 (N_13847,N_13609,N_13726);
xor U13848 (N_13848,N_13613,N_13605);
and U13849 (N_13849,N_13735,N_13752);
xor U13850 (N_13850,N_13655,N_13685);
xnor U13851 (N_13851,N_13750,N_13640);
nand U13852 (N_13852,N_13710,N_13689);
and U13853 (N_13853,N_13702,N_13629);
xor U13854 (N_13854,N_13734,N_13694);
and U13855 (N_13855,N_13720,N_13655);
and U13856 (N_13856,N_13753,N_13693);
xor U13857 (N_13857,N_13718,N_13723);
xor U13858 (N_13858,N_13653,N_13611);
xor U13859 (N_13859,N_13634,N_13671);
or U13860 (N_13860,N_13641,N_13749);
and U13861 (N_13861,N_13643,N_13621);
xnor U13862 (N_13862,N_13607,N_13714);
or U13863 (N_13863,N_13683,N_13752);
nor U13864 (N_13864,N_13671,N_13620);
nand U13865 (N_13865,N_13699,N_13728);
and U13866 (N_13866,N_13713,N_13714);
and U13867 (N_13867,N_13730,N_13736);
nor U13868 (N_13868,N_13736,N_13746);
and U13869 (N_13869,N_13644,N_13756);
or U13870 (N_13870,N_13697,N_13623);
and U13871 (N_13871,N_13715,N_13601);
nand U13872 (N_13872,N_13639,N_13601);
xnor U13873 (N_13873,N_13705,N_13658);
or U13874 (N_13874,N_13729,N_13665);
nor U13875 (N_13875,N_13607,N_13665);
nand U13876 (N_13876,N_13620,N_13711);
nand U13877 (N_13877,N_13681,N_13708);
xor U13878 (N_13878,N_13730,N_13647);
nor U13879 (N_13879,N_13682,N_13721);
nand U13880 (N_13880,N_13633,N_13680);
nand U13881 (N_13881,N_13629,N_13699);
and U13882 (N_13882,N_13738,N_13647);
and U13883 (N_13883,N_13602,N_13636);
xor U13884 (N_13884,N_13658,N_13691);
xnor U13885 (N_13885,N_13704,N_13697);
xor U13886 (N_13886,N_13700,N_13640);
nand U13887 (N_13887,N_13682,N_13726);
or U13888 (N_13888,N_13715,N_13615);
or U13889 (N_13889,N_13714,N_13643);
nand U13890 (N_13890,N_13606,N_13717);
nor U13891 (N_13891,N_13656,N_13666);
xnor U13892 (N_13892,N_13725,N_13697);
and U13893 (N_13893,N_13711,N_13603);
xnor U13894 (N_13894,N_13633,N_13612);
nor U13895 (N_13895,N_13663,N_13728);
nand U13896 (N_13896,N_13734,N_13638);
nor U13897 (N_13897,N_13607,N_13748);
or U13898 (N_13898,N_13742,N_13600);
or U13899 (N_13899,N_13661,N_13719);
or U13900 (N_13900,N_13741,N_13656);
or U13901 (N_13901,N_13618,N_13739);
nor U13902 (N_13902,N_13746,N_13743);
or U13903 (N_13903,N_13746,N_13639);
and U13904 (N_13904,N_13748,N_13669);
or U13905 (N_13905,N_13686,N_13713);
nor U13906 (N_13906,N_13615,N_13722);
or U13907 (N_13907,N_13718,N_13651);
and U13908 (N_13908,N_13616,N_13728);
nand U13909 (N_13909,N_13700,N_13731);
nand U13910 (N_13910,N_13736,N_13749);
xor U13911 (N_13911,N_13611,N_13701);
nand U13912 (N_13912,N_13705,N_13624);
xor U13913 (N_13913,N_13662,N_13716);
or U13914 (N_13914,N_13663,N_13717);
and U13915 (N_13915,N_13654,N_13710);
nor U13916 (N_13916,N_13642,N_13734);
or U13917 (N_13917,N_13619,N_13675);
and U13918 (N_13918,N_13735,N_13630);
and U13919 (N_13919,N_13642,N_13747);
nand U13920 (N_13920,N_13845,N_13840);
or U13921 (N_13921,N_13804,N_13793);
nand U13922 (N_13922,N_13792,N_13770);
or U13923 (N_13923,N_13786,N_13876);
nand U13924 (N_13924,N_13900,N_13869);
xnor U13925 (N_13925,N_13892,N_13831);
nand U13926 (N_13926,N_13916,N_13797);
nand U13927 (N_13927,N_13824,N_13885);
and U13928 (N_13928,N_13861,N_13838);
or U13929 (N_13929,N_13846,N_13810);
and U13930 (N_13930,N_13774,N_13827);
xor U13931 (N_13931,N_13908,N_13798);
nand U13932 (N_13932,N_13785,N_13794);
or U13933 (N_13933,N_13800,N_13820);
or U13934 (N_13934,N_13802,N_13782);
nand U13935 (N_13935,N_13821,N_13765);
nand U13936 (N_13936,N_13805,N_13829);
nand U13937 (N_13937,N_13807,N_13855);
or U13938 (N_13938,N_13812,N_13907);
nand U13939 (N_13939,N_13780,N_13883);
and U13940 (N_13940,N_13849,N_13760);
or U13941 (N_13941,N_13769,N_13790);
nand U13942 (N_13942,N_13880,N_13814);
and U13943 (N_13943,N_13872,N_13826);
nor U13944 (N_13944,N_13902,N_13816);
and U13945 (N_13945,N_13813,N_13918);
nand U13946 (N_13946,N_13832,N_13776);
nand U13947 (N_13947,N_13778,N_13862);
or U13948 (N_13948,N_13766,N_13773);
nor U13949 (N_13949,N_13775,N_13823);
nand U13950 (N_13950,N_13895,N_13799);
xor U13951 (N_13951,N_13904,N_13866);
or U13952 (N_13952,N_13839,N_13762);
nor U13953 (N_13953,N_13897,N_13871);
nand U13954 (N_13954,N_13905,N_13859);
nor U13955 (N_13955,N_13764,N_13864);
or U13956 (N_13956,N_13777,N_13819);
xor U13957 (N_13957,N_13772,N_13914);
and U13958 (N_13958,N_13847,N_13853);
nor U13959 (N_13959,N_13867,N_13860);
xor U13960 (N_13960,N_13913,N_13811);
nor U13961 (N_13961,N_13910,N_13806);
nor U13962 (N_13962,N_13868,N_13779);
xor U13963 (N_13963,N_13808,N_13768);
nand U13964 (N_13964,N_13801,N_13865);
xor U13965 (N_13965,N_13852,N_13771);
and U13966 (N_13966,N_13884,N_13899);
nand U13967 (N_13967,N_13815,N_13873);
or U13968 (N_13968,N_13834,N_13877);
or U13969 (N_13969,N_13888,N_13791);
and U13970 (N_13970,N_13919,N_13881);
nand U13971 (N_13971,N_13903,N_13917);
nor U13972 (N_13972,N_13788,N_13874);
and U13973 (N_13973,N_13842,N_13878);
nor U13974 (N_13974,N_13822,N_13896);
nand U13975 (N_13975,N_13795,N_13784);
nor U13976 (N_13976,N_13889,N_13893);
nand U13977 (N_13977,N_13843,N_13817);
or U13978 (N_13978,N_13854,N_13879);
xnor U13979 (N_13979,N_13870,N_13890);
xnor U13980 (N_13980,N_13858,N_13828);
or U13981 (N_13981,N_13850,N_13763);
nand U13982 (N_13982,N_13886,N_13851);
and U13983 (N_13983,N_13901,N_13898);
nand U13984 (N_13984,N_13887,N_13837);
or U13985 (N_13985,N_13848,N_13856);
and U13986 (N_13986,N_13796,N_13803);
or U13987 (N_13987,N_13767,N_13915);
nand U13988 (N_13988,N_13789,N_13830);
and U13989 (N_13989,N_13891,N_13809);
nor U13990 (N_13990,N_13761,N_13911);
xnor U13991 (N_13991,N_13863,N_13912);
nand U13992 (N_13992,N_13841,N_13882);
nand U13993 (N_13993,N_13844,N_13875);
or U13994 (N_13994,N_13787,N_13906);
and U13995 (N_13995,N_13894,N_13835);
nor U13996 (N_13996,N_13825,N_13909);
and U13997 (N_13997,N_13833,N_13857);
nor U13998 (N_13998,N_13818,N_13783);
and U13999 (N_13999,N_13781,N_13836);
xnor U14000 (N_14000,N_13853,N_13762);
or U14001 (N_14001,N_13857,N_13917);
and U14002 (N_14002,N_13855,N_13898);
xnor U14003 (N_14003,N_13847,N_13859);
xor U14004 (N_14004,N_13889,N_13839);
and U14005 (N_14005,N_13774,N_13787);
nand U14006 (N_14006,N_13837,N_13803);
or U14007 (N_14007,N_13787,N_13879);
xnor U14008 (N_14008,N_13794,N_13865);
xnor U14009 (N_14009,N_13871,N_13821);
or U14010 (N_14010,N_13879,N_13899);
nor U14011 (N_14011,N_13893,N_13782);
nor U14012 (N_14012,N_13887,N_13776);
and U14013 (N_14013,N_13880,N_13861);
nand U14014 (N_14014,N_13868,N_13902);
nor U14015 (N_14015,N_13882,N_13768);
and U14016 (N_14016,N_13833,N_13809);
nor U14017 (N_14017,N_13836,N_13916);
xnor U14018 (N_14018,N_13834,N_13794);
and U14019 (N_14019,N_13863,N_13804);
nand U14020 (N_14020,N_13864,N_13901);
nand U14021 (N_14021,N_13801,N_13896);
nand U14022 (N_14022,N_13816,N_13808);
nand U14023 (N_14023,N_13855,N_13881);
xor U14024 (N_14024,N_13766,N_13839);
xor U14025 (N_14025,N_13845,N_13804);
or U14026 (N_14026,N_13870,N_13820);
and U14027 (N_14027,N_13771,N_13833);
and U14028 (N_14028,N_13803,N_13875);
and U14029 (N_14029,N_13811,N_13919);
or U14030 (N_14030,N_13846,N_13819);
and U14031 (N_14031,N_13762,N_13821);
nand U14032 (N_14032,N_13813,N_13838);
or U14033 (N_14033,N_13894,N_13831);
xor U14034 (N_14034,N_13907,N_13795);
or U14035 (N_14035,N_13804,N_13848);
nor U14036 (N_14036,N_13876,N_13828);
xor U14037 (N_14037,N_13890,N_13789);
nand U14038 (N_14038,N_13841,N_13760);
nand U14039 (N_14039,N_13901,N_13866);
nand U14040 (N_14040,N_13843,N_13893);
nand U14041 (N_14041,N_13872,N_13833);
and U14042 (N_14042,N_13799,N_13781);
or U14043 (N_14043,N_13886,N_13826);
and U14044 (N_14044,N_13855,N_13867);
or U14045 (N_14045,N_13765,N_13841);
or U14046 (N_14046,N_13790,N_13802);
or U14047 (N_14047,N_13865,N_13787);
and U14048 (N_14048,N_13806,N_13770);
nor U14049 (N_14049,N_13806,N_13816);
and U14050 (N_14050,N_13762,N_13823);
xnor U14051 (N_14051,N_13915,N_13895);
nor U14052 (N_14052,N_13789,N_13898);
and U14053 (N_14053,N_13880,N_13903);
or U14054 (N_14054,N_13915,N_13777);
nor U14055 (N_14055,N_13825,N_13806);
or U14056 (N_14056,N_13899,N_13902);
nor U14057 (N_14057,N_13900,N_13786);
nor U14058 (N_14058,N_13768,N_13806);
nand U14059 (N_14059,N_13857,N_13888);
and U14060 (N_14060,N_13809,N_13849);
and U14061 (N_14061,N_13831,N_13908);
nor U14062 (N_14062,N_13811,N_13813);
or U14063 (N_14063,N_13832,N_13834);
nor U14064 (N_14064,N_13912,N_13839);
nand U14065 (N_14065,N_13788,N_13832);
nor U14066 (N_14066,N_13840,N_13781);
xnor U14067 (N_14067,N_13903,N_13800);
xor U14068 (N_14068,N_13770,N_13862);
and U14069 (N_14069,N_13835,N_13775);
and U14070 (N_14070,N_13776,N_13911);
nor U14071 (N_14071,N_13813,N_13830);
xor U14072 (N_14072,N_13858,N_13873);
and U14073 (N_14073,N_13874,N_13817);
nand U14074 (N_14074,N_13833,N_13810);
nor U14075 (N_14075,N_13907,N_13886);
xor U14076 (N_14076,N_13829,N_13862);
or U14077 (N_14077,N_13838,N_13831);
nand U14078 (N_14078,N_13768,N_13885);
and U14079 (N_14079,N_13856,N_13888);
or U14080 (N_14080,N_13998,N_13986);
or U14081 (N_14081,N_14055,N_14046);
xor U14082 (N_14082,N_13990,N_13993);
nand U14083 (N_14083,N_13992,N_14005);
nand U14084 (N_14084,N_13931,N_13967);
and U14085 (N_14085,N_13977,N_14030);
nand U14086 (N_14086,N_13988,N_13972);
nand U14087 (N_14087,N_14036,N_13980);
nor U14088 (N_14088,N_14037,N_14031);
xnor U14089 (N_14089,N_14026,N_14052);
xnor U14090 (N_14090,N_14050,N_14072);
and U14091 (N_14091,N_14061,N_13947);
and U14092 (N_14092,N_14003,N_13973);
and U14093 (N_14093,N_13983,N_14075);
xnor U14094 (N_14094,N_14073,N_13978);
xnor U14095 (N_14095,N_13937,N_14014);
nor U14096 (N_14096,N_14000,N_14007);
or U14097 (N_14097,N_14045,N_14028);
xor U14098 (N_14098,N_14048,N_13969);
nand U14099 (N_14099,N_14006,N_14067);
nand U14100 (N_14100,N_14018,N_13960);
nand U14101 (N_14101,N_13965,N_13925);
nor U14102 (N_14102,N_14011,N_14034);
xor U14103 (N_14103,N_13957,N_14001);
nor U14104 (N_14104,N_13975,N_14059);
xnor U14105 (N_14105,N_13933,N_13964);
xnor U14106 (N_14106,N_14049,N_14077);
and U14107 (N_14107,N_13970,N_13951);
xor U14108 (N_14108,N_13971,N_13929);
xnor U14109 (N_14109,N_13942,N_14040);
nor U14110 (N_14110,N_13943,N_13921);
or U14111 (N_14111,N_13999,N_14066);
or U14112 (N_14112,N_14070,N_14008);
nand U14113 (N_14113,N_14009,N_14013);
xor U14114 (N_14114,N_14039,N_14032);
nand U14115 (N_14115,N_13995,N_14064);
xnor U14116 (N_14116,N_13981,N_13923);
or U14117 (N_14117,N_14012,N_14060);
nand U14118 (N_14118,N_13982,N_14053);
xor U14119 (N_14119,N_13991,N_14042);
and U14120 (N_14120,N_13966,N_14038);
or U14121 (N_14121,N_14063,N_13920);
or U14122 (N_14122,N_13935,N_13939);
nand U14123 (N_14123,N_14019,N_13932);
nor U14124 (N_14124,N_13940,N_14068);
and U14125 (N_14125,N_13944,N_13989);
and U14126 (N_14126,N_13930,N_14071);
or U14127 (N_14127,N_14079,N_14010);
nand U14128 (N_14128,N_14078,N_14004);
xor U14129 (N_14129,N_13946,N_14074);
xor U14130 (N_14130,N_14002,N_13955);
and U14131 (N_14131,N_13994,N_13962);
or U14132 (N_14132,N_14027,N_14076);
nand U14133 (N_14133,N_13949,N_13997);
nand U14134 (N_14134,N_13985,N_14025);
and U14135 (N_14135,N_13987,N_14054);
nand U14136 (N_14136,N_13938,N_13996);
nor U14137 (N_14137,N_13956,N_14017);
and U14138 (N_14138,N_14029,N_14062);
xnor U14139 (N_14139,N_14016,N_13934);
nor U14140 (N_14140,N_13945,N_14020);
xor U14141 (N_14141,N_13941,N_13968);
nand U14142 (N_14142,N_14065,N_13954);
nor U14143 (N_14143,N_13950,N_13926);
nor U14144 (N_14144,N_14033,N_13961);
or U14145 (N_14145,N_14024,N_14043);
nor U14146 (N_14146,N_13952,N_14057);
and U14147 (N_14147,N_13924,N_14044);
and U14148 (N_14148,N_13927,N_13936);
nand U14149 (N_14149,N_14035,N_14041);
nand U14150 (N_14150,N_14015,N_13922);
nor U14151 (N_14151,N_14022,N_14069);
nor U14152 (N_14152,N_13958,N_13974);
xnor U14153 (N_14153,N_13979,N_13976);
or U14154 (N_14154,N_14023,N_14021);
nor U14155 (N_14155,N_14056,N_13948);
and U14156 (N_14156,N_13928,N_13959);
and U14157 (N_14157,N_13984,N_14047);
nand U14158 (N_14158,N_14051,N_13963);
or U14159 (N_14159,N_14058,N_13953);
or U14160 (N_14160,N_13958,N_13969);
nor U14161 (N_14161,N_13940,N_14013);
or U14162 (N_14162,N_14071,N_14067);
or U14163 (N_14163,N_14014,N_13929);
xor U14164 (N_14164,N_14014,N_13995);
or U14165 (N_14165,N_14068,N_13930);
xor U14166 (N_14166,N_14015,N_13960);
xor U14167 (N_14167,N_13939,N_13929);
nand U14168 (N_14168,N_14028,N_14041);
xnor U14169 (N_14169,N_13984,N_13952);
or U14170 (N_14170,N_13968,N_14078);
xnor U14171 (N_14171,N_13987,N_13972);
or U14172 (N_14172,N_14072,N_14041);
nor U14173 (N_14173,N_13974,N_13975);
xor U14174 (N_14174,N_13971,N_13932);
or U14175 (N_14175,N_14051,N_14071);
nand U14176 (N_14176,N_14075,N_14056);
xnor U14177 (N_14177,N_14016,N_13929);
nand U14178 (N_14178,N_14070,N_13956);
and U14179 (N_14179,N_13933,N_14044);
or U14180 (N_14180,N_13933,N_13992);
and U14181 (N_14181,N_13929,N_13952);
nand U14182 (N_14182,N_14014,N_13983);
nor U14183 (N_14183,N_13986,N_13963);
nor U14184 (N_14184,N_13961,N_14044);
and U14185 (N_14185,N_14004,N_13930);
xnor U14186 (N_14186,N_13927,N_13994);
nor U14187 (N_14187,N_13943,N_14048);
or U14188 (N_14188,N_14047,N_13956);
xor U14189 (N_14189,N_14043,N_14019);
xor U14190 (N_14190,N_13973,N_14047);
or U14191 (N_14191,N_13970,N_13962);
xor U14192 (N_14192,N_14008,N_14049);
nand U14193 (N_14193,N_14079,N_13937);
and U14194 (N_14194,N_14058,N_13965);
nand U14195 (N_14195,N_13934,N_14014);
nand U14196 (N_14196,N_14034,N_13973);
nand U14197 (N_14197,N_14062,N_13929);
nor U14198 (N_14198,N_13940,N_14051);
nor U14199 (N_14199,N_13950,N_14054);
nand U14200 (N_14200,N_14063,N_13981);
and U14201 (N_14201,N_13972,N_13938);
or U14202 (N_14202,N_13972,N_13976);
nand U14203 (N_14203,N_14003,N_14032);
nor U14204 (N_14204,N_13966,N_13993);
or U14205 (N_14205,N_13951,N_13973);
nor U14206 (N_14206,N_14079,N_14019);
and U14207 (N_14207,N_13991,N_14027);
or U14208 (N_14208,N_14078,N_13922);
and U14209 (N_14209,N_14012,N_14010);
or U14210 (N_14210,N_14037,N_13967);
nor U14211 (N_14211,N_13929,N_13926);
or U14212 (N_14212,N_13959,N_13981);
and U14213 (N_14213,N_14030,N_13991);
and U14214 (N_14214,N_13960,N_14047);
nor U14215 (N_14215,N_13952,N_13978);
or U14216 (N_14216,N_13950,N_13953);
and U14217 (N_14217,N_14045,N_13999);
xnor U14218 (N_14218,N_14006,N_13973);
nor U14219 (N_14219,N_13930,N_14052);
and U14220 (N_14220,N_13986,N_13954);
nor U14221 (N_14221,N_13997,N_14006);
nor U14222 (N_14222,N_13950,N_14003);
or U14223 (N_14223,N_13932,N_13952);
and U14224 (N_14224,N_14018,N_13926);
nand U14225 (N_14225,N_14022,N_14050);
or U14226 (N_14226,N_14029,N_14063);
and U14227 (N_14227,N_13968,N_14000);
and U14228 (N_14228,N_13973,N_14053);
xor U14229 (N_14229,N_14007,N_14079);
and U14230 (N_14230,N_13930,N_13972);
xor U14231 (N_14231,N_14079,N_14001);
xnor U14232 (N_14232,N_14006,N_14044);
nand U14233 (N_14233,N_14023,N_13983);
xnor U14234 (N_14234,N_14032,N_13982);
or U14235 (N_14235,N_14060,N_13931);
and U14236 (N_14236,N_13954,N_14049);
and U14237 (N_14237,N_13949,N_13922);
nand U14238 (N_14238,N_14073,N_13985);
and U14239 (N_14239,N_14046,N_13925);
nand U14240 (N_14240,N_14206,N_14157);
or U14241 (N_14241,N_14091,N_14171);
xor U14242 (N_14242,N_14092,N_14232);
xor U14243 (N_14243,N_14177,N_14194);
xnor U14244 (N_14244,N_14097,N_14188);
nand U14245 (N_14245,N_14161,N_14183);
or U14246 (N_14246,N_14208,N_14237);
and U14247 (N_14247,N_14176,N_14081);
and U14248 (N_14248,N_14121,N_14129);
or U14249 (N_14249,N_14198,N_14219);
xor U14250 (N_14250,N_14185,N_14104);
and U14251 (N_14251,N_14186,N_14153);
and U14252 (N_14252,N_14196,N_14202);
nor U14253 (N_14253,N_14162,N_14150);
or U14254 (N_14254,N_14133,N_14170);
nor U14255 (N_14255,N_14166,N_14090);
nor U14256 (N_14256,N_14189,N_14199);
and U14257 (N_14257,N_14229,N_14149);
and U14258 (N_14258,N_14126,N_14107);
or U14259 (N_14259,N_14220,N_14167);
xnor U14260 (N_14260,N_14106,N_14168);
and U14261 (N_14261,N_14083,N_14098);
nor U14262 (N_14262,N_14156,N_14148);
nor U14263 (N_14263,N_14099,N_14154);
xor U14264 (N_14264,N_14127,N_14197);
nor U14265 (N_14265,N_14173,N_14226);
or U14266 (N_14266,N_14190,N_14163);
or U14267 (N_14267,N_14096,N_14215);
and U14268 (N_14268,N_14214,N_14120);
and U14269 (N_14269,N_14174,N_14239);
nor U14270 (N_14270,N_14087,N_14200);
or U14271 (N_14271,N_14184,N_14141);
and U14272 (N_14272,N_14180,N_14195);
or U14273 (N_14273,N_14193,N_14134);
xnor U14274 (N_14274,N_14088,N_14136);
nor U14275 (N_14275,N_14231,N_14212);
nand U14276 (N_14276,N_14085,N_14109);
or U14277 (N_14277,N_14105,N_14110);
xor U14278 (N_14278,N_14086,N_14221);
and U14279 (N_14279,N_14236,N_14155);
xor U14280 (N_14280,N_14178,N_14207);
nand U14281 (N_14281,N_14204,N_14125);
or U14282 (N_14282,N_14138,N_14179);
nand U14283 (N_14283,N_14228,N_14146);
xor U14284 (N_14284,N_14147,N_14172);
or U14285 (N_14285,N_14094,N_14131);
xnor U14286 (N_14286,N_14211,N_14080);
nand U14287 (N_14287,N_14235,N_14139);
nor U14288 (N_14288,N_14218,N_14140);
nand U14289 (N_14289,N_14192,N_14113);
xnor U14290 (N_14290,N_14114,N_14234);
nor U14291 (N_14291,N_14095,N_14213);
or U14292 (N_14292,N_14209,N_14123);
nor U14293 (N_14293,N_14227,N_14160);
xnor U14294 (N_14294,N_14108,N_14143);
nand U14295 (N_14295,N_14223,N_14159);
and U14296 (N_14296,N_14158,N_14082);
xnor U14297 (N_14297,N_14205,N_14137);
nand U14298 (N_14298,N_14128,N_14175);
nand U14299 (N_14299,N_14201,N_14210);
nor U14300 (N_14300,N_14164,N_14135);
and U14301 (N_14301,N_14115,N_14238);
nor U14302 (N_14302,N_14117,N_14233);
nand U14303 (N_14303,N_14118,N_14122);
xor U14304 (N_14304,N_14181,N_14124);
nor U14305 (N_14305,N_14119,N_14116);
or U14306 (N_14306,N_14132,N_14144);
nor U14307 (N_14307,N_14089,N_14101);
nand U14308 (N_14308,N_14142,N_14112);
or U14309 (N_14309,N_14169,N_14225);
and U14310 (N_14310,N_14151,N_14187);
nand U14311 (N_14311,N_14145,N_14217);
or U14312 (N_14312,N_14103,N_14203);
nor U14313 (N_14313,N_14230,N_14111);
nand U14314 (N_14314,N_14165,N_14152);
xnor U14315 (N_14315,N_14102,N_14182);
nor U14316 (N_14316,N_14100,N_14224);
and U14317 (N_14317,N_14216,N_14222);
or U14318 (N_14318,N_14084,N_14130);
and U14319 (N_14319,N_14191,N_14093);
nor U14320 (N_14320,N_14155,N_14136);
and U14321 (N_14321,N_14089,N_14204);
nand U14322 (N_14322,N_14156,N_14129);
xor U14323 (N_14323,N_14236,N_14159);
or U14324 (N_14324,N_14125,N_14173);
nand U14325 (N_14325,N_14182,N_14171);
nand U14326 (N_14326,N_14217,N_14238);
or U14327 (N_14327,N_14199,N_14131);
nor U14328 (N_14328,N_14111,N_14173);
or U14329 (N_14329,N_14225,N_14146);
xnor U14330 (N_14330,N_14205,N_14190);
xor U14331 (N_14331,N_14192,N_14097);
or U14332 (N_14332,N_14196,N_14112);
nor U14333 (N_14333,N_14080,N_14104);
nor U14334 (N_14334,N_14151,N_14116);
nor U14335 (N_14335,N_14211,N_14173);
and U14336 (N_14336,N_14230,N_14229);
nor U14337 (N_14337,N_14156,N_14203);
nor U14338 (N_14338,N_14222,N_14160);
nand U14339 (N_14339,N_14099,N_14085);
nand U14340 (N_14340,N_14172,N_14099);
or U14341 (N_14341,N_14212,N_14184);
nor U14342 (N_14342,N_14092,N_14115);
xor U14343 (N_14343,N_14214,N_14199);
nor U14344 (N_14344,N_14192,N_14162);
or U14345 (N_14345,N_14168,N_14130);
nor U14346 (N_14346,N_14194,N_14216);
nor U14347 (N_14347,N_14100,N_14087);
nor U14348 (N_14348,N_14181,N_14205);
nand U14349 (N_14349,N_14191,N_14104);
or U14350 (N_14350,N_14153,N_14199);
xor U14351 (N_14351,N_14209,N_14235);
or U14352 (N_14352,N_14145,N_14172);
nand U14353 (N_14353,N_14124,N_14215);
or U14354 (N_14354,N_14167,N_14080);
or U14355 (N_14355,N_14154,N_14123);
xor U14356 (N_14356,N_14131,N_14133);
nor U14357 (N_14357,N_14094,N_14151);
or U14358 (N_14358,N_14182,N_14176);
xnor U14359 (N_14359,N_14230,N_14095);
nor U14360 (N_14360,N_14205,N_14090);
and U14361 (N_14361,N_14208,N_14190);
nand U14362 (N_14362,N_14108,N_14137);
or U14363 (N_14363,N_14124,N_14184);
or U14364 (N_14364,N_14140,N_14183);
or U14365 (N_14365,N_14132,N_14166);
or U14366 (N_14366,N_14082,N_14145);
nor U14367 (N_14367,N_14210,N_14083);
xnor U14368 (N_14368,N_14174,N_14125);
xnor U14369 (N_14369,N_14130,N_14233);
or U14370 (N_14370,N_14204,N_14213);
nor U14371 (N_14371,N_14191,N_14236);
xor U14372 (N_14372,N_14216,N_14160);
nand U14373 (N_14373,N_14129,N_14082);
and U14374 (N_14374,N_14221,N_14226);
nand U14375 (N_14375,N_14186,N_14127);
and U14376 (N_14376,N_14085,N_14168);
nand U14377 (N_14377,N_14153,N_14206);
nor U14378 (N_14378,N_14105,N_14141);
nor U14379 (N_14379,N_14137,N_14138);
xor U14380 (N_14380,N_14166,N_14097);
nor U14381 (N_14381,N_14223,N_14153);
nor U14382 (N_14382,N_14224,N_14211);
and U14383 (N_14383,N_14224,N_14101);
nor U14384 (N_14384,N_14093,N_14182);
or U14385 (N_14385,N_14173,N_14104);
nand U14386 (N_14386,N_14185,N_14161);
or U14387 (N_14387,N_14234,N_14112);
and U14388 (N_14388,N_14226,N_14138);
xnor U14389 (N_14389,N_14141,N_14103);
nand U14390 (N_14390,N_14181,N_14163);
or U14391 (N_14391,N_14098,N_14229);
and U14392 (N_14392,N_14234,N_14107);
nor U14393 (N_14393,N_14184,N_14136);
nor U14394 (N_14394,N_14192,N_14081);
or U14395 (N_14395,N_14145,N_14221);
xor U14396 (N_14396,N_14232,N_14093);
nand U14397 (N_14397,N_14108,N_14081);
xnor U14398 (N_14398,N_14196,N_14134);
nor U14399 (N_14399,N_14136,N_14145);
nor U14400 (N_14400,N_14258,N_14316);
or U14401 (N_14401,N_14296,N_14274);
nor U14402 (N_14402,N_14251,N_14328);
xor U14403 (N_14403,N_14397,N_14326);
xnor U14404 (N_14404,N_14351,N_14343);
and U14405 (N_14405,N_14312,N_14279);
xnor U14406 (N_14406,N_14369,N_14333);
and U14407 (N_14407,N_14280,N_14273);
nand U14408 (N_14408,N_14385,N_14281);
xnor U14409 (N_14409,N_14345,N_14347);
nand U14410 (N_14410,N_14303,N_14348);
and U14411 (N_14411,N_14310,N_14388);
and U14412 (N_14412,N_14276,N_14295);
nor U14413 (N_14413,N_14387,N_14382);
and U14414 (N_14414,N_14356,N_14308);
xnor U14415 (N_14415,N_14318,N_14257);
nand U14416 (N_14416,N_14291,N_14275);
xnor U14417 (N_14417,N_14357,N_14313);
nor U14418 (N_14418,N_14371,N_14393);
or U14419 (N_14419,N_14241,N_14368);
nand U14420 (N_14420,N_14277,N_14346);
nor U14421 (N_14421,N_14358,N_14390);
xnor U14422 (N_14422,N_14248,N_14319);
nand U14423 (N_14423,N_14270,N_14256);
or U14424 (N_14424,N_14323,N_14289);
and U14425 (N_14425,N_14342,N_14355);
nand U14426 (N_14426,N_14362,N_14272);
or U14427 (N_14427,N_14396,N_14250);
xor U14428 (N_14428,N_14389,N_14324);
nand U14429 (N_14429,N_14361,N_14314);
or U14430 (N_14430,N_14302,N_14288);
nand U14431 (N_14431,N_14254,N_14386);
xnor U14432 (N_14432,N_14244,N_14309);
and U14433 (N_14433,N_14311,N_14378);
and U14434 (N_14434,N_14344,N_14354);
xor U14435 (N_14435,N_14394,N_14320);
nor U14436 (N_14436,N_14304,N_14242);
and U14437 (N_14437,N_14322,N_14359);
nor U14438 (N_14438,N_14262,N_14253);
and U14439 (N_14439,N_14332,N_14383);
or U14440 (N_14440,N_14325,N_14297);
xnor U14441 (N_14441,N_14301,N_14375);
xnor U14442 (N_14442,N_14271,N_14287);
and U14443 (N_14443,N_14300,N_14374);
nor U14444 (N_14444,N_14370,N_14266);
nand U14445 (N_14445,N_14399,N_14284);
xnor U14446 (N_14446,N_14264,N_14364);
or U14447 (N_14447,N_14376,N_14350);
and U14448 (N_14448,N_14373,N_14377);
nand U14449 (N_14449,N_14384,N_14372);
or U14450 (N_14450,N_14391,N_14349);
xor U14451 (N_14451,N_14380,N_14298);
or U14452 (N_14452,N_14240,N_14247);
xor U14453 (N_14453,N_14363,N_14306);
or U14454 (N_14454,N_14249,N_14243);
nor U14455 (N_14455,N_14285,N_14299);
and U14456 (N_14456,N_14268,N_14398);
nor U14457 (N_14457,N_14341,N_14269);
nand U14458 (N_14458,N_14327,N_14246);
nor U14459 (N_14459,N_14365,N_14282);
and U14460 (N_14460,N_14263,N_14353);
or U14461 (N_14461,N_14330,N_14307);
nor U14462 (N_14462,N_14267,N_14252);
and U14463 (N_14463,N_14283,N_14367);
or U14464 (N_14464,N_14352,N_14360);
nand U14465 (N_14465,N_14294,N_14338);
or U14466 (N_14466,N_14337,N_14339);
xor U14467 (N_14467,N_14329,N_14331);
nand U14468 (N_14468,N_14379,N_14292);
nor U14469 (N_14469,N_14315,N_14260);
xnor U14470 (N_14470,N_14317,N_14381);
nor U14471 (N_14471,N_14265,N_14255);
xor U14472 (N_14472,N_14245,N_14395);
nor U14473 (N_14473,N_14334,N_14340);
nor U14474 (N_14474,N_14278,N_14335);
nand U14475 (N_14475,N_14336,N_14305);
nor U14476 (N_14476,N_14321,N_14366);
nand U14477 (N_14477,N_14290,N_14259);
nand U14478 (N_14478,N_14261,N_14293);
nor U14479 (N_14479,N_14286,N_14392);
xor U14480 (N_14480,N_14310,N_14272);
nand U14481 (N_14481,N_14297,N_14256);
or U14482 (N_14482,N_14358,N_14365);
nor U14483 (N_14483,N_14311,N_14348);
nor U14484 (N_14484,N_14283,N_14377);
or U14485 (N_14485,N_14363,N_14380);
nor U14486 (N_14486,N_14391,N_14329);
or U14487 (N_14487,N_14288,N_14306);
and U14488 (N_14488,N_14331,N_14294);
or U14489 (N_14489,N_14257,N_14340);
nand U14490 (N_14490,N_14398,N_14312);
xor U14491 (N_14491,N_14380,N_14320);
nand U14492 (N_14492,N_14345,N_14314);
nor U14493 (N_14493,N_14331,N_14254);
xor U14494 (N_14494,N_14331,N_14313);
and U14495 (N_14495,N_14282,N_14397);
and U14496 (N_14496,N_14288,N_14323);
nand U14497 (N_14497,N_14363,N_14368);
xor U14498 (N_14498,N_14326,N_14303);
or U14499 (N_14499,N_14255,N_14349);
nor U14500 (N_14500,N_14347,N_14302);
or U14501 (N_14501,N_14265,N_14372);
nand U14502 (N_14502,N_14323,N_14240);
or U14503 (N_14503,N_14398,N_14348);
xnor U14504 (N_14504,N_14316,N_14341);
nor U14505 (N_14505,N_14298,N_14300);
nand U14506 (N_14506,N_14372,N_14318);
xnor U14507 (N_14507,N_14372,N_14373);
xor U14508 (N_14508,N_14362,N_14382);
and U14509 (N_14509,N_14331,N_14270);
or U14510 (N_14510,N_14317,N_14298);
or U14511 (N_14511,N_14355,N_14387);
nand U14512 (N_14512,N_14241,N_14298);
nor U14513 (N_14513,N_14266,N_14330);
and U14514 (N_14514,N_14387,N_14274);
xor U14515 (N_14515,N_14307,N_14305);
xnor U14516 (N_14516,N_14257,N_14269);
nand U14517 (N_14517,N_14252,N_14284);
nor U14518 (N_14518,N_14279,N_14378);
nand U14519 (N_14519,N_14390,N_14395);
nand U14520 (N_14520,N_14263,N_14288);
or U14521 (N_14521,N_14358,N_14347);
xnor U14522 (N_14522,N_14364,N_14327);
or U14523 (N_14523,N_14362,N_14289);
nor U14524 (N_14524,N_14339,N_14262);
or U14525 (N_14525,N_14260,N_14290);
or U14526 (N_14526,N_14264,N_14291);
or U14527 (N_14527,N_14298,N_14259);
and U14528 (N_14528,N_14361,N_14358);
nand U14529 (N_14529,N_14379,N_14332);
and U14530 (N_14530,N_14245,N_14316);
or U14531 (N_14531,N_14321,N_14287);
and U14532 (N_14532,N_14307,N_14265);
or U14533 (N_14533,N_14358,N_14394);
nand U14534 (N_14534,N_14281,N_14273);
nand U14535 (N_14535,N_14321,N_14274);
or U14536 (N_14536,N_14373,N_14360);
and U14537 (N_14537,N_14315,N_14324);
xor U14538 (N_14538,N_14358,N_14375);
nor U14539 (N_14539,N_14335,N_14351);
nor U14540 (N_14540,N_14303,N_14306);
xnor U14541 (N_14541,N_14275,N_14268);
nand U14542 (N_14542,N_14308,N_14330);
and U14543 (N_14543,N_14276,N_14350);
and U14544 (N_14544,N_14368,N_14291);
nand U14545 (N_14545,N_14360,N_14377);
and U14546 (N_14546,N_14391,N_14263);
nand U14547 (N_14547,N_14246,N_14268);
nand U14548 (N_14548,N_14383,N_14359);
and U14549 (N_14549,N_14375,N_14398);
nor U14550 (N_14550,N_14243,N_14312);
xnor U14551 (N_14551,N_14321,N_14340);
nor U14552 (N_14552,N_14367,N_14333);
nand U14553 (N_14553,N_14366,N_14256);
nor U14554 (N_14554,N_14374,N_14378);
xor U14555 (N_14555,N_14331,N_14278);
xnor U14556 (N_14556,N_14255,N_14292);
nand U14557 (N_14557,N_14378,N_14337);
nand U14558 (N_14558,N_14291,N_14391);
nor U14559 (N_14559,N_14280,N_14379);
or U14560 (N_14560,N_14557,N_14488);
and U14561 (N_14561,N_14512,N_14481);
nand U14562 (N_14562,N_14539,N_14521);
or U14563 (N_14563,N_14545,N_14415);
xnor U14564 (N_14564,N_14434,N_14503);
xor U14565 (N_14565,N_14422,N_14445);
xor U14566 (N_14566,N_14556,N_14437);
nand U14567 (N_14567,N_14526,N_14507);
xor U14568 (N_14568,N_14458,N_14485);
nand U14569 (N_14569,N_14454,N_14551);
xnor U14570 (N_14570,N_14559,N_14531);
nor U14571 (N_14571,N_14524,N_14471);
and U14572 (N_14572,N_14495,N_14509);
nand U14573 (N_14573,N_14427,N_14476);
nand U14574 (N_14574,N_14525,N_14423);
and U14575 (N_14575,N_14520,N_14497);
nand U14576 (N_14576,N_14455,N_14494);
xnor U14577 (N_14577,N_14461,N_14440);
xnor U14578 (N_14578,N_14530,N_14433);
xor U14579 (N_14579,N_14432,N_14428);
xnor U14580 (N_14580,N_14438,N_14414);
and U14581 (N_14581,N_14532,N_14550);
and U14582 (N_14582,N_14417,N_14547);
and U14583 (N_14583,N_14538,N_14413);
nor U14584 (N_14584,N_14493,N_14470);
xor U14585 (N_14585,N_14500,N_14552);
and U14586 (N_14586,N_14502,N_14534);
and U14587 (N_14587,N_14501,N_14468);
and U14588 (N_14588,N_14449,N_14439);
and U14589 (N_14589,N_14490,N_14451);
nor U14590 (N_14590,N_14477,N_14448);
or U14591 (N_14591,N_14518,N_14456);
or U14592 (N_14592,N_14523,N_14499);
nor U14593 (N_14593,N_14441,N_14425);
nor U14594 (N_14594,N_14412,N_14489);
nand U14595 (N_14595,N_14513,N_14549);
nor U14596 (N_14596,N_14486,N_14558);
and U14597 (N_14597,N_14540,N_14464);
and U14598 (N_14598,N_14491,N_14444);
or U14599 (N_14599,N_14517,N_14403);
nand U14600 (N_14600,N_14407,N_14527);
nor U14601 (N_14601,N_14515,N_14400);
or U14602 (N_14602,N_14528,N_14429);
nor U14603 (N_14603,N_14506,N_14410);
nor U14604 (N_14604,N_14514,N_14483);
or U14605 (N_14605,N_14548,N_14555);
xnor U14606 (N_14606,N_14478,N_14504);
nor U14607 (N_14607,N_14474,N_14430);
nor U14608 (N_14608,N_14541,N_14505);
nor U14609 (N_14609,N_14463,N_14411);
xnor U14610 (N_14610,N_14453,N_14409);
and U14611 (N_14611,N_14492,N_14416);
and U14612 (N_14612,N_14450,N_14544);
or U14613 (N_14613,N_14508,N_14510);
xor U14614 (N_14614,N_14462,N_14546);
nand U14615 (N_14615,N_14472,N_14402);
and U14616 (N_14616,N_14479,N_14447);
and U14617 (N_14617,N_14473,N_14542);
nor U14618 (N_14618,N_14484,N_14406);
or U14619 (N_14619,N_14424,N_14419);
or U14620 (N_14620,N_14535,N_14543);
or U14621 (N_14621,N_14446,N_14460);
and U14622 (N_14622,N_14436,N_14519);
and U14623 (N_14623,N_14420,N_14553);
nor U14624 (N_14624,N_14435,N_14457);
and U14625 (N_14625,N_14480,N_14487);
or U14626 (N_14626,N_14404,N_14496);
or U14627 (N_14627,N_14469,N_14537);
xor U14628 (N_14628,N_14405,N_14421);
xor U14629 (N_14629,N_14475,N_14431);
nor U14630 (N_14630,N_14498,N_14533);
or U14631 (N_14631,N_14467,N_14443);
nor U14632 (N_14632,N_14442,N_14452);
nor U14633 (N_14633,N_14482,N_14465);
and U14634 (N_14634,N_14459,N_14466);
and U14635 (N_14635,N_14529,N_14426);
xor U14636 (N_14636,N_14554,N_14516);
nor U14637 (N_14637,N_14536,N_14522);
or U14638 (N_14638,N_14401,N_14408);
and U14639 (N_14639,N_14418,N_14511);
or U14640 (N_14640,N_14429,N_14527);
nand U14641 (N_14641,N_14537,N_14553);
and U14642 (N_14642,N_14442,N_14435);
or U14643 (N_14643,N_14451,N_14549);
nor U14644 (N_14644,N_14541,N_14409);
nor U14645 (N_14645,N_14439,N_14511);
and U14646 (N_14646,N_14405,N_14531);
or U14647 (N_14647,N_14532,N_14519);
nand U14648 (N_14648,N_14408,N_14537);
or U14649 (N_14649,N_14541,N_14493);
and U14650 (N_14650,N_14532,N_14529);
or U14651 (N_14651,N_14521,N_14555);
nand U14652 (N_14652,N_14474,N_14515);
nor U14653 (N_14653,N_14444,N_14537);
or U14654 (N_14654,N_14540,N_14461);
nor U14655 (N_14655,N_14445,N_14557);
and U14656 (N_14656,N_14444,N_14433);
xor U14657 (N_14657,N_14488,N_14449);
and U14658 (N_14658,N_14521,N_14474);
xor U14659 (N_14659,N_14520,N_14506);
or U14660 (N_14660,N_14456,N_14441);
nor U14661 (N_14661,N_14544,N_14426);
or U14662 (N_14662,N_14456,N_14527);
or U14663 (N_14663,N_14558,N_14546);
xor U14664 (N_14664,N_14447,N_14417);
nand U14665 (N_14665,N_14430,N_14519);
xnor U14666 (N_14666,N_14414,N_14441);
or U14667 (N_14667,N_14528,N_14461);
xor U14668 (N_14668,N_14547,N_14409);
or U14669 (N_14669,N_14541,N_14548);
and U14670 (N_14670,N_14449,N_14534);
and U14671 (N_14671,N_14490,N_14429);
nand U14672 (N_14672,N_14495,N_14504);
nor U14673 (N_14673,N_14415,N_14484);
nor U14674 (N_14674,N_14531,N_14472);
and U14675 (N_14675,N_14476,N_14504);
or U14676 (N_14676,N_14410,N_14432);
xor U14677 (N_14677,N_14499,N_14483);
and U14678 (N_14678,N_14429,N_14439);
and U14679 (N_14679,N_14479,N_14417);
and U14680 (N_14680,N_14441,N_14424);
and U14681 (N_14681,N_14520,N_14433);
xnor U14682 (N_14682,N_14486,N_14441);
and U14683 (N_14683,N_14519,N_14401);
nor U14684 (N_14684,N_14473,N_14556);
and U14685 (N_14685,N_14532,N_14487);
and U14686 (N_14686,N_14550,N_14545);
nand U14687 (N_14687,N_14433,N_14402);
xor U14688 (N_14688,N_14457,N_14483);
or U14689 (N_14689,N_14414,N_14470);
and U14690 (N_14690,N_14493,N_14468);
nor U14691 (N_14691,N_14509,N_14467);
xor U14692 (N_14692,N_14556,N_14513);
and U14693 (N_14693,N_14444,N_14438);
nand U14694 (N_14694,N_14445,N_14512);
nor U14695 (N_14695,N_14489,N_14520);
xor U14696 (N_14696,N_14450,N_14493);
and U14697 (N_14697,N_14505,N_14449);
or U14698 (N_14698,N_14415,N_14460);
nand U14699 (N_14699,N_14445,N_14542);
nand U14700 (N_14700,N_14421,N_14546);
and U14701 (N_14701,N_14424,N_14501);
or U14702 (N_14702,N_14403,N_14499);
and U14703 (N_14703,N_14427,N_14545);
xor U14704 (N_14704,N_14506,N_14441);
or U14705 (N_14705,N_14520,N_14455);
or U14706 (N_14706,N_14510,N_14494);
nand U14707 (N_14707,N_14515,N_14490);
nor U14708 (N_14708,N_14426,N_14424);
xor U14709 (N_14709,N_14457,N_14491);
nand U14710 (N_14710,N_14546,N_14450);
nand U14711 (N_14711,N_14504,N_14532);
nand U14712 (N_14712,N_14437,N_14527);
xnor U14713 (N_14713,N_14462,N_14412);
nor U14714 (N_14714,N_14518,N_14433);
nor U14715 (N_14715,N_14487,N_14438);
or U14716 (N_14716,N_14536,N_14537);
xor U14717 (N_14717,N_14525,N_14494);
and U14718 (N_14718,N_14462,N_14531);
nand U14719 (N_14719,N_14455,N_14420);
or U14720 (N_14720,N_14680,N_14588);
xor U14721 (N_14721,N_14631,N_14619);
xor U14722 (N_14722,N_14703,N_14614);
or U14723 (N_14723,N_14692,N_14686);
or U14724 (N_14724,N_14570,N_14673);
and U14725 (N_14725,N_14636,N_14685);
nand U14726 (N_14726,N_14564,N_14629);
nor U14727 (N_14727,N_14700,N_14571);
or U14728 (N_14728,N_14602,N_14618);
nand U14729 (N_14729,N_14649,N_14663);
nor U14730 (N_14730,N_14682,N_14711);
nor U14731 (N_14731,N_14590,N_14671);
nor U14732 (N_14732,N_14643,N_14639);
and U14733 (N_14733,N_14578,N_14708);
or U14734 (N_14734,N_14664,N_14581);
or U14735 (N_14735,N_14652,N_14647);
nor U14736 (N_14736,N_14665,N_14698);
or U14737 (N_14737,N_14568,N_14583);
nor U14738 (N_14738,N_14599,N_14580);
nor U14739 (N_14739,N_14715,N_14697);
xnor U14740 (N_14740,N_14689,N_14702);
nor U14741 (N_14741,N_14696,N_14677);
or U14742 (N_14742,N_14625,N_14662);
nor U14743 (N_14743,N_14562,N_14718);
nand U14744 (N_14744,N_14667,N_14596);
or U14745 (N_14745,N_14710,N_14719);
nor U14746 (N_14746,N_14582,N_14575);
xor U14747 (N_14747,N_14579,N_14617);
nor U14748 (N_14748,N_14714,N_14585);
nor U14749 (N_14749,N_14632,N_14678);
and U14750 (N_14750,N_14569,N_14656);
nor U14751 (N_14751,N_14597,N_14572);
nand U14752 (N_14752,N_14563,N_14676);
xnor U14753 (N_14753,N_14594,N_14699);
or U14754 (N_14754,N_14712,N_14717);
nand U14755 (N_14755,N_14616,N_14603);
xor U14756 (N_14756,N_14679,N_14574);
or U14757 (N_14757,N_14684,N_14670);
xnor U14758 (N_14758,N_14620,N_14660);
or U14759 (N_14759,N_14567,N_14648);
and U14760 (N_14760,N_14604,N_14630);
or U14761 (N_14761,N_14638,N_14654);
xnor U14762 (N_14762,N_14668,N_14659);
xor U14763 (N_14763,N_14576,N_14691);
and U14764 (N_14764,N_14657,N_14693);
or U14765 (N_14765,N_14709,N_14566);
xor U14766 (N_14766,N_14624,N_14607);
and U14767 (N_14767,N_14612,N_14672);
and U14768 (N_14768,N_14586,N_14600);
nand U14769 (N_14769,N_14611,N_14633);
and U14770 (N_14770,N_14705,N_14695);
nor U14771 (N_14771,N_14621,N_14650);
nor U14772 (N_14772,N_14615,N_14593);
nor U14773 (N_14773,N_14589,N_14669);
or U14774 (N_14774,N_14661,N_14688);
and U14775 (N_14775,N_14622,N_14584);
nand U14776 (N_14776,N_14561,N_14646);
nand U14777 (N_14777,N_14675,N_14606);
and U14778 (N_14778,N_14713,N_14626);
nand U14779 (N_14779,N_14644,N_14634);
xor U14780 (N_14780,N_14627,N_14577);
or U14781 (N_14781,N_14666,N_14706);
or U14782 (N_14782,N_14704,N_14707);
or U14783 (N_14783,N_14645,N_14674);
or U14784 (N_14784,N_14658,N_14587);
nor U14785 (N_14785,N_14655,N_14608);
xor U14786 (N_14786,N_14641,N_14601);
and U14787 (N_14787,N_14637,N_14628);
nand U14788 (N_14788,N_14605,N_14591);
nand U14789 (N_14789,N_14681,N_14653);
or U14790 (N_14790,N_14573,N_14716);
or U14791 (N_14791,N_14640,N_14701);
or U14792 (N_14792,N_14635,N_14687);
nand U14793 (N_14793,N_14623,N_14613);
and U14794 (N_14794,N_14694,N_14565);
and U14795 (N_14795,N_14690,N_14592);
or U14796 (N_14796,N_14651,N_14642);
xnor U14797 (N_14797,N_14610,N_14609);
and U14798 (N_14798,N_14560,N_14598);
or U14799 (N_14799,N_14683,N_14595);
nand U14800 (N_14800,N_14633,N_14706);
nor U14801 (N_14801,N_14711,N_14709);
xnor U14802 (N_14802,N_14597,N_14671);
xor U14803 (N_14803,N_14661,N_14669);
nor U14804 (N_14804,N_14653,N_14696);
and U14805 (N_14805,N_14648,N_14601);
and U14806 (N_14806,N_14598,N_14616);
or U14807 (N_14807,N_14575,N_14604);
nor U14808 (N_14808,N_14596,N_14615);
xnor U14809 (N_14809,N_14708,N_14629);
xor U14810 (N_14810,N_14671,N_14630);
nor U14811 (N_14811,N_14657,N_14664);
nand U14812 (N_14812,N_14671,N_14708);
nor U14813 (N_14813,N_14693,N_14700);
or U14814 (N_14814,N_14566,N_14581);
or U14815 (N_14815,N_14717,N_14622);
or U14816 (N_14816,N_14674,N_14617);
and U14817 (N_14817,N_14664,N_14623);
xor U14818 (N_14818,N_14677,N_14639);
and U14819 (N_14819,N_14618,N_14631);
or U14820 (N_14820,N_14600,N_14661);
or U14821 (N_14821,N_14627,N_14673);
and U14822 (N_14822,N_14590,N_14561);
or U14823 (N_14823,N_14653,N_14571);
nand U14824 (N_14824,N_14647,N_14637);
and U14825 (N_14825,N_14669,N_14610);
nand U14826 (N_14826,N_14618,N_14629);
xnor U14827 (N_14827,N_14647,N_14604);
or U14828 (N_14828,N_14683,N_14634);
and U14829 (N_14829,N_14657,N_14696);
nand U14830 (N_14830,N_14585,N_14685);
xnor U14831 (N_14831,N_14565,N_14681);
nand U14832 (N_14832,N_14604,N_14609);
nor U14833 (N_14833,N_14653,N_14607);
xor U14834 (N_14834,N_14579,N_14608);
nor U14835 (N_14835,N_14692,N_14647);
and U14836 (N_14836,N_14614,N_14642);
or U14837 (N_14837,N_14711,N_14671);
and U14838 (N_14838,N_14704,N_14642);
nand U14839 (N_14839,N_14625,N_14710);
nand U14840 (N_14840,N_14619,N_14583);
or U14841 (N_14841,N_14615,N_14647);
nand U14842 (N_14842,N_14719,N_14690);
or U14843 (N_14843,N_14636,N_14691);
and U14844 (N_14844,N_14572,N_14665);
or U14845 (N_14845,N_14681,N_14689);
and U14846 (N_14846,N_14639,N_14699);
xor U14847 (N_14847,N_14718,N_14618);
and U14848 (N_14848,N_14693,N_14562);
nand U14849 (N_14849,N_14692,N_14637);
and U14850 (N_14850,N_14645,N_14656);
or U14851 (N_14851,N_14695,N_14570);
nand U14852 (N_14852,N_14583,N_14656);
and U14853 (N_14853,N_14597,N_14570);
nor U14854 (N_14854,N_14616,N_14715);
and U14855 (N_14855,N_14599,N_14581);
xor U14856 (N_14856,N_14576,N_14655);
nor U14857 (N_14857,N_14695,N_14676);
nor U14858 (N_14858,N_14598,N_14610);
or U14859 (N_14859,N_14565,N_14579);
and U14860 (N_14860,N_14571,N_14636);
xnor U14861 (N_14861,N_14686,N_14625);
nand U14862 (N_14862,N_14657,N_14638);
and U14863 (N_14863,N_14617,N_14577);
nor U14864 (N_14864,N_14705,N_14594);
xnor U14865 (N_14865,N_14565,N_14677);
xnor U14866 (N_14866,N_14646,N_14587);
nor U14867 (N_14867,N_14632,N_14609);
nor U14868 (N_14868,N_14608,N_14705);
xnor U14869 (N_14869,N_14584,N_14623);
or U14870 (N_14870,N_14596,N_14608);
nand U14871 (N_14871,N_14707,N_14699);
and U14872 (N_14872,N_14628,N_14663);
and U14873 (N_14873,N_14701,N_14707);
nand U14874 (N_14874,N_14718,N_14693);
nand U14875 (N_14875,N_14605,N_14583);
or U14876 (N_14876,N_14612,N_14677);
or U14877 (N_14877,N_14663,N_14599);
or U14878 (N_14878,N_14680,N_14714);
nor U14879 (N_14879,N_14621,N_14569);
nor U14880 (N_14880,N_14738,N_14821);
xnor U14881 (N_14881,N_14816,N_14751);
xnor U14882 (N_14882,N_14830,N_14809);
or U14883 (N_14883,N_14775,N_14745);
nand U14884 (N_14884,N_14862,N_14755);
nand U14885 (N_14885,N_14824,N_14831);
and U14886 (N_14886,N_14833,N_14864);
and U14887 (N_14887,N_14777,N_14754);
and U14888 (N_14888,N_14844,N_14740);
or U14889 (N_14889,N_14855,N_14759);
xnor U14890 (N_14890,N_14868,N_14849);
nand U14891 (N_14891,N_14869,N_14765);
nand U14892 (N_14892,N_14865,N_14763);
xnor U14893 (N_14893,N_14805,N_14877);
or U14894 (N_14894,N_14787,N_14792);
xnor U14895 (N_14895,N_14747,N_14720);
and U14896 (N_14896,N_14825,N_14814);
or U14897 (N_14897,N_14871,N_14803);
nand U14898 (N_14898,N_14790,N_14737);
xor U14899 (N_14899,N_14772,N_14863);
nand U14900 (N_14900,N_14807,N_14750);
or U14901 (N_14901,N_14776,N_14866);
and U14902 (N_14902,N_14749,N_14723);
xor U14903 (N_14903,N_14734,N_14732);
nand U14904 (N_14904,N_14843,N_14736);
and U14905 (N_14905,N_14794,N_14757);
and U14906 (N_14906,N_14832,N_14857);
xnor U14907 (N_14907,N_14852,N_14822);
and U14908 (N_14908,N_14823,N_14768);
nand U14909 (N_14909,N_14743,N_14742);
nand U14910 (N_14910,N_14771,N_14836);
and U14911 (N_14911,N_14834,N_14806);
xor U14912 (N_14912,N_14724,N_14813);
and U14913 (N_14913,N_14756,N_14791);
nand U14914 (N_14914,N_14785,N_14876);
nor U14915 (N_14915,N_14827,N_14867);
nand U14916 (N_14916,N_14727,N_14878);
nand U14917 (N_14917,N_14829,N_14762);
nand U14918 (N_14918,N_14782,N_14860);
xnor U14919 (N_14919,N_14808,N_14845);
nor U14920 (N_14920,N_14797,N_14722);
or U14921 (N_14921,N_14744,N_14850);
nor U14922 (N_14922,N_14766,N_14815);
or U14923 (N_14923,N_14870,N_14798);
or U14924 (N_14924,N_14841,N_14802);
nor U14925 (N_14925,N_14826,N_14801);
nor U14926 (N_14926,N_14856,N_14793);
nand U14927 (N_14927,N_14858,N_14764);
nor U14928 (N_14928,N_14835,N_14781);
nor U14929 (N_14929,N_14861,N_14872);
or U14930 (N_14930,N_14770,N_14767);
xnor U14931 (N_14931,N_14859,N_14739);
and U14932 (N_14932,N_14774,N_14758);
and U14933 (N_14933,N_14840,N_14753);
or U14934 (N_14934,N_14788,N_14819);
xor U14935 (N_14935,N_14741,N_14847);
nor U14936 (N_14936,N_14726,N_14760);
or U14937 (N_14937,N_14800,N_14789);
xnor U14938 (N_14938,N_14804,N_14853);
nor U14939 (N_14939,N_14799,N_14731);
nor U14940 (N_14940,N_14851,N_14879);
and U14941 (N_14941,N_14773,N_14735);
or U14942 (N_14942,N_14796,N_14780);
nand U14943 (N_14943,N_14846,N_14779);
or U14944 (N_14944,N_14784,N_14818);
and U14945 (N_14945,N_14786,N_14875);
and U14946 (N_14946,N_14778,N_14842);
nand U14947 (N_14947,N_14761,N_14728);
nand U14948 (N_14948,N_14873,N_14874);
xnor U14949 (N_14949,N_14795,N_14729);
xnor U14950 (N_14950,N_14810,N_14828);
and U14951 (N_14951,N_14820,N_14838);
nor U14952 (N_14952,N_14752,N_14848);
nand U14953 (N_14953,N_14817,N_14839);
nor U14954 (N_14954,N_14812,N_14854);
or U14955 (N_14955,N_14725,N_14837);
xnor U14956 (N_14956,N_14733,N_14748);
nand U14957 (N_14957,N_14769,N_14746);
nand U14958 (N_14958,N_14811,N_14721);
nor U14959 (N_14959,N_14730,N_14783);
and U14960 (N_14960,N_14863,N_14832);
nand U14961 (N_14961,N_14848,N_14870);
nor U14962 (N_14962,N_14753,N_14805);
nand U14963 (N_14963,N_14850,N_14786);
nand U14964 (N_14964,N_14769,N_14862);
or U14965 (N_14965,N_14738,N_14822);
nand U14966 (N_14966,N_14835,N_14833);
nand U14967 (N_14967,N_14817,N_14828);
xnor U14968 (N_14968,N_14817,N_14794);
and U14969 (N_14969,N_14739,N_14811);
nor U14970 (N_14970,N_14752,N_14776);
nor U14971 (N_14971,N_14769,N_14825);
and U14972 (N_14972,N_14872,N_14808);
xnor U14973 (N_14973,N_14770,N_14769);
or U14974 (N_14974,N_14757,N_14777);
and U14975 (N_14975,N_14827,N_14754);
nand U14976 (N_14976,N_14777,N_14854);
or U14977 (N_14977,N_14846,N_14720);
nor U14978 (N_14978,N_14746,N_14805);
nand U14979 (N_14979,N_14836,N_14797);
or U14980 (N_14980,N_14879,N_14771);
or U14981 (N_14981,N_14869,N_14777);
nor U14982 (N_14982,N_14742,N_14780);
xnor U14983 (N_14983,N_14866,N_14752);
nor U14984 (N_14984,N_14861,N_14868);
nand U14985 (N_14985,N_14865,N_14757);
xnor U14986 (N_14986,N_14804,N_14797);
and U14987 (N_14987,N_14749,N_14801);
or U14988 (N_14988,N_14735,N_14781);
or U14989 (N_14989,N_14754,N_14815);
nand U14990 (N_14990,N_14801,N_14823);
or U14991 (N_14991,N_14811,N_14785);
or U14992 (N_14992,N_14779,N_14830);
nor U14993 (N_14993,N_14859,N_14854);
xnor U14994 (N_14994,N_14757,N_14721);
nor U14995 (N_14995,N_14732,N_14792);
and U14996 (N_14996,N_14810,N_14815);
nor U14997 (N_14997,N_14750,N_14759);
or U14998 (N_14998,N_14784,N_14750);
nor U14999 (N_14999,N_14773,N_14850);
nand U15000 (N_15000,N_14789,N_14775);
and U15001 (N_15001,N_14732,N_14766);
xnor U15002 (N_15002,N_14800,N_14757);
or U15003 (N_15003,N_14814,N_14847);
or U15004 (N_15004,N_14740,N_14759);
nand U15005 (N_15005,N_14821,N_14878);
or U15006 (N_15006,N_14787,N_14865);
nor U15007 (N_15007,N_14869,N_14726);
nor U15008 (N_15008,N_14836,N_14721);
or U15009 (N_15009,N_14841,N_14758);
nor U15010 (N_15010,N_14785,N_14803);
xnor U15011 (N_15011,N_14846,N_14816);
xnor U15012 (N_15012,N_14756,N_14812);
nor U15013 (N_15013,N_14745,N_14853);
and U15014 (N_15014,N_14865,N_14870);
xnor U15015 (N_15015,N_14728,N_14731);
nand U15016 (N_15016,N_14833,N_14848);
nand U15017 (N_15017,N_14828,N_14827);
nand U15018 (N_15018,N_14809,N_14775);
or U15019 (N_15019,N_14851,N_14776);
nor U15020 (N_15020,N_14722,N_14738);
or U15021 (N_15021,N_14751,N_14835);
and U15022 (N_15022,N_14758,N_14844);
or U15023 (N_15023,N_14813,N_14859);
nand U15024 (N_15024,N_14738,N_14772);
xnor U15025 (N_15025,N_14729,N_14841);
xor U15026 (N_15026,N_14784,N_14832);
xor U15027 (N_15027,N_14796,N_14799);
nand U15028 (N_15028,N_14756,N_14855);
or U15029 (N_15029,N_14779,N_14820);
and U15030 (N_15030,N_14766,N_14819);
nor U15031 (N_15031,N_14846,N_14787);
and U15032 (N_15032,N_14736,N_14859);
and U15033 (N_15033,N_14837,N_14755);
or U15034 (N_15034,N_14733,N_14761);
nor U15035 (N_15035,N_14845,N_14721);
and U15036 (N_15036,N_14723,N_14867);
nand U15037 (N_15037,N_14839,N_14826);
xnor U15038 (N_15038,N_14771,N_14736);
xnor U15039 (N_15039,N_14835,N_14792);
nor U15040 (N_15040,N_14887,N_15039);
and U15041 (N_15041,N_14989,N_15032);
xor U15042 (N_15042,N_14931,N_15006);
nand U15043 (N_15043,N_14995,N_14913);
nand U15044 (N_15044,N_14891,N_14990);
nand U15045 (N_15045,N_14934,N_14881);
or U15046 (N_15046,N_14986,N_15014);
or U15047 (N_15047,N_14912,N_15000);
xnor U15048 (N_15048,N_14978,N_14972);
or U15049 (N_15049,N_15024,N_15010);
and U15050 (N_15050,N_14946,N_14938);
xor U15051 (N_15051,N_14927,N_14994);
xnor U15052 (N_15052,N_14922,N_15022);
nand U15053 (N_15053,N_15003,N_14999);
xnor U15054 (N_15054,N_15035,N_15015);
and U15055 (N_15055,N_14958,N_14925);
or U15056 (N_15056,N_14955,N_14949);
nor U15057 (N_15057,N_14880,N_14899);
nor U15058 (N_15058,N_14945,N_14983);
xor U15059 (N_15059,N_14906,N_14971);
or U15060 (N_15060,N_14884,N_15038);
xnor U15061 (N_15061,N_14905,N_15019);
or U15062 (N_15062,N_14897,N_14997);
nand U15063 (N_15063,N_14982,N_14892);
xor U15064 (N_15064,N_14943,N_14885);
nand U15065 (N_15065,N_15020,N_14962);
xor U15066 (N_15066,N_14967,N_14993);
nor U15067 (N_15067,N_14957,N_14920);
nor U15068 (N_15068,N_14987,N_14919);
nor U15069 (N_15069,N_14902,N_14903);
nand U15070 (N_15070,N_15004,N_15030);
nand U15071 (N_15071,N_14965,N_14923);
nand U15072 (N_15072,N_14896,N_14947);
or U15073 (N_15073,N_14939,N_14954);
nand U15074 (N_15074,N_15001,N_15028);
and U15075 (N_15075,N_14904,N_14964);
or U15076 (N_15076,N_14911,N_15002);
xnor U15077 (N_15077,N_14936,N_14952);
nor U15078 (N_15078,N_15036,N_14966);
or U15079 (N_15079,N_14914,N_14969);
xor U15080 (N_15080,N_14948,N_14998);
or U15081 (N_15081,N_15008,N_14981);
xnor U15082 (N_15082,N_14980,N_14932);
or U15083 (N_15083,N_14973,N_15016);
and U15084 (N_15084,N_14890,N_14907);
nor U15085 (N_15085,N_15009,N_14960);
nor U15086 (N_15086,N_15037,N_14956);
or U15087 (N_15087,N_14895,N_14910);
or U15088 (N_15088,N_14928,N_14886);
and U15089 (N_15089,N_14942,N_14883);
or U15090 (N_15090,N_14889,N_14894);
and U15091 (N_15091,N_14926,N_14963);
xnor U15092 (N_15092,N_14900,N_15029);
and U15093 (N_15093,N_14970,N_14898);
or U15094 (N_15094,N_14968,N_14916);
and U15095 (N_15095,N_15021,N_14941);
and U15096 (N_15096,N_14901,N_14933);
or U15097 (N_15097,N_14930,N_14996);
xnor U15098 (N_15098,N_14924,N_15031);
or U15099 (N_15099,N_14959,N_14888);
nand U15100 (N_15100,N_14893,N_14940);
and U15101 (N_15101,N_14929,N_14984);
nand U15102 (N_15102,N_15005,N_14992);
nor U15103 (N_15103,N_15027,N_15012);
or U15104 (N_15104,N_14953,N_15023);
and U15105 (N_15105,N_15018,N_14976);
xor U15106 (N_15106,N_14951,N_14937);
nor U15107 (N_15107,N_14935,N_14961);
xnor U15108 (N_15108,N_15017,N_14915);
xnor U15109 (N_15109,N_14975,N_14944);
and U15110 (N_15110,N_14988,N_15007);
nand U15111 (N_15111,N_15026,N_15025);
nor U15112 (N_15112,N_15034,N_14977);
and U15113 (N_15113,N_14917,N_15033);
and U15114 (N_15114,N_15013,N_14974);
nand U15115 (N_15115,N_14950,N_14882);
nor U15116 (N_15116,N_14908,N_15011);
nand U15117 (N_15117,N_14918,N_14985);
nand U15118 (N_15118,N_14909,N_14991);
nor U15119 (N_15119,N_14979,N_14921);
and U15120 (N_15120,N_14950,N_14889);
xnor U15121 (N_15121,N_14882,N_14957);
and U15122 (N_15122,N_14988,N_14981);
nor U15123 (N_15123,N_14933,N_14946);
or U15124 (N_15124,N_14911,N_14905);
nand U15125 (N_15125,N_14883,N_14887);
and U15126 (N_15126,N_14958,N_14938);
and U15127 (N_15127,N_14976,N_14924);
or U15128 (N_15128,N_14909,N_14992);
and U15129 (N_15129,N_15011,N_14992);
and U15130 (N_15130,N_14967,N_14880);
or U15131 (N_15131,N_14930,N_14927);
and U15132 (N_15132,N_14928,N_14896);
and U15133 (N_15133,N_14940,N_14977);
or U15134 (N_15134,N_14909,N_14997);
xnor U15135 (N_15135,N_15003,N_14934);
xor U15136 (N_15136,N_14985,N_14984);
nand U15137 (N_15137,N_14979,N_14944);
nand U15138 (N_15138,N_14990,N_14906);
xor U15139 (N_15139,N_14886,N_14963);
or U15140 (N_15140,N_14883,N_14937);
xnor U15141 (N_15141,N_14923,N_15022);
nor U15142 (N_15142,N_14900,N_14927);
nand U15143 (N_15143,N_14882,N_14904);
or U15144 (N_15144,N_14989,N_14993);
and U15145 (N_15145,N_14919,N_14948);
nor U15146 (N_15146,N_14931,N_14950);
or U15147 (N_15147,N_15037,N_14955);
nor U15148 (N_15148,N_14908,N_14885);
nand U15149 (N_15149,N_14985,N_15018);
nor U15150 (N_15150,N_14932,N_14952);
nor U15151 (N_15151,N_14965,N_14948);
nor U15152 (N_15152,N_14991,N_14952);
nor U15153 (N_15153,N_14997,N_14967);
nor U15154 (N_15154,N_14922,N_14989);
xnor U15155 (N_15155,N_14930,N_15008);
and U15156 (N_15156,N_14955,N_15015);
or U15157 (N_15157,N_15009,N_15010);
and U15158 (N_15158,N_15015,N_15016);
nand U15159 (N_15159,N_14915,N_14901);
xor U15160 (N_15160,N_15015,N_15019);
nand U15161 (N_15161,N_15006,N_14885);
or U15162 (N_15162,N_14948,N_14985);
and U15163 (N_15163,N_14924,N_14986);
nand U15164 (N_15164,N_14996,N_14955);
nand U15165 (N_15165,N_15016,N_14983);
or U15166 (N_15166,N_15025,N_14977);
nor U15167 (N_15167,N_14907,N_14971);
nand U15168 (N_15168,N_14926,N_15033);
and U15169 (N_15169,N_15016,N_14901);
and U15170 (N_15170,N_14985,N_14908);
nor U15171 (N_15171,N_14973,N_14931);
nor U15172 (N_15172,N_14951,N_15030);
nand U15173 (N_15173,N_14967,N_14881);
or U15174 (N_15174,N_14947,N_14953);
xor U15175 (N_15175,N_14968,N_14922);
and U15176 (N_15176,N_14896,N_14924);
nor U15177 (N_15177,N_14925,N_14977);
xor U15178 (N_15178,N_14923,N_14995);
and U15179 (N_15179,N_14928,N_14964);
nor U15180 (N_15180,N_14919,N_14915);
or U15181 (N_15181,N_14939,N_14932);
nand U15182 (N_15182,N_14955,N_14975);
or U15183 (N_15183,N_14987,N_14904);
nor U15184 (N_15184,N_15015,N_14945);
xor U15185 (N_15185,N_15035,N_14988);
nor U15186 (N_15186,N_14980,N_14969);
xor U15187 (N_15187,N_14886,N_15008);
nand U15188 (N_15188,N_14907,N_14996);
and U15189 (N_15189,N_15030,N_14977);
xor U15190 (N_15190,N_15008,N_15025);
or U15191 (N_15191,N_15012,N_14990);
and U15192 (N_15192,N_14977,N_14907);
xnor U15193 (N_15193,N_14881,N_14922);
or U15194 (N_15194,N_14941,N_14974);
nor U15195 (N_15195,N_14935,N_15032);
or U15196 (N_15196,N_15008,N_14972);
nor U15197 (N_15197,N_14897,N_14925);
or U15198 (N_15198,N_14901,N_14965);
xnor U15199 (N_15199,N_15005,N_14926);
and U15200 (N_15200,N_15056,N_15069);
nor U15201 (N_15201,N_15085,N_15132);
and U15202 (N_15202,N_15109,N_15175);
or U15203 (N_15203,N_15139,N_15179);
nand U15204 (N_15204,N_15187,N_15077);
xor U15205 (N_15205,N_15090,N_15197);
nand U15206 (N_15206,N_15159,N_15119);
xnor U15207 (N_15207,N_15093,N_15165);
xor U15208 (N_15208,N_15078,N_15071);
and U15209 (N_15209,N_15082,N_15100);
nand U15210 (N_15210,N_15174,N_15063);
nand U15211 (N_15211,N_15150,N_15134);
nor U15212 (N_15212,N_15041,N_15108);
nor U15213 (N_15213,N_15199,N_15182);
nand U15214 (N_15214,N_15146,N_15044);
nor U15215 (N_15215,N_15130,N_15147);
or U15216 (N_15216,N_15181,N_15194);
and U15217 (N_15217,N_15042,N_15114);
nand U15218 (N_15218,N_15178,N_15050);
nor U15219 (N_15219,N_15047,N_15158);
or U15220 (N_15220,N_15127,N_15117);
and U15221 (N_15221,N_15048,N_15155);
nor U15222 (N_15222,N_15188,N_15148);
and U15223 (N_15223,N_15123,N_15052);
xnor U15224 (N_15224,N_15040,N_15136);
nor U15225 (N_15225,N_15133,N_15166);
xnor U15226 (N_15226,N_15060,N_15170);
nand U15227 (N_15227,N_15157,N_15124);
nor U15228 (N_15228,N_15092,N_15125);
nand U15229 (N_15229,N_15081,N_15099);
nor U15230 (N_15230,N_15137,N_15111);
nand U15231 (N_15231,N_15173,N_15152);
nand U15232 (N_15232,N_15183,N_15054);
or U15233 (N_15233,N_15043,N_15172);
nand U15234 (N_15234,N_15186,N_15189);
xor U15235 (N_15235,N_15107,N_15084);
nand U15236 (N_15236,N_15129,N_15121);
and U15237 (N_15237,N_15167,N_15191);
and U15238 (N_15238,N_15154,N_15110);
nand U15239 (N_15239,N_15074,N_15196);
nand U15240 (N_15240,N_15120,N_15102);
and U15241 (N_15241,N_15195,N_15138);
or U15242 (N_15242,N_15091,N_15051);
xor U15243 (N_15243,N_15104,N_15087);
and U15244 (N_15244,N_15103,N_15122);
xor U15245 (N_15245,N_15067,N_15145);
nor U15246 (N_15246,N_15094,N_15143);
nand U15247 (N_15247,N_15112,N_15079);
nand U15248 (N_15248,N_15068,N_15177);
or U15249 (N_15249,N_15126,N_15180);
nor U15250 (N_15250,N_15062,N_15171);
nor U15251 (N_15251,N_15151,N_15176);
nor U15252 (N_15252,N_15080,N_15089);
xor U15253 (N_15253,N_15131,N_15190);
xor U15254 (N_15254,N_15163,N_15113);
nor U15255 (N_15255,N_15073,N_15193);
xor U15256 (N_15256,N_15061,N_15192);
or U15257 (N_15257,N_15198,N_15164);
or U15258 (N_15258,N_15064,N_15115);
and U15259 (N_15259,N_15098,N_15184);
xor U15260 (N_15260,N_15160,N_15140);
nor U15261 (N_15261,N_15095,N_15053);
and U15262 (N_15262,N_15141,N_15070);
nor U15263 (N_15263,N_15116,N_15144);
or U15264 (N_15264,N_15066,N_15083);
and U15265 (N_15265,N_15156,N_15169);
nand U15266 (N_15266,N_15161,N_15168);
xor U15267 (N_15267,N_15065,N_15162);
nor U15268 (N_15268,N_15153,N_15059);
nor U15269 (N_15269,N_15045,N_15118);
nor U15270 (N_15270,N_15142,N_15046);
xnor U15271 (N_15271,N_15149,N_15106);
and U15272 (N_15272,N_15105,N_15096);
or U15273 (N_15273,N_15076,N_15185);
xor U15274 (N_15274,N_15101,N_15072);
and U15275 (N_15275,N_15135,N_15088);
or U15276 (N_15276,N_15055,N_15128);
or U15277 (N_15277,N_15097,N_15058);
or U15278 (N_15278,N_15057,N_15049);
nand U15279 (N_15279,N_15075,N_15086);
xnor U15280 (N_15280,N_15186,N_15147);
nor U15281 (N_15281,N_15075,N_15193);
nor U15282 (N_15282,N_15193,N_15040);
xor U15283 (N_15283,N_15045,N_15091);
or U15284 (N_15284,N_15097,N_15170);
xnor U15285 (N_15285,N_15171,N_15094);
nand U15286 (N_15286,N_15052,N_15154);
nor U15287 (N_15287,N_15180,N_15087);
nor U15288 (N_15288,N_15088,N_15148);
nor U15289 (N_15289,N_15150,N_15131);
nand U15290 (N_15290,N_15174,N_15152);
or U15291 (N_15291,N_15112,N_15052);
and U15292 (N_15292,N_15045,N_15051);
and U15293 (N_15293,N_15177,N_15181);
nand U15294 (N_15294,N_15046,N_15193);
or U15295 (N_15295,N_15167,N_15119);
nor U15296 (N_15296,N_15042,N_15072);
nand U15297 (N_15297,N_15064,N_15043);
nand U15298 (N_15298,N_15088,N_15066);
xor U15299 (N_15299,N_15140,N_15091);
nor U15300 (N_15300,N_15093,N_15100);
xnor U15301 (N_15301,N_15056,N_15170);
and U15302 (N_15302,N_15174,N_15116);
xnor U15303 (N_15303,N_15185,N_15115);
nand U15304 (N_15304,N_15165,N_15159);
nand U15305 (N_15305,N_15172,N_15118);
or U15306 (N_15306,N_15163,N_15072);
or U15307 (N_15307,N_15109,N_15156);
or U15308 (N_15308,N_15173,N_15110);
xnor U15309 (N_15309,N_15191,N_15047);
or U15310 (N_15310,N_15068,N_15122);
and U15311 (N_15311,N_15079,N_15196);
nand U15312 (N_15312,N_15104,N_15130);
xnor U15313 (N_15313,N_15068,N_15073);
xor U15314 (N_15314,N_15119,N_15168);
nand U15315 (N_15315,N_15185,N_15136);
nor U15316 (N_15316,N_15185,N_15057);
nand U15317 (N_15317,N_15105,N_15050);
or U15318 (N_15318,N_15100,N_15119);
nor U15319 (N_15319,N_15052,N_15124);
and U15320 (N_15320,N_15050,N_15042);
xnor U15321 (N_15321,N_15162,N_15079);
and U15322 (N_15322,N_15151,N_15080);
and U15323 (N_15323,N_15173,N_15179);
or U15324 (N_15324,N_15144,N_15163);
or U15325 (N_15325,N_15108,N_15186);
xor U15326 (N_15326,N_15162,N_15121);
and U15327 (N_15327,N_15049,N_15151);
xnor U15328 (N_15328,N_15070,N_15184);
nor U15329 (N_15329,N_15160,N_15149);
and U15330 (N_15330,N_15051,N_15154);
or U15331 (N_15331,N_15133,N_15096);
and U15332 (N_15332,N_15155,N_15127);
nor U15333 (N_15333,N_15159,N_15055);
nor U15334 (N_15334,N_15186,N_15110);
or U15335 (N_15335,N_15117,N_15152);
and U15336 (N_15336,N_15160,N_15094);
or U15337 (N_15337,N_15134,N_15082);
or U15338 (N_15338,N_15107,N_15067);
and U15339 (N_15339,N_15173,N_15071);
nor U15340 (N_15340,N_15145,N_15170);
and U15341 (N_15341,N_15057,N_15180);
xor U15342 (N_15342,N_15178,N_15129);
nand U15343 (N_15343,N_15046,N_15188);
or U15344 (N_15344,N_15194,N_15152);
nor U15345 (N_15345,N_15138,N_15082);
and U15346 (N_15346,N_15109,N_15108);
xor U15347 (N_15347,N_15163,N_15185);
nand U15348 (N_15348,N_15194,N_15189);
or U15349 (N_15349,N_15097,N_15057);
xnor U15350 (N_15350,N_15149,N_15096);
nor U15351 (N_15351,N_15141,N_15154);
xor U15352 (N_15352,N_15128,N_15085);
nand U15353 (N_15353,N_15129,N_15103);
nand U15354 (N_15354,N_15048,N_15129);
nor U15355 (N_15355,N_15051,N_15098);
and U15356 (N_15356,N_15112,N_15181);
xor U15357 (N_15357,N_15069,N_15161);
or U15358 (N_15358,N_15162,N_15198);
or U15359 (N_15359,N_15198,N_15113);
nor U15360 (N_15360,N_15254,N_15287);
nand U15361 (N_15361,N_15313,N_15256);
or U15362 (N_15362,N_15317,N_15329);
or U15363 (N_15363,N_15326,N_15239);
or U15364 (N_15364,N_15301,N_15358);
nand U15365 (N_15365,N_15248,N_15316);
nand U15366 (N_15366,N_15359,N_15200);
xor U15367 (N_15367,N_15344,N_15240);
xor U15368 (N_15368,N_15349,N_15201);
nand U15369 (N_15369,N_15230,N_15224);
nand U15370 (N_15370,N_15289,N_15333);
nor U15371 (N_15371,N_15261,N_15241);
or U15372 (N_15372,N_15236,N_15281);
nor U15373 (N_15373,N_15343,N_15304);
or U15374 (N_15374,N_15257,N_15214);
or U15375 (N_15375,N_15271,N_15314);
and U15376 (N_15376,N_15217,N_15250);
nor U15377 (N_15377,N_15235,N_15307);
xnor U15378 (N_15378,N_15219,N_15288);
xnor U15379 (N_15379,N_15290,N_15232);
or U15380 (N_15380,N_15345,N_15267);
nand U15381 (N_15381,N_15223,N_15296);
or U15382 (N_15382,N_15251,N_15341);
or U15383 (N_15383,N_15202,N_15286);
xnor U15384 (N_15384,N_15342,N_15302);
xor U15385 (N_15385,N_15243,N_15218);
nor U15386 (N_15386,N_15348,N_15300);
nand U15387 (N_15387,N_15221,N_15279);
xor U15388 (N_15388,N_15322,N_15228);
nand U15389 (N_15389,N_15208,N_15244);
xor U15390 (N_15390,N_15350,N_15278);
nand U15391 (N_15391,N_15211,N_15245);
xor U15392 (N_15392,N_15310,N_15273);
nor U15393 (N_15393,N_15233,N_15357);
or U15394 (N_15394,N_15203,N_15274);
xnor U15395 (N_15395,N_15294,N_15249);
and U15396 (N_15396,N_15353,N_15298);
or U15397 (N_15397,N_15285,N_15325);
nor U15398 (N_15398,N_15283,N_15258);
nor U15399 (N_15399,N_15204,N_15277);
nand U15400 (N_15400,N_15297,N_15226);
nor U15401 (N_15401,N_15276,N_15265);
or U15402 (N_15402,N_15275,N_15242);
nor U15403 (N_15403,N_15334,N_15324);
xor U15404 (N_15404,N_15282,N_15262);
xnor U15405 (N_15405,N_15321,N_15237);
or U15406 (N_15406,N_15253,N_15319);
nand U15407 (N_15407,N_15227,N_15337);
nor U15408 (N_15408,N_15209,N_15260);
nand U15409 (N_15409,N_15303,N_15330);
nand U15410 (N_15410,N_15340,N_15293);
and U15411 (N_15411,N_15263,N_15323);
nand U15412 (N_15412,N_15335,N_15354);
and U15413 (N_15413,N_15247,N_15234);
nor U15414 (N_15414,N_15306,N_15331);
nand U15415 (N_15415,N_15339,N_15222);
nand U15416 (N_15416,N_15338,N_15205);
xnor U15417 (N_15417,N_15212,N_15272);
or U15418 (N_15418,N_15246,N_15320);
nor U15419 (N_15419,N_15327,N_15280);
and U15420 (N_15420,N_15231,N_15206);
nand U15421 (N_15421,N_15291,N_15238);
nand U15422 (N_15422,N_15336,N_15346);
nor U15423 (N_15423,N_15215,N_15355);
or U15424 (N_15424,N_15229,N_15352);
and U15425 (N_15425,N_15351,N_15347);
and U15426 (N_15426,N_15213,N_15356);
nor U15427 (N_15427,N_15259,N_15315);
xnor U15428 (N_15428,N_15225,N_15270);
xor U15429 (N_15429,N_15207,N_15308);
nand U15430 (N_15430,N_15268,N_15266);
or U15431 (N_15431,N_15299,N_15305);
nand U15432 (N_15432,N_15311,N_15312);
nand U15433 (N_15433,N_15210,N_15264);
or U15434 (N_15434,N_15328,N_15332);
nor U15435 (N_15435,N_15295,N_15220);
nor U15436 (N_15436,N_15284,N_15318);
xor U15437 (N_15437,N_15292,N_15255);
nand U15438 (N_15438,N_15252,N_15269);
and U15439 (N_15439,N_15309,N_15216);
nor U15440 (N_15440,N_15263,N_15288);
or U15441 (N_15441,N_15336,N_15318);
nand U15442 (N_15442,N_15331,N_15241);
and U15443 (N_15443,N_15265,N_15252);
and U15444 (N_15444,N_15337,N_15256);
and U15445 (N_15445,N_15218,N_15297);
or U15446 (N_15446,N_15216,N_15226);
nand U15447 (N_15447,N_15342,N_15329);
nor U15448 (N_15448,N_15243,N_15211);
nor U15449 (N_15449,N_15213,N_15302);
nand U15450 (N_15450,N_15306,N_15268);
nor U15451 (N_15451,N_15319,N_15226);
xnor U15452 (N_15452,N_15358,N_15276);
nor U15453 (N_15453,N_15350,N_15210);
nor U15454 (N_15454,N_15244,N_15240);
nor U15455 (N_15455,N_15326,N_15253);
xor U15456 (N_15456,N_15340,N_15290);
xnor U15457 (N_15457,N_15230,N_15342);
xnor U15458 (N_15458,N_15239,N_15296);
or U15459 (N_15459,N_15291,N_15208);
nand U15460 (N_15460,N_15340,N_15355);
and U15461 (N_15461,N_15286,N_15236);
and U15462 (N_15462,N_15324,N_15323);
nand U15463 (N_15463,N_15336,N_15347);
xor U15464 (N_15464,N_15286,N_15203);
or U15465 (N_15465,N_15253,N_15337);
nand U15466 (N_15466,N_15318,N_15202);
xor U15467 (N_15467,N_15348,N_15325);
or U15468 (N_15468,N_15319,N_15222);
nor U15469 (N_15469,N_15303,N_15233);
and U15470 (N_15470,N_15294,N_15237);
or U15471 (N_15471,N_15299,N_15255);
nor U15472 (N_15472,N_15350,N_15216);
nor U15473 (N_15473,N_15231,N_15247);
and U15474 (N_15474,N_15202,N_15273);
and U15475 (N_15475,N_15342,N_15327);
nand U15476 (N_15476,N_15285,N_15275);
and U15477 (N_15477,N_15295,N_15311);
or U15478 (N_15478,N_15333,N_15306);
nand U15479 (N_15479,N_15340,N_15246);
or U15480 (N_15480,N_15303,N_15209);
and U15481 (N_15481,N_15286,N_15271);
xor U15482 (N_15482,N_15349,N_15204);
nand U15483 (N_15483,N_15346,N_15222);
nor U15484 (N_15484,N_15250,N_15206);
nand U15485 (N_15485,N_15252,N_15221);
and U15486 (N_15486,N_15327,N_15274);
or U15487 (N_15487,N_15349,N_15209);
xnor U15488 (N_15488,N_15302,N_15222);
xor U15489 (N_15489,N_15249,N_15340);
or U15490 (N_15490,N_15229,N_15323);
xnor U15491 (N_15491,N_15324,N_15317);
or U15492 (N_15492,N_15225,N_15262);
or U15493 (N_15493,N_15352,N_15269);
and U15494 (N_15494,N_15326,N_15292);
nor U15495 (N_15495,N_15312,N_15300);
nor U15496 (N_15496,N_15327,N_15303);
and U15497 (N_15497,N_15297,N_15295);
nor U15498 (N_15498,N_15229,N_15216);
nor U15499 (N_15499,N_15220,N_15276);
nor U15500 (N_15500,N_15342,N_15236);
and U15501 (N_15501,N_15348,N_15205);
xor U15502 (N_15502,N_15284,N_15313);
nand U15503 (N_15503,N_15311,N_15304);
nand U15504 (N_15504,N_15297,N_15261);
or U15505 (N_15505,N_15265,N_15309);
nor U15506 (N_15506,N_15233,N_15247);
and U15507 (N_15507,N_15207,N_15246);
nand U15508 (N_15508,N_15303,N_15286);
xor U15509 (N_15509,N_15291,N_15247);
nand U15510 (N_15510,N_15272,N_15283);
nand U15511 (N_15511,N_15265,N_15227);
xor U15512 (N_15512,N_15224,N_15220);
or U15513 (N_15513,N_15208,N_15212);
and U15514 (N_15514,N_15342,N_15309);
and U15515 (N_15515,N_15220,N_15300);
nor U15516 (N_15516,N_15340,N_15348);
xnor U15517 (N_15517,N_15215,N_15258);
or U15518 (N_15518,N_15222,N_15326);
xor U15519 (N_15519,N_15290,N_15272);
and U15520 (N_15520,N_15499,N_15456);
nand U15521 (N_15521,N_15360,N_15408);
and U15522 (N_15522,N_15392,N_15422);
xor U15523 (N_15523,N_15469,N_15470);
nand U15524 (N_15524,N_15486,N_15425);
nand U15525 (N_15525,N_15375,N_15516);
nor U15526 (N_15526,N_15447,N_15517);
xnor U15527 (N_15527,N_15501,N_15439);
xor U15528 (N_15528,N_15423,N_15380);
nor U15529 (N_15529,N_15513,N_15403);
nand U15530 (N_15530,N_15485,N_15378);
or U15531 (N_15531,N_15479,N_15490);
nand U15532 (N_15532,N_15473,N_15399);
xnor U15533 (N_15533,N_15420,N_15453);
and U15534 (N_15534,N_15460,N_15498);
nor U15535 (N_15535,N_15371,N_15481);
nand U15536 (N_15536,N_15494,N_15471);
nor U15537 (N_15537,N_15396,N_15434);
and U15538 (N_15538,N_15383,N_15372);
and U15539 (N_15539,N_15386,N_15376);
xnor U15540 (N_15540,N_15418,N_15433);
xor U15541 (N_15541,N_15487,N_15368);
nor U15542 (N_15542,N_15363,N_15437);
nand U15543 (N_15543,N_15455,N_15413);
xnor U15544 (N_15544,N_15493,N_15509);
xnor U15545 (N_15545,N_15404,N_15365);
nand U15546 (N_15546,N_15429,N_15377);
or U15547 (N_15547,N_15384,N_15388);
nor U15548 (N_15548,N_15482,N_15489);
nand U15549 (N_15549,N_15458,N_15477);
xor U15550 (N_15550,N_15491,N_15454);
nor U15551 (N_15551,N_15385,N_15367);
or U15552 (N_15552,N_15512,N_15478);
nand U15553 (N_15553,N_15411,N_15450);
or U15554 (N_15554,N_15506,N_15467);
xnor U15555 (N_15555,N_15510,N_15515);
nand U15556 (N_15556,N_15381,N_15504);
and U15557 (N_15557,N_15448,N_15427);
xnor U15558 (N_15558,N_15415,N_15410);
and U15559 (N_15559,N_15511,N_15503);
xnor U15560 (N_15560,N_15374,N_15519);
nand U15561 (N_15561,N_15430,N_15514);
nand U15562 (N_15562,N_15397,N_15406);
and U15563 (N_15563,N_15438,N_15435);
nor U15564 (N_15564,N_15441,N_15366);
or U15565 (N_15565,N_15462,N_15496);
or U15566 (N_15566,N_15364,N_15446);
nor U15567 (N_15567,N_15472,N_15445);
xnor U15568 (N_15568,N_15407,N_15390);
nor U15569 (N_15569,N_15484,N_15443);
xor U15570 (N_15570,N_15409,N_15497);
and U15571 (N_15571,N_15432,N_15436);
nor U15572 (N_15572,N_15492,N_15505);
nor U15573 (N_15573,N_15459,N_15463);
nand U15574 (N_15574,N_15476,N_15465);
xor U15575 (N_15575,N_15468,N_15419);
nand U15576 (N_15576,N_15393,N_15461);
nor U15577 (N_15577,N_15480,N_15398);
and U15578 (N_15578,N_15387,N_15449);
nand U15579 (N_15579,N_15424,N_15369);
nor U15580 (N_15580,N_15466,N_15444);
xnor U15581 (N_15581,N_15395,N_15373);
nand U15582 (N_15582,N_15421,N_15488);
xnor U15583 (N_15583,N_15428,N_15400);
nand U15584 (N_15584,N_15389,N_15405);
nand U15585 (N_15585,N_15379,N_15426);
nor U15586 (N_15586,N_15495,N_15475);
or U15587 (N_15587,N_15451,N_15464);
and U15588 (N_15588,N_15440,N_15382);
xnor U15589 (N_15589,N_15394,N_15414);
or U15590 (N_15590,N_15474,N_15508);
xor U15591 (N_15591,N_15417,N_15412);
nor U15592 (N_15592,N_15452,N_15431);
and U15593 (N_15593,N_15457,N_15507);
and U15594 (N_15594,N_15370,N_15362);
or U15595 (N_15595,N_15442,N_15500);
and U15596 (N_15596,N_15416,N_15391);
or U15597 (N_15597,N_15361,N_15518);
nand U15598 (N_15598,N_15483,N_15402);
nor U15599 (N_15599,N_15401,N_15502);
nand U15600 (N_15600,N_15398,N_15466);
nor U15601 (N_15601,N_15485,N_15495);
nor U15602 (N_15602,N_15392,N_15368);
nor U15603 (N_15603,N_15490,N_15488);
nor U15604 (N_15604,N_15464,N_15418);
nor U15605 (N_15605,N_15474,N_15463);
xnor U15606 (N_15606,N_15361,N_15504);
nand U15607 (N_15607,N_15496,N_15452);
nand U15608 (N_15608,N_15461,N_15423);
or U15609 (N_15609,N_15388,N_15370);
nor U15610 (N_15610,N_15448,N_15414);
nor U15611 (N_15611,N_15422,N_15405);
and U15612 (N_15612,N_15476,N_15496);
or U15613 (N_15613,N_15435,N_15361);
nand U15614 (N_15614,N_15492,N_15498);
and U15615 (N_15615,N_15371,N_15478);
xor U15616 (N_15616,N_15428,N_15435);
nand U15617 (N_15617,N_15457,N_15512);
or U15618 (N_15618,N_15373,N_15409);
xnor U15619 (N_15619,N_15424,N_15435);
or U15620 (N_15620,N_15419,N_15382);
and U15621 (N_15621,N_15399,N_15516);
or U15622 (N_15622,N_15443,N_15449);
or U15623 (N_15623,N_15512,N_15410);
and U15624 (N_15624,N_15391,N_15515);
nand U15625 (N_15625,N_15377,N_15439);
nand U15626 (N_15626,N_15505,N_15451);
xnor U15627 (N_15627,N_15391,N_15378);
and U15628 (N_15628,N_15500,N_15437);
and U15629 (N_15629,N_15384,N_15440);
nand U15630 (N_15630,N_15364,N_15480);
xor U15631 (N_15631,N_15393,N_15443);
or U15632 (N_15632,N_15492,N_15501);
nand U15633 (N_15633,N_15366,N_15360);
nor U15634 (N_15634,N_15463,N_15384);
xor U15635 (N_15635,N_15439,N_15489);
xor U15636 (N_15636,N_15487,N_15403);
nand U15637 (N_15637,N_15440,N_15371);
and U15638 (N_15638,N_15491,N_15362);
nor U15639 (N_15639,N_15394,N_15436);
nand U15640 (N_15640,N_15498,N_15501);
xnor U15641 (N_15641,N_15513,N_15481);
and U15642 (N_15642,N_15491,N_15397);
nand U15643 (N_15643,N_15478,N_15460);
or U15644 (N_15644,N_15458,N_15486);
and U15645 (N_15645,N_15392,N_15400);
xor U15646 (N_15646,N_15460,N_15383);
nand U15647 (N_15647,N_15388,N_15385);
or U15648 (N_15648,N_15445,N_15442);
xor U15649 (N_15649,N_15413,N_15454);
nor U15650 (N_15650,N_15470,N_15472);
or U15651 (N_15651,N_15468,N_15375);
nor U15652 (N_15652,N_15475,N_15389);
nand U15653 (N_15653,N_15469,N_15484);
or U15654 (N_15654,N_15475,N_15463);
and U15655 (N_15655,N_15378,N_15363);
and U15656 (N_15656,N_15376,N_15469);
or U15657 (N_15657,N_15400,N_15426);
xnor U15658 (N_15658,N_15468,N_15436);
and U15659 (N_15659,N_15487,N_15395);
xnor U15660 (N_15660,N_15512,N_15507);
nand U15661 (N_15661,N_15418,N_15398);
or U15662 (N_15662,N_15517,N_15409);
xnor U15663 (N_15663,N_15376,N_15516);
nand U15664 (N_15664,N_15387,N_15479);
nor U15665 (N_15665,N_15457,N_15419);
and U15666 (N_15666,N_15454,N_15373);
nor U15667 (N_15667,N_15381,N_15388);
nand U15668 (N_15668,N_15368,N_15376);
or U15669 (N_15669,N_15447,N_15420);
nand U15670 (N_15670,N_15452,N_15383);
nor U15671 (N_15671,N_15391,N_15465);
xnor U15672 (N_15672,N_15498,N_15473);
or U15673 (N_15673,N_15467,N_15401);
xnor U15674 (N_15674,N_15449,N_15382);
and U15675 (N_15675,N_15393,N_15399);
nand U15676 (N_15676,N_15369,N_15400);
nor U15677 (N_15677,N_15496,N_15379);
or U15678 (N_15678,N_15438,N_15517);
nand U15679 (N_15679,N_15396,N_15467);
or U15680 (N_15680,N_15647,N_15653);
or U15681 (N_15681,N_15670,N_15537);
and U15682 (N_15682,N_15623,N_15579);
nor U15683 (N_15683,N_15550,N_15568);
nor U15684 (N_15684,N_15671,N_15551);
nor U15685 (N_15685,N_15588,N_15565);
and U15686 (N_15686,N_15669,N_15608);
or U15687 (N_15687,N_15650,N_15627);
or U15688 (N_15688,N_15635,N_15609);
and U15689 (N_15689,N_15555,N_15530);
nand U15690 (N_15690,N_15592,N_15668);
or U15691 (N_15691,N_15590,N_15628);
and U15692 (N_15692,N_15634,N_15545);
xor U15693 (N_15693,N_15667,N_15656);
nor U15694 (N_15694,N_15672,N_15642);
nand U15695 (N_15695,N_15646,N_15576);
xnor U15696 (N_15696,N_15649,N_15524);
and U15697 (N_15697,N_15613,N_15595);
and U15698 (N_15698,N_15677,N_15658);
and U15699 (N_15699,N_15578,N_15601);
and U15700 (N_15700,N_15631,N_15533);
and U15701 (N_15701,N_15525,N_15539);
and U15702 (N_15702,N_15639,N_15603);
nor U15703 (N_15703,N_15641,N_15552);
xnor U15704 (N_15704,N_15665,N_15549);
or U15705 (N_15705,N_15541,N_15597);
and U15706 (N_15706,N_15643,N_15547);
or U15707 (N_15707,N_15558,N_15527);
or U15708 (N_15708,N_15598,N_15632);
xor U15709 (N_15709,N_15559,N_15618);
nor U15710 (N_15710,N_15625,N_15678);
or U15711 (N_15711,N_15544,N_15538);
and U15712 (N_15712,N_15575,N_15536);
xor U15713 (N_15713,N_15633,N_15528);
and U15714 (N_15714,N_15562,N_15619);
nand U15715 (N_15715,N_15583,N_15580);
nor U15716 (N_15716,N_15617,N_15660);
and U15717 (N_15717,N_15651,N_15676);
and U15718 (N_15718,N_15620,N_15548);
or U15719 (N_15719,N_15546,N_15584);
or U15720 (N_15720,N_15679,N_15574);
nand U15721 (N_15721,N_15630,N_15564);
nor U15722 (N_15722,N_15520,N_15523);
nor U15723 (N_15723,N_15593,N_15573);
nor U15724 (N_15724,N_15581,N_15654);
nand U15725 (N_15725,N_15589,N_15621);
or U15726 (N_15726,N_15610,N_15605);
or U15727 (N_15727,N_15553,N_15594);
xnor U15728 (N_15728,N_15535,N_15532);
and U15729 (N_15729,N_15529,N_15560);
or U15730 (N_15730,N_15612,N_15615);
and U15731 (N_15731,N_15582,N_15540);
and U15732 (N_15732,N_15543,N_15640);
and U15733 (N_15733,N_15648,N_15569);
xnor U15734 (N_15734,N_15542,N_15596);
or U15735 (N_15735,N_15534,N_15563);
nand U15736 (N_15736,N_15659,N_15591);
and U15737 (N_15737,N_15662,N_15616);
xor U15738 (N_15738,N_15664,N_15561);
or U15739 (N_15739,N_15566,N_15636);
nand U15740 (N_15740,N_15526,N_15663);
and U15741 (N_15741,N_15614,N_15661);
and U15742 (N_15742,N_15522,N_15666);
and U15743 (N_15743,N_15556,N_15607);
nor U15744 (N_15744,N_15602,N_15570);
and U15745 (N_15745,N_15673,N_15638);
nor U15746 (N_15746,N_15587,N_15572);
nand U15747 (N_15747,N_15622,N_15624);
or U15748 (N_15748,N_15585,N_15611);
and U15749 (N_15749,N_15637,N_15674);
and U15750 (N_15750,N_15557,N_15577);
and U15751 (N_15751,N_15645,N_15531);
or U15752 (N_15752,N_15600,N_15521);
and U15753 (N_15753,N_15606,N_15567);
nand U15754 (N_15754,N_15644,N_15586);
nor U15755 (N_15755,N_15629,N_15604);
or U15756 (N_15756,N_15599,N_15571);
and U15757 (N_15757,N_15657,N_15626);
nor U15758 (N_15758,N_15554,N_15652);
and U15759 (N_15759,N_15675,N_15655);
nand U15760 (N_15760,N_15662,N_15672);
nor U15761 (N_15761,N_15586,N_15604);
nand U15762 (N_15762,N_15651,N_15623);
or U15763 (N_15763,N_15669,N_15626);
nor U15764 (N_15764,N_15549,N_15590);
nand U15765 (N_15765,N_15620,N_15656);
xor U15766 (N_15766,N_15657,N_15612);
or U15767 (N_15767,N_15605,N_15669);
xnor U15768 (N_15768,N_15668,N_15539);
nand U15769 (N_15769,N_15600,N_15524);
xor U15770 (N_15770,N_15551,N_15657);
nor U15771 (N_15771,N_15599,N_15678);
xor U15772 (N_15772,N_15610,N_15649);
xnor U15773 (N_15773,N_15568,N_15633);
and U15774 (N_15774,N_15623,N_15570);
nor U15775 (N_15775,N_15574,N_15642);
and U15776 (N_15776,N_15646,N_15618);
nor U15777 (N_15777,N_15620,N_15556);
or U15778 (N_15778,N_15579,N_15588);
nor U15779 (N_15779,N_15533,N_15587);
xnor U15780 (N_15780,N_15589,N_15655);
nand U15781 (N_15781,N_15628,N_15579);
xnor U15782 (N_15782,N_15586,N_15527);
nor U15783 (N_15783,N_15628,N_15653);
nor U15784 (N_15784,N_15590,N_15653);
nor U15785 (N_15785,N_15620,N_15582);
xor U15786 (N_15786,N_15588,N_15647);
or U15787 (N_15787,N_15603,N_15597);
or U15788 (N_15788,N_15624,N_15653);
xnor U15789 (N_15789,N_15671,N_15587);
xnor U15790 (N_15790,N_15550,N_15620);
nor U15791 (N_15791,N_15624,N_15677);
nor U15792 (N_15792,N_15618,N_15650);
nor U15793 (N_15793,N_15664,N_15553);
nor U15794 (N_15794,N_15600,N_15566);
and U15795 (N_15795,N_15591,N_15638);
nand U15796 (N_15796,N_15627,N_15575);
nor U15797 (N_15797,N_15638,N_15575);
xnor U15798 (N_15798,N_15608,N_15644);
nand U15799 (N_15799,N_15542,N_15646);
nor U15800 (N_15800,N_15535,N_15602);
xnor U15801 (N_15801,N_15567,N_15621);
nand U15802 (N_15802,N_15609,N_15663);
xor U15803 (N_15803,N_15538,N_15672);
nor U15804 (N_15804,N_15631,N_15561);
nand U15805 (N_15805,N_15625,N_15575);
nor U15806 (N_15806,N_15610,N_15647);
or U15807 (N_15807,N_15671,N_15673);
nor U15808 (N_15808,N_15527,N_15638);
and U15809 (N_15809,N_15613,N_15561);
xor U15810 (N_15810,N_15619,N_15603);
nand U15811 (N_15811,N_15669,N_15544);
nand U15812 (N_15812,N_15533,N_15676);
nor U15813 (N_15813,N_15594,N_15624);
nand U15814 (N_15814,N_15674,N_15678);
nand U15815 (N_15815,N_15638,N_15534);
xnor U15816 (N_15816,N_15563,N_15531);
nand U15817 (N_15817,N_15543,N_15678);
nand U15818 (N_15818,N_15544,N_15650);
nor U15819 (N_15819,N_15595,N_15612);
or U15820 (N_15820,N_15616,N_15636);
xnor U15821 (N_15821,N_15601,N_15639);
xnor U15822 (N_15822,N_15652,N_15618);
nor U15823 (N_15823,N_15575,N_15607);
nand U15824 (N_15824,N_15535,N_15537);
and U15825 (N_15825,N_15576,N_15562);
nand U15826 (N_15826,N_15587,N_15635);
nor U15827 (N_15827,N_15593,N_15604);
or U15828 (N_15828,N_15676,N_15546);
or U15829 (N_15829,N_15595,N_15590);
and U15830 (N_15830,N_15528,N_15606);
nor U15831 (N_15831,N_15636,N_15656);
nor U15832 (N_15832,N_15603,N_15636);
and U15833 (N_15833,N_15531,N_15607);
nand U15834 (N_15834,N_15537,N_15528);
xor U15835 (N_15835,N_15591,N_15597);
xor U15836 (N_15836,N_15634,N_15599);
nor U15837 (N_15837,N_15673,N_15602);
or U15838 (N_15838,N_15568,N_15527);
xnor U15839 (N_15839,N_15609,N_15600);
xor U15840 (N_15840,N_15680,N_15714);
nand U15841 (N_15841,N_15784,N_15740);
xor U15842 (N_15842,N_15819,N_15753);
nand U15843 (N_15843,N_15718,N_15737);
xnor U15844 (N_15844,N_15754,N_15704);
nand U15845 (N_15845,N_15774,N_15726);
or U15846 (N_15846,N_15722,N_15729);
and U15847 (N_15847,N_15821,N_15822);
nand U15848 (N_15848,N_15776,N_15743);
and U15849 (N_15849,N_15684,N_15758);
and U15850 (N_15850,N_15744,N_15763);
or U15851 (N_15851,N_15793,N_15810);
xor U15852 (N_15852,N_15792,N_15688);
nand U15853 (N_15853,N_15800,N_15804);
or U15854 (N_15854,N_15707,N_15789);
or U15855 (N_15855,N_15765,N_15723);
or U15856 (N_15856,N_15709,N_15690);
or U15857 (N_15857,N_15833,N_15694);
nor U15858 (N_15858,N_15731,N_15782);
xnor U15859 (N_15859,N_15686,N_15733);
xor U15860 (N_15860,N_15735,N_15755);
xor U15861 (N_15861,N_15805,N_15682);
and U15862 (N_15862,N_15697,N_15770);
and U15863 (N_15863,N_15826,N_15780);
xor U15864 (N_15864,N_15681,N_15706);
xnor U15865 (N_15865,N_15728,N_15752);
nor U15866 (N_15866,N_15708,N_15785);
and U15867 (N_15867,N_15716,N_15698);
nor U15868 (N_15868,N_15803,N_15831);
or U15869 (N_15869,N_15795,N_15699);
or U15870 (N_15870,N_15683,N_15832);
and U15871 (N_15871,N_15787,N_15788);
xnor U15872 (N_15872,N_15835,N_15693);
or U15873 (N_15873,N_15809,N_15823);
xor U15874 (N_15874,N_15739,N_15692);
nand U15875 (N_15875,N_15830,N_15724);
xor U15876 (N_15876,N_15719,N_15838);
or U15877 (N_15877,N_15815,N_15705);
nor U15878 (N_15878,N_15814,N_15839);
xnor U15879 (N_15879,N_15797,N_15757);
xnor U15880 (N_15880,N_15691,N_15772);
or U15881 (N_15881,N_15813,N_15818);
xor U15882 (N_15882,N_15759,N_15713);
xnor U15883 (N_15883,N_15746,N_15736);
xnor U15884 (N_15884,N_15715,N_15790);
and U15885 (N_15885,N_15764,N_15796);
nor U15886 (N_15886,N_15687,N_15837);
and U15887 (N_15887,N_15689,N_15773);
nand U15888 (N_15888,N_15730,N_15750);
nand U15889 (N_15889,N_15742,N_15771);
and U15890 (N_15890,N_15766,N_15747);
nand U15891 (N_15891,N_15762,N_15768);
or U15892 (N_15892,N_15783,N_15756);
and U15893 (N_15893,N_15828,N_15761);
nand U15894 (N_15894,N_15751,N_15760);
and U15895 (N_15895,N_15791,N_15827);
and U15896 (N_15896,N_15801,N_15700);
xnor U15897 (N_15897,N_15727,N_15717);
nor U15898 (N_15898,N_15685,N_15775);
or U15899 (N_15899,N_15806,N_15695);
nand U15900 (N_15900,N_15703,N_15808);
nand U15901 (N_15901,N_15829,N_15817);
nand U15902 (N_15902,N_15799,N_15834);
xor U15903 (N_15903,N_15712,N_15767);
nor U15904 (N_15904,N_15824,N_15778);
nor U15905 (N_15905,N_15721,N_15781);
and U15906 (N_15906,N_15696,N_15802);
nor U15907 (N_15907,N_15836,N_15725);
xor U15908 (N_15908,N_15816,N_15798);
or U15909 (N_15909,N_15749,N_15820);
or U15910 (N_15910,N_15812,N_15720);
nand U15911 (N_15911,N_15701,N_15734);
or U15912 (N_15912,N_15710,N_15769);
or U15913 (N_15913,N_15741,N_15745);
nand U15914 (N_15914,N_15748,N_15811);
nor U15915 (N_15915,N_15794,N_15807);
and U15916 (N_15916,N_15732,N_15702);
xnor U15917 (N_15917,N_15738,N_15779);
or U15918 (N_15918,N_15777,N_15825);
xor U15919 (N_15919,N_15711,N_15786);
xnor U15920 (N_15920,N_15724,N_15772);
or U15921 (N_15921,N_15684,N_15805);
nand U15922 (N_15922,N_15717,N_15797);
xor U15923 (N_15923,N_15772,N_15725);
nor U15924 (N_15924,N_15762,N_15733);
nand U15925 (N_15925,N_15804,N_15832);
xor U15926 (N_15926,N_15739,N_15722);
or U15927 (N_15927,N_15807,N_15816);
nor U15928 (N_15928,N_15779,N_15823);
nor U15929 (N_15929,N_15781,N_15821);
xnor U15930 (N_15930,N_15742,N_15830);
nand U15931 (N_15931,N_15810,N_15704);
nand U15932 (N_15932,N_15704,N_15696);
nor U15933 (N_15933,N_15773,N_15683);
nor U15934 (N_15934,N_15696,N_15712);
nor U15935 (N_15935,N_15753,N_15791);
or U15936 (N_15936,N_15778,N_15787);
nand U15937 (N_15937,N_15803,N_15728);
or U15938 (N_15938,N_15702,N_15696);
nand U15939 (N_15939,N_15720,N_15777);
and U15940 (N_15940,N_15801,N_15751);
or U15941 (N_15941,N_15713,N_15710);
or U15942 (N_15942,N_15752,N_15739);
xnor U15943 (N_15943,N_15696,N_15778);
xor U15944 (N_15944,N_15779,N_15698);
nor U15945 (N_15945,N_15812,N_15838);
or U15946 (N_15946,N_15758,N_15761);
and U15947 (N_15947,N_15818,N_15765);
and U15948 (N_15948,N_15796,N_15808);
or U15949 (N_15949,N_15703,N_15771);
or U15950 (N_15950,N_15805,N_15782);
nor U15951 (N_15951,N_15733,N_15716);
nor U15952 (N_15952,N_15687,N_15806);
xnor U15953 (N_15953,N_15826,N_15702);
and U15954 (N_15954,N_15724,N_15797);
or U15955 (N_15955,N_15824,N_15783);
nand U15956 (N_15956,N_15808,N_15780);
nand U15957 (N_15957,N_15704,N_15735);
nor U15958 (N_15958,N_15682,N_15698);
xnor U15959 (N_15959,N_15743,N_15692);
and U15960 (N_15960,N_15808,N_15719);
and U15961 (N_15961,N_15801,N_15809);
nand U15962 (N_15962,N_15742,N_15699);
or U15963 (N_15963,N_15695,N_15797);
and U15964 (N_15964,N_15777,N_15753);
or U15965 (N_15965,N_15703,N_15690);
xnor U15966 (N_15966,N_15818,N_15809);
or U15967 (N_15967,N_15726,N_15685);
nand U15968 (N_15968,N_15830,N_15744);
and U15969 (N_15969,N_15837,N_15750);
nand U15970 (N_15970,N_15836,N_15812);
or U15971 (N_15971,N_15755,N_15765);
or U15972 (N_15972,N_15745,N_15780);
xor U15973 (N_15973,N_15800,N_15821);
xor U15974 (N_15974,N_15826,N_15714);
or U15975 (N_15975,N_15740,N_15715);
xor U15976 (N_15976,N_15764,N_15833);
or U15977 (N_15977,N_15793,N_15689);
nand U15978 (N_15978,N_15799,N_15777);
or U15979 (N_15979,N_15709,N_15698);
or U15980 (N_15980,N_15731,N_15828);
nor U15981 (N_15981,N_15835,N_15724);
xor U15982 (N_15982,N_15735,N_15727);
and U15983 (N_15983,N_15816,N_15826);
or U15984 (N_15984,N_15800,N_15809);
nand U15985 (N_15985,N_15821,N_15794);
nor U15986 (N_15986,N_15824,N_15757);
xnor U15987 (N_15987,N_15708,N_15813);
nor U15988 (N_15988,N_15742,N_15686);
nor U15989 (N_15989,N_15680,N_15802);
and U15990 (N_15990,N_15717,N_15770);
nand U15991 (N_15991,N_15750,N_15726);
or U15992 (N_15992,N_15788,N_15756);
nor U15993 (N_15993,N_15795,N_15717);
or U15994 (N_15994,N_15713,N_15764);
nor U15995 (N_15995,N_15697,N_15681);
nand U15996 (N_15996,N_15696,N_15835);
or U15997 (N_15997,N_15709,N_15754);
and U15998 (N_15998,N_15771,N_15839);
and U15999 (N_15999,N_15760,N_15741);
or U16000 (N_16000,N_15911,N_15970);
nand U16001 (N_16001,N_15876,N_15968);
nand U16002 (N_16002,N_15844,N_15973);
or U16003 (N_16003,N_15870,N_15916);
nor U16004 (N_16004,N_15993,N_15977);
xnor U16005 (N_16005,N_15902,N_15941);
xnor U16006 (N_16006,N_15983,N_15913);
xor U16007 (N_16007,N_15855,N_15953);
xnor U16008 (N_16008,N_15900,N_15928);
or U16009 (N_16009,N_15960,N_15965);
or U16010 (N_16010,N_15975,N_15853);
or U16011 (N_16011,N_15852,N_15978);
or U16012 (N_16012,N_15950,N_15894);
xnor U16013 (N_16013,N_15860,N_15964);
xor U16014 (N_16014,N_15985,N_15895);
or U16015 (N_16015,N_15847,N_15871);
or U16016 (N_16016,N_15869,N_15962);
nor U16017 (N_16017,N_15969,N_15859);
nand U16018 (N_16018,N_15972,N_15868);
or U16019 (N_16019,N_15920,N_15882);
nand U16020 (N_16020,N_15863,N_15927);
or U16021 (N_16021,N_15939,N_15990);
nand U16022 (N_16022,N_15872,N_15888);
nor U16023 (N_16023,N_15959,N_15932);
nand U16024 (N_16024,N_15843,N_15942);
nor U16025 (N_16025,N_15848,N_15922);
and U16026 (N_16026,N_15849,N_15933);
nand U16027 (N_16027,N_15884,N_15886);
and U16028 (N_16028,N_15906,N_15845);
or U16029 (N_16029,N_15867,N_15981);
xor U16030 (N_16030,N_15999,N_15861);
or U16031 (N_16031,N_15952,N_15944);
xnor U16032 (N_16032,N_15992,N_15877);
xnor U16033 (N_16033,N_15976,N_15926);
and U16034 (N_16034,N_15866,N_15919);
and U16035 (N_16035,N_15908,N_15974);
or U16036 (N_16036,N_15946,N_15857);
nor U16037 (N_16037,N_15892,N_15929);
and U16038 (N_16038,N_15930,N_15874);
xnor U16039 (N_16039,N_15923,N_15945);
nand U16040 (N_16040,N_15955,N_15910);
and U16041 (N_16041,N_15889,N_15984);
xor U16042 (N_16042,N_15914,N_15988);
xor U16043 (N_16043,N_15865,N_15846);
or U16044 (N_16044,N_15898,N_15947);
nand U16045 (N_16045,N_15873,N_15891);
or U16046 (N_16046,N_15948,N_15904);
or U16047 (N_16047,N_15934,N_15841);
xnor U16048 (N_16048,N_15951,N_15921);
xor U16049 (N_16049,N_15980,N_15971);
xnor U16050 (N_16050,N_15901,N_15840);
nor U16051 (N_16051,N_15851,N_15903);
or U16052 (N_16052,N_15887,N_15905);
nor U16053 (N_16053,N_15850,N_15938);
xnor U16054 (N_16054,N_15979,N_15967);
and U16055 (N_16055,N_15896,N_15996);
and U16056 (N_16056,N_15924,N_15864);
nand U16057 (N_16057,N_15912,N_15879);
xor U16058 (N_16058,N_15925,N_15995);
or U16059 (N_16059,N_15935,N_15994);
or U16060 (N_16060,N_15883,N_15949);
or U16061 (N_16061,N_15880,N_15907);
nand U16062 (N_16062,N_15957,N_15897);
or U16063 (N_16063,N_15966,N_15991);
nor U16064 (N_16064,N_15854,N_15899);
nand U16065 (N_16065,N_15856,N_15881);
nor U16066 (N_16066,N_15842,N_15986);
or U16067 (N_16067,N_15998,N_15936);
and U16068 (N_16068,N_15875,N_15890);
and U16069 (N_16069,N_15982,N_15940);
nand U16070 (N_16070,N_15943,N_15997);
nor U16071 (N_16071,N_15989,N_15954);
and U16072 (N_16072,N_15885,N_15937);
nor U16073 (N_16073,N_15893,N_15878);
xor U16074 (N_16074,N_15956,N_15987);
or U16075 (N_16075,N_15963,N_15909);
nor U16076 (N_16076,N_15862,N_15931);
and U16077 (N_16077,N_15961,N_15958);
or U16078 (N_16078,N_15915,N_15858);
nand U16079 (N_16079,N_15918,N_15917);
or U16080 (N_16080,N_15861,N_15978);
or U16081 (N_16081,N_15986,N_15918);
nor U16082 (N_16082,N_15892,N_15969);
and U16083 (N_16083,N_15973,N_15995);
and U16084 (N_16084,N_15868,N_15899);
and U16085 (N_16085,N_15975,N_15852);
or U16086 (N_16086,N_15858,N_15904);
or U16087 (N_16087,N_15997,N_15978);
nor U16088 (N_16088,N_15994,N_15892);
nand U16089 (N_16089,N_15951,N_15909);
nor U16090 (N_16090,N_15867,N_15877);
nand U16091 (N_16091,N_15859,N_15856);
and U16092 (N_16092,N_15975,N_15929);
or U16093 (N_16093,N_15976,N_15998);
and U16094 (N_16094,N_15994,N_15898);
nand U16095 (N_16095,N_15865,N_15860);
or U16096 (N_16096,N_15865,N_15899);
nand U16097 (N_16097,N_15887,N_15875);
xor U16098 (N_16098,N_15966,N_15927);
nand U16099 (N_16099,N_15914,N_15885);
nor U16100 (N_16100,N_15958,N_15926);
or U16101 (N_16101,N_15843,N_15902);
xor U16102 (N_16102,N_15965,N_15877);
nor U16103 (N_16103,N_15913,N_15995);
nand U16104 (N_16104,N_15842,N_15965);
nor U16105 (N_16105,N_15944,N_15987);
nand U16106 (N_16106,N_15922,N_15876);
and U16107 (N_16107,N_15880,N_15926);
or U16108 (N_16108,N_15975,N_15994);
or U16109 (N_16109,N_15906,N_15879);
and U16110 (N_16110,N_15899,N_15945);
nand U16111 (N_16111,N_15934,N_15848);
xor U16112 (N_16112,N_15924,N_15929);
nor U16113 (N_16113,N_15898,N_15972);
or U16114 (N_16114,N_15862,N_15935);
xnor U16115 (N_16115,N_15874,N_15974);
nand U16116 (N_16116,N_15909,N_15911);
nor U16117 (N_16117,N_15907,N_15955);
xnor U16118 (N_16118,N_15847,N_15972);
or U16119 (N_16119,N_15985,N_15846);
nand U16120 (N_16120,N_15962,N_15943);
or U16121 (N_16121,N_15896,N_15902);
nor U16122 (N_16122,N_15953,N_15908);
xnor U16123 (N_16123,N_15866,N_15992);
xnor U16124 (N_16124,N_15843,N_15973);
and U16125 (N_16125,N_15873,N_15945);
or U16126 (N_16126,N_15976,N_15906);
or U16127 (N_16127,N_15849,N_15907);
and U16128 (N_16128,N_15879,N_15859);
or U16129 (N_16129,N_15976,N_15866);
nand U16130 (N_16130,N_15890,N_15948);
and U16131 (N_16131,N_15846,N_15916);
nor U16132 (N_16132,N_15846,N_15844);
and U16133 (N_16133,N_15982,N_15953);
nand U16134 (N_16134,N_15857,N_15999);
or U16135 (N_16135,N_15922,N_15910);
and U16136 (N_16136,N_15864,N_15907);
xnor U16137 (N_16137,N_15915,N_15905);
and U16138 (N_16138,N_15946,N_15968);
xnor U16139 (N_16139,N_15990,N_15843);
nand U16140 (N_16140,N_15933,N_15894);
xnor U16141 (N_16141,N_15841,N_15987);
or U16142 (N_16142,N_15946,N_15911);
or U16143 (N_16143,N_15844,N_15908);
nand U16144 (N_16144,N_15894,N_15884);
or U16145 (N_16145,N_15992,N_15959);
nand U16146 (N_16146,N_15933,N_15893);
or U16147 (N_16147,N_15973,N_15880);
xnor U16148 (N_16148,N_15948,N_15963);
or U16149 (N_16149,N_15901,N_15911);
nor U16150 (N_16150,N_15896,N_15994);
nor U16151 (N_16151,N_15865,N_15916);
or U16152 (N_16152,N_15953,N_15865);
or U16153 (N_16153,N_15922,N_15885);
or U16154 (N_16154,N_15985,N_15997);
and U16155 (N_16155,N_15869,N_15860);
nor U16156 (N_16156,N_15938,N_15934);
nand U16157 (N_16157,N_15989,N_15967);
nor U16158 (N_16158,N_15941,N_15992);
and U16159 (N_16159,N_15910,N_15963);
or U16160 (N_16160,N_16130,N_16115);
and U16161 (N_16161,N_16109,N_16000);
nand U16162 (N_16162,N_16137,N_16028);
xnor U16163 (N_16163,N_16027,N_16108);
xor U16164 (N_16164,N_16141,N_16129);
or U16165 (N_16165,N_16003,N_16045);
nor U16166 (N_16166,N_16062,N_16106);
nor U16167 (N_16167,N_16042,N_16075);
and U16168 (N_16168,N_16071,N_16127);
and U16169 (N_16169,N_16128,N_16155);
xor U16170 (N_16170,N_16002,N_16123);
xor U16171 (N_16171,N_16012,N_16124);
nand U16172 (N_16172,N_16135,N_16030);
and U16173 (N_16173,N_16011,N_16097);
nand U16174 (N_16174,N_16121,N_16138);
xnor U16175 (N_16175,N_16026,N_16089);
nand U16176 (N_16176,N_16020,N_16100);
nor U16177 (N_16177,N_16080,N_16052);
nor U16178 (N_16178,N_16139,N_16152);
xnor U16179 (N_16179,N_16081,N_16043);
nor U16180 (N_16180,N_16046,N_16051);
and U16181 (N_16181,N_16018,N_16093);
nand U16182 (N_16182,N_16107,N_16008);
and U16183 (N_16183,N_16092,N_16038);
xor U16184 (N_16184,N_16060,N_16058);
or U16185 (N_16185,N_16063,N_16035);
or U16186 (N_16186,N_16113,N_16001);
xor U16187 (N_16187,N_16024,N_16087);
or U16188 (N_16188,N_16104,N_16007);
nand U16189 (N_16189,N_16053,N_16077);
nand U16190 (N_16190,N_16009,N_16049);
or U16191 (N_16191,N_16034,N_16016);
and U16192 (N_16192,N_16103,N_16022);
nor U16193 (N_16193,N_16091,N_16023);
or U16194 (N_16194,N_16118,N_16116);
nand U16195 (N_16195,N_16096,N_16144);
and U16196 (N_16196,N_16082,N_16067);
and U16197 (N_16197,N_16010,N_16122);
nor U16198 (N_16198,N_16140,N_16094);
xor U16199 (N_16199,N_16095,N_16147);
and U16200 (N_16200,N_16061,N_16076);
nor U16201 (N_16201,N_16054,N_16031);
and U16202 (N_16202,N_16134,N_16132);
nor U16203 (N_16203,N_16072,N_16083);
and U16204 (N_16204,N_16117,N_16150);
nor U16205 (N_16205,N_16146,N_16085);
and U16206 (N_16206,N_16056,N_16125);
nor U16207 (N_16207,N_16069,N_16044);
xor U16208 (N_16208,N_16073,N_16143);
or U16209 (N_16209,N_16057,N_16157);
xnor U16210 (N_16210,N_16017,N_16154);
nor U16211 (N_16211,N_16102,N_16032);
xor U16212 (N_16212,N_16112,N_16047);
xor U16213 (N_16213,N_16004,N_16156);
nand U16214 (N_16214,N_16055,N_16105);
or U16215 (N_16215,N_16066,N_16159);
nand U16216 (N_16216,N_16015,N_16084);
nand U16217 (N_16217,N_16033,N_16021);
nand U16218 (N_16218,N_16114,N_16153);
nand U16219 (N_16219,N_16111,N_16101);
and U16220 (N_16220,N_16151,N_16119);
nor U16221 (N_16221,N_16039,N_16098);
nor U16222 (N_16222,N_16090,N_16088);
nand U16223 (N_16223,N_16037,N_16025);
xor U16224 (N_16224,N_16065,N_16120);
and U16225 (N_16225,N_16041,N_16145);
xnor U16226 (N_16226,N_16131,N_16064);
nand U16227 (N_16227,N_16005,N_16099);
and U16228 (N_16228,N_16149,N_16086);
nand U16229 (N_16229,N_16040,N_16079);
nor U16230 (N_16230,N_16048,N_16136);
nor U16231 (N_16231,N_16078,N_16110);
nand U16232 (N_16232,N_16068,N_16133);
xor U16233 (N_16233,N_16019,N_16036);
and U16234 (N_16234,N_16050,N_16142);
or U16235 (N_16235,N_16148,N_16126);
nor U16236 (N_16236,N_16014,N_16029);
nand U16237 (N_16237,N_16158,N_16006);
nor U16238 (N_16238,N_16013,N_16070);
or U16239 (N_16239,N_16074,N_16059);
and U16240 (N_16240,N_16112,N_16070);
xnor U16241 (N_16241,N_16082,N_16000);
or U16242 (N_16242,N_16080,N_16024);
and U16243 (N_16243,N_16101,N_16097);
nor U16244 (N_16244,N_16151,N_16130);
nor U16245 (N_16245,N_16046,N_16059);
xor U16246 (N_16246,N_16118,N_16096);
xor U16247 (N_16247,N_16090,N_16092);
xor U16248 (N_16248,N_16017,N_16058);
nand U16249 (N_16249,N_16115,N_16034);
nand U16250 (N_16250,N_16038,N_16067);
or U16251 (N_16251,N_16097,N_16014);
and U16252 (N_16252,N_16024,N_16152);
xnor U16253 (N_16253,N_16083,N_16082);
nand U16254 (N_16254,N_16032,N_16135);
nand U16255 (N_16255,N_16147,N_16068);
nand U16256 (N_16256,N_16096,N_16136);
nand U16257 (N_16257,N_16122,N_16025);
xnor U16258 (N_16258,N_16113,N_16143);
or U16259 (N_16259,N_16095,N_16068);
and U16260 (N_16260,N_16033,N_16038);
nor U16261 (N_16261,N_16077,N_16001);
xor U16262 (N_16262,N_16124,N_16020);
or U16263 (N_16263,N_16039,N_16113);
nand U16264 (N_16264,N_16100,N_16051);
nor U16265 (N_16265,N_16079,N_16058);
xnor U16266 (N_16266,N_16021,N_16000);
nand U16267 (N_16267,N_16144,N_16099);
or U16268 (N_16268,N_16113,N_16096);
xnor U16269 (N_16269,N_16038,N_16151);
or U16270 (N_16270,N_16007,N_16064);
nand U16271 (N_16271,N_16059,N_16047);
or U16272 (N_16272,N_16012,N_16106);
or U16273 (N_16273,N_16118,N_16014);
xnor U16274 (N_16274,N_16104,N_16100);
and U16275 (N_16275,N_16105,N_16024);
nand U16276 (N_16276,N_16065,N_16071);
nor U16277 (N_16277,N_16148,N_16013);
nor U16278 (N_16278,N_16063,N_16013);
and U16279 (N_16279,N_16003,N_16080);
nand U16280 (N_16280,N_16100,N_16060);
xnor U16281 (N_16281,N_16083,N_16129);
xor U16282 (N_16282,N_16111,N_16059);
xnor U16283 (N_16283,N_16053,N_16015);
nor U16284 (N_16284,N_16101,N_16026);
and U16285 (N_16285,N_16034,N_16078);
xnor U16286 (N_16286,N_16103,N_16019);
nand U16287 (N_16287,N_16058,N_16032);
nand U16288 (N_16288,N_16078,N_16151);
xor U16289 (N_16289,N_16106,N_16038);
nand U16290 (N_16290,N_16122,N_16058);
or U16291 (N_16291,N_16013,N_16096);
or U16292 (N_16292,N_16092,N_16151);
and U16293 (N_16293,N_16029,N_16099);
and U16294 (N_16294,N_16083,N_16145);
or U16295 (N_16295,N_16140,N_16092);
xor U16296 (N_16296,N_16000,N_16132);
or U16297 (N_16297,N_16099,N_16011);
or U16298 (N_16298,N_16087,N_16005);
nand U16299 (N_16299,N_16130,N_16041);
xor U16300 (N_16300,N_16032,N_16107);
xnor U16301 (N_16301,N_16051,N_16126);
nand U16302 (N_16302,N_16037,N_16155);
xor U16303 (N_16303,N_16128,N_16061);
and U16304 (N_16304,N_16080,N_16040);
nor U16305 (N_16305,N_16151,N_16004);
nor U16306 (N_16306,N_16151,N_16061);
nand U16307 (N_16307,N_16092,N_16102);
or U16308 (N_16308,N_16047,N_16033);
and U16309 (N_16309,N_16144,N_16052);
nand U16310 (N_16310,N_16121,N_16004);
xor U16311 (N_16311,N_16077,N_16091);
nand U16312 (N_16312,N_16053,N_16004);
nand U16313 (N_16313,N_16028,N_16136);
nand U16314 (N_16314,N_16132,N_16039);
or U16315 (N_16315,N_16002,N_16046);
nand U16316 (N_16316,N_16039,N_16057);
nand U16317 (N_16317,N_16118,N_16090);
nand U16318 (N_16318,N_16015,N_16058);
xor U16319 (N_16319,N_16128,N_16000);
nor U16320 (N_16320,N_16199,N_16200);
xnor U16321 (N_16321,N_16259,N_16202);
nor U16322 (N_16322,N_16168,N_16162);
and U16323 (N_16323,N_16184,N_16305);
xnor U16324 (N_16324,N_16232,N_16255);
nor U16325 (N_16325,N_16211,N_16175);
and U16326 (N_16326,N_16312,N_16256);
nand U16327 (N_16327,N_16169,N_16237);
nor U16328 (N_16328,N_16313,N_16223);
xor U16329 (N_16329,N_16174,N_16236);
or U16330 (N_16330,N_16285,N_16178);
or U16331 (N_16331,N_16274,N_16183);
nor U16332 (N_16332,N_16300,N_16282);
xnor U16333 (N_16333,N_16231,N_16176);
xnor U16334 (N_16334,N_16230,N_16311);
or U16335 (N_16335,N_16227,N_16217);
or U16336 (N_16336,N_16319,N_16238);
or U16337 (N_16337,N_16318,N_16278);
nand U16338 (N_16338,N_16161,N_16197);
nor U16339 (N_16339,N_16204,N_16276);
nand U16340 (N_16340,N_16171,N_16273);
or U16341 (N_16341,N_16265,N_16242);
nor U16342 (N_16342,N_16304,N_16293);
nor U16343 (N_16343,N_16166,N_16193);
xnor U16344 (N_16344,N_16264,N_16291);
or U16345 (N_16345,N_16247,N_16233);
nand U16346 (N_16346,N_16210,N_16206);
or U16347 (N_16347,N_16270,N_16296);
nand U16348 (N_16348,N_16287,N_16167);
xor U16349 (N_16349,N_16295,N_16198);
and U16350 (N_16350,N_16267,N_16194);
xnor U16351 (N_16351,N_16219,N_16288);
nor U16352 (N_16352,N_16249,N_16252);
or U16353 (N_16353,N_16209,N_16299);
nand U16354 (N_16354,N_16315,N_16173);
nand U16355 (N_16355,N_16261,N_16165);
and U16356 (N_16356,N_16213,N_16281);
or U16357 (N_16357,N_16228,N_16316);
nand U16358 (N_16358,N_16308,N_16235);
nor U16359 (N_16359,N_16286,N_16272);
nand U16360 (N_16360,N_16181,N_16292);
nand U16361 (N_16361,N_16203,N_16170);
nand U16362 (N_16362,N_16241,N_16279);
xnor U16363 (N_16363,N_16257,N_16254);
and U16364 (N_16364,N_16244,N_16275);
xnor U16365 (N_16365,N_16240,N_16283);
xnor U16366 (N_16366,N_16212,N_16268);
nand U16367 (N_16367,N_16163,N_16207);
or U16368 (N_16368,N_16185,N_16306);
and U16369 (N_16369,N_16195,N_16191);
xor U16370 (N_16370,N_16208,N_16298);
nor U16371 (N_16371,N_16239,N_16269);
nor U16372 (N_16372,N_16243,N_16224);
xor U16373 (N_16373,N_16205,N_16303);
and U16374 (N_16374,N_16192,N_16218);
nand U16375 (N_16375,N_16301,N_16215);
nand U16376 (N_16376,N_16297,N_16221);
and U16377 (N_16377,N_16309,N_16289);
xnor U16378 (N_16378,N_16177,N_16307);
and U16379 (N_16379,N_16234,N_16190);
nand U16380 (N_16380,N_16196,N_16310);
xnor U16381 (N_16381,N_16260,N_16188);
nand U16382 (N_16382,N_16189,N_16245);
and U16383 (N_16383,N_16271,N_16263);
or U16384 (N_16384,N_16284,N_16248);
or U16385 (N_16385,N_16186,N_16180);
nand U16386 (N_16386,N_16160,N_16182);
nor U16387 (N_16387,N_16246,N_16251);
nor U16388 (N_16388,N_16314,N_16294);
nand U16389 (N_16389,N_16172,N_16214);
xor U16390 (N_16390,N_16253,N_16225);
or U16391 (N_16391,N_16229,N_16164);
nand U16392 (N_16392,N_16290,N_16280);
and U16393 (N_16393,N_16222,N_16277);
nand U16394 (N_16394,N_16226,N_16220);
xor U16395 (N_16395,N_16258,N_16179);
or U16396 (N_16396,N_16266,N_16201);
xor U16397 (N_16397,N_16262,N_16317);
nor U16398 (N_16398,N_16250,N_16216);
and U16399 (N_16399,N_16302,N_16187);
nor U16400 (N_16400,N_16227,N_16182);
nor U16401 (N_16401,N_16263,N_16202);
xor U16402 (N_16402,N_16180,N_16317);
or U16403 (N_16403,N_16291,N_16184);
or U16404 (N_16404,N_16197,N_16227);
and U16405 (N_16405,N_16266,N_16241);
nor U16406 (N_16406,N_16179,N_16196);
xnor U16407 (N_16407,N_16315,N_16257);
xnor U16408 (N_16408,N_16226,N_16314);
and U16409 (N_16409,N_16277,N_16244);
and U16410 (N_16410,N_16288,N_16199);
nand U16411 (N_16411,N_16236,N_16179);
and U16412 (N_16412,N_16222,N_16315);
and U16413 (N_16413,N_16180,N_16189);
and U16414 (N_16414,N_16209,N_16289);
nand U16415 (N_16415,N_16227,N_16255);
nand U16416 (N_16416,N_16216,N_16241);
nor U16417 (N_16417,N_16203,N_16269);
or U16418 (N_16418,N_16265,N_16246);
xnor U16419 (N_16419,N_16280,N_16167);
nor U16420 (N_16420,N_16256,N_16253);
or U16421 (N_16421,N_16231,N_16161);
and U16422 (N_16422,N_16193,N_16312);
nand U16423 (N_16423,N_16162,N_16294);
nand U16424 (N_16424,N_16269,N_16229);
nand U16425 (N_16425,N_16280,N_16303);
or U16426 (N_16426,N_16221,N_16286);
nand U16427 (N_16427,N_16283,N_16214);
nor U16428 (N_16428,N_16304,N_16240);
nand U16429 (N_16429,N_16180,N_16179);
nor U16430 (N_16430,N_16208,N_16300);
or U16431 (N_16431,N_16281,N_16225);
xor U16432 (N_16432,N_16216,N_16227);
xor U16433 (N_16433,N_16279,N_16173);
nor U16434 (N_16434,N_16203,N_16184);
and U16435 (N_16435,N_16310,N_16235);
and U16436 (N_16436,N_16188,N_16242);
or U16437 (N_16437,N_16300,N_16173);
xor U16438 (N_16438,N_16211,N_16162);
nand U16439 (N_16439,N_16168,N_16284);
or U16440 (N_16440,N_16312,N_16262);
xor U16441 (N_16441,N_16230,N_16253);
xnor U16442 (N_16442,N_16238,N_16247);
nand U16443 (N_16443,N_16196,N_16216);
and U16444 (N_16444,N_16319,N_16165);
and U16445 (N_16445,N_16182,N_16301);
or U16446 (N_16446,N_16300,N_16248);
or U16447 (N_16447,N_16277,N_16295);
nand U16448 (N_16448,N_16193,N_16235);
or U16449 (N_16449,N_16182,N_16310);
nand U16450 (N_16450,N_16187,N_16308);
or U16451 (N_16451,N_16276,N_16265);
xor U16452 (N_16452,N_16275,N_16216);
nand U16453 (N_16453,N_16240,N_16292);
nand U16454 (N_16454,N_16291,N_16169);
and U16455 (N_16455,N_16260,N_16293);
nor U16456 (N_16456,N_16267,N_16179);
nand U16457 (N_16457,N_16241,N_16298);
xor U16458 (N_16458,N_16238,N_16268);
or U16459 (N_16459,N_16244,N_16310);
nor U16460 (N_16460,N_16179,N_16189);
or U16461 (N_16461,N_16248,N_16260);
xor U16462 (N_16462,N_16273,N_16163);
and U16463 (N_16463,N_16316,N_16200);
nand U16464 (N_16464,N_16183,N_16206);
nand U16465 (N_16465,N_16256,N_16187);
nand U16466 (N_16466,N_16161,N_16315);
or U16467 (N_16467,N_16249,N_16309);
and U16468 (N_16468,N_16310,N_16281);
xnor U16469 (N_16469,N_16178,N_16199);
and U16470 (N_16470,N_16311,N_16246);
and U16471 (N_16471,N_16174,N_16214);
xor U16472 (N_16472,N_16287,N_16251);
nand U16473 (N_16473,N_16204,N_16313);
or U16474 (N_16474,N_16167,N_16209);
xnor U16475 (N_16475,N_16202,N_16225);
or U16476 (N_16476,N_16260,N_16291);
xnor U16477 (N_16477,N_16300,N_16262);
or U16478 (N_16478,N_16318,N_16247);
nand U16479 (N_16479,N_16227,N_16177);
nor U16480 (N_16480,N_16393,N_16342);
nor U16481 (N_16481,N_16375,N_16357);
xnor U16482 (N_16482,N_16413,N_16432);
xnor U16483 (N_16483,N_16441,N_16479);
xnor U16484 (N_16484,N_16386,N_16349);
and U16485 (N_16485,N_16424,N_16425);
nor U16486 (N_16486,N_16325,N_16336);
and U16487 (N_16487,N_16411,N_16348);
nor U16488 (N_16488,N_16380,N_16414);
nor U16489 (N_16489,N_16396,N_16446);
nand U16490 (N_16490,N_16454,N_16382);
nand U16491 (N_16491,N_16407,N_16324);
and U16492 (N_16492,N_16395,N_16459);
xor U16493 (N_16493,N_16404,N_16340);
and U16494 (N_16494,N_16360,N_16335);
nor U16495 (N_16495,N_16328,N_16326);
xnor U16496 (N_16496,N_16439,N_16457);
nor U16497 (N_16497,N_16369,N_16381);
nand U16498 (N_16498,N_16376,N_16426);
or U16499 (N_16499,N_16433,N_16472);
and U16500 (N_16500,N_16379,N_16378);
and U16501 (N_16501,N_16430,N_16387);
and U16502 (N_16502,N_16400,N_16374);
and U16503 (N_16503,N_16391,N_16420);
nand U16504 (N_16504,N_16397,N_16416);
or U16505 (N_16505,N_16428,N_16410);
or U16506 (N_16506,N_16474,N_16398);
nor U16507 (N_16507,N_16465,N_16394);
xor U16508 (N_16508,N_16355,N_16384);
or U16509 (N_16509,N_16419,N_16361);
or U16510 (N_16510,N_16356,N_16385);
xnor U16511 (N_16511,N_16403,N_16339);
xor U16512 (N_16512,N_16467,N_16445);
or U16513 (N_16513,N_16329,N_16346);
nor U16514 (N_16514,N_16405,N_16471);
and U16515 (N_16515,N_16322,N_16427);
or U16516 (N_16516,N_16388,N_16370);
or U16517 (N_16517,N_16418,N_16417);
xor U16518 (N_16518,N_16351,N_16408);
nor U16519 (N_16519,N_16367,N_16451);
and U16520 (N_16520,N_16347,N_16429);
or U16521 (N_16521,N_16452,N_16473);
nand U16522 (N_16522,N_16358,N_16449);
and U16523 (N_16523,N_16475,N_16354);
nand U16524 (N_16524,N_16353,N_16442);
and U16525 (N_16525,N_16331,N_16458);
and U16526 (N_16526,N_16401,N_16437);
xnor U16527 (N_16527,N_16438,N_16434);
or U16528 (N_16528,N_16476,N_16444);
xor U16529 (N_16529,N_16320,N_16462);
xor U16530 (N_16530,N_16455,N_16364);
nor U16531 (N_16531,N_16362,N_16383);
nor U16532 (N_16532,N_16443,N_16321);
nand U16533 (N_16533,N_16423,N_16453);
nand U16534 (N_16534,N_16345,N_16344);
nand U16535 (N_16535,N_16366,N_16341);
xnor U16536 (N_16536,N_16460,N_16371);
nor U16537 (N_16537,N_16338,N_16402);
xor U16538 (N_16538,N_16440,N_16415);
or U16539 (N_16539,N_16435,N_16334);
and U16540 (N_16540,N_16447,N_16470);
nand U16541 (N_16541,N_16332,N_16390);
or U16542 (N_16542,N_16365,N_16327);
nand U16543 (N_16543,N_16466,N_16477);
and U16544 (N_16544,N_16464,N_16409);
xor U16545 (N_16545,N_16421,N_16350);
or U16546 (N_16546,N_16343,N_16461);
or U16547 (N_16547,N_16412,N_16406);
and U16548 (N_16548,N_16389,N_16363);
xnor U16549 (N_16549,N_16478,N_16323);
nor U16550 (N_16550,N_16469,N_16436);
and U16551 (N_16551,N_16368,N_16422);
nor U16552 (N_16552,N_16372,N_16359);
and U16553 (N_16553,N_16468,N_16463);
and U16554 (N_16554,N_16399,N_16377);
xor U16555 (N_16555,N_16450,N_16431);
and U16556 (N_16556,N_16392,N_16333);
and U16557 (N_16557,N_16330,N_16337);
nand U16558 (N_16558,N_16352,N_16373);
and U16559 (N_16559,N_16456,N_16448);
xnor U16560 (N_16560,N_16462,N_16418);
and U16561 (N_16561,N_16474,N_16394);
nor U16562 (N_16562,N_16457,N_16443);
nor U16563 (N_16563,N_16391,N_16462);
xor U16564 (N_16564,N_16444,N_16396);
nand U16565 (N_16565,N_16423,N_16370);
nand U16566 (N_16566,N_16412,N_16363);
nand U16567 (N_16567,N_16413,N_16441);
nor U16568 (N_16568,N_16366,N_16372);
or U16569 (N_16569,N_16345,N_16351);
nor U16570 (N_16570,N_16469,N_16356);
or U16571 (N_16571,N_16376,N_16410);
nand U16572 (N_16572,N_16440,N_16471);
xor U16573 (N_16573,N_16320,N_16331);
xor U16574 (N_16574,N_16417,N_16468);
nor U16575 (N_16575,N_16325,N_16467);
and U16576 (N_16576,N_16451,N_16383);
nand U16577 (N_16577,N_16367,N_16338);
nor U16578 (N_16578,N_16378,N_16358);
nand U16579 (N_16579,N_16377,N_16338);
xor U16580 (N_16580,N_16432,N_16329);
nand U16581 (N_16581,N_16477,N_16377);
or U16582 (N_16582,N_16449,N_16375);
nor U16583 (N_16583,N_16345,N_16428);
and U16584 (N_16584,N_16421,N_16349);
nand U16585 (N_16585,N_16455,N_16450);
or U16586 (N_16586,N_16402,N_16478);
nand U16587 (N_16587,N_16435,N_16374);
nor U16588 (N_16588,N_16460,N_16455);
or U16589 (N_16589,N_16356,N_16345);
nand U16590 (N_16590,N_16462,N_16363);
and U16591 (N_16591,N_16344,N_16369);
or U16592 (N_16592,N_16346,N_16416);
xor U16593 (N_16593,N_16459,N_16327);
nand U16594 (N_16594,N_16413,N_16479);
nor U16595 (N_16595,N_16372,N_16444);
nor U16596 (N_16596,N_16332,N_16443);
or U16597 (N_16597,N_16450,N_16412);
and U16598 (N_16598,N_16378,N_16376);
xnor U16599 (N_16599,N_16380,N_16340);
and U16600 (N_16600,N_16350,N_16384);
and U16601 (N_16601,N_16330,N_16401);
nor U16602 (N_16602,N_16327,N_16340);
nor U16603 (N_16603,N_16332,N_16396);
and U16604 (N_16604,N_16414,N_16384);
and U16605 (N_16605,N_16462,N_16361);
xnor U16606 (N_16606,N_16460,N_16396);
nor U16607 (N_16607,N_16472,N_16360);
xor U16608 (N_16608,N_16441,N_16366);
or U16609 (N_16609,N_16381,N_16352);
or U16610 (N_16610,N_16354,N_16356);
xor U16611 (N_16611,N_16428,N_16471);
and U16612 (N_16612,N_16406,N_16376);
xor U16613 (N_16613,N_16384,N_16323);
and U16614 (N_16614,N_16448,N_16432);
xnor U16615 (N_16615,N_16446,N_16322);
or U16616 (N_16616,N_16475,N_16327);
xnor U16617 (N_16617,N_16405,N_16344);
and U16618 (N_16618,N_16423,N_16415);
or U16619 (N_16619,N_16342,N_16394);
and U16620 (N_16620,N_16328,N_16430);
or U16621 (N_16621,N_16358,N_16397);
xnor U16622 (N_16622,N_16457,N_16453);
and U16623 (N_16623,N_16392,N_16439);
nor U16624 (N_16624,N_16414,N_16375);
nand U16625 (N_16625,N_16350,N_16342);
or U16626 (N_16626,N_16390,N_16479);
nand U16627 (N_16627,N_16323,N_16341);
nand U16628 (N_16628,N_16466,N_16467);
xor U16629 (N_16629,N_16437,N_16322);
nand U16630 (N_16630,N_16442,N_16373);
xor U16631 (N_16631,N_16412,N_16459);
nand U16632 (N_16632,N_16468,N_16429);
xnor U16633 (N_16633,N_16320,N_16373);
and U16634 (N_16634,N_16459,N_16466);
or U16635 (N_16635,N_16359,N_16366);
nand U16636 (N_16636,N_16416,N_16444);
and U16637 (N_16637,N_16459,N_16323);
nand U16638 (N_16638,N_16328,N_16346);
or U16639 (N_16639,N_16389,N_16431);
nor U16640 (N_16640,N_16623,N_16541);
nand U16641 (N_16641,N_16481,N_16510);
or U16642 (N_16642,N_16587,N_16483);
or U16643 (N_16643,N_16611,N_16598);
and U16644 (N_16644,N_16637,N_16572);
nor U16645 (N_16645,N_16584,N_16561);
or U16646 (N_16646,N_16488,N_16624);
xnor U16647 (N_16647,N_16616,N_16563);
nand U16648 (N_16648,N_16582,N_16524);
xnor U16649 (N_16649,N_16580,N_16634);
or U16650 (N_16650,N_16608,N_16631);
nand U16651 (N_16651,N_16602,N_16539);
xnor U16652 (N_16652,N_16540,N_16530);
nand U16653 (N_16653,N_16484,N_16621);
nor U16654 (N_16654,N_16565,N_16523);
nor U16655 (N_16655,N_16490,N_16542);
nand U16656 (N_16656,N_16566,N_16562);
or U16657 (N_16657,N_16569,N_16532);
xnor U16658 (N_16658,N_16609,N_16491);
and U16659 (N_16659,N_16589,N_16633);
xnor U16660 (N_16660,N_16612,N_16525);
nand U16661 (N_16661,N_16546,N_16513);
or U16662 (N_16662,N_16489,N_16570);
or U16663 (N_16663,N_16578,N_16617);
nand U16664 (N_16664,N_16629,N_16554);
and U16665 (N_16665,N_16552,N_16636);
xnor U16666 (N_16666,N_16596,N_16494);
nor U16667 (N_16667,N_16568,N_16529);
or U16668 (N_16668,N_16545,N_16620);
nand U16669 (N_16669,N_16543,N_16625);
nor U16670 (N_16670,N_16507,N_16506);
nand U16671 (N_16671,N_16607,N_16597);
xor U16672 (N_16672,N_16614,N_16590);
and U16673 (N_16673,N_16618,N_16533);
nand U16674 (N_16674,N_16535,N_16610);
or U16675 (N_16675,N_16586,N_16601);
nand U16676 (N_16676,N_16505,N_16503);
nand U16677 (N_16677,N_16560,N_16514);
or U16678 (N_16678,N_16551,N_16604);
nor U16679 (N_16679,N_16579,N_16512);
and U16680 (N_16680,N_16504,N_16564);
or U16681 (N_16681,N_16583,N_16613);
and U16682 (N_16682,N_16549,N_16509);
and U16683 (N_16683,N_16559,N_16515);
or U16684 (N_16684,N_16526,N_16627);
nand U16685 (N_16685,N_16577,N_16605);
and U16686 (N_16686,N_16594,N_16606);
nor U16687 (N_16687,N_16635,N_16518);
xnor U16688 (N_16688,N_16585,N_16521);
or U16689 (N_16689,N_16638,N_16499);
xnor U16690 (N_16690,N_16573,N_16544);
and U16691 (N_16691,N_16557,N_16599);
and U16692 (N_16692,N_16622,N_16520);
nor U16693 (N_16693,N_16528,N_16511);
and U16694 (N_16694,N_16496,N_16516);
and U16695 (N_16695,N_16547,N_16500);
xnor U16696 (N_16696,N_16498,N_16630);
and U16697 (N_16697,N_16501,N_16576);
nand U16698 (N_16698,N_16522,N_16619);
and U16699 (N_16699,N_16493,N_16567);
nor U16700 (N_16700,N_16592,N_16508);
and U16701 (N_16701,N_16639,N_16555);
nand U16702 (N_16702,N_16527,N_16497);
xnor U16703 (N_16703,N_16603,N_16574);
nand U16704 (N_16704,N_16593,N_16575);
nor U16705 (N_16705,N_16519,N_16492);
nand U16706 (N_16706,N_16480,N_16517);
nor U16707 (N_16707,N_16534,N_16553);
nor U16708 (N_16708,N_16571,N_16550);
or U16709 (N_16709,N_16626,N_16588);
or U16710 (N_16710,N_16600,N_16615);
or U16711 (N_16711,N_16482,N_16632);
xnor U16712 (N_16712,N_16595,N_16495);
or U16713 (N_16713,N_16486,N_16531);
xor U16714 (N_16714,N_16548,N_16537);
or U16715 (N_16715,N_16591,N_16538);
nor U16716 (N_16716,N_16502,N_16536);
and U16717 (N_16717,N_16558,N_16581);
xnor U16718 (N_16718,N_16487,N_16556);
or U16719 (N_16719,N_16628,N_16485);
and U16720 (N_16720,N_16590,N_16497);
nand U16721 (N_16721,N_16597,N_16559);
xnor U16722 (N_16722,N_16607,N_16593);
xnor U16723 (N_16723,N_16615,N_16552);
nor U16724 (N_16724,N_16592,N_16617);
or U16725 (N_16725,N_16548,N_16530);
nand U16726 (N_16726,N_16598,N_16526);
nand U16727 (N_16727,N_16589,N_16527);
xnor U16728 (N_16728,N_16625,N_16604);
and U16729 (N_16729,N_16598,N_16639);
nand U16730 (N_16730,N_16499,N_16550);
nor U16731 (N_16731,N_16610,N_16626);
or U16732 (N_16732,N_16505,N_16578);
or U16733 (N_16733,N_16524,N_16521);
or U16734 (N_16734,N_16586,N_16573);
nand U16735 (N_16735,N_16566,N_16610);
xor U16736 (N_16736,N_16568,N_16554);
or U16737 (N_16737,N_16624,N_16638);
nand U16738 (N_16738,N_16595,N_16625);
nand U16739 (N_16739,N_16576,N_16495);
xor U16740 (N_16740,N_16488,N_16536);
xor U16741 (N_16741,N_16582,N_16558);
xor U16742 (N_16742,N_16504,N_16604);
nand U16743 (N_16743,N_16558,N_16639);
or U16744 (N_16744,N_16572,N_16567);
or U16745 (N_16745,N_16596,N_16553);
xnor U16746 (N_16746,N_16506,N_16524);
xnor U16747 (N_16747,N_16529,N_16506);
or U16748 (N_16748,N_16607,N_16491);
nand U16749 (N_16749,N_16497,N_16570);
nor U16750 (N_16750,N_16556,N_16566);
nand U16751 (N_16751,N_16619,N_16598);
nor U16752 (N_16752,N_16567,N_16486);
nand U16753 (N_16753,N_16487,N_16494);
nand U16754 (N_16754,N_16627,N_16552);
xor U16755 (N_16755,N_16577,N_16571);
or U16756 (N_16756,N_16498,N_16500);
nand U16757 (N_16757,N_16538,N_16580);
nor U16758 (N_16758,N_16617,N_16549);
nand U16759 (N_16759,N_16594,N_16508);
or U16760 (N_16760,N_16569,N_16638);
nor U16761 (N_16761,N_16582,N_16638);
nor U16762 (N_16762,N_16635,N_16544);
and U16763 (N_16763,N_16507,N_16628);
xor U16764 (N_16764,N_16590,N_16507);
xnor U16765 (N_16765,N_16546,N_16492);
nand U16766 (N_16766,N_16636,N_16522);
xor U16767 (N_16767,N_16619,N_16611);
or U16768 (N_16768,N_16503,N_16494);
or U16769 (N_16769,N_16498,N_16502);
nand U16770 (N_16770,N_16628,N_16538);
nand U16771 (N_16771,N_16540,N_16485);
and U16772 (N_16772,N_16554,N_16538);
nor U16773 (N_16773,N_16502,N_16609);
nand U16774 (N_16774,N_16602,N_16615);
nor U16775 (N_16775,N_16627,N_16553);
nand U16776 (N_16776,N_16635,N_16631);
nand U16777 (N_16777,N_16541,N_16581);
nand U16778 (N_16778,N_16534,N_16570);
xnor U16779 (N_16779,N_16610,N_16634);
nor U16780 (N_16780,N_16515,N_16555);
or U16781 (N_16781,N_16481,N_16579);
nor U16782 (N_16782,N_16572,N_16609);
nor U16783 (N_16783,N_16634,N_16618);
nor U16784 (N_16784,N_16547,N_16635);
and U16785 (N_16785,N_16574,N_16506);
xor U16786 (N_16786,N_16629,N_16515);
nor U16787 (N_16787,N_16536,N_16484);
nor U16788 (N_16788,N_16492,N_16559);
or U16789 (N_16789,N_16624,N_16547);
xnor U16790 (N_16790,N_16566,N_16528);
or U16791 (N_16791,N_16520,N_16509);
nand U16792 (N_16792,N_16598,N_16538);
and U16793 (N_16793,N_16592,N_16502);
and U16794 (N_16794,N_16521,N_16494);
nand U16795 (N_16795,N_16591,N_16624);
and U16796 (N_16796,N_16592,N_16504);
and U16797 (N_16797,N_16569,N_16524);
or U16798 (N_16798,N_16529,N_16517);
and U16799 (N_16799,N_16482,N_16548);
nand U16800 (N_16800,N_16649,N_16730);
nor U16801 (N_16801,N_16647,N_16791);
xor U16802 (N_16802,N_16675,N_16793);
xnor U16803 (N_16803,N_16714,N_16657);
and U16804 (N_16804,N_16758,N_16690);
and U16805 (N_16805,N_16781,N_16694);
and U16806 (N_16806,N_16787,N_16754);
or U16807 (N_16807,N_16679,N_16670);
xor U16808 (N_16808,N_16705,N_16764);
nand U16809 (N_16809,N_16671,N_16742);
nor U16810 (N_16810,N_16662,N_16652);
and U16811 (N_16811,N_16646,N_16772);
nand U16812 (N_16812,N_16777,N_16704);
nor U16813 (N_16813,N_16729,N_16760);
nand U16814 (N_16814,N_16737,N_16786);
xnor U16815 (N_16815,N_16677,N_16695);
or U16816 (N_16816,N_16718,N_16715);
and U16817 (N_16817,N_16792,N_16667);
xnor U16818 (N_16818,N_16698,N_16726);
nor U16819 (N_16819,N_16684,N_16768);
or U16820 (N_16820,N_16683,N_16798);
and U16821 (N_16821,N_16733,N_16753);
nor U16822 (N_16822,N_16750,N_16748);
nand U16823 (N_16823,N_16776,N_16680);
nor U16824 (N_16824,N_16645,N_16672);
nand U16825 (N_16825,N_16736,N_16743);
nand U16826 (N_16826,N_16745,N_16659);
or U16827 (N_16827,N_16713,N_16767);
or U16828 (N_16828,N_16644,N_16785);
nand U16829 (N_16829,N_16681,N_16719);
xnor U16830 (N_16830,N_16725,N_16751);
nor U16831 (N_16831,N_16693,N_16707);
or U16832 (N_16832,N_16642,N_16674);
nor U16833 (N_16833,N_16689,N_16727);
xnor U16834 (N_16834,N_16685,N_16789);
nor U16835 (N_16835,N_16778,N_16716);
and U16836 (N_16836,N_16722,N_16796);
xnor U16837 (N_16837,N_16773,N_16752);
nand U16838 (N_16838,N_16676,N_16782);
nand U16839 (N_16839,N_16757,N_16660);
and U16840 (N_16840,N_16643,N_16756);
and U16841 (N_16841,N_16720,N_16653);
and U16842 (N_16842,N_16711,N_16759);
nand U16843 (N_16843,N_16721,N_16666);
or U16844 (N_16844,N_16700,N_16774);
nand U16845 (N_16845,N_16784,N_16769);
xnor U16846 (N_16846,N_16740,N_16738);
nand U16847 (N_16847,N_16797,N_16708);
xnor U16848 (N_16848,N_16651,N_16661);
and U16849 (N_16849,N_16795,N_16664);
and U16850 (N_16850,N_16678,N_16744);
xor U16851 (N_16851,N_16691,N_16766);
and U16852 (N_16852,N_16702,N_16741);
nor U16853 (N_16853,N_16663,N_16731);
or U16854 (N_16854,N_16739,N_16710);
xor U16855 (N_16855,N_16656,N_16723);
or U16856 (N_16856,N_16701,N_16790);
nor U16857 (N_16857,N_16775,N_16779);
nor U16858 (N_16858,N_16697,N_16709);
or U16859 (N_16859,N_16735,N_16706);
or U16860 (N_16860,N_16640,N_16762);
nor U16861 (N_16861,N_16771,N_16692);
xnor U16862 (N_16862,N_16765,N_16712);
nor U16863 (N_16863,N_16699,N_16682);
nor U16864 (N_16864,N_16717,N_16770);
or U16865 (N_16865,N_16780,N_16761);
or U16866 (N_16866,N_16788,N_16650);
nand U16867 (N_16867,N_16673,N_16783);
or U16868 (N_16868,N_16668,N_16669);
xor U16869 (N_16869,N_16665,N_16658);
nand U16870 (N_16870,N_16724,N_16654);
and U16871 (N_16871,N_16749,N_16688);
nand U16872 (N_16872,N_16696,N_16687);
nand U16873 (N_16873,N_16641,N_16728);
nor U16874 (N_16874,N_16755,N_16794);
nand U16875 (N_16875,N_16686,N_16746);
nor U16876 (N_16876,N_16732,N_16799);
nand U16877 (N_16877,N_16747,N_16734);
nor U16878 (N_16878,N_16648,N_16703);
and U16879 (N_16879,N_16655,N_16763);
or U16880 (N_16880,N_16768,N_16767);
nand U16881 (N_16881,N_16715,N_16676);
or U16882 (N_16882,N_16729,N_16732);
and U16883 (N_16883,N_16719,N_16657);
or U16884 (N_16884,N_16640,N_16755);
or U16885 (N_16885,N_16713,N_16676);
and U16886 (N_16886,N_16731,N_16697);
or U16887 (N_16887,N_16706,N_16695);
nand U16888 (N_16888,N_16783,N_16696);
nor U16889 (N_16889,N_16669,N_16773);
nor U16890 (N_16890,N_16752,N_16782);
and U16891 (N_16891,N_16692,N_16707);
nand U16892 (N_16892,N_16760,N_16744);
and U16893 (N_16893,N_16650,N_16672);
or U16894 (N_16894,N_16739,N_16751);
nor U16895 (N_16895,N_16730,N_16750);
or U16896 (N_16896,N_16774,N_16681);
nand U16897 (N_16897,N_16712,N_16734);
and U16898 (N_16898,N_16701,N_16719);
or U16899 (N_16899,N_16651,N_16663);
and U16900 (N_16900,N_16659,N_16774);
xor U16901 (N_16901,N_16711,N_16658);
nor U16902 (N_16902,N_16702,N_16747);
and U16903 (N_16903,N_16698,N_16706);
xor U16904 (N_16904,N_16684,N_16723);
xor U16905 (N_16905,N_16798,N_16766);
nor U16906 (N_16906,N_16642,N_16792);
nor U16907 (N_16907,N_16707,N_16750);
or U16908 (N_16908,N_16709,N_16661);
xnor U16909 (N_16909,N_16712,N_16691);
and U16910 (N_16910,N_16767,N_16695);
xor U16911 (N_16911,N_16753,N_16773);
xnor U16912 (N_16912,N_16799,N_16755);
or U16913 (N_16913,N_16727,N_16690);
or U16914 (N_16914,N_16652,N_16725);
and U16915 (N_16915,N_16662,N_16791);
and U16916 (N_16916,N_16678,N_16764);
nor U16917 (N_16917,N_16744,N_16738);
nand U16918 (N_16918,N_16767,N_16722);
nor U16919 (N_16919,N_16771,N_16688);
nand U16920 (N_16920,N_16766,N_16659);
and U16921 (N_16921,N_16733,N_16697);
and U16922 (N_16922,N_16774,N_16648);
nand U16923 (N_16923,N_16789,N_16694);
and U16924 (N_16924,N_16710,N_16735);
and U16925 (N_16925,N_16708,N_16715);
nand U16926 (N_16926,N_16669,N_16730);
nand U16927 (N_16927,N_16681,N_16687);
nand U16928 (N_16928,N_16678,N_16688);
nor U16929 (N_16929,N_16770,N_16735);
nand U16930 (N_16930,N_16793,N_16752);
nor U16931 (N_16931,N_16772,N_16770);
nand U16932 (N_16932,N_16748,N_16768);
and U16933 (N_16933,N_16721,N_16732);
and U16934 (N_16934,N_16782,N_16683);
nand U16935 (N_16935,N_16654,N_16714);
or U16936 (N_16936,N_16762,N_16739);
or U16937 (N_16937,N_16688,N_16777);
xnor U16938 (N_16938,N_16724,N_16649);
and U16939 (N_16939,N_16669,N_16657);
or U16940 (N_16940,N_16747,N_16658);
xnor U16941 (N_16941,N_16651,N_16799);
nand U16942 (N_16942,N_16703,N_16770);
or U16943 (N_16943,N_16644,N_16727);
nor U16944 (N_16944,N_16783,N_16709);
nor U16945 (N_16945,N_16770,N_16734);
nand U16946 (N_16946,N_16721,N_16789);
or U16947 (N_16947,N_16650,N_16727);
nor U16948 (N_16948,N_16799,N_16653);
xnor U16949 (N_16949,N_16785,N_16757);
and U16950 (N_16950,N_16684,N_16642);
nor U16951 (N_16951,N_16794,N_16714);
and U16952 (N_16952,N_16752,N_16775);
xor U16953 (N_16953,N_16728,N_16766);
xnor U16954 (N_16954,N_16789,N_16760);
or U16955 (N_16955,N_16658,N_16657);
or U16956 (N_16956,N_16667,N_16691);
or U16957 (N_16957,N_16776,N_16675);
and U16958 (N_16958,N_16647,N_16692);
and U16959 (N_16959,N_16728,N_16774);
and U16960 (N_16960,N_16935,N_16954);
nor U16961 (N_16961,N_16848,N_16822);
or U16962 (N_16962,N_16886,N_16811);
and U16963 (N_16963,N_16933,N_16882);
nand U16964 (N_16964,N_16813,N_16930);
and U16965 (N_16965,N_16948,N_16911);
nor U16966 (N_16966,N_16940,N_16898);
or U16967 (N_16967,N_16836,N_16835);
nor U16968 (N_16968,N_16870,N_16864);
xor U16969 (N_16969,N_16901,N_16957);
and U16970 (N_16970,N_16927,N_16907);
nand U16971 (N_16971,N_16863,N_16847);
nor U16972 (N_16972,N_16902,N_16910);
and U16973 (N_16973,N_16939,N_16909);
or U16974 (N_16974,N_16956,N_16936);
nand U16975 (N_16975,N_16887,N_16873);
and U16976 (N_16976,N_16819,N_16807);
nand U16977 (N_16977,N_16913,N_16867);
nor U16978 (N_16978,N_16820,N_16818);
and U16979 (N_16979,N_16938,N_16841);
nor U16980 (N_16980,N_16879,N_16843);
xnor U16981 (N_16981,N_16949,N_16832);
nand U16982 (N_16982,N_16850,N_16888);
xnor U16983 (N_16983,N_16905,N_16906);
xor U16984 (N_16984,N_16868,N_16830);
nand U16985 (N_16985,N_16885,N_16849);
nand U16986 (N_16986,N_16871,N_16881);
or U16987 (N_16987,N_16800,N_16853);
or U16988 (N_16988,N_16892,N_16904);
xnor U16989 (N_16989,N_16840,N_16896);
and U16990 (N_16990,N_16923,N_16953);
and U16991 (N_16991,N_16816,N_16918);
and U16992 (N_16992,N_16903,N_16883);
nand U16993 (N_16993,N_16947,N_16890);
xnor U16994 (N_16994,N_16893,N_16854);
and U16995 (N_16995,N_16929,N_16937);
nor U16996 (N_16996,N_16814,N_16812);
or U16997 (N_16997,N_16931,N_16869);
and U16998 (N_16998,N_16915,N_16926);
xnor U16999 (N_16999,N_16861,N_16874);
nor U17000 (N_17000,N_16922,N_16808);
and U17001 (N_17001,N_16838,N_16855);
or U17002 (N_17002,N_16803,N_16859);
and U17003 (N_17003,N_16846,N_16959);
nor U17004 (N_17004,N_16875,N_16815);
xor U17005 (N_17005,N_16851,N_16942);
or U17006 (N_17006,N_16834,N_16857);
and U17007 (N_17007,N_16884,N_16845);
nand U17008 (N_17008,N_16878,N_16920);
nand U17009 (N_17009,N_16856,N_16829);
xor U17010 (N_17010,N_16862,N_16865);
and U17011 (N_17011,N_16943,N_16806);
nor U17012 (N_17012,N_16925,N_16833);
and U17013 (N_17013,N_16919,N_16950);
nor U17014 (N_17014,N_16952,N_16889);
and U17015 (N_17015,N_16928,N_16821);
xor U17016 (N_17016,N_16916,N_16858);
xor U17017 (N_17017,N_16955,N_16932);
nor U17018 (N_17018,N_16945,N_16917);
or U17019 (N_17019,N_16852,N_16891);
xnor U17020 (N_17020,N_16877,N_16866);
and U17021 (N_17021,N_16880,N_16827);
or U17022 (N_17022,N_16946,N_16908);
nand U17023 (N_17023,N_16899,N_16921);
xnor U17024 (N_17024,N_16839,N_16824);
nor U17025 (N_17025,N_16831,N_16900);
or U17026 (N_17026,N_16801,N_16944);
nand U17027 (N_17027,N_16895,N_16897);
or U17028 (N_17028,N_16941,N_16872);
nor U17029 (N_17029,N_16951,N_16912);
xnor U17030 (N_17030,N_16817,N_16809);
and U17031 (N_17031,N_16810,N_16837);
or U17032 (N_17032,N_16805,N_16825);
or U17033 (N_17033,N_16924,N_16934);
and U17034 (N_17034,N_16914,N_16804);
and U17035 (N_17035,N_16894,N_16802);
xor U17036 (N_17036,N_16828,N_16826);
nor U17037 (N_17037,N_16860,N_16842);
or U17038 (N_17038,N_16876,N_16958);
nand U17039 (N_17039,N_16844,N_16823);
and U17040 (N_17040,N_16895,N_16950);
or U17041 (N_17041,N_16887,N_16825);
nor U17042 (N_17042,N_16931,N_16914);
or U17043 (N_17043,N_16879,N_16827);
xor U17044 (N_17044,N_16876,N_16808);
xnor U17045 (N_17045,N_16844,N_16818);
xnor U17046 (N_17046,N_16805,N_16911);
xor U17047 (N_17047,N_16808,N_16891);
nor U17048 (N_17048,N_16821,N_16805);
nand U17049 (N_17049,N_16915,N_16816);
nor U17050 (N_17050,N_16913,N_16944);
or U17051 (N_17051,N_16943,N_16836);
xnor U17052 (N_17052,N_16908,N_16928);
nor U17053 (N_17053,N_16959,N_16805);
xor U17054 (N_17054,N_16922,N_16950);
nor U17055 (N_17055,N_16863,N_16835);
nand U17056 (N_17056,N_16950,N_16906);
nand U17057 (N_17057,N_16875,N_16907);
xor U17058 (N_17058,N_16814,N_16824);
or U17059 (N_17059,N_16842,N_16867);
nor U17060 (N_17060,N_16929,N_16827);
or U17061 (N_17061,N_16836,N_16938);
nor U17062 (N_17062,N_16882,N_16890);
and U17063 (N_17063,N_16888,N_16920);
nor U17064 (N_17064,N_16867,N_16818);
nand U17065 (N_17065,N_16887,N_16813);
or U17066 (N_17066,N_16838,N_16949);
nor U17067 (N_17067,N_16881,N_16911);
and U17068 (N_17068,N_16873,N_16928);
nand U17069 (N_17069,N_16917,N_16883);
and U17070 (N_17070,N_16809,N_16850);
xor U17071 (N_17071,N_16954,N_16864);
nand U17072 (N_17072,N_16852,N_16929);
nor U17073 (N_17073,N_16856,N_16890);
or U17074 (N_17074,N_16842,N_16824);
nor U17075 (N_17075,N_16897,N_16851);
and U17076 (N_17076,N_16916,N_16937);
xnor U17077 (N_17077,N_16944,N_16956);
or U17078 (N_17078,N_16830,N_16842);
nor U17079 (N_17079,N_16902,N_16934);
nand U17080 (N_17080,N_16852,N_16883);
xor U17081 (N_17081,N_16807,N_16839);
and U17082 (N_17082,N_16938,N_16945);
and U17083 (N_17083,N_16841,N_16906);
nor U17084 (N_17084,N_16878,N_16811);
nor U17085 (N_17085,N_16908,N_16916);
xor U17086 (N_17086,N_16922,N_16810);
nor U17087 (N_17087,N_16837,N_16901);
nor U17088 (N_17088,N_16836,N_16807);
nand U17089 (N_17089,N_16808,N_16945);
and U17090 (N_17090,N_16908,N_16947);
nand U17091 (N_17091,N_16858,N_16839);
nor U17092 (N_17092,N_16856,N_16842);
nand U17093 (N_17093,N_16958,N_16807);
nor U17094 (N_17094,N_16928,N_16943);
nand U17095 (N_17095,N_16829,N_16957);
or U17096 (N_17096,N_16812,N_16888);
or U17097 (N_17097,N_16804,N_16835);
nor U17098 (N_17098,N_16805,N_16915);
xor U17099 (N_17099,N_16948,N_16914);
and U17100 (N_17100,N_16859,N_16822);
or U17101 (N_17101,N_16881,N_16926);
or U17102 (N_17102,N_16822,N_16808);
nand U17103 (N_17103,N_16898,N_16957);
or U17104 (N_17104,N_16941,N_16846);
and U17105 (N_17105,N_16859,N_16853);
nor U17106 (N_17106,N_16831,N_16824);
nor U17107 (N_17107,N_16839,N_16853);
and U17108 (N_17108,N_16857,N_16827);
xnor U17109 (N_17109,N_16881,N_16936);
xor U17110 (N_17110,N_16835,N_16806);
and U17111 (N_17111,N_16818,N_16908);
nor U17112 (N_17112,N_16944,N_16843);
xnor U17113 (N_17113,N_16925,N_16872);
nor U17114 (N_17114,N_16915,N_16866);
nor U17115 (N_17115,N_16863,N_16884);
nand U17116 (N_17116,N_16890,N_16933);
xor U17117 (N_17117,N_16813,N_16919);
nand U17118 (N_17118,N_16939,N_16848);
nand U17119 (N_17119,N_16819,N_16865);
xnor U17120 (N_17120,N_16996,N_17044);
nor U17121 (N_17121,N_17114,N_17059);
or U17122 (N_17122,N_17010,N_17111);
nor U17123 (N_17123,N_17066,N_17116);
or U17124 (N_17124,N_17039,N_17004);
nor U17125 (N_17125,N_17074,N_17043);
nand U17126 (N_17126,N_16989,N_16967);
and U17127 (N_17127,N_16962,N_16994);
and U17128 (N_17128,N_17050,N_17042);
or U17129 (N_17129,N_17073,N_17086);
or U17130 (N_17130,N_16984,N_17077);
nand U17131 (N_17131,N_17033,N_17089);
and U17132 (N_17132,N_17037,N_17031);
nand U17133 (N_17133,N_16990,N_17081);
nand U17134 (N_17134,N_17021,N_17094);
and U17135 (N_17135,N_17075,N_17061);
and U17136 (N_17136,N_17102,N_17062);
and U17137 (N_17137,N_16993,N_17014);
nand U17138 (N_17138,N_17057,N_17012);
or U17139 (N_17139,N_17065,N_17008);
nand U17140 (N_17140,N_17001,N_16997);
nand U17141 (N_17141,N_17119,N_17015);
and U17142 (N_17142,N_17090,N_17003);
and U17143 (N_17143,N_17082,N_17006);
and U17144 (N_17144,N_17052,N_17105);
and U17145 (N_17145,N_17005,N_17067);
nor U17146 (N_17146,N_17013,N_17106);
and U17147 (N_17147,N_17071,N_17099);
and U17148 (N_17148,N_17007,N_16999);
and U17149 (N_17149,N_17040,N_16966);
xor U17150 (N_17150,N_17097,N_16983);
nand U17151 (N_17151,N_16976,N_16965);
nor U17152 (N_17152,N_17038,N_17104);
or U17153 (N_17153,N_17023,N_17109);
nand U17154 (N_17154,N_17095,N_17103);
and U17155 (N_17155,N_16968,N_17088);
xor U17156 (N_17156,N_17063,N_17055);
or U17157 (N_17157,N_17058,N_16960);
and U17158 (N_17158,N_17064,N_17087);
nand U17159 (N_17159,N_17049,N_16981);
xnor U17160 (N_17160,N_17002,N_17026);
xnor U17161 (N_17161,N_17072,N_17076);
or U17162 (N_17162,N_17027,N_17020);
xnor U17163 (N_17163,N_17011,N_17115);
or U17164 (N_17164,N_16988,N_16970);
nand U17165 (N_17165,N_16985,N_16980);
and U17166 (N_17166,N_16995,N_16978);
or U17167 (N_17167,N_17112,N_17069);
or U17168 (N_17168,N_16974,N_16964);
and U17169 (N_17169,N_16986,N_17035);
and U17170 (N_17170,N_16992,N_17117);
nor U17171 (N_17171,N_17100,N_16969);
or U17172 (N_17172,N_17022,N_17048);
and U17173 (N_17173,N_17017,N_17018);
nor U17174 (N_17174,N_17110,N_17034);
xor U17175 (N_17175,N_17098,N_17030);
and U17176 (N_17176,N_17080,N_17084);
nand U17177 (N_17177,N_16987,N_16977);
or U17178 (N_17178,N_16998,N_17047);
xor U17179 (N_17179,N_16979,N_17036);
and U17180 (N_17180,N_17113,N_17032);
or U17181 (N_17181,N_17107,N_17028);
or U17182 (N_17182,N_16991,N_17108);
xor U17183 (N_17183,N_17068,N_17085);
and U17184 (N_17184,N_17118,N_17009);
or U17185 (N_17185,N_17041,N_17046);
xor U17186 (N_17186,N_17016,N_16972);
nand U17187 (N_17187,N_17092,N_17060);
and U17188 (N_17188,N_16961,N_17025);
xor U17189 (N_17189,N_16971,N_17078);
xor U17190 (N_17190,N_17029,N_17053);
nand U17191 (N_17191,N_17019,N_17051);
and U17192 (N_17192,N_17093,N_17000);
nand U17193 (N_17193,N_17091,N_17054);
nand U17194 (N_17194,N_17024,N_16982);
xnor U17195 (N_17195,N_17056,N_17083);
and U17196 (N_17196,N_17096,N_16973);
nand U17197 (N_17197,N_17045,N_16975);
and U17198 (N_17198,N_16963,N_17070);
xnor U17199 (N_17199,N_17079,N_17101);
xor U17200 (N_17200,N_16979,N_17079);
nand U17201 (N_17201,N_17018,N_17083);
nand U17202 (N_17202,N_17049,N_16989);
or U17203 (N_17203,N_17002,N_17103);
and U17204 (N_17204,N_17086,N_17043);
xor U17205 (N_17205,N_17110,N_17019);
xnor U17206 (N_17206,N_17045,N_17061);
or U17207 (N_17207,N_17101,N_17094);
or U17208 (N_17208,N_16973,N_17117);
nand U17209 (N_17209,N_16974,N_17012);
or U17210 (N_17210,N_17093,N_17047);
xor U17211 (N_17211,N_16970,N_17029);
nand U17212 (N_17212,N_17118,N_17057);
nand U17213 (N_17213,N_17037,N_17008);
nand U17214 (N_17214,N_16995,N_17065);
nand U17215 (N_17215,N_17117,N_17043);
xnor U17216 (N_17216,N_17029,N_17012);
nor U17217 (N_17217,N_17031,N_17052);
and U17218 (N_17218,N_16977,N_17066);
or U17219 (N_17219,N_16967,N_16983);
xnor U17220 (N_17220,N_17070,N_17110);
or U17221 (N_17221,N_17102,N_17114);
and U17222 (N_17222,N_16980,N_17114);
nor U17223 (N_17223,N_17027,N_17054);
or U17224 (N_17224,N_17011,N_17116);
xnor U17225 (N_17225,N_17065,N_16999);
or U17226 (N_17226,N_17061,N_17087);
or U17227 (N_17227,N_17102,N_16977);
nand U17228 (N_17228,N_16985,N_17110);
or U17229 (N_17229,N_17097,N_17111);
or U17230 (N_17230,N_16980,N_17035);
nor U17231 (N_17231,N_17105,N_17113);
xnor U17232 (N_17232,N_16998,N_17053);
xnor U17233 (N_17233,N_17010,N_17064);
nand U17234 (N_17234,N_17055,N_16984);
nand U17235 (N_17235,N_16987,N_16996);
or U17236 (N_17236,N_17084,N_17076);
nor U17237 (N_17237,N_17095,N_17075);
xnor U17238 (N_17238,N_17119,N_17045);
nand U17239 (N_17239,N_17057,N_17074);
xor U17240 (N_17240,N_17041,N_17062);
nand U17241 (N_17241,N_17106,N_17103);
and U17242 (N_17242,N_17066,N_16993);
or U17243 (N_17243,N_17013,N_17022);
nor U17244 (N_17244,N_17083,N_16980);
and U17245 (N_17245,N_17006,N_17043);
and U17246 (N_17246,N_16990,N_17082);
xor U17247 (N_17247,N_16970,N_17032);
or U17248 (N_17248,N_17022,N_17064);
or U17249 (N_17249,N_17036,N_16982);
and U17250 (N_17250,N_16990,N_17044);
and U17251 (N_17251,N_16971,N_17021);
or U17252 (N_17252,N_17068,N_17088);
and U17253 (N_17253,N_17074,N_17069);
nand U17254 (N_17254,N_17104,N_17001);
nor U17255 (N_17255,N_17101,N_17015);
xnor U17256 (N_17256,N_17026,N_17053);
and U17257 (N_17257,N_16990,N_16999);
xor U17258 (N_17258,N_17065,N_16969);
or U17259 (N_17259,N_16983,N_17053);
xor U17260 (N_17260,N_17027,N_17083);
xnor U17261 (N_17261,N_17063,N_16984);
or U17262 (N_17262,N_16996,N_16995);
nand U17263 (N_17263,N_17100,N_17065);
nand U17264 (N_17264,N_17094,N_17010);
nor U17265 (N_17265,N_17019,N_17118);
and U17266 (N_17266,N_16976,N_17092);
and U17267 (N_17267,N_17103,N_17076);
nor U17268 (N_17268,N_17009,N_17034);
and U17269 (N_17269,N_17020,N_17019);
nor U17270 (N_17270,N_17097,N_17071);
and U17271 (N_17271,N_17053,N_17002);
and U17272 (N_17272,N_16993,N_16961);
nand U17273 (N_17273,N_17053,N_17062);
nand U17274 (N_17274,N_17057,N_17060);
or U17275 (N_17275,N_17073,N_16966);
nor U17276 (N_17276,N_16987,N_17041);
nand U17277 (N_17277,N_17023,N_17118);
and U17278 (N_17278,N_16993,N_16990);
xor U17279 (N_17279,N_17074,N_16983);
and U17280 (N_17280,N_17271,N_17277);
and U17281 (N_17281,N_17264,N_17128);
nand U17282 (N_17282,N_17265,N_17208);
nand U17283 (N_17283,N_17240,N_17153);
xnor U17284 (N_17284,N_17256,N_17231);
xnor U17285 (N_17285,N_17195,N_17201);
or U17286 (N_17286,N_17272,N_17234);
and U17287 (N_17287,N_17155,N_17172);
or U17288 (N_17288,N_17185,N_17204);
and U17289 (N_17289,N_17138,N_17224);
and U17290 (N_17290,N_17170,N_17164);
nor U17291 (N_17291,N_17205,N_17179);
and U17292 (N_17292,N_17122,N_17151);
or U17293 (N_17293,N_17216,N_17140);
nand U17294 (N_17294,N_17182,N_17142);
nand U17295 (N_17295,N_17166,N_17251);
nand U17296 (N_17296,N_17167,N_17202);
or U17297 (N_17297,N_17220,N_17243);
nor U17298 (N_17298,N_17219,N_17181);
nor U17299 (N_17299,N_17269,N_17248);
nor U17300 (N_17300,N_17250,N_17214);
nand U17301 (N_17301,N_17120,N_17160);
xnor U17302 (N_17302,N_17154,N_17156);
or U17303 (N_17303,N_17162,N_17244);
and U17304 (N_17304,N_17130,N_17279);
or U17305 (N_17305,N_17133,N_17126);
or U17306 (N_17306,N_17207,N_17124);
xnor U17307 (N_17307,N_17253,N_17139);
and U17308 (N_17308,N_17157,N_17144);
or U17309 (N_17309,N_17146,N_17178);
or U17310 (N_17310,N_17136,N_17218);
and U17311 (N_17311,N_17236,N_17221);
and U17312 (N_17312,N_17127,N_17262);
nand U17313 (N_17313,N_17203,N_17230);
and U17314 (N_17314,N_17276,N_17275);
xnor U17315 (N_17315,N_17237,N_17238);
nor U17316 (N_17316,N_17158,N_17186);
and U17317 (N_17317,N_17169,N_17193);
nor U17318 (N_17318,N_17239,N_17165);
and U17319 (N_17319,N_17267,N_17147);
nand U17320 (N_17320,N_17227,N_17266);
nor U17321 (N_17321,N_17190,N_17171);
and U17322 (N_17322,N_17273,N_17168);
nor U17323 (N_17323,N_17192,N_17255);
nor U17324 (N_17324,N_17226,N_17206);
nor U17325 (N_17325,N_17197,N_17247);
xor U17326 (N_17326,N_17199,N_17233);
or U17327 (N_17327,N_17261,N_17232);
nand U17328 (N_17328,N_17198,N_17215);
or U17329 (N_17329,N_17246,N_17184);
and U17330 (N_17330,N_17163,N_17173);
and U17331 (N_17331,N_17148,N_17252);
or U17332 (N_17332,N_17141,N_17210);
xor U17333 (N_17333,N_17209,N_17228);
nand U17334 (N_17334,N_17242,N_17191);
and U17335 (N_17335,N_17121,N_17212);
and U17336 (N_17336,N_17225,N_17260);
or U17337 (N_17337,N_17145,N_17143);
xor U17338 (N_17338,N_17176,N_17200);
or U17339 (N_17339,N_17152,N_17196);
or U17340 (N_17340,N_17188,N_17263);
nand U17341 (N_17341,N_17134,N_17268);
xor U17342 (N_17342,N_17161,N_17180);
or U17343 (N_17343,N_17257,N_17129);
nor U17344 (N_17344,N_17229,N_17258);
nand U17345 (N_17345,N_17241,N_17274);
nor U17346 (N_17346,N_17123,N_17194);
xor U17347 (N_17347,N_17235,N_17249);
nand U17348 (N_17348,N_17189,N_17149);
and U17349 (N_17349,N_17150,N_17174);
xor U17350 (N_17350,N_17159,N_17278);
and U17351 (N_17351,N_17175,N_17245);
and U17352 (N_17352,N_17187,N_17177);
and U17353 (N_17353,N_17217,N_17254);
and U17354 (N_17354,N_17125,N_17135);
xnor U17355 (N_17355,N_17183,N_17131);
nor U17356 (N_17356,N_17137,N_17213);
xnor U17357 (N_17357,N_17132,N_17211);
or U17358 (N_17358,N_17270,N_17223);
nand U17359 (N_17359,N_17222,N_17259);
and U17360 (N_17360,N_17162,N_17137);
and U17361 (N_17361,N_17251,N_17171);
nand U17362 (N_17362,N_17171,N_17200);
or U17363 (N_17363,N_17208,N_17256);
nor U17364 (N_17364,N_17156,N_17195);
and U17365 (N_17365,N_17249,N_17160);
and U17366 (N_17366,N_17223,N_17232);
nand U17367 (N_17367,N_17229,N_17262);
or U17368 (N_17368,N_17264,N_17138);
nor U17369 (N_17369,N_17278,N_17276);
nor U17370 (N_17370,N_17228,N_17170);
and U17371 (N_17371,N_17273,N_17212);
and U17372 (N_17372,N_17128,N_17189);
nand U17373 (N_17373,N_17198,N_17196);
and U17374 (N_17374,N_17141,N_17189);
and U17375 (N_17375,N_17179,N_17184);
and U17376 (N_17376,N_17140,N_17132);
nand U17377 (N_17377,N_17163,N_17241);
nor U17378 (N_17378,N_17139,N_17195);
or U17379 (N_17379,N_17241,N_17186);
nand U17380 (N_17380,N_17215,N_17162);
or U17381 (N_17381,N_17257,N_17143);
nand U17382 (N_17382,N_17242,N_17144);
nor U17383 (N_17383,N_17140,N_17238);
or U17384 (N_17384,N_17157,N_17225);
xor U17385 (N_17385,N_17242,N_17243);
or U17386 (N_17386,N_17142,N_17176);
or U17387 (N_17387,N_17253,N_17160);
nor U17388 (N_17388,N_17209,N_17276);
nor U17389 (N_17389,N_17214,N_17136);
xor U17390 (N_17390,N_17207,N_17269);
or U17391 (N_17391,N_17268,N_17184);
nor U17392 (N_17392,N_17167,N_17124);
nor U17393 (N_17393,N_17192,N_17216);
nor U17394 (N_17394,N_17157,N_17138);
or U17395 (N_17395,N_17130,N_17158);
nor U17396 (N_17396,N_17155,N_17269);
xnor U17397 (N_17397,N_17187,N_17179);
or U17398 (N_17398,N_17237,N_17220);
nand U17399 (N_17399,N_17177,N_17176);
nor U17400 (N_17400,N_17126,N_17258);
xor U17401 (N_17401,N_17199,N_17269);
nor U17402 (N_17402,N_17171,N_17151);
and U17403 (N_17403,N_17137,N_17255);
or U17404 (N_17404,N_17142,N_17159);
and U17405 (N_17405,N_17168,N_17238);
nor U17406 (N_17406,N_17232,N_17216);
nand U17407 (N_17407,N_17251,N_17210);
nor U17408 (N_17408,N_17222,N_17245);
xor U17409 (N_17409,N_17122,N_17264);
or U17410 (N_17410,N_17225,N_17165);
nor U17411 (N_17411,N_17141,N_17173);
nand U17412 (N_17412,N_17220,N_17279);
nor U17413 (N_17413,N_17227,N_17123);
nor U17414 (N_17414,N_17227,N_17132);
nor U17415 (N_17415,N_17268,N_17148);
and U17416 (N_17416,N_17233,N_17227);
nand U17417 (N_17417,N_17224,N_17269);
nand U17418 (N_17418,N_17263,N_17179);
or U17419 (N_17419,N_17159,N_17201);
xnor U17420 (N_17420,N_17230,N_17246);
xnor U17421 (N_17421,N_17124,N_17274);
and U17422 (N_17422,N_17275,N_17218);
and U17423 (N_17423,N_17191,N_17278);
nor U17424 (N_17424,N_17182,N_17189);
nor U17425 (N_17425,N_17182,N_17228);
nand U17426 (N_17426,N_17148,N_17130);
nor U17427 (N_17427,N_17138,N_17189);
or U17428 (N_17428,N_17176,N_17226);
or U17429 (N_17429,N_17259,N_17256);
nor U17430 (N_17430,N_17193,N_17137);
nor U17431 (N_17431,N_17249,N_17124);
or U17432 (N_17432,N_17172,N_17175);
and U17433 (N_17433,N_17131,N_17218);
and U17434 (N_17434,N_17215,N_17257);
nand U17435 (N_17435,N_17218,N_17123);
nand U17436 (N_17436,N_17122,N_17202);
nor U17437 (N_17437,N_17179,N_17149);
and U17438 (N_17438,N_17212,N_17192);
xor U17439 (N_17439,N_17159,N_17239);
nand U17440 (N_17440,N_17371,N_17303);
or U17441 (N_17441,N_17329,N_17335);
nand U17442 (N_17442,N_17432,N_17295);
or U17443 (N_17443,N_17377,N_17393);
or U17444 (N_17444,N_17418,N_17289);
nor U17445 (N_17445,N_17394,N_17398);
or U17446 (N_17446,N_17438,N_17286);
nand U17447 (N_17447,N_17357,N_17334);
nand U17448 (N_17448,N_17387,N_17378);
nand U17449 (N_17449,N_17317,N_17422);
nand U17450 (N_17450,N_17296,N_17281);
and U17451 (N_17451,N_17380,N_17374);
or U17452 (N_17452,N_17407,N_17320);
nand U17453 (N_17453,N_17395,N_17353);
nand U17454 (N_17454,N_17341,N_17330);
nor U17455 (N_17455,N_17434,N_17345);
xnor U17456 (N_17456,N_17304,N_17437);
xnor U17457 (N_17457,N_17429,N_17340);
xor U17458 (N_17458,N_17337,N_17417);
xnor U17459 (N_17459,N_17376,N_17409);
xnor U17460 (N_17460,N_17372,N_17397);
nand U17461 (N_17461,N_17413,N_17318);
xor U17462 (N_17462,N_17389,N_17391);
xnor U17463 (N_17463,N_17399,N_17435);
nand U17464 (N_17464,N_17412,N_17368);
and U17465 (N_17465,N_17439,N_17410);
xnor U17466 (N_17466,N_17373,N_17332);
nand U17467 (N_17467,N_17382,N_17293);
or U17468 (N_17468,N_17356,N_17323);
or U17469 (N_17469,N_17348,N_17384);
or U17470 (N_17470,N_17350,N_17426);
xnor U17471 (N_17471,N_17363,N_17362);
nand U17472 (N_17472,N_17331,N_17325);
or U17473 (N_17473,N_17369,N_17321);
nor U17474 (N_17474,N_17347,N_17421);
nor U17475 (N_17475,N_17388,N_17346);
and U17476 (N_17476,N_17354,N_17342);
and U17477 (N_17477,N_17411,N_17360);
nand U17478 (N_17478,N_17338,N_17367);
or U17479 (N_17479,N_17327,N_17308);
xnor U17480 (N_17480,N_17358,N_17401);
xnor U17481 (N_17481,N_17381,N_17386);
xnor U17482 (N_17482,N_17285,N_17291);
xnor U17483 (N_17483,N_17425,N_17299);
xnor U17484 (N_17484,N_17352,N_17280);
nor U17485 (N_17485,N_17297,N_17423);
xnor U17486 (N_17486,N_17290,N_17316);
or U17487 (N_17487,N_17405,N_17349);
nor U17488 (N_17488,N_17314,N_17390);
xor U17489 (N_17489,N_17305,N_17416);
nand U17490 (N_17490,N_17312,N_17403);
and U17491 (N_17491,N_17336,N_17375);
nand U17492 (N_17492,N_17370,N_17402);
xor U17493 (N_17493,N_17292,N_17315);
nor U17494 (N_17494,N_17379,N_17288);
xnor U17495 (N_17495,N_17400,N_17351);
xor U17496 (N_17496,N_17319,N_17283);
nor U17497 (N_17497,N_17326,N_17428);
nor U17498 (N_17498,N_17436,N_17424);
nand U17499 (N_17499,N_17408,N_17344);
nand U17500 (N_17500,N_17300,N_17383);
xnor U17501 (N_17501,N_17359,N_17406);
and U17502 (N_17502,N_17311,N_17298);
xor U17503 (N_17503,N_17430,N_17301);
nor U17504 (N_17504,N_17287,N_17282);
or U17505 (N_17505,N_17420,N_17309);
or U17506 (N_17506,N_17415,N_17284);
nor U17507 (N_17507,N_17333,N_17433);
xor U17508 (N_17508,N_17302,N_17404);
xor U17509 (N_17509,N_17385,N_17427);
or U17510 (N_17510,N_17328,N_17366);
and U17511 (N_17511,N_17324,N_17414);
and U17512 (N_17512,N_17310,N_17365);
nor U17513 (N_17513,N_17392,N_17364);
xnor U17514 (N_17514,N_17306,N_17431);
xnor U17515 (N_17515,N_17396,N_17313);
xor U17516 (N_17516,N_17307,N_17294);
nand U17517 (N_17517,N_17339,N_17361);
nor U17518 (N_17518,N_17322,N_17343);
and U17519 (N_17519,N_17419,N_17355);
or U17520 (N_17520,N_17435,N_17414);
and U17521 (N_17521,N_17344,N_17374);
and U17522 (N_17522,N_17290,N_17327);
nand U17523 (N_17523,N_17350,N_17308);
nand U17524 (N_17524,N_17339,N_17300);
xnor U17525 (N_17525,N_17329,N_17437);
and U17526 (N_17526,N_17292,N_17404);
and U17527 (N_17527,N_17429,N_17380);
nand U17528 (N_17528,N_17353,N_17348);
or U17529 (N_17529,N_17406,N_17404);
nor U17530 (N_17530,N_17336,N_17432);
nor U17531 (N_17531,N_17317,N_17385);
xnor U17532 (N_17532,N_17406,N_17412);
nand U17533 (N_17533,N_17301,N_17377);
xor U17534 (N_17534,N_17430,N_17351);
xor U17535 (N_17535,N_17368,N_17347);
and U17536 (N_17536,N_17366,N_17290);
nand U17537 (N_17537,N_17346,N_17329);
nor U17538 (N_17538,N_17322,N_17375);
or U17539 (N_17539,N_17411,N_17396);
nor U17540 (N_17540,N_17337,N_17395);
or U17541 (N_17541,N_17371,N_17401);
and U17542 (N_17542,N_17392,N_17399);
and U17543 (N_17543,N_17313,N_17364);
nand U17544 (N_17544,N_17426,N_17303);
nand U17545 (N_17545,N_17422,N_17351);
xnor U17546 (N_17546,N_17354,N_17403);
or U17547 (N_17547,N_17401,N_17336);
nor U17548 (N_17548,N_17433,N_17298);
nor U17549 (N_17549,N_17357,N_17305);
nor U17550 (N_17550,N_17371,N_17368);
and U17551 (N_17551,N_17424,N_17352);
nor U17552 (N_17552,N_17422,N_17346);
and U17553 (N_17553,N_17374,N_17354);
or U17554 (N_17554,N_17376,N_17402);
xor U17555 (N_17555,N_17377,N_17420);
nor U17556 (N_17556,N_17390,N_17339);
and U17557 (N_17557,N_17361,N_17420);
nor U17558 (N_17558,N_17376,N_17318);
xor U17559 (N_17559,N_17291,N_17360);
nor U17560 (N_17560,N_17419,N_17303);
or U17561 (N_17561,N_17360,N_17345);
and U17562 (N_17562,N_17308,N_17299);
nand U17563 (N_17563,N_17286,N_17422);
nand U17564 (N_17564,N_17432,N_17385);
nor U17565 (N_17565,N_17435,N_17339);
or U17566 (N_17566,N_17362,N_17354);
or U17567 (N_17567,N_17313,N_17333);
or U17568 (N_17568,N_17426,N_17348);
xnor U17569 (N_17569,N_17410,N_17340);
nand U17570 (N_17570,N_17356,N_17326);
nor U17571 (N_17571,N_17400,N_17295);
nand U17572 (N_17572,N_17365,N_17388);
or U17573 (N_17573,N_17290,N_17293);
xor U17574 (N_17574,N_17287,N_17315);
and U17575 (N_17575,N_17373,N_17288);
xor U17576 (N_17576,N_17319,N_17420);
or U17577 (N_17577,N_17342,N_17282);
xnor U17578 (N_17578,N_17405,N_17384);
or U17579 (N_17579,N_17439,N_17417);
or U17580 (N_17580,N_17433,N_17299);
xor U17581 (N_17581,N_17431,N_17285);
or U17582 (N_17582,N_17290,N_17320);
nor U17583 (N_17583,N_17436,N_17326);
and U17584 (N_17584,N_17394,N_17397);
and U17585 (N_17585,N_17438,N_17362);
and U17586 (N_17586,N_17339,N_17353);
nand U17587 (N_17587,N_17404,N_17331);
and U17588 (N_17588,N_17402,N_17396);
nor U17589 (N_17589,N_17355,N_17424);
or U17590 (N_17590,N_17305,N_17316);
nor U17591 (N_17591,N_17296,N_17345);
xor U17592 (N_17592,N_17310,N_17313);
nand U17593 (N_17593,N_17342,N_17413);
or U17594 (N_17594,N_17395,N_17306);
nor U17595 (N_17595,N_17312,N_17340);
or U17596 (N_17596,N_17399,N_17340);
nor U17597 (N_17597,N_17422,N_17393);
nand U17598 (N_17598,N_17410,N_17345);
nand U17599 (N_17599,N_17392,N_17318);
nor U17600 (N_17600,N_17572,N_17502);
and U17601 (N_17601,N_17577,N_17472);
xor U17602 (N_17602,N_17445,N_17529);
or U17603 (N_17603,N_17453,N_17480);
nand U17604 (N_17604,N_17581,N_17525);
or U17605 (N_17605,N_17508,N_17509);
and U17606 (N_17606,N_17542,N_17588);
nand U17607 (N_17607,N_17555,N_17573);
or U17608 (N_17608,N_17452,N_17496);
nor U17609 (N_17609,N_17544,N_17597);
or U17610 (N_17610,N_17457,N_17510);
xor U17611 (N_17611,N_17536,N_17540);
and U17612 (N_17612,N_17578,N_17467);
nand U17613 (N_17613,N_17460,N_17517);
nor U17614 (N_17614,N_17596,N_17538);
nor U17615 (N_17615,N_17490,N_17575);
nand U17616 (N_17616,N_17507,N_17491);
and U17617 (N_17617,N_17527,N_17455);
nor U17618 (N_17618,N_17591,N_17478);
and U17619 (N_17619,N_17474,N_17513);
xor U17620 (N_17620,N_17493,N_17459);
or U17621 (N_17621,N_17488,N_17515);
nor U17622 (N_17622,N_17458,N_17442);
or U17623 (N_17623,N_17470,N_17454);
nand U17624 (N_17624,N_17516,N_17558);
or U17625 (N_17625,N_17504,N_17528);
xor U17626 (N_17626,N_17522,N_17567);
xnor U17627 (N_17627,N_17543,N_17506);
and U17628 (N_17628,N_17585,N_17565);
nand U17629 (N_17629,N_17589,N_17551);
xnor U17630 (N_17630,N_17500,N_17594);
and U17631 (N_17631,N_17449,N_17448);
and U17632 (N_17632,N_17590,N_17479);
xnor U17633 (N_17633,N_17463,N_17599);
xor U17634 (N_17634,N_17560,N_17440);
nor U17635 (N_17635,N_17566,N_17532);
xnor U17636 (N_17636,N_17571,N_17563);
nor U17637 (N_17637,N_17530,N_17446);
xor U17638 (N_17638,N_17557,N_17464);
nand U17639 (N_17639,N_17546,N_17564);
nor U17640 (N_17640,N_17511,N_17524);
xor U17641 (N_17641,N_17518,N_17537);
and U17642 (N_17642,N_17486,N_17451);
xor U17643 (N_17643,N_17444,N_17497);
nor U17644 (N_17644,N_17568,N_17547);
nand U17645 (N_17645,N_17576,N_17570);
and U17646 (N_17646,N_17554,N_17450);
and U17647 (N_17647,N_17512,N_17489);
nor U17648 (N_17648,N_17461,N_17531);
or U17649 (N_17649,N_17443,N_17465);
xor U17650 (N_17650,N_17477,N_17521);
xor U17651 (N_17651,N_17494,N_17476);
xor U17652 (N_17652,N_17447,N_17485);
or U17653 (N_17653,N_17535,N_17498);
nor U17654 (N_17654,N_17481,N_17556);
nor U17655 (N_17655,N_17505,N_17492);
and U17656 (N_17656,N_17559,N_17482);
nor U17657 (N_17657,N_17523,N_17595);
xnor U17658 (N_17658,N_17514,N_17562);
nand U17659 (N_17659,N_17548,N_17499);
or U17660 (N_17660,N_17471,N_17533);
nor U17661 (N_17661,N_17469,N_17466);
nand U17662 (N_17662,N_17520,N_17441);
or U17663 (N_17663,N_17501,N_17593);
and U17664 (N_17664,N_17462,N_17468);
xnor U17665 (N_17665,N_17519,N_17586);
and U17666 (N_17666,N_17553,N_17545);
xor U17667 (N_17667,N_17574,N_17475);
or U17668 (N_17668,N_17583,N_17483);
nand U17669 (N_17669,N_17487,N_17473);
and U17670 (N_17670,N_17456,N_17539);
xor U17671 (N_17671,N_17541,N_17561);
nand U17672 (N_17672,N_17569,N_17584);
nand U17673 (N_17673,N_17579,N_17552);
nand U17674 (N_17674,N_17587,N_17592);
nand U17675 (N_17675,N_17550,N_17582);
nand U17676 (N_17676,N_17580,N_17526);
or U17677 (N_17677,N_17484,N_17503);
xnor U17678 (N_17678,N_17598,N_17534);
and U17679 (N_17679,N_17549,N_17495);
xor U17680 (N_17680,N_17542,N_17549);
or U17681 (N_17681,N_17569,N_17538);
nor U17682 (N_17682,N_17574,N_17454);
and U17683 (N_17683,N_17480,N_17476);
nand U17684 (N_17684,N_17441,N_17575);
nor U17685 (N_17685,N_17541,N_17553);
nor U17686 (N_17686,N_17578,N_17470);
nand U17687 (N_17687,N_17478,N_17473);
and U17688 (N_17688,N_17450,N_17474);
xor U17689 (N_17689,N_17448,N_17557);
and U17690 (N_17690,N_17519,N_17485);
xor U17691 (N_17691,N_17471,N_17538);
and U17692 (N_17692,N_17529,N_17480);
and U17693 (N_17693,N_17467,N_17552);
xor U17694 (N_17694,N_17559,N_17537);
nand U17695 (N_17695,N_17567,N_17549);
or U17696 (N_17696,N_17510,N_17596);
and U17697 (N_17697,N_17595,N_17561);
or U17698 (N_17698,N_17568,N_17577);
xnor U17699 (N_17699,N_17452,N_17442);
or U17700 (N_17700,N_17535,N_17509);
xor U17701 (N_17701,N_17570,N_17516);
nor U17702 (N_17702,N_17452,N_17475);
and U17703 (N_17703,N_17463,N_17536);
xor U17704 (N_17704,N_17509,N_17555);
xnor U17705 (N_17705,N_17529,N_17582);
nor U17706 (N_17706,N_17564,N_17453);
xnor U17707 (N_17707,N_17454,N_17598);
or U17708 (N_17708,N_17499,N_17457);
nor U17709 (N_17709,N_17590,N_17531);
nor U17710 (N_17710,N_17503,N_17580);
xnor U17711 (N_17711,N_17593,N_17503);
nand U17712 (N_17712,N_17481,N_17533);
nor U17713 (N_17713,N_17540,N_17488);
or U17714 (N_17714,N_17492,N_17525);
or U17715 (N_17715,N_17487,N_17579);
nand U17716 (N_17716,N_17499,N_17547);
nor U17717 (N_17717,N_17481,N_17518);
xnor U17718 (N_17718,N_17483,N_17524);
and U17719 (N_17719,N_17571,N_17539);
xor U17720 (N_17720,N_17524,N_17486);
xor U17721 (N_17721,N_17480,N_17565);
xor U17722 (N_17722,N_17561,N_17523);
nand U17723 (N_17723,N_17487,N_17481);
and U17724 (N_17724,N_17530,N_17559);
nor U17725 (N_17725,N_17469,N_17579);
and U17726 (N_17726,N_17577,N_17518);
nand U17727 (N_17727,N_17479,N_17524);
or U17728 (N_17728,N_17447,N_17559);
and U17729 (N_17729,N_17524,N_17538);
or U17730 (N_17730,N_17483,N_17594);
or U17731 (N_17731,N_17537,N_17451);
and U17732 (N_17732,N_17469,N_17529);
nor U17733 (N_17733,N_17580,N_17449);
nor U17734 (N_17734,N_17540,N_17443);
xor U17735 (N_17735,N_17551,N_17563);
xor U17736 (N_17736,N_17481,N_17590);
nor U17737 (N_17737,N_17573,N_17506);
or U17738 (N_17738,N_17457,N_17462);
nor U17739 (N_17739,N_17493,N_17598);
xor U17740 (N_17740,N_17575,N_17487);
nor U17741 (N_17741,N_17598,N_17510);
or U17742 (N_17742,N_17446,N_17553);
nor U17743 (N_17743,N_17578,N_17456);
and U17744 (N_17744,N_17530,N_17570);
xnor U17745 (N_17745,N_17473,N_17559);
xnor U17746 (N_17746,N_17463,N_17469);
nor U17747 (N_17747,N_17567,N_17547);
nand U17748 (N_17748,N_17514,N_17579);
nor U17749 (N_17749,N_17484,N_17474);
xnor U17750 (N_17750,N_17526,N_17532);
nand U17751 (N_17751,N_17444,N_17454);
xor U17752 (N_17752,N_17493,N_17478);
xnor U17753 (N_17753,N_17571,N_17503);
or U17754 (N_17754,N_17445,N_17584);
xor U17755 (N_17755,N_17539,N_17560);
nand U17756 (N_17756,N_17570,N_17441);
nand U17757 (N_17757,N_17511,N_17510);
nor U17758 (N_17758,N_17570,N_17460);
xor U17759 (N_17759,N_17473,N_17445);
xor U17760 (N_17760,N_17719,N_17604);
or U17761 (N_17761,N_17702,N_17676);
nand U17762 (N_17762,N_17696,N_17661);
xor U17763 (N_17763,N_17623,N_17669);
and U17764 (N_17764,N_17624,N_17641);
and U17765 (N_17765,N_17745,N_17618);
xnor U17766 (N_17766,N_17734,N_17673);
nor U17767 (N_17767,N_17628,N_17667);
and U17768 (N_17768,N_17698,N_17680);
nor U17769 (N_17769,N_17655,N_17678);
nor U17770 (N_17770,N_17755,N_17674);
nand U17771 (N_17771,N_17621,N_17646);
xnor U17772 (N_17772,N_17640,N_17751);
or U17773 (N_17773,N_17607,N_17701);
xor U17774 (N_17774,N_17620,N_17649);
nor U17775 (N_17775,N_17718,N_17602);
or U17776 (N_17776,N_17601,N_17697);
xor U17777 (N_17777,N_17611,N_17738);
or U17778 (N_17778,N_17730,N_17662);
nor U17779 (N_17779,N_17677,N_17672);
and U17780 (N_17780,N_17693,N_17668);
xor U17781 (N_17781,N_17622,N_17748);
and U17782 (N_17782,N_17631,N_17694);
or U17783 (N_17783,N_17685,N_17713);
nor U17784 (N_17784,N_17653,N_17758);
or U17785 (N_17785,N_17705,N_17615);
or U17786 (N_17786,N_17651,N_17639);
xnor U17787 (N_17787,N_17675,N_17626);
xor U17788 (N_17788,N_17741,N_17715);
nor U17789 (N_17789,N_17629,N_17689);
nor U17790 (N_17790,N_17703,N_17635);
xnor U17791 (N_17791,N_17744,N_17603);
xnor U17792 (N_17792,N_17728,N_17656);
xnor U17793 (N_17793,N_17636,N_17643);
nor U17794 (N_17794,N_17746,N_17700);
nand U17795 (N_17795,N_17756,N_17743);
nand U17796 (N_17796,N_17707,N_17690);
nor U17797 (N_17797,N_17658,N_17613);
or U17798 (N_17798,N_17616,N_17752);
nor U17799 (N_17799,N_17648,N_17633);
nand U17800 (N_17800,N_17609,N_17660);
nor U17801 (N_17801,N_17654,N_17722);
nand U17802 (N_17802,N_17724,N_17638);
and U17803 (N_17803,N_17731,N_17757);
and U17804 (N_17804,N_17632,N_17606);
or U17805 (N_17805,N_17735,N_17681);
xor U17806 (N_17806,N_17671,N_17686);
nand U17807 (N_17807,N_17650,N_17617);
xor U17808 (N_17808,N_17727,N_17634);
nand U17809 (N_17809,N_17706,N_17747);
nand U17810 (N_17810,N_17692,N_17647);
nor U17811 (N_17811,N_17625,N_17630);
xor U17812 (N_17812,N_17708,N_17659);
nand U17813 (N_17813,N_17753,N_17600);
or U17814 (N_17814,N_17726,N_17644);
nand U17815 (N_17815,N_17704,N_17712);
xnor U17816 (N_17816,N_17645,N_17714);
xnor U17817 (N_17817,N_17666,N_17736);
nand U17818 (N_17818,N_17683,N_17754);
xnor U17819 (N_17819,N_17688,N_17740);
xnor U17820 (N_17820,N_17614,N_17642);
or U17821 (N_17821,N_17652,N_17721);
or U17822 (N_17822,N_17716,N_17657);
and U17823 (N_17823,N_17739,N_17663);
nor U17824 (N_17824,N_17695,N_17750);
nor U17825 (N_17825,N_17709,N_17749);
xor U17826 (N_17826,N_17717,N_17665);
nand U17827 (N_17827,N_17733,N_17737);
and U17828 (N_17828,N_17619,N_17742);
nor U17829 (N_17829,N_17691,N_17605);
nand U17830 (N_17830,N_17610,N_17608);
or U17831 (N_17831,N_17612,N_17679);
xnor U17832 (N_17832,N_17637,N_17627);
xor U17833 (N_17833,N_17699,N_17759);
nor U17834 (N_17834,N_17720,N_17729);
nand U17835 (N_17835,N_17711,N_17725);
nor U17836 (N_17836,N_17710,N_17684);
nor U17837 (N_17837,N_17723,N_17670);
or U17838 (N_17838,N_17732,N_17682);
and U17839 (N_17839,N_17687,N_17664);
and U17840 (N_17840,N_17738,N_17731);
and U17841 (N_17841,N_17721,N_17719);
and U17842 (N_17842,N_17707,N_17600);
or U17843 (N_17843,N_17758,N_17685);
and U17844 (N_17844,N_17756,N_17723);
or U17845 (N_17845,N_17678,N_17696);
or U17846 (N_17846,N_17671,N_17657);
and U17847 (N_17847,N_17684,N_17656);
xor U17848 (N_17848,N_17673,N_17606);
and U17849 (N_17849,N_17652,N_17720);
and U17850 (N_17850,N_17640,N_17629);
and U17851 (N_17851,N_17690,N_17703);
xor U17852 (N_17852,N_17758,N_17661);
and U17853 (N_17853,N_17701,N_17703);
nand U17854 (N_17854,N_17622,N_17712);
and U17855 (N_17855,N_17627,N_17663);
xnor U17856 (N_17856,N_17667,N_17646);
nor U17857 (N_17857,N_17620,N_17701);
or U17858 (N_17858,N_17675,N_17678);
and U17859 (N_17859,N_17618,N_17703);
nand U17860 (N_17860,N_17686,N_17730);
nand U17861 (N_17861,N_17603,N_17683);
nand U17862 (N_17862,N_17608,N_17697);
xor U17863 (N_17863,N_17660,N_17622);
xor U17864 (N_17864,N_17622,N_17676);
nor U17865 (N_17865,N_17617,N_17713);
xor U17866 (N_17866,N_17601,N_17734);
nand U17867 (N_17867,N_17631,N_17685);
and U17868 (N_17868,N_17667,N_17714);
nand U17869 (N_17869,N_17720,N_17653);
or U17870 (N_17870,N_17738,N_17756);
nor U17871 (N_17871,N_17749,N_17706);
nor U17872 (N_17872,N_17737,N_17699);
nand U17873 (N_17873,N_17759,N_17618);
and U17874 (N_17874,N_17621,N_17693);
xnor U17875 (N_17875,N_17625,N_17704);
or U17876 (N_17876,N_17624,N_17630);
nand U17877 (N_17877,N_17652,N_17682);
or U17878 (N_17878,N_17652,N_17710);
or U17879 (N_17879,N_17732,N_17621);
nor U17880 (N_17880,N_17628,N_17686);
nand U17881 (N_17881,N_17657,N_17746);
or U17882 (N_17882,N_17615,N_17748);
nand U17883 (N_17883,N_17702,N_17656);
nor U17884 (N_17884,N_17679,N_17725);
and U17885 (N_17885,N_17663,N_17632);
nand U17886 (N_17886,N_17700,N_17712);
nor U17887 (N_17887,N_17689,N_17697);
or U17888 (N_17888,N_17661,N_17606);
and U17889 (N_17889,N_17673,N_17749);
xnor U17890 (N_17890,N_17759,N_17747);
nor U17891 (N_17891,N_17717,N_17603);
or U17892 (N_17892,N_17653,N_17724);
xnor U17893 (N_17893,N_17658,N_17708);
and U17894 (N_17894,N_17715,N_17600);
nand U17895 (N_17895,N_17716,N_17666);
and U17896 (N_17896,N_17679,N_17672);
xnor U17897 (N_17897,N_17644,N_17623);
nor U17898 (N_17898,N_17637,N_17744);
or U17899 (N_17899,N_17667,N_17606);
or U17900 (N_17900,N_17623,N_17671);
xnor U17901 (N_17901,N_17735,N_17632);
xnor U17902 (N_17902,N_17744,N_17606);
nand U17903 (N_17903,N_17747,N_17623);
and U17904 (N_17904,N_17666,N_17705);
xor U17905 (N_17905,N_17751,N_17710);
nor U17906 (N_17906,N_17749,N_17711);
and U17907 (N_17907,N_17642,N_17669);
and U17908 (N_17908,N_17692,N_17678);
and U17909 (N_17909,N_17714,N_17753);
and U17910 (N_17910,N_17675,N_17663);
nor U17911 (N_17911,N_17736,N_17724);
nand U17912 (N_17912,N_17699,N_17669);
or U17913 (N_17913,N_17712,N_17648);
xor U17914 (N_17914,N_17715,N_17703);
and U17915 (N_17915,N_17651,N_17655);
and U17916 (N_17916,N_17751,N_17753);
nor U17917 (N_17917,N_17676,N_17726);
or U17918 (N_17918,N_17616,N_17715);
or U17919 (N_17919,N_17604,N_17651);
xnor U17920 (N_17920,N_17914,N_17776);
or U17921 (N_17921,N_17867,N_17772);
or U17922 (N_17922,N_17899,N_17805);
and U17923 (N_17923,N_17795,N_17840);
and U17924 (N_17924,N_17808,N_17855);
and U17925 (N_17925,N_17880,N_17900);
xor U17926 (N_17926,N_17858,N_17768);
nand U17927 (N_17927,N_17910,N_17783);
nand U17928 (N_17928,N_17796,N_17777);
xnor U17929 (N_17929,N_17835,N_17807);
nor U17930 (N_17930,N_17890,N_17761);
nand U17931 (N_17931,N_17903,N_17888);
and U17932 (N_17932,N_17820,N_17852);
xor U17933 (N_17933,N_17764,N_17894);
nor U17934 (N_17934,N_17862,N_17865);
nand U17935 (N_17935,N_17819,N_17875);
xnor U17936 (N_17936,N_17773,N_17872);
or U17937 (N_17937,N_17789,N_17871);
nor U17938 (N_17938,N_17901,N_17848);
nor U17939 (N_17939,N_17834,N_17780);
nor U17940 (N_17940,N_17821,N_17895);
and U17941 (N_17941,N_17787,N_17916);
nand U17942 (N_17942,N_17866,N_17778);
and U17943 (N_17943,N_17896,N_17849);
xnor U17944 (N_17944,N_17817,N_17878);
or U17945 (N_17945,N_17803,N_17830);
and U17946 (N_17946,N_17767,N_17881);
and U17947 (N_17947,N_17831,N_17909);
and U17948 (N_17948,N_17873,N_17863);
nor U17949 (N_17949,N_17814,N_17763);
nand U17950 (N_17950,N_17799,N_17847);
xnor U17951 (N_17951,N_17824,N_17774);
and U17952 (N_17952,N_17775,N_17887);
xor U17953 (N_17953,N_17892,N_17845);
xor U17954 (N_17954,N_17846,N_17853);
or U17955 (N_17955,N_17809,N_17859);
or U17956 (N_17956,N_17785,N_17870);
xnor U17957 (N_17957,N_17826,N_17850);
nor U17958 (N_17958,N_17802,N_17765);
xor U17959 (N_17959,N_17917,N_17829);
nor U17960 (N_17960,N_17770,N_17883);
and U17961 (N_17961,N_17898,N_17836);
xnor U17962 (N_17962,N_17915,N_17891);
nor U17963 (N_17963,N_17860,N_17794);
nor U17964 (N_17964,N_17893,N_17804);
or U17965 (N_17965,N_17879,N_17864);
nor U17966 (N_17966,N_17885,N_17791);
xor U17967 (N_17967,N_17912,N_17902);
nand U17968 (N_17968,N_17919,N_17818);
xor U17969 (N_17969,N_17877,N_17766);
nand U17970 (N_17970,N_17854,N_17868);
and U17971 (N_17971,N_17813,N_17907);
and U17972 (N_17972,N_17806,N_17779);
and U17973 (N_17973,N_17843,N_17838);
nor U17974 (N_17974,N_17913,N_17839);
or U17975 (N_17975,N_17889,N_17832);
or U17976 (N_17976,N_17801,N_17797);
xor U17977 (N_17977,N_17786,N_17788);
xor U17978 (N_17978,N_17897,N_17781);
xor U17979 (N_17979,N_17822,N_17782);
and U17980 (N_17980,N_17884,N_17790);
and U17981 (N_17981,N_17861,N_17810);
or U17982 (N_17982,N_17816,N_17825);
and U17983 (N_17983,N_17911,N_17771);
and U17984 (N_17984,N_17833,N_17857);
and U17985 (N_17985,N_17841,N_17869);
or U17986 (N_17986,N_17798,N_17874);
nor U17987 (N_17987,N_17828,N_17918);
nand U17988 (N_17988,N_17823,N_17886);
or U17989 (N_17989,N_17760,N_17792);
nor U17990 (N_17990,N_17851,N_17815);
or U17991 (N_17991,N_17856,N_17812);
xor U17992 (N_17992,N_17837,N_17827);
nor U17993 (N_17993,N_17844,N_17906);
and U17994 (N_17994,N_17905,N_17762);
xnor U17995 (N_17995,N_17908,N_17811);
or U17996 (N_17996,N_17800,N_17793);
xor U17997 (N_17997,N_17876,N_17904);
nand U17998 (N_17998,N_17769,N_17784);
nor U17999 (N_17999,N_17882,N_17842);
xnor U18000 (N_18000,N_17908,N_17871);
or U18001 (N_18001,N_17840,N_17766);
or U18002 (N_18002,N_17860,N_17829);
xnor U18003 (N_18003,N_17798,N_17915);
nand U18004 (N_18004,N_17829,N_17767);
and U18005 (N_18005,N_17805,N_17813);
nor U18006 (N_18006,N_17833,N_17822);
nand U18007 (N_18007,N_17904,N_17771);
or U18008 (N_18008,N_17761,N_17885);
nor U18009 (N_18009,N_17910,N_17851);
nand U18010 (N_18010,N_17901,N_17809);
or U18011 (N_18011,N_17898,N_17880);
nor U18012 (N_18012,N_17776,N_17768);
nor U18013 (N_18013,N_17833,N_17878);
or U18014 (N_18014,N_17822,N_17872);
nor U18015 (N_18015,N_17786,N_17912);
nand U18016 (N_18016,N_17866,N_17769);
xor U18017 (N_18017,N_17798,N_17863);
nand U18018 (N_18018,N_17851,N_17797);
nor U18019 (N_18019,N_17795,N_17780);
nor U18020 (N_18020,N_17831,N_17762);
and U18021 (N_18021,N_17888,N_17883);
nor U18022 (N_18022,N_17911,N_17823);
xnor U18023 (N_18023,N_17887,N_17815);
nand U18024 (N_18024,N_17810,N_17839);
nand U18025 (N_18025,N_17816,N_17789);
or U18026 (N_18026,N_17885,N_17845);
and U18027 (N_18027,N_17894,N_17774);
nand U18028 (N_18028,N_17856,N_17889);
and U18029 (N_18029,N_17867,N_17761);
nand U18030 (N_18030,N_17829,N_17814);
and U18031 (N_18031,N_17851,N_17911);
nor U18032 (N_18032,N_17818,N_17852);
nand U18033 (N_18033,N_17907,N_17816);
nand U18034 (N_18034,N_17828,N_17807);
nand U18035 (N_18035,N_17779,N_17902);
or U18036 (N_18036,N_17867,N_17833);
xor U18037 (N_18037,N_17821,N_17860);
xnor U18038 (N_18038,N_17820,N_17850);
xnor U18039 (N_18039,N_17833,N_17792);
nand U18040 (N_18040,N_17812,N_17810);
nand U18041 (N_18041,N_17839,N_17773);
nor U18042 (N_18042,N_17833,N_17858);
xnor U18043 (N_18043,N_17761,N_17806);
and U18044 (N_18044,N_17854,N_17875);
xor U18045 (N_18045,N_17873,N_17821);
and U18046 (N_18046,N_17822,N_17873);
xor U18047 (N_18047,N_17794,N_17897);
xor U18048 (N_18048,N_17841,N_17804);
xor U18049 (N_18049,N_17851,N_17885);
nand U18050 (N_18050,N_17807,N_17862);
xor U18051 (N_18051,N_17797,N_17909);
and U18052 (N_18052,N_17822,N_17763);
or U18053 (N_18053,N_17764,N_17830);
nor U18054 (N_18054,N_17904,N_17761);
or U18055 (N_18055,N_17790,N_17842);
xnor U18056 (N_18056,N_17790,N_17828);
and U18057 (N_18057,N_17911,N_17901);
nand U18058 (N_18058,N_17769,N_17805);
or U18059 (N_18059,N_17771,N_17798);
nand U18060 (N_18060,N_17825,N_17840);
nand U18061 (N_18061,N_17789,N_17895);
and U18062 (N_18062,N_17828,N_17765);
nor U18063 (N_18063,N_17896,N_17780);
nor U18064 (N_18064,N_17873,N_17772);
and U18065 (N_18065,N_17835,N_17776);
and U18066 (N_18066,N_17767,N_17868);
or U18067 (N_18067,N_17809,N_17788);
nand U18068 (N_18068,N_17877,N_17776);
and U18069 (N_18069,N_17839,N_17797);
nor U18070 (N_18070,N_17896,N_17769);
nor U18071 (N_18071,N_17839,N_17915);
and U18072 (N_18072,N_17881,N_17783);
nor U18073 (N_18073,N_17905,N_17801);
nor U18074 (N_18074,N_17783,N_17816);
and U18075 (N_18075,N_17813,N_17895);
or U18076 (N_18076,N_17798,N_17866);
and U18077 (N_18077,N_17825,N_17823);
and U18078 (N_18078,N_17909,N_17815);
or U18079 (N_18079,N_17919,N_17779);
nor U18080 (N_18080,N_17958,N_18012);
nor U18081 (N_18081,N_18025,N_18003);
and U18082 (N_18082,N_18058,N_18021);
xnor U18083 (N_18083,N_17946,N_18076);
nor U18084 (N_18084,N_17985,N_18020);
xnor U18085 (N_18085,N_17997,N_17967);
or U18086 (N_18086,N_17936,N_17925);
or U18087 (N_18087,N_17930,N_17952);
nor U18088 (N_18088,N_18030,N_17949);
and U18089 (N_18089,N_18029,N_17940);
nand U18090 (N_18090,N_18049,N_18052);
nand U18091 (N_18091,N_18041,N_17968);
nand U18092 (N_18092,N_18018,N_17923);
or U18093 (N_18093,N_18002,N_17992);
and U18094 (N_18094,N_17947,N_18038);
and U18095 (N_18095,N_17957,N_17933);
xor U18096 (N_18096,N_18053,N_17945);
nor U18097 (N_18097,N_17970,N_18051);
and U18098 (N_18098,N_17964,N_17963);
and U18099 (N_18099,N_18063,N_18036);
and U18100 (N_18100,N_17995,N_18026);
or U18101 (N_18101,N_17960,N_18023);
xor U18102 (N_18102,N_18048,N_18060);
nor U18103 (N_18103,N_18014,N_18004);
xor U18104 (N_18104,N_18019,N_17984);
nor U18105 (N_18105,N_17969,N_18042);
xnor U18106 (N_18106,N_18079,N_17961);
nor U18107 (N_18107,N_17932,N_18006);
nand U18108 (N_18108,N_18070,N_18069);
or U18109 (N_18109,N_18043,N_18062);
nor U18110 (N_18110,N_18039,N_17924);
nor U18111 (N_18111,N_18075,N_17935);
and U18112 (N_18112,N_18037,N_17953);
xnor U18113 (N_18113,N_17966,N_17942);
nand U18114 (N_18114,N_18068,N_17978);
nor U18115 (N_18115,N_17980,N_17929);
nand U18116 (N_18116,N_17938,N_17962);
nand U18117 (N_18117,N_18010,N_18045);
nand U18118 (N_18118,N_17937,N_18000);
nor U18119 (N_18119,N_18040,N_18007);
nor U18120 (N_18120,N_18071,N_18054);
nand U18121 (N_18121,N_18044,N_17979);
or U18122 (N_18122,N_17921,N_17993);
nand U18123 (N_18123,N_17926,N_18047);
and U18124 (N_18124,N_18032,N_18066);
nand U18125 (N_18125,N_17934,N_18067);
nand U18126 (N_18126,N_17941,N_17955);
and U18127 (N_18127,N_17971,N_18055);
or U18128 (N_18128,N_18024,N_18001);
xor U18129 (N_18129,N_17983,N_18064);
nand U18130 (N_18130,N_17999,N_18017);
and U18131 (N_18131,N_17986,N_17928);
and U18132 (N_18132,N_17972,N_18008);
or U18133 (N_18133,N_17991,N_18016);
nor U18134 (N_18134,N_18013,N_18035);
and U18135 (N_18135,N_18065,N_18074);
xor U18136 (N_18136,N_17944,N_18072);
nand U18137 (N_18137,N_17975,N_18050);
xor U18138 (N_18138,N_17954,N_17927);
xor U18139 (N_18139,N_17951,N_18027);
xnor U18140 (N_18140,N_18061,N_18073);
nand U18141 (N_18141,N_17982,N_17998);
and U18142 (N_18142,N_18028,N_18057);
nor U18143 (N_18143,N_17981,N_17931);
nor U18144 (N_18144,N_17987,N_18078);
and U18145 (N_18145,N_17922,N_17920);
and U18146 (N_18146,N_18009,N_17989);
or U18147 (N_18147,N_18015,N_17994);
or U18148 (N_18148,N_18022,N_18059);
or U18149 (N_18149,N_17948,N_17988);
nor U18150 (N_18150,N_18056,N_17965);
nand U18151 (N_18151,N_17943,N_18011);
or U18152 (N_18152,N_18046,N_17974);
or U18153 (N_18153,N_18005,N_17959);
nor U18154 (N_18154,N_18033,N_18031);
nand U18155 (N_18155,N_17990,N_17956);
xnor U18156 (N_18156,N_17939,N_18034);
or U18157 (N_18157,N_17950,N_18077);
xnor U18158 (N_18158,N_17976,N_17996);
nor U18159 (N_18159,N_17973,N_17977);
and U18160 (N_18160,N_17955,N_18048);
xnor U18161 (N_18161,N_17968,N_18016);
xnor U18162 (N_18162,N_18064,N_18001);
xor U18163 (N_18163,N_17998,N_18035);
and U18164 (N_18164,N_17974,N_17997);
and U18165 (N_18165,N_17943,N_18061);
nor U18166 (N_18166,N_18078,N_18066);
and U18167 (N_18167,N_17958,N_18070);
or U18168 (N_18168,N_17956,N_17936);
or U18169 (N_18169,N_17971,N_18063);
or U18170 (N_18170,N_17986,N_18066);
xnor U18171 (N_18171,N_17946,N_18025);
nand U18172 (N_18172,N_17991,N_17978);
and U18173 (N_18173,N_17934,N_17941);
xnor U18174 (N_18174,N_18066,N_18025);
or U18175 (N_18175,N_17950,N_18065);
nand U18176 (N_18176,N_18043,N_17959);
nand U18177 (N_18177,N_18023,N_17981);
or U18178 (N_18178,N_18039,N_17999);
nor U18179 (N_18179,N_17994,N_18058);
xnor U18180 (N_18180,N_18007,N_18035);
and U18181 (N_18181,N_18046,N_17940);
or U18182 (N_18182,N_17937,N_18037);
nor U18183 (N_18183,N_17979,N_17935);
and U18184 (N_18184,N_18007,N_18032);
and U18185 (N_18185,N_17933,N_17977);
xor U18186 (N_18186,N_18072,N_18027);
xnor U18187 (N_18187,N_18009,N_17935);
nor U18188 (N_18188,N_17949,N_17955);
and U18189 (N_18189,N_18019,N_17995);
xor U18190 (N_18190,N_17992,N_17952);
and U18191 (N_18191,N_18007,N_18031);
or U18192 (N_18192,N_17931,N_18062);
nand U18193 (N_18193,N_17941,N_17995);
and U18194 (N_18194,N_18033,N_17942);
nor U18195 (N_18195,N_18031,N_17991);
nand U18196 (N_18196,N_18075,N_18040);
or U18197 (N_18197,N_18072,N_17942);
or U18198 (N_18198,N_17958,N_17989);
nand U18199 (N_18199,N_17922,N_18036);
nor U18200 (N_18200,N_18012,N_17976);
or U18201 (N_18201,N_18055,N_18035);
or U18202 (N_18202,N_18007,N_18074);
xor U18203 (N_18203,N_18006,N_17926);
xnor U18204 (N_18204,N_17924,N_17934);
nor U18205 (N_18205,N_17937,N_17957);
or U18206 (N_18206,N_18006,N_17935);
nand U18207 (N_18207,N_18059,N_17944);
nor U18208 (N_18208,N_17996,N_17998);
nor U18209 (N_18209,N_18006,N_17996);
xor U18210 (N_18210,N_17968,N_17999);
nand U18211 (N_18211,N_17964,N_17976);
xnor U18212 (N_18212,N_18008,N_17981);
nand U18213 (N_18213,N_17957,N_18072);
and U18214 (N_18214,N_18051,N_18039);
or U18215 (N_18215,N_17930,N_18078);
or U18216 (N_18216,N_17933,N_17943);
nor U18217 (N_18217,N_17964,N_17980);
and U18218 (N_18218,N_17994,N_18000);
or U18219 (N_18219,N_17976,N_17989);
xnor U18220 (N_18220,N_17926,N_18025);
nor U18221 (N_18221,N_17995,N_18033);
nor U18222 (N_18222,N_17945,N_17983);
nor U18223 (N_18223,N_17984,N_18067);
or U18224 (N_18224,N_17934,N_18058);
or U18225 (N_18225,N_17963,N_17943);
xnor U18226 (N_18226,N_18004,N_17992);
xor U18227 (N_18227,N_18007,N_18048);
nand U18228 (N_18228,N_17947,N_17982);
nand U18229 (N_18229,N_17937,N_18002);
nor U18230 (N_18230,N_17989,N_18020);
xor U18231 (N_18231,N_17972,N_18078);
xor U18232 (N_18232,N_18035,N_18008);
nand U18233 (N_18233,N_18044,N_18045);
and U18234 (N_18234,N_18075,N_18051);
nand U18235 (N_18235,N_18054,N_18010);
and U18236 (N_18236,N_17941,N_17952);
nand U18237 (N_18237,N_17957,N_17999);
xor U18238 (N_18238,N_18053,N_17999);
xnor U18239 (N_18239,N_17939,N_18012);
nand U18240 (N_18240,N_18163,N_18088);
nor U18241 (N_18241,N_18232,N_18092);
nand U18242 (N_18242,N_18168,N_18237);
xor U18243 (N_18243,N_18233,N_18124);
xnor U18244 (N_18244,N_18118,N_18089);
or U18245 (N_18245,N_18167,N_18186);
nand U18246 (N_18246,N_18132,N_18174);
nor U18247 (N_18247,N_18086,N_18109);
xnor U18248 (N_18248,N_18166,N_18111);
nor U18249 (N_18249,N_18221,N_18189);
nand U18250 (N_18250,N_18103,N_18145);
nor U18251 (N_18251,N_18129,N_18213);
nor U18252 (N_18252,N_18101,N_18217);
or U18253 (N_18253,N_18117,N_18087);
or U18254 (N_18254,N_18203,N_18164);
or U18255 (N_18255,N_18238,N_18114);
or U18256 (N_18256,N_18219,N_18106);
xnor U18257 (N_18257,N_18160,N_18119);
and U18258 (N_18258,N_18093,N_18141);
nor U18259 (N_18259,N_18094,N_18159);
nand U18260 (N_18260,N_18229,N_18150);
nor U18261 (N_18261,N_18140,N_18107);
nor U18262 (N_18262,N_18112,N_18157);
xnor U18263 (N_18263,N_18175,N_18134);
or U18264 (N_18264,N_18153,N_18155);
and U18265 (N_18265,N_18080,N_18161);
or U18266 (N_18266,N_18211,N_18130);
nor U18267 (N_18267,N_18196,N_18147);
and U18268 (N_18268,N_18225,N_18165);
or U18269 (N_18269,N_18183,N_18182);
nand U18270 (N_18270,N_18235,N_18181);
nand U18271 (N_18271,N_18122,N_18102);
or U18272 (N_18272,N_18091,N_18226);
nand U18273 (N_18273,N_18179,N_18202);
or U18274 (N_18274,N_18146,N_18172);
nand U18275 (N_18275,N_18144,N_18227);
nor U18276 (N_18276,N_18208,N_18131);
nor U18277 (N_18277,N_18192,N_18239);
nor U18278 (N_18278,N_18199,N_18082);
and U18279 (N_18279,N_18188,N_18123);
nor U18280 (N_18280,N_18204,N_18215);
or U18281 (N_18281,N_18162,N_18185);
nand U18282 (N_18282,N_18184,N_18095);
xor U18283 (N_18283,N_18170,N_18214);
nor U18284 (N_18284,N_18205,N_18126);
nand U18285 (N_18285,N_18152,N_18190);
nor U18286 (N_18286,N_18169,N_18154);
and U18287 (N_18287,N_18084,N_18137);
or U18288 (N_18288,N_18139,N_18231);
xnor U18289 (N_18289,N_18136,N_18135);
or U18290 (N_18290,N_18223,N_18197);
and U18291 (N_18291,N_18104,N_18187);
and U18292 (N_18292,N_18090,N_18220);
xor U18293 (N_18293,N_18120,N_18230);
xnor U18294 (N_18294,N_18236,N_18216);
and U18295 (N_18295,N_18178,N_18201);
xnor U18296 (N_18296,N_18206,N_18194);
and U18297 (N_18297,N_18171,N_18083);
nand U18298 (N_18298,N_18098,N_18099);
and U18299 (N_18299,N_18096,N_18097);
nor U18300 (N_18300,N_18200,N_18193);
nor U18301 (N_18301,N_18133,N_18151);
xnor U18302 (N_18302,N_18228,N_18212);
nor U18303 (N_18303,N_18156,N_18148);
nor U18304 (N_18304,N_18113,N_18100);
xnor U18305 (N_18305,N_18195,N_18085);
xnor U18306 (N_18306,N_18110,N_18149);
nand U18307 (N_18307,N_18108,N_18224);
nor U18308 (N_18308,N_18180,N_18218);
xnor U18309 (N_18309,N_18143,N_18198);
and U18310 (N_18310,N_18128,N_18191);
or U18311 (N_18311,N_18105,N_18173);
nand U18312 (N_18312,N_18210,N_18234);
nand U18313 (N_18313,N_18158,N_18125);
nor U18314 (N_18314,N_18116,N_18115);
and U18315 (N_18315,N_18207,N_18127);
nor U18316 (N_18316,N_18177,N_18081);
xor U18317 (N_18317,N_18138,N_18121);
or U18318 (N_18318,N_18142,N_18176);
xor U18319 (N_18319,N_18222,N_18209);
nor U18320 (N_18320,N_18171,N_18133);
nand U18321 (N_18321,N_18186,N_18088);
nand U18322 (N_18322,N_18199,N_18222);
xnor U18323 (N_18323,N_18177,N_18187);
nor U18324 (N_18324,N_18195,N_18082);
or U18325 (N_18325,N_18080,N_18136);
and U18326 (N_18326,N_18117,N_18198);
xor U18327 (N_18327,N_18087,N_18113);
or U18328 (N_18328,N_18223,N_18205);
and U18329 (N_18329,N_18149,N_18238);
nor U18330 (N_18330,N_18214,N_18144);
nand U18331 (N_18331,N_18140,N_18194);
and U18332 (N_18332,N_18167,N_18228);
and U18333 (N_18333,N_18235,N_18195);
nand U18334 (N_18334,N_18132,N_18109);
nor U18335 (N_18335,N_18101,N_18108);
xor U18336 (N_18336,N_18124,N_18119);
nor U18337 (N_18337,N_18147,N_18139);
or U18338 (N_18338,N_18140,N_18112);
nand U18339 (N_18339,N_18229,N_18224);
xnor U18340 (N_18340,N_18204,N_18097);
or U18341 (N_18341,N_18143,N_18189);
xor U18342 (N_18342,N_18092,N_18131);
nand U18343 (N_18343,N_18109,N_18177);
nor U18344 (N_18344,N_18115,N_18100);
nor U18345 (N_18345,N_18093,N_18201);
xnor U18346 (N_18346,N_18150,N_18202);
xnor U18347 (N_18347,N_18149,N_18128);
and U18348 (N_18348,N_18142,N_18229);
nor U18349 (N_18349,N_18187,N_18167);
and U18350 (N_18350,N_18092,N_18190);
and U18351 (N_18351,N_18113,N_18196);
nor U18352 (N_18352,N_18189,N_18099);
and U18353 (N_18353,N_18176,N_18098);
and U18354 (N_18354,N_18132,N_18093);
xor U18355 (N_18355,N_18135,N_18162);
nand U18356 (N_18356,N_18115,N_18090);
nand U18357 (N_18357,N_18218,N_18191);
nand U18358 (N_18358,N_18146,N_18137);
xor U18359 (N_18359,N_18131,N_18158);
nor U18360 (N_18360,N_18150,N_18110);
xor U18361 (N_18361,N_18164,N_18120);
nand U18362 (N_18362,N_18231,N_18239);
nor U18363 (N_18363,N_18186,N_18092);
and U18364 (N_18364,N_18125,N_18187);
xor U18365 (N_18365,N_18145,N_18099);
nand U18366 (N_18366,N_18152,N_18131);
or U18367 (N_18367,N_18172,N_18221);
or U18368 (N_18368,N_18095,N_18150);
nor U18369 (N_18369,N_18139,N_18190);
xor U18370 (N_18370,N_18114,N_18109);
nand U18371 (N_18371,N_18173,N_18186);
or U18372 (N_18372,N_18149,N_18232);
and U18373 (N_18373,N_18207,N_18189);
and U18374 (N_18374,N_18158,N_18093);
and U18375 (N_18375,N_18216,N_18104);
or U18376 (N_18376,N_18200,N_18223);
xor U18377 (N_18377,N_18126,N_18163);
nor U18378 (N_18378,N_18226,N_18155);
xor U18379 (N_18379,N_18161,N_18083);
xor U18380 (N_18380,N_18089,N_18100);
nand U18381 (N_18381,N_18108,N_18128);
nor U18382 (N_18382,N_18170,N_18229);
nor U18383 (N_18383,N_18094,N_18123);
nand U18384 (N_18384,N_18151,N_18142);
or U18385 (N_18385,N_18198,N_18235);
and U18386 (N_18386,N_18173,N_18089);
nor U18387 (N_18387,N_18123,N_18095);
and U18388 (N_18388,N_18231,N_18134);
and U18389 (N_18389,N_18222,N_18203);
and U18390 (N_18390,N_18189,N_18081);
and U18391 (N_18391,N_18170,N_18092);
nand U18392 (N_18392,N_18154,N_18147);
or U18393 (N_18393,N_18216,N_18169);
nand U18394 (N_18394,N_18203,N_18092);
nand U18395 (N_18395,N_18147,N_18138);
nor U18396 (N_18396,N_18139,N_18205);
nor U18397 (N_18397,N_18141,N_18132);
nand U18398 (N_18398,N_18170,N_18227);
nand U18399 (N_18399,N_18102,N_18094);
nand U18400 (N_18400,N_18342,N_18305);
or U18401 (N_18401,N_18343,N_18287);
nor U18402 (N_18402,N_18397,N_18340);
nand U18403 (N_18403,N_18244,N_18331);
and U18404 (N_18404,N_18281,N_18316);
nand U18405 (N_18405,N_18393,N_18285);
xnor U18406 (N_18406,N_18248,N_18251);
nand U18407 (N_18407,N_18260,N_18278);
and U18408 (N_18408,N_18346,N_18321);
or U18409 (N_18409,N_18280,N_18390);
or U18410 (N_18410,N_18338,N_18257);
or U18411 (N_18411,N_18362,N_18290);
nand U18412 (N_18412,N_18303,N_18368);
and U18413 (N_18413,N_18386,N_18242);
nand U18414 (N_18414,N_18322,N_18375);
xnor U18415 (N_18415,N_18376,N_18345);
and U18416 (N_18416,N_18330,N_18337);
nor U18417 (N_18417,N_18319,N_18279);
xor U18418 (N_18418,N_18306,N_18336);
nand U18419 (N_18419,N_18344,N_18275);
nand U18420 (N_18420,N_18364,N_18254);
or U18421 (N_18421,N_18387,N_18325);
xor U18422 (N_18422,N_18284,N_18385);
or U18423 (N_18423,N_18332,N_18311);
nand U18424 (N_18424,N_18371,N_18291);
or U18425 (N_18425,N_18264,N_18252);
xor U18426 (N_18426,N_18380,N_18259);
and U18427 (N_18427,N_18266,N_18367);
xor U18428 (N_18428,N_18297,N_18274);
xnor U18429 (N_18429,N_18392,N_18333);
nor U18430 (N_18430,N_18261,N_18292);
nor U18431 (N_18431,N_18369,N_18396);
or U18432 (N_18432,N_18370,N_18341);
xor U18433 (N_18433,N_18263,N_18398);
and U18434 (N_18434,N_18272,N_18366);
or U18435 (N_18435,N_18379,N_18293);
nand U18436 (N_18436,N_18327,N_18283);
nand U18437 (N_18437,N_18247,N_18240);
or U18438 (N_18438,N_18276,N_18383);
or U18439 (N_18439,N_18348,N_18391);
xor U18440 (N_18440,N_18350,N_18246);
xnor U18441 (N_18441,N_18310,N_18381);
and U18442 (N_18442,N_18289,N_18324);
nor U18443 (N_18443,N_18241,N_18268);
nor U18444 (N_18444,N_18250,N_18378);
nor U18445 (N_18445,N_18315,N_18394);
nor U18446 (N_18446,N_18355,N_18365);
and U18447 (N_18447,N_18295,N_18351);
nor U18448 (N_18448,N_18389,N_18294);
nand U18449 (N_18449,N_18271,N_18357);
and U18450 (N_18450,N_18384,N_18258);
and U18451 (N_18451,N_18313,N_18270);
nor U18452 (N_18452,N_18300,N_18356);
nor U18453 (N_18453,N_18363,N_18395);
nor U18454 (N_18454,N_18269,N_18388);
or U18455 (N_18455,N_18323,N_18317);
nand U18456 (N_18456,N_18359,N_18358);
nand U18457 (N_18457,N_18301,N_18299);
or U18458 (N_18458,N_18334,N_18328);
nor U18459 (N_18459,N_18372,N_18382);
nand U18460 (N_18460,N_18326,N_18373);
nand U18461 (N_18461,N_18349,N_18353);
nor U18462 (N_18462,N_18298,N_18320);
nor U18463 (N_18463,N_18352,N_18256);
or U18464 (N_18464,N_18318,N_18354);
or U18465 (N_18465,N_18339,N_18347);
xnor U18466 (N_18466,N_18308,N_18267);
nand U18467 (N_18467,N_18302,N_18253);
or U18468 (N_18468,N_18399,N_18277);
xor U18469 (N_18469,N_18245,N_18309);
or U18470 (N_18470,N_18360,N_18329);
nand U18471 (N_18471,N_18361,N_18249);
and U18472 (N_18472,N_18377,N_18243);
nand U18473 (N_18473,N_18255,N_18314);
xnor U18474 (N_18474,N_18288,N_18265);
and U18475 (N_18475,N_18312,N_18273);
nand U18476 (N_18476,N_18335,N_18304);
nand U18477 (N_18477,N_18307,N_18262);
and U18478 (N_18478,N_18286,N_18296);
xnor U18479 (N_18479,N_18374,N_18282);
xnor U18480 (N_18480,N_18393,N_18356);
and U18481 (N_18481,N_18352,N_18336);
and U18482 (N_18482,N_18393,N_18302);
or U18483 (N_18483,N_18357,N_18380);
or U18484 (N_18484,N_18364,N_18359);
xnor U18485 (N_18485,N_18301,N_18342);
nor U18486 (N_18486,N_18385,N_18370);
nand U18487 (N_18487,N_18347,N_18294);
or U18488 (N_18488,N_18398,N_18355);
nor U18489 (N_18489,N_18355,N_18256);
or U18490 (N_18490,N_18323,N_18352);
or U18491 (N_18491,N_18297,N_18385);
nand U18492 (N_18492,N_18376,N_18295);
or U18493 (N_18493,N_18258,N_18377);
or U18494 (N_18494,N_18297,N_18308);
xnor U18495 (N_18495,N_18395,N_18399);
xor U18496 (N_18496,N_18379,N_18280);
nor U18497 (N_18497,N_18368,N_18265);
nand U18498 (N_18498,N_18340,N_18278);
nor U18499 (N_18499,N_18351,N_18343);
nor U18500 (N_18500,N_18285,N_18308);
xnor U18501 (N_18501,N_18331,N_18376);
nor U18502 (N_18502,N_18395,N_18277);
xor U18503 (N_18503,N_18366,N_18286);
xor U18504 (N_18504,N_18332,N_18262);
or U18505 (N_18505,N_18314,N_18320);
nor U18506 (N_18506,N_18369,N_18368);
or U18507 (N_18507,N_18368,N_18329);
xnor U18508 (N_18508,N_18244,N_18392);
and U18509 (N_18509,N_18367,N_18391);
nor U18510 (N_18510,N_18268,N_18339);
and U18511 (N_18511,N_18269,N_18357);
nand U18512 (N_18512,N_18241,N_18395);
xor U18513 (N_18513,N_18356,N_18278);
or U18514 (N_18514,N_18278,N_18322);
and U18515 (N_18515,N_18255,N_18332);
and U18516 (N_18516,N_18338,N_18299);
nor U18517 (N_18517,N_18389,N_18247);
nand U18518 (N_18518,N_18266,N_18291);
or U18519 (N_18519,N_18280,N_18285);
or U18520 (N_18520,N_18376,N_18347);
nand U18521 (N_18521,N_18284,N_18281);
or U18522 (N_18522,N_18296,N_18302);
nor U18523 (N_18523,N_18316,N_18350);
nor U18524 (N_18524,N_18319,N_18320);
xor U18525 (N_18525,N_18245,N_18353);
nand U18526 (N_18526,N_18305,N_18352);
and U18527 (N_18527,N_18373,N_18299);
nand U18528 (N_18528,N_18369,N_18282);
and U18529 (N_18529,N_18349,N_18321);
or U18530 (N_18530,N_18334,N_18337);
or U18531 (N_18531,N_18261,N_18289);
nand U18532 (N_18532,N_18373,N_18388);
or U18533 (N_18533,N_18382,N_18290);
nand U18534 (N_18534,N_18322,N_18330);
and U18535 (N_18535,N_18241,N_18243);
nor U18536 (N_18536,N_18396,N_18377);
or U18537 (N_18537,N_18284,N_18349);
or U18538 (N_18538,N_18350,N_18378);
nand U18539 (N_18539,N_18305,N_18394);
or U18540 (N_18540,N_18306,N_18313);
nor U18541 (N_18541,N_18366,N_18377);
or U18542 (N_18542,N_18259,N_18280);
nor U18543 (N_18543,N_18307,N_18315);
xnor U18544 (N_18544,N_18350,N_18368);
or U18545 (N_18545,N_18396,N_18326);
and U18546 (N_18546,N_18364,N_18290);
nand U18547 (N_18547,N_18365,N_18393);
and U18548 (N_18548,N_18395,N_18285);
or U18549 (N_18549,N_18270,N_18290);
xnor U18550 (N_18550,N_18291,N_18348);
xnor U18551 (N_18551,N_18355,N_18263);
and U18552 (N_18552,N_18335,N_18330);
xor U18553 (N_18553,N_18295,N_18253);
and U18554 (N_18554,N_18341,N_18349);
xnor U18555 (N_18555,N_18318,N_18390);
nor U18556 (N_18556,N_18336,N_18375);
nand U18557 (N_18557,N_18284,N_18294);
nor U18558 (N_18558,N_18326,N_18249);
or U18559 (N_18559,N_18278,N_18248);
or U18560 (N_18560,N_18520,N_18424);
nor U18561 (N_18561,N_18553,N_18433);
nor U18562 (N_18562,N_18530,N_18437);
nand U18563 (N_18563,N_18442,N_18533);
or U18564 (N_18564,N_18488,N_18508);
nor U18565 (N_18565,N_18401,N_18532);
nor U18566 (N_18566,N_18494,N_18458);
nor U18567 (N_18567,N_18501,N_18426);
nor U18568 (N_18568,N_18413,N_18486);
or U18569 (N_18569,N_18429,N_18545);
nor U18570 (N_18570,N_18435,N_18524);
or U18571 (N_18571,N_18521,N_18474);
and U18572 (N_18572,N_18403,N_18446);
nand U18573 (N_18573,N_18452,N_18402);
nor U18574 (N_18574,N_18469,N_18544);
xor U18575 (N_18575,N_18484,N_18473);
and U18576 (N_18576,N_18536,N_18415);
nand U18577 (N_18577,N_18542,N_18518);
or U18578 (N_18578,N_18491,N_18467);
xor U18579 (N_18579,N_18511,N_18465);
xnor U18580 (N_18580,N_18460,N_18557);
nand U18581 (N_18581,N_18490,N_18555);
nor U18582 (N_18582,N_18483,N_18480);
nor U18583 (N_18583,N_18522,N_18495);
and U18584 (N_18584,N_18512,N_18552);
nand U18585 (N_18585,N_18478,N_18422);
or U18586 (N_18586,N_18550,N_18427);
xor U18587 (N_18587,N_18510,N_18447);
nor U18588 (N_18588,N_18537,N_18517);
nor U18589 (N_18589,N_18493,N_18459);
xor U18590 (N_18590,N_18481,N_18534);
nor U18591 (N_18591,N_18472,N_18408);
nor U18592 (N_18592,N_18436,N_18500);
and U18593 (N_18593,N_18453,N_18538);
nand U18594 (N_18594,N_18464,N_18513);
xor U18595 (N_18595,N_18431,N_18412);
and U18596 (N_18596,N_18423,N_18461);
nand U18597 (N_18597,N_18438,N_18556);
nand U18598 (N_18598,N_18425,N_18502);
nor U18599 (N_18599,N_18514,N_18479);
xnor U18600 (N_18600,N_18531,N_18439);
xnor U18601 (N_18601,N_18516,N_18410);
xnor U18602 (N_18602,N_18441,N_18466);
nand U18603 (N_18603,N_18462,N_18509);
xnor U18604 (N_18604,N_18525,N_18539);
xnor U18605 (N_18605,N_18418,N_18499);
nor U18606 (N_18606,N_18476,N_18430);
nand U18607 (N_18607,N_18409,N_18405);
or U18608 (N_18608,N_18507,N_18443);
and U18609 (N_18609,N_18440,N_18457);
and U18610 (N_18610,N_18449,N_18420);
nand U18611 (N_18611,N_18463,N_18541);
and U18612 (N_18612,N_18489,N_18468);
xnor U18613 (N_18613,N_18451,N_18496);
nand U18614 (N_18614,N_18543,N_18548);
nor U18615 (N_18615,N_18498,N_18471);
nor U18616 (N_18616,N_18400,N_18527);
nor U18617 (N_18617,N_18419,N_18515);
nor U18618 (N_18618,N_18421,N_18519);
and U18619 (N_18619,N_18540,N_18404);
nor U18620 (N_18620,N_18432,N_18434);
and U18621 (N_18621,N_18414,N_18428);
nor U18622 (N_18622,N_18448,N_18455);
or U18623 (N_18623,N_18475,N_18417);
nor U18624 (N_18624,N_18547,N_18492);
and U18625 (N_18625,N_18497,N_18445);
nand U18626 (N_18626,N_18456,N_18482);
nor U18627 (N_18627,N_18529,N_18407);
nor U18628 (N_18628,N_18526,N_18549);
xnor U18629 (N_18629,N_18487,N_18416);
nor U18630 (N_18630,N_18406,N_18470);
or U18631 (N_18631,N_18444,N_18503);
nor U18632 (N_18632,N_18454,N_18546);
nor U18633 (N_18633,N_18485,N_18558);
and U18634 (N_18634,N_18559,N_18506);
and U18635 (N_18635,N_18504,N_18450);
xnor U18636 (N_18636,N_18528,N_18554);
nand U18637 (N_18637,N_18551,N_18505);
nor U18638 (N_18638,N_18411,N_18535);
nor U18639 (N_18639,N_18523,N_18477);
nand U18640 (N_18640,N_18488,N_18423);
nor U18641 (N_18641,N_18419,N_18514);
and U18642 (N_18642,N_18482,N_18433);
xor U18643 (N_18643,N_18418,N_18530);
nand U18644 (N_18644,N_18489,N_18539);
xor U18645 (N_18645,N_18465,N_18510);
nor U18646 (N_18646,N_18558,N_18415);
xnor U18647 (N_18647,N_18476,N_18473);
nor U18648 (N_18648,N_18525,N_18548);
or U18649 (N_18649,N_18421,N_18558);
nor U18650 (N_18650,N_18528,N_18409);
and U18651 (N_18651,N_18459,N_18432);
nand U18652 (N_18652,N_18428,N_18557);
or U18653 (N_18653,N_18489,N_18450);
nor U18654 (N_18654,N_18483,N_18469);
nor U18655 (N_18655,N_18504,N_18464);
or U18656 (N_18656,N_18523,N_18534);
xnor U18657 (N_18657,N_18441,N_18418);
nand U18658 (N_18658,N_18457,N_18513);
and U18659 (N_18659,N_18464,N_18427);
or U18660 (N_18660,N_18535,N_18539);
or U18661 (N_18661,N_18553,N_18403);
nor U18662 (N_18662,N_18486,N_18448);
xnor U18663 (N_18663,N_18411,N_18468);
nor U18664 (N_18664,N_18545,N_18412);
and U18665 (N_18665,N_18460,N_18414);
nand U18666 (N_18666,N_18547,N_18419);
nor U18667 (N_18667,N_18450,N_18414);
nor U18668 (N_18668,N_18502,N_18538);
nand U18669 (N_18669,N_18454,N_18525);
nand U18670 (N_18670,N_18426,N_18455);
or U18671 (N_18671,N_18491,N_18511);
xnor U18672 (N_18672,N_18422,N_18554);
xnor U18673 (N_18673,N_18508,N_18497);
and U18674 (N_18674,N_18536,N_18480);
xor U18675 (N_18675,N_18498,N_18470);
nor U18676 (N_18676,N_18559,N_18525);
nand U18677 (N_18677,N_18455,N_18446);
nand U18678 (N_18678,N_18522,N_18438);
or U18679 (N_18679,N_18485,N_18495);
xnor U18680 (N_18680,N_18457,N_18519);
and U18681 (N_18681,N_18491,N_18404);
or U18682 (N_18682,N_18407,N_18468);
or U18683 (N_18683,N_18432,N_18408);
nand U18684 (N_18684,N_18462,N_18502);
or U18685 (N_18685,N_18517,N_18488);
xnor U18686 (N_18686,N_18472,N_18535);
xor U18687 (N_18687,N_18457,N_18430);
nand U18688 (N_18688,N_18442,N_18437);
or U18689 (N_18689,N_18480,N_18429);
and U18690 (N_18690,N_18517,N_18413);
or U18691 (N_18691,N_18433,N_18452);
and U18692 (N_18692,N_18541,N_18534);
nand U18693 (N_18693,N_18411,N_18403);
nand U18694 (N_18694,N_18524,N_18512);
xnor U18695 (N_18695,N_18553,N_18549);
xnor U18696 (N_18696,N_18417,N_18541);
nand U18697 (N_18697,N_18462,N_18470);
nor U18698 (N_18698,N_18540,N_18490);
nand U18699 (N_18699,N_18526,N_18439);
and U18700 (N_18700,N_18480,N_18549);
nor U18701 (N_18701,N_18503,N_18425);
xor U18702 (N_18702,N_18535,N_18529);
xor U18703 (N_18703,N_18445,N_18559);
xnor U18704 (N_18704,N_18458,N_18408);
nor U18705 (N_18705,N_18538,N_18512);
xnor U18706 (N_18706,N_18492,N_18439);
nor U18707 (N_18707,N_18536,N_18436);
nor U18708 (N_18708,N_18468,N_18426);
and U18709 (N_18709,N_18553,N_18404);
xnor U18710 (N_18710,N_18454,N_18533);
nor U18711 (N_18711,N_18517,N_18532);
and U18712 (N_18712,N_18559,N_18537);
nor U18713 (N_18713,N_18502,N_18535);
nor U18714 (N_18714,N_18480,N_18514);
nand U18715 (N_18715,N_18525,N_18467);
nand U18716 (N_18716,N_18431,N_18458);
nand U18717 (N_18717,N_18518,N_18413);
nor U18718 (N_18718,N_18427,N_18518);
nor U18719 (N_18719,N_18524,N_18523);
xnor U18720 (N_18720,N_18678,N_18569);
or U18721 (N_18721,N_18717,N_18658);
nand U18722 (N_18722,N_18666,N_18711);
and U18723 (N_18723,N_18576,N_18644);
xor U18724 (N_18724,N_18682,N_18680);
and U18725 (N_18725,N_18607,N_18700);
nand U18726 (N_18726,N_18625,N_18573);
or U18727 (N_18727,N_18656,N_18636);
xor U18728 (N_18728,N_18697,N_18568);
and U18729 (N_18729,N_18595,N_18616);
and U18730 (N_18730,N_18591,N_18604);
or U18731 (N_18731,N_18713,N_18574);
nor U18732 (N_18732,N_18686,N_18602);
and U18733 (N_18733,N_18619,N_18598);
or U18734 (N_18734,N_18630,N_18694);
nor U18735 (N_18735,N_18706,N_18719);
or U18736 (N_18736,N_18632,N_18642);
nand U18737 (N_18737,N_18652,N_18605);
or U18738 (N_18738,N_18701,N_18703);
nor U18739 (N_18739,N_18673,N_18661);
nor U18740 (N_18740,N_18640,N_18690);
nand U18741 (N_18741,N_18611,N_18663);
nand U18742 (N_18742,N_18597,N_18578);
xnor U18743 (N_18743,N_18708,N_18621);
and U18744 (N_18744,N_18638,N_18583);
and U18745 (N_18745,N_18702,N_18592);
nor U18746 (N_18746,N_18715,N_18596);
or U18747 (N_18747,N_18571,N_18565);
nor U18748 (N_18748,N_18566,N_18693);
xor U18749 (N_18749,N_18675,N_18631);
and U18750 (N_18750,N_18589,N_18651);
xnor U18751 (N_18751,N_18584,N_18635);
or U18752 (N_18752,N_18660,N_18648);
xnor U18753 (N_18753,N_18710,N_18582);
xor U18754 (N_18754,N_18714,N_18696);
xnor U18755 (N_18755,N_18609,N_18691);
nor U18756 (N_18756,N_18615,N_18688);
and U18757 (N_18757,N_18575,N_18590);
or U18758 (N_18758,N_18683,N_18643);
nand U18759 (N_18759,N_18587,N_18664);
or U18760 (N_18760,N_18679,N_18685);
or U18761 (N_18761,N_18671,N_18601);
nand U18762 (N_18762,N_18639,N_18654);
nand U18763 (N_18763,N_18709,N_18624);
or U18764 (N_18764,N_18672,N_18646);
nor U18765 (N_18765,N_18704,N_18674);
nor U18766 (N_18766,N_18695,N_18716);
and U18767 (N_18767,N_18562,N_18699);
xor U18768 (N_18768,N_18599,N_18603);
nand U18769 (N_18769,N_18641,N_18705);
nor U18770 (N_18770,N_18689,N_18614);
and U18771 (N_18771,N_18626,N_18655);
or U18772 (N_18772,N_18620,N_18677);
and U18773 (N_18773,N_18588,N_18662);
nand U18774 (N_18774,N_18561,N_18667);
and U18775 (N_18775,N_18628,N_18634);
nand U18776 (N_18776,N_18618,N_18637);
nor U18777 (N_18777,N_18600,N_18612);
and U18778 (N_18778,N_18687,N_18567);
xnor U18779 (N_18779,N_18572,N_18563);
nor U18780 (N_18780,N_18606,N_18594);
nor U18781 (N_18781,N_18579,N_18627);
nand U18782 (N_18782,N_18681,N_18608);
xnor U18783 (N_18783,N_18613,N_18585);
and U18784 (N_18784,N_18617,N_18629);
or U18785 (N_18785,N_18560,N_18698);
and U18786 (N_18786,N_18593,N_18684);
nor U18787 (N_18787,N_18712,N_18610);
and U18788 (N_18788,N_18633,N_18718);
and U18789 (N_18789,N_18650,N_18659);
nor U18790 (N_18790,N_18692,N_18623);
and U18791 (N_18791,N_18581,N_18577);
xor U18792 (N_18792,N_18570,N_18649);
nand U18793 (N_18793,N_18653,N_18668);
xnor U18794 (N_18794,N_18564,N_18586);
nand U18795 (N_18795,N_18707,N_18669);
xnor U18796 (N_18796,N_18647,N_18580);
and U18797 (N_18797,N_18676,N_18665);
xor U18798 (N_18798,N_18657,N_18670);
or U18799 (N_18799,N_18645,N_18622);
xnor U18800 (N_18800,N_18624,N_18707);
nand U18801 (N_18801,N_18708,N_18611);
nor U18802 (N_18802,N_18591,N_18584);
nor U18803 (N_18803,N_18694,N_18672);
or U18804 (N_18804,N_18700,N_18683);
nand U18805 (N_18805,N_18709,N_18574);
and U18806 (N_18806,N_18663,N_18592);
nand U18807 (N_18807,N_18716,N_18719);
nand U18808 (N_18808,N_18588,N_18679);
nand U18809 (N_18809,N_18589,N_18613);
or U18810 (N_18810,N_18705,N_18665);
nor U18811 (N_18811,N_18568,N_18698);
nand U18812 (N_18812,N_18602,N_18667);
and U18813 (N_18813,N_18699,N_18629);
nor U18814 (N_18814,N_18629,N_18561);
xnor U18815 (N_18815,N_18706,N_18603);
or U18816 (N_18816,N_18638,N_18594);
or U18817 (N_18817,N_18710,N_18692);
and U18818 (N_18818,N_18690,N_18663);
or U18819 (N_18819,N_18719,N_18571);
nor U18820 (N_18820,N_18642,N_18705);
nand U18821 (N_18821,N_18604,N_18594);
and U18822 (N_18822,N_18704,N_18699);
nor U18823 (N_18823,N_18589,N_18579);
nor U18824 (N_18824,N_18561,N_18659);
and U18825 (N_18825,N_18714,N_18610);
or U18826 (N_18826,N_18717,N_18605);
or U18827 (N_18827,N_18669,N_18668);
and U18828 (N_18828,N_18719,N_18578);
or U18829 (N_18829,N_18587,N_18666);
or U18830 (N_18830,N_18687,N_18606);
and U18831 (N_18831,N_18612,N_18573);
nand U18832 (N_18832,N_18617,N_18649);
and U18833 (N_18833,N_18710,N_18668);
nand U18834 (N_18834,N_18669,N_18591);
nor U18835 (N_18835,N_18629,N_18718);
nor U18836 (N_18836,N_18633,N_18588);
and U18837 (N_18837,N_18639,N_18668);
nor U18838 (N_18838,N_18707,N_18700);
xor U18839 (N_18839,N_18717,N_18674);
nor U18840 (N_18840,N_18645,N_18601);
nand U18841 (N_18841,N_18626,N_18712);
xnor U18842 (N_18842,N_18657,N_18694);
or U18843 (N_18843,N_18719,N_18576);
or U18844 (N_18844,N_18568,N_18601);
nor U18845 (N_18845,N_18703,N_18674);
nand U18846 (N_18846,N_18641,N_18699);
or U18847 (N_18847,N_18593,N_18691);
nor U18848 (N_18848,N_18681,N_18631);
xor U18849 (N_18849,N_18633,N_18641);
xnor U18850 (N_18850,N_18658,N_18645);
and U18851 (N_18851,N_18576,N_18612);
or U18852 (N_18852,N_18567,N_18689);
xnor U18853 (N_18853,N_18595,N_18599);
and U18854 (N_18854,N_18604,N_18689);
xor U18855 (N_18855,N_18613,N_18583);
or U18856 (N_18856,N_18678,N_18590);
xnor U18857 (N_18857,N_18616,N_18564);
xor U18858 (N_18858,N_18680,N_18710);
xnor U18859 (N_18859,N_18704,N_18562);
nor U18860 (N_18860,N_18565,N_18605);
and U18861 (N_18861,N_18620,N_18610);
or U18862 (N_18862,N_18575,N_18643);
nand U18863 (N_18863,N_18641,N_18685);
or U18864 (N_18864,N_18704,N_18676);
or U18865 (N_18865,N_18672,N_18701);
or U18866 (N_18866,N_18701,N_18580);
nand U18867 (N_18867,N_18622,N_18576);
xnor U18868 (N_18868,N_18578,N_18576);
nor U18869 (N_18869,N_18709,N_18612);
xor U18870 (N_18870,N_18689,N_18607);
nand U18871 (N_18871,N_18672,N_18697);
or U18872 (N_18872,N_18700,N_18682);
or U18873 (N_18873,N_18571,N_18587);
and U18874 (N_18874,N_18654,N_18711);
or U18875 (N_18875,N_18675,N_18684);
xnor U18876 (N_18876,N_18560,N_18676);
and U18877 (N_18877,N_18686,N_18683);
nor U18878 (N_18878,N_18684,N_18677);
nor U18879 (N_18879,N_18672,N_18594);
nor U18880 (N_18880,N_18808,N_18812);
and U18881 (N_18881,N_18787,N_18863);
nor U18882 (N_18882,N_18839,N_18872);
nand U18883 (N_18883,N_18758,N_18725);
xor U18884 (N_18884,N_18753,N_18746);
xor U18885 (N_18885,N_18771,N_18747);
xor U18886 (N_18886,N_18790,N_18735);
and U18887 (N_18887,N_18760,N_18806);
nor U18888 (N_18888,N_18728,N_18737);
or U18889 (N_18889,N_18794,N_18843);
and U18890 (N_18890,N_18866,N_18763);
nand U18891 (N_18891,N_18798,N_18785);
nor U18892 (N_18892,N_18727,N_18765);
or U18893 (N_18893,N_18722,N_18743);
and U18894 (N_18894,N_18802,N_18836);
or U18895 (N_18895,N_18804,N_18830);
nand U18896 (N_18896,N_18762,N_18814);
nand U18897 (N_18897,N_18878,N_18849);
nor U18898 (N_18898,N_18869,N_18871);
nand U18899 (N_18899,N_18870,N_18831);
nor U18900 (N_18900,N_18773,N_18741);
nand U18901 (N_18901,N_18826,N_18770);
and U18902 (N_18902,N_18797,N_18769);
and U18903 (N_18903,N_18755,N_18852);
or U18904 (N_18904,N_18840,N_18823);
or U18905 (N_18905,N_18857,N_18854);
nor U18906 (N_18906,N_18759,N_18739);
xor U18907 (N_18907,N_18767,N_18850);
and U18908 (N_18908,N_18782,N_18800);
or U18909 (N_18909,N_18845,N_18732);
xor U18910 (N_18910,N_18786,N_18721);
nand U18911 (N_18911,N_18818,N_18780);
and U18912 (N_18912,N_18734,N_18875);
xor U18913 (N_18913,N_18811,N_18768);
nand U18914 (N_18914,N_18778,N_18873);
nor U18915 (N_18915,N_18820,N_18807);
nor U18916 (N_18916,N_18766,N_18748);
xnor U18917 (N_18917,N_18856,N_18847);
xnor U18918 (N_18918,N_18874,N_18777);
xnor U18919 (N_18919,N_18775,N_18877);
nor U18920 (N_18920,N_18783,N_18835);
and U18921 (N_18921,N_18729,N_18825);
or U18922 (N_18922,N_18796,N_18761);
nand U18923 (N_18923,N_18861,N_18744);
nand U18924 (N_18924,N_18738,N_18832);
nor U18925 (N_18925,N_18859,N_18865);
and U18926 (N_18926,N_18833,N_18801);
and U18927 (N_18927,N_18844,N_18779);
nand U18928 (N_18928,N_18803,N_18858);
nor U18929 (N_18929,N_18730,N_18822);
xor U18930 (N_18930,N_18816,N_18819);
or U18931 (N_18931,N_18784,N_18726);
nor U18932 (N_18932,N_18772,N_18757);
nor U18933 (N_18933,N_18828,N_18723);
nand U18934 (N_18934,N_18838,N_18751);
xnor U18935 (N_18935,N_18754,N_18842);
or U18936 (N_18936,N_18862,N_18810);
or U18937 (N_18937,N_18799,N_18740);
and U18938 (N_18938,N_18792,N_18837);
nor U18939 (N_18939,N_18867,N_18736);
xnor U18940 (N_18940,N_18829,N_18750);
nand U18941 (N_18941,N_18791,N_18821);
or U18942 (N_18942,N_18776,N_18813);
xnor U18943 (N_18943,N_18749,N_18809);
and U18944 (N_18944,N_18855,N_18868);
and U18945 (N_18945,N_18724,N_18817);
and U18946 (N_18946,N_18851,N_18795);
xnor U18947 (N_18947,N_18756,N_18793);
nor U18948 (N_18948,N_18745,N_18848);
nand U18949 (N_18949,N_18824,N_18731);
or U18950 (N_18950,N_18815,N_18853);
and U18951 (N_18951,N_18841,N_18827);
and U18952 (N_18952,N_18876,N_18846);
nor U18953 (N_18953,N_18774,N_18781);
and U18954 (N_18954,N_18720,N_18860);
or U18955 (N_18955,N_18788,N_18879);
or U18956 (N_18956,N_18789,N_18864);
nor U18957 (N_18957,N_18834,N_18752);
or U18958 (N_18958,N_18742,N_18805);
nor U18959 (N_18959,N_18764,N_18733);
or U18960 (N_18960,N_18821,N_18849);
and U18961 (N_18961,N_18748,N_18749);
nand U18962 (N_18962,N_18749,N_18728);
nor U18963 (N_18963,N_18864,N_18800);
or U18964 (N_18964,N_18772,N_18791);
xor U18965 (N_18965,N_18787,N_18811);
nand U18966 (N_18966,N_18795,N_18776);
xnor U18967 (N_18967,N_18865,N_18792);
nor U18968 (N_18968,N_18764,N_18866);
xnor U18969 (N_18969,N_18786,N_18835);
and U18970 (N_18970,N_18843,N_18727);
and U18971 (N_18971,N_18827,N_18859);
xor U18972 (N_18972,N_18761,N_18822);
xor U18973 (N_18973,N_18721,N_18774);
and U18974 (N_18974,N_18769,N_18755);
or U18975 (N_18975,N_18832,N_18765);
nand U18976 (N_18976,N_18779,N_18858);
and U18977 (N_18977,N_18824,N_18801);
and U18978 (N_18978,N_18799,N_18832);
nor U18979 (N_18979,N_18748,N_18822);
nand U18980 (N_18980,N_18798,N_18770);
and U18981 (N_18981,N_18761,N_18741);
or U18982 (N_18982,N_18856,N_18793);
xor U18983 (N_18983,N_18766,N_18780);
and U18984 (N_18984,N_18849,N_18759);
xor U18985 (N_18985,N_18784,N_18799);
and U18986 (N_18986,N_18823,N_18831);
nor U18987 (N_18987,N_18856,N_18855);
or U18988 (N_18988,N_18827,N_18816);
and U18989 (N_18989,N_18839,N_18803);
or U18990 (N_18990,N_18878,N_18866);
nor U18991 (N_18991,N_18834,N_18873);
nand U18992 (N_18992,N_18822,N_18756);
nor U18993 (N_18993,N_18824,N_18724);
or U18994 (N_18994,N_18787,N_18868);
nor U18995 (N_18995,N_18802,N_18834);
or U18996 (N_18996,N_18860,N_18848);
nor U18997 (N_18997,N_18786,N_18813);
xnor U18998 (N_18998,N_18862,N_18774);
nor U18999 (N_18999,N_18734,N_18837);
nor U19000 (N_19000,N_18845,N_18784);
nor U19001 (N_19001,N_18725,N_18768);
or U19002 (N_19002,N_18738,N_18726);
and U19003 (N_19003,N_18798,N_18814);
nor U19004 (N_19004,N_18758,N_18840);
and U19005 (N_19005,N_18837,N_18847);
and U19006 (N_19006,N_18814,N_18724);
or U19007 (N_19007,N_18838,N_18750);
xnor U19008 (N_19008,N_18868,N_18862);
nand U19009 (N_19009,N_18842,N_18822);
nor U19010 (N_19010,N_18840,N_18878);
nand U19011 (N_19011,N_18829,N_18809);
nand U19012 (N_19012,N_18762,N_18793);
and U19013 (N_19013,N_18825,N_18848);
xor U19014 (N_19014,N_18764,N_18856);
and U19015 (N_19015,N_18851,N_18726);
xor U19016 (N_19016,N_18747,N_18868);
or U19017 (N_19017,N_18759,N_18805);
or U19018 (N_19018,N_18762,N_18854);
and U19019 (N_19019,N_18777,N_18759);
or U19020 (N_19020,N_18726,N_18857);
and U19021 (N_19021,N_18763,N_18852);
nor U19022 (N_19022,N_18786,N_18841);
and U19023 (N_19023,N_18739,N_18842);
nor U19024 (N_19024,N_18777,N_18840);
or U19025 (N_19025,N_18869,N_18841);
and U19026 (N_19026,N_18743,N_18795);
nand U19027 (N_19027,N_18842,N_18845);
and U19028 (N_19028,N_18842,N_18859);
xor U19029 (N_19029,N_18861,N_18777);
nand U19030 (N_19030,N_18758,N_18768);
nor U19031 (N_19031,N_18767,N_18725);
and U19032 (N_19032,N_18836,N_18799);
or U19033 (N_19033,N_18731,N_18721);
nor U19034 (N_19034,N_18828,N_18743);
and U19035 (N_19035,N_18793,N_18737);
nor U19036 (N_19036,N_18823,N_18739);
nor U19037 (N_19037,N_18755,N_18803);
nor U19038 (N_19038,N_18831,N_18840);
and U19039 (N_19039,N_18816,N_18849);
nand U19040 (N_19040,N_18880,N_18930);
or U19041 (N_19041,N_18926,N_18934);
and U19042 (N_19042,N_18935,N_18972);
nor U19043 (N_19043,N_18938,N_18893);
nor U19044 (N_19044,N_18923,N_18950);
nand U19045 (N_19045,N_18920,N_18936);
xnor U19046 (N_19046,N_18987,N_18957);
nand U19047 (N_19047,N_18925,N_18974);
and U19048 (N_19048,N_18988,N_19028);
nand U19049 (N_19049,N_18929,N_18958);
xor U19050 (N_19050,N_18921,N_18952);
xnor U19051 (N_19051,N_18889,N_18986);
and U19052 (N_19052,N_18985,N_18981);
or U19053 (N_19053,N_19008,N_18907);
nand U19054 (N_19054,N_19026,N_18970);
or U19055 (N_19055,N_18931,N_18960);
or U19056 (N_19056,N_18975,N_18997);
nand U19057 (N_19057,N_18977,N_18899);
or U19058 (N_19058,N_18906,N_18881);
nand U19059 (N_19059,N_18976,N_18979);
nand U19060 (N_19060,N_19037,N_18946);
xor U19061 (N_19061,N_19038,N_18910);
nand U19062 (N_19062,N_18883,N_19015);
xnor U19063 (N_19063,N_19010,N_19002);
nand U19064 (N_19064,N_18983,N_18953);
or U19065 (N_19065,N_19019,N_18944);
and U19066 (N_19066,N_18890,N_18994);
nand U19067 (N_19067,N_19003,N_18888);
nand U19068 (N_19068,N_18941,N_19034);
and U19069 (N_19069,N_18965,N_19025);
xor U19070 (N_19070,N_19020,N_18966);
or U19071 (N_19071,N_19004,N_18991);
nand U19072 (N_19072,N_18905,N_19012);
or U19073 (N_19073,N_18927,N_19013);
nand U19074 (N_19074,N_18917,N_18971);
xnor U19075 (N_19075,N_18891,N_18898);
xnor U19076 (N_19076,N_19023,N_18908);
nand U19077 (N_19077,N_18999,N_18992);
xnor U19078 (N_19078,N_19036,N_19006);
nor U19079 (N_19079,N_19001,N_18990);
nand U19080 (N_19080,N_19016,N_19007);
nand U19081 (N_19081,N_19024,N_18933);
xor U19082 (N_19082,N_18904,N_18900);
xnor U19083 (N_19083,N_18964,N_18998);
and U19084 (N_19084,N_18968,N_18911);
xor U19085 (N_19085,N_18980,N_18951);
xnor U19086 (N_19086,N_18909,N_18897);
or U19087 (N_19087,N_18945,N_18943);
or U19088 (N_19088,N_18892,N_18959);
and U19089 (N_19089,N_18993,N_18969);
or U19090 (N_19090,N_18894,N_19005);
and U19091 (N_19091,N_18887,N_18996);
and U19092 (N_19092,N_18942,N_18896);
and U19093 (N_19093,N_18922,N_18995);
or U19094 (N_19094,N_18963,N_18884);
or U19095 (N_19095,N_18895,N_19022);
or U19096 (N_19096,N_18961,N_18902);
or U19097 (N_19097,N_18928,N_18956);
nor U19098 (N_19098,N_18932,N_18914);
nand U19099 (N_19099,N_18919,N_18947);
nor U19100 (N_19100,N_18903,N_18967);
and U19101 (N_19101,N_18973,N_18918);
and U19102 (N_19102,N_19027,N_18916);
xor U19103 (N_19103,N_19039,N_18912);
or U19104 (N_19104,N_18948,N_18924);
xor U19105 (N_19105,N_19018,N_19032);
and U19106 (N_19106,N_19031,N_19035);
or U19107 (N_19107,N_19009,N_18915);
nand U19108 (N_19108,N_19014,N_18885);
or U19109 (N_19109,N_19011,N_18984);
xnor U19110 (N_19110,N_18982,N_18882);
xor U19111 (N_19111,N_18955,N_18886);
nor U19112 (N_19112,N_19017,N_18989);
or U19113 (N_19113,N_18939,N_18901);
nor U19114 (N_19114,N_19029,N_19030);
or U19115 (N_19115,N_18954,N_18978);
or U19116 (N_19116,N_19000,N_18913);
and U19117 (N_19117,N_18962,N_18940);
and U19118 (N_19118,N_19021,N_18949);
or U19119 (N_19119,N_18937,N_19033);
nor U19120 (N_19120,N_19028,N_18915);
xor U19121 (N_19121,N_18884,N_18989);
nor U19122 (N_19122,N_18901,N_18883);
nor U19123 (N_19123,N_18912,N_18946);
or U19124 (N_19124,N_18931,N_18969);
nor U19125 (N_19125,N_18959,N_18917);
and U19126 (N_19126,N_18992,N_18926);
nor U19127 (N_19127,N_19031,N_18881);
xor U19128 (N_19128,N_18919,N_18966);
nand U19129 (N_19129,N_18945,N_19019);
nand U19130 (N_19130,N_18900,N_18927);
xnor U19131 (N_19131,N_18882,N_19016);
nor U19132 (N_19132,N_18936,N_18894);
xnor U19133 (N_19133,N_18987,N_19017);
nand U19134 (N_19134,N_18904,N_18916);
xor U19135 (N_19135,N_18886,N_18913);
and U19136 (N_19136,N_18923,N_18991);
and U19137 (N_19137,N_19005,N_18893);
or U19138 (N_19138,N_18887,N_18941);
and U19139 (N_19139,N_18963,N_18902);
nand U19140 (N_19140,N_18918,N_18896);
and U19141 (N_19141,N_18913,N_18927);
nand U19142 (N_19142,N_18892,N_18940);
nor U19143 (N_19143,N_18952,N_18900);
nor U19144 (N_19144,N_18952,N_19022);
nor U19145 (N_19145,N_18956,N_19015);
nor U19146 (N_19146,N_19025,N_19021);
or U19147 (N_19147,N_18950,N_18905);
xnor U19148 (N_19148,N_18924,N_18906);
xnor U19149 (N_19149,N_18906,N_18969);
and U19150 (N_19150,N_18969,N_18919);
and U19151 (N_19151,N_18953,N_18995);
and U19152 (N_19152,N_18917,N_19023);
or U19153 (N_19153,N_18914,N_18952);
or U19154 (N_19154,N_18940,N_18936);
nor U19155 (N_19155,N_18889,N_18943);
nand U19156 (N_19156,N_18979,N_18893);
nor U19157 (N_19157,N_18893,N_18963);
nor U19158 (N_19158,N_19038,N_18880);
nor U19159 (N_19159,N_18996,N_18954);
or U19160 (N_19160,N_18983,N_18930);
nor U19161 (N_19161,N_18963,N_18936);
nand U19162 (N_19162,N_19021,N_18906);
nand U19163 (N_19163,N_18939,N_18917);
nor U19164 (N_19164,N_18906,N_18882);
or U19165 (N_19165,N_19002,N_19028);
and U19166 (N_19166,N_18964,N_18992);
or U19167 (N_19167,N_19017,N_18885);
nand U19168 (N_19168,N_19021,N_18914);
nor U19169 (N_19169,N_18997,N_18942);
nand U19170 (N_19170,N_19022,N_19025);
and U19171 (N_19171,N_18941,N_18903);
nor U19172 (N_19172,N_18897,N_19030);
and U19173 (N_19173,N_18894,N_18971);
and U19174 (N_19174,N_18899,N_19025);
nand U19175 (N_19175,N_18969,N_18933);
xnor U19176 (N_19176,N_18982,N_19018);
and U19177 (N_19177,N_18977,N_19039);
nand U19178 (N_19178,N_18898,N_18910);
nor U19179 (N_19179,N_18904,N_19035);
xnor U19180 (N_19180,N_18979,N_18999);
or U19181 (N_19181,N_18931,N_19036);
nand U19182 (N_19182,N_18887,N_19013);
or U19183 (N_19183,N_19008,N_18896);
nor U19184 (N_19184,N_18929,N_19008);
or U19185 (N_19185,N_18880,N_18989);
nand U19186 (N_19186,N_18932,N_18976);
or U19187 (N_19187,N_19017,N_18953);
and U19188 (N_19188,N_18903,N_19025);
xor U19189 (N_19189,N_19018,N_19010);
nand U19190 (N_19190,N_19008,N_18959);
xor U19191 (N_19191,N_18881,N_19006);
or U19192 (N_19192,N_18924,N_19012);
xor U19193 (N_19193,N_18917,N_18921);
xnor U19194 (N_19194,N_18994,N_19023);
and U19195 (N_19195,N_18958,N_18910);
nand U19196 (N_19196,N_19009,N_19022);
and U19197 (N_19197,N_19007,N_18890);
and U19198 (N_19198,N_18903,N_18895);
and U19199 (N_19199,N_18984,N_18961);
and U19200 (N_19200,N_19093,N_19117);
and U19201 (N_19201,N_19172,N_19195);
and U19202 (N_19202,N_19052,N_19105);
and U19203 (N_19203,N_19078,N_19061);
xnor U19204 (N_19204,N_19095,N_19196);
nor U19205 (N_19205,N_19171,N_19167);
nor U19206 (N_19206,N_19118,N_19136);
nor U19207 (N_19207,N_19109,N_19113);
or U19208 (N_19208,N_19069,N_19180);
and U19209 (N_19209,N_19150,N_19125);
or U19210 (N_19210,N_19175,N_19141);
nand U19211 (N_19211,N_19074,N_19126);
nor U19212 (N_19212,N_19155,N_19191);
and U19213 (N_19213,N_19197,N_19144);
and U19214 (N_19214,N_19173,N_19084);
nor U19215 (N_19215,N_19177,N_19193);
nor U19216 (N_19216,N_19176,N_19154);
xor U19217 (N_19217,N_19156,N_19116);
nor U19218 (N_19218,N_19070,N_19045);
and U19219 (N_19219,N_19063,N_19168);
or U19220 (N_19220,N_19146,N_19164);
or U19221 (N_19221,N_19137,N_19131);
or U19222 (N_19222,N_19089,N_19130);
xnor U19223 (N_19223,N_19088,N_19111);
or U19224 (N_19224,N_19099,N_19096);
nor U19225 (N_19225,N_19056,N_19148);
or U19226 (N_19226,N_19059,N_19139);
nor U19227 (N_19227,N_19067,N_19047);
nand U19228 (N_19228,N_19182,N_19066);
nor U19229 (N_19229,N_19120,N_19153);
and U19230 (N_19230,N_19040,N_19127);
xnor U19231 (N_19231,N_19194,N_19138);
or U19232 (N_19232,N_19190,N_19103);
xnor U19233 (N_19233,N_19149,N_19179);
nor U19234 (N_19234,N_19152,N_19049);
or U19235 (N_19235,N_19188,N_19134);
or U19236 (N_19236,N_19170,N_19142);
xor U19237 (N_19237,N_19097,N_19083);
or U19238 (N_19238,N_19145,N_19062);
or U19239 (N_19239,N_19077,N_19058);
xnor U19240 (N_19240,N_19124,N_19053);
nand U19241 (N_19241,N_19107,N_19114);
and U19242 (N_19242,N_19080,N_19187);
nand U19243 (N_19243,N_19108,N_19046);
xor U19244 (N_19244,N_19199,N_19106);
and U19245 (N_19245,N_19165,N_19178);
nor U19246 (N_19246,N_19132,N_19184);
or U19247 (N_19247,N_19082,N_19169);
and U19248 (N_19248,N_19041,N_19163);
nor U19249 (N_19249,N_19166,N_19051);
xnor U19250 (N_19250,N_19123,N_19189);
nor U19251 (N_19251,N_19048,N_19174);
nor U19252 (N_19252,N_19147,N_19151);
or U19253 (N_19253,N_19057,N_19181);
and U19254 (N_19254,N_19086,N_19094);
nor U19255 (N_19255,N_19186,N_19085);
and U19256 (N_19256,N_19087,N_19104);
and U19257 (N_19257,N_19101,N_19112);
xor U19258 (N_19258,N_19162,N_19133);
and U19259 (N_19259,N_19050,N_19055);
and U19260 (N_19260,N_19079,N_19140);
xnor U19261 (N_19261,N_19198,N_19185);
nor U19262 (N_19262,N_19064,N_19143);
nor U19263 (N_19263,N_19091,N_19060);
nand U19264 (N_19264,N_19158,N_19073);
nor U19265 (N_19265,N_19128,N_19115);
nand U19266 (N_19266,N_19122,N_19121);
nor U19267 (N_19267,N_19090,N_19072);
nor U19268 (N_19268,N_19161,N_19068);
nor U19269 (N_19269,N_19054,N_19160);
or U19270 (N_19270,N_19043,N_19065);
xor U19271 (N_19271,N_19081,N_19135);
xnor U19272 (N_19272,N_19092,N_19157);
or U19273 (N_19273,N_19100,N_19071);
xor U19274 (N_19274,N_19102,N_19119);
nand U19275 (N_19275,N_19042,N_19192);
nand U19276 (N_19276,N_19129,N_19183);
or U19277 (N_19277,N_19075,N_19044);
xor U19278 (N_19278,N_19098,N_19159);
nand U19279 (N_19279,N_19110,N_19076);
and U19280 (N_19280,N_19149,N_19116);
nand U19281 (N_19281,N_19187,N_19184);
xor U19282 (N_19282,N_19100,N_19183);
nor U19283 (N_19283,N_19099,N_19149);
nor U19284 (N_19284,N_19092,N_19119);
and U19285 (N_19285,N_19071,N_19087);
and U19286 (N_19286,N_19129,N_19174);
and U19287 (N_19287,N_19056,N_19184);
nor U19288 (N_19288,N_19061,N_19157);
and U19289 (N_19289,N_19042,N_19173);
or U19290 (N_19290,N_19187,N_19166);
nand U19291 (N_19291,N_19138,N_19050);
or U19292 (N_19292,N_19086,N_19110);
and U19293 (N_19293,N_19081,N_19073);
and U19294 (N_19294,N_19116,N_19070);
or U19295 (N_19295,N_19075,N_19090);
nor U19296 (N_19296,N_19079,N_19109);
nand U19297 (N_19297,N_19167,N_19147);
nand U19298 (N_19298,N_19062,N_19104);
nor U19299 (N_19299,N_19150,N_19151);
xor U19300 (N_19300,N_19128,N_19150);
nand U19301 (N_19301,N_19069,N_19192);
or U19302 (N_19302,N_19042,N_19100);
nand U19303 (N_19303,N_19192,N_19158);
and U19304 (N_19304,N_19108,N_19195);
nor U19305 (N_19305,N_19143,N_19118);
xnor U19306 (N_19306,N_19059,N_19078);
nand U19307 (N_19307,N_19110,N_19096);
or U19308 (N_19308,N_19062,N_19147);
nor U19309 (N_19309,N_19101,N_19042);
and U19310 (N_19310,N_19199,N_19067);
and U19311 (N_19311,N_19171,N_19087);
nand U19312 (N_19312,N_19189,N_19186);
and U19313 (N_19313,N_19136,N_19067);
xnor U19314 (N_19314,N_19044,N_19179);
nor U19315 (N_19315,N_19055,N_19051);
and U19316 (N_19316,N_19132,N_19113);
nand U19317 (N_19317,N_19153,N_19188);
or U19318 (N_19318,N_19188,N_19165);
nand U19319 (N_19319,N_19112,N_19058);
and U19320 (N_19320,N_19129,N_19080);
and U19321 (N_19321,N_19182,N_19191);
and U19322 (N_19322,N_19130,N_19057);
and U19323 (N_19323,N_19047,N_19091);
or U19324 (N_19324,N_19116,N_19086);
nand U19325 (N_19325,N_19068,N_19175);
nand U19326 (N_19326,N_19180,N_19172);
nand U19327 (N_19327,N_19072,N_19075);
and U19328 (N_19328,N_19191,N_19095);
nor U19329 (N_19329,N_19138,N_19190);
nand U19330 (N_19330,N_19101,N_19106);
nor U19331 (N_19331,N_19163,N_19073);
and U19332 (N_19332,N_19091,N_19138);
xor U19333 (N_19333,N_19076,N_19092);
and U19334 (N_19334,N_19075,N_19135);
xnor U19335 (N_19335,N_19046,N_19182);
and U19336 (N_19336,N_19089,N_19055);
nand U19337 (N_19337,N_19058,N_19090);
xor U19338 (N_19338,N_19057,N_19172);
and U19339 (N_19339,N_19157,N_19186);
nand U19340 (N_19340,N_19098,N_19185);
nand U19341 (N_19341,N_19057,N_19199);
xnor U19342 (N_19342,N_19165,N_19083);
nor U19343 (N_19343,N_19045,N_19111);
nor U19344 (N_19344,N_19161,N_19166);
xnor U19345 (N_19345,N_19153,N_19142);
nand U19346 (N_19346,N_19178,N_19103);
xnor U19347 (N_19347,N_19123,N_19081);
and U19348 (N_19348,N_19069,N_19104);
nor U19349 (N_19349,N_19092,N_19087);
and U19350 (N_19350,N_19111,N_19120);
xor U19351 (N_19351,N_19146,N_19061);
nand U19352 (N_19352,N_19135,N_19078);
nor U19353 (N_19353,N_19185,N_19175);
nor U19354 (N_19354,N_19051,N_19068);
nand U19355 (N_19355,N_19081,N_19182);
xnor U19356 (N_19356,N_19135,N_19045);
or U19357 (N_19357,N_19160,N_19092);
and U19358 (N_19358,N_19111,N_19181);
and U19359 (N_19359,N_19073,N_19129);
nand U19360 (N_19360,N_19302,N_19201);
xnor U19361 (N_19361,N_19281,N_19222);
or U19362 (N_19362,N_19290,N_19348);
or U19363 (N_19363,N_19349,N_19326);
and U19364 (N_19364,N_19214,N_19252);
nor U19365 (N_19365,N_19221,N_19200);
xnor U19366 (N_19366,N_19242,N_19213);
or U19367 (N_19367,N_19299,N_19257);
nor U19368 (N_19368,N_19263,N_19323);
nand U19369 (N_19369,N_19311,N_19205);
nand U19370 (N_19370,N_19286,N_19235);
nand U19371 (N_19371,N_19340,N_19225);
nor U19372 (N_19372,N_19271,N_19224);
xor U19373 (N_19373,N_19218,N_19246);
xnor U19374 (N_19374,N_19353,N_19301);
nand U19375 (N_19375,N_19317,N_19313);
nor U19376 (N_19376,N_19335,N_19328);
and U19377 (N_19377,N_19244,N_19256);
nand U19378 (N_19378,N_19356,N_19274);
xor U19379 (N_19379,N_19273,N_19337);
or U19380 (N_19380,N_19260,N_19261);
and U19381 (N_19381,N_19347,N_19240);
xnor U19382 (N_19382,N_19230,N_19316);
nor U19383 (N_19383,N_19231,N_19278);
and U19384 (N_19384,N_19283,N_19219);
nor U19385 (N_19385,N_19314,N_19354);
nand U19386 (N_19386,N_19295,N_19220);
or U19387 (N_19387,N_19296,N_19289);
or U19388 (N_19388,N_19344,N_19331);
and U19389 (N_19389,N_19282,N_19357);
nor U19390 (N_19390,N_19208,N_19312);
nand U19391 (N_19391,N_19203,N_19236);
or U19392 (N_19392,N_19292,N_19322);
or U19393 (N_19393,N_19265,N_19234);
nor U19394 (N_19394,N_19300,N_19209);
and U19395 (N_19395,N_19215,N_19321);
nand U19396 (N_19396,N_19298,N_19207);
nor U19397 (N_19397,N_19249,N_19206);
and U19398 (N_19398,N_19287,N_19343);
nor U19399 (N_19399,N_19336,N_19284);
xor U19400 (N_19400,N_19254,N_19232);
nand U19401 (N_19401,N_19293,N_19248);
or U19402 (N_19402,N_19303,N_19294);
or U19403 (N_19403,N_19251,N_19346);
nor U19404 (N_19404,N_19266,N_19358);
nor U19405 (N_19405,N_19239,N_19329);
or U19406 (N_19406,N_19210,N_19342);
or U19407 (N_19407,N_19226,N_19279);
xor U19408 (N_19408,N_19307,N_19351);
nand U19409 (N_19409,N_19217,N_19268);
nor U19410 (N_19410,N_19228,N_19276);
nor U19411 (N_19411,N_19325,N_19238);
and U19412 (N_19412,N_19237,N_19275);
nor U19413 (N_19413,N_19332,N_19309);
or U19414 (N_19414,N_19330,N_19269);
xor U19415 (N_19415,N_19280,N_19359);
nand U19416 (N_19416,N_19233,N_19288);
or U19417 (N_19417,N_19315,N_19339);
or U19418 (N_19418,N_19319,N_19270);
and U19419 (N_19419,N_19255,N_19334);
or U19420 (N_19420,N_19247,N_19350);
xnor U19421 (N_19421,N_19310,N_19291);
and U19422 (N_19422,N_19223,N_19241);
nor U19423 (N_19423,N_19264,N_19285);
or U19424 (N_19424,N_19250,N_19306);
and U19425 (N_19425,N_19333,N_19211);
nand U19426 (N_19426,N_19320,N_19229);
xnor U19427 (N_19427,N_19324,N_19227);
and U19428 (N_19428,N_19308,N_19341);
xnor U19429 (N_19429,N_19297,N_19305);
and U19430 (N_19430,N_19262,N_19355);
nor U19431 (N_19431,N_19212,N_19338);
nor U19432 (N_19432,N_19259,N_19258);
and U19433 (N_19433,N_19253,N_19345);
nand U19434 (N_19434,N_19327,N_19318);
nand U19435 (N_19435,N_19202,N_19304);
nor U19436 (N_19436,N_19245,N_19267);
and U19437 (N_19437,N_19352,N_19277);
and U19438 (N_19438,N_19216,N_19272);
nor U19439 (N_19439,N_19243,N_19204);
or U19440 (N_19440,N_19251,N_19350);
xor U19441 (N_19441,N_19214,N_19335);
or U19442 (N_19442,N_19288,N_19324);
nand U19443 (N_19443,N_19207,N_19340);
or U19444 (N_19444,N_19255,N_19305);
or U19445 (N_19445,N_19243,N_19289);
and U19446 (N_19446,N_19231,N_19233);
nor U19447 (N_19447,N_19252,N_19317);
nor U19448 (N_19448,N_19319,N_19303);
xor U19449 (N_19449,N_19231,N_19322);
or U19450 (N_19450,N_19271,N_19338);
and U19451 (N_19451,N_19203,N_19357);
or U19452 (N_19452,N_19293,N_19294);
or U19453 (N_19453,N_19209,N_19231);
nor U19454 (N_19454,N_19236,N_19346);
xor U19455 (N_19455,N_19207,N_19316);
xor U19456 (N_19456,N_19265,N_19317);
and U19457 (N_19457,N_19292,N_19305);
or U19458 (N_19458,N_19286,N_19231);
or U19459 (N_19459,N_19253,N_19225);
nor U19460 (N_19460,N_19231,N_19351);
and U19461 (N_19461,N_19283,N_19272);
and U19462 (N_19462,N_19230,N_19277);
xnor U19463 (N_19463,N_19244,N_19227);
xnor U19464 (N_19464,N_19201,N_19329);
and U19465 (N_19465,N_19208,N_19277);
xnor U19466 (N_19466,N_19356,N_19343);
nand U19467 (N_19467,N_19315,N_19313);
nor U19468 (N_19468,N_19295,N_19253);
nor U19469 (N_19469,N_19268,N_19308);
or U19470 (N_19470,N_19200,N_19223);
or U19471 (N_19471,N_19221,N_19283);
nor U19472 (N_19472,N_19251,N_19264);
and U19473 (N_19473,N_19214,N_19217);
or U19474 (N_19474,N_19275,N_19302);
and U19475 (N_19475,N_19338,N_19207);
xor U19476 (N_19476,N_19326,N_19278);
nor U19477 (N_19477,N_19297,N_19246);
and U19478 (N_19478,N_19304,N_19277);
nand U19479 (N_19479,N_19219,N_19261);
xor U19480 (N_19480,N_19202,N_19283);
or U19481 (N_19481,N_19283,N_19304);
nand U19482 (N_19482,N_19295,N_19241);
and U19483 (N_19483,N_19348,N_19325);
nor U19484 (N_19484,N_19269,N_19290);
and U19485 (N_19485,N_19221,N_19355);
xnor U19486 (N_19486,N_19211,N_19249);
nor U19487 (N_19487,N_19302,N_19340);
nor U19488 (N_19488,N_19343,N_19286);
and U19489 (N_19489,N_19326,N_19205);
and U19490 (N_19490,N_19322,N_19334);
or U19491 (N_19491,N_19221,N_19325);
and U19492 (N_19492,N_19276,N_19335);
nand U19493 (N_19493,N_19225,N_19335);
xor U19494 (N_19494,N_19308,N_19263);
or U19495 (N_19495,N_19341,N_19318);
xor U19496 (N_19496,N_19231,N_19305);
nand U19497 (N_19497,N_19296,N_19339);
xor U19498 (N_19498,N_19203,N_19332);
or U19499 (N_19499,N_19355,N_19354);
nand U19500 (N_19500,N_19294,N_19349);
and U19501 (N_19501,N_19204,N_19271);
or U19502 (N_19502,N_19252,N_19323);
or U19503 (N_19503,N_19238,N_19346);
xnor U19504 (N_19504,N_19300,N_19249);
and U19505 (N_19505,N_19268,N_19240);
or U19506 (N_19506,N_19279,N_19221);
or U19507 (N_19507,N_19204,N_19343);
nor U19508 (N_19508,N_19359,N_19316);
and U19509 (N_19509,N_19256,N_19298);
or U19510 (N_19510,N_19253,N_19316);
xnor U19511 (N_19511,N_19270,N_19254);
and U19512 (N_19512,N_19288,N_19220);
and U19513 (N_19513,N_19235,N_19255);
or U19514 (N_19514,N_19343,N_19346);
nand U19515 (N_19515,N_19292,N_19320);
nor U19516 (N_19516,N_19236,N_19327);
and U19517 (N_19517,N_19268,N_19327);
and U19518 (N_19518,N_19340,N_19206);
nand U19519 (N_19519,N_19288,N_19201);
xor U19520 (N_19520,N_19452,N_19412);
nor U19521 (N_19521,N_19395,N_19508);
nor U19522 (N_19522,N_19469,N_19378);
and U19523 (N_19523,N_19511,N_19403);
nor U19524 (N_19524,N_19515,N_19392);
nand U19525 (N_19525,N_19411,N_19492);
nand U19526 (N_19526,N_19414,N_19502);
nor U19527 (N_19527,N_19361,N_19484);
or U19528 (N_19528,N_19510,N_19471);
nand U19529 (N_19529,N_19419,N_19498);
nand U19530 (N_19530,N_19420,N_19401);
and U19531 (N_19531,N_19387,N_19404);
nand U19532 (N_19532,N_19421,N_19388);
and U19533 (N_19533,N_19390,N_19424);
xnor U19534 (N_19534,N_19481,N_19438);
xnor U19535 (N_19535,N_19485,N_19369);
xor U19536 (N_19536,N_19407,N_19391);
nand U19537 (N_19537,N_19368,N_19457);
and U19538 (N_19538,N_19431,N_19425);
nor U19539 (N_19539,N_19429,N_19422);
nor U19540 (N_19540,N_19513,N_19427);
xor U19541 (N_19541,N_19413,N_19479);
nand U19542 (N_19542,N_19493,N_19463);
nand U19543 (N_19543,N_19494,N_19491);
and U19544 (N_19544,N_19423,N_19503);
and U19545 (N_19545,N_19468,N_19461);
nand U19546 (N_19546,N_19384,N_19379);
nand U19547 (N_19547,N_19495,N_19381);
and U19548 (N_19548,N_19377,N_19478);
nor U19549 (N_19549,N_19464,N_19446);
nor U19550 (N_19550,N_19505,N_19436);
and U19551 (N_19551,N_19439,N_19454);
or U19552 (N_19552,N_19486,N_19488);
xnor U19553 (N_19553,N_19458,N_19451);
xnor U19554 (N_19554,N_19405,N_19385);
xnor U19555 (N_19555,N_19473,N_19466);
nand U19556 (N_19556,N_19509,N_19383);
nor U19557 (N_19557,N_19393,N_19363);
nand U19558 (N_19558,N_19366,N_19415);
and U19559 (N_19559,N_19443,N_19465);
or U19560 (N_19560,N_19449,N_19367);
nand U19561 (N_19561,N_19455,N_19459);
nor U19562 (N_19562,N_19482,N_19389);
or U19563 (N_19563,N_19432,N_19374);
nand U19564 (N_19564,N_19496,N_19402);
and U19565 (N_19565,N_19408,N_19472);
xor U19566 (N_19566,N_19376,N_19428);
xor U19567 (N_19567,N_19364,N_19409);
nand U19568 (N_19568,N_19433,N_19506);
and U19569 (N_19569,N_19489,N_19410);
nor U19570 (N_19570,N_19518,N_19483);
nor U19571 (N_19571,N_19448,N_19430);
xnor U19572 (N_19572,N_19440,N_19477);
and U19573 (N_19573,N_19514,N_19399);
nor U19574 (N_19574,N_19417,N_19370);
nor U19575 (N_19575,N_19400,N_19397);
nand U19576 (N_19576,N_19434,N_19375);
xor U19577 (N_19577,N_19362,N_19437);
and U19578 (N_19578,N_19456,N_19490);
nor U19579 (N_19579,N_19373,N_19426);
xnor U19580 (N_19580,N_19445,N_19418);
or U19581 (N_19581,N_19504,N_19453);
nand U19582 (N_19582,N_19516,N_19444);
nand U19583 (N_19583,N_19460,N_19474);
and U19584 (N_19584,N_19476,N_19450);
and U19585 (N_19585,N_19416,N_19398);
or U19586 (N_19586,N_19441,N_19365);
xor U19587 (N_19587,N_19467,N_19380);
nand U19588 (N_19588,N_19499,N_19501);
and U19589 (N_19589,N_19372,N_19442);
nand U19590 (N_19590,N_19406,N_19517);
or U19591 (N_19591,N_19386,N_19360);
nand U19592 (N_19592,N_19462,N_19512);
and U19593 (N_19593,N_19396,N_19487);
xnor U19594 (N_19594,N_19435,N_19519);
nand U19595 (N_19595,N_19497,N_19371);
nand U19596 (N_19596,N_19447,N_19480);
or U19597 (N_19597,N_19507,N_19475);
and U19598 (N_19598,N_19500,N_19382);
nand U19599 (N_19599,N_19394,N_19470);
xor U19600 (N_19600,N_19433,N_19509);
xnor U19601 (N_19601,N_19393,N_19409);
xor U19602 (N_19602,N_19511,N_19385);
xnor U19603 (N_19603,N_19418,N_19405);
xnor U19604 (N_19604,N_19493,N_19518);
xor U19605 (N_19605,N_19501,N_19428);
or U19606 (N_19606,N_19394,N_19397);
or U19607 (N_19607,N_19516,N_19367);
and U19608 (N_19608,N_19478,N_19502);
and U19609 (N_19609,N_19491,N_19514);
nand U19610 (N_19610,N_19489,N_19373);
nand U19611 (N_19611,N_19361,N_19376);
and U19612 (N_19612,N_19388,N_19483);
nand U19613 (N_19613,N_19448,N_19480);
and U19614 (N_19614,N_19424,N_19501);
and U19615 (N_19615,N_19394,N_19440);
and U19616 (N_19616,N_19472,N_19518);
nand U19617 (N_19617,N_19373,N_19416);
xor U19618 (N_19618,N_19388,N_19406);
nor U19619 (N_19619,N_19399,N_19452);
xor U19620 (N_19620,N_19455,N_19499);
or U19621 (N_19621,N_19462,N_19422);
xnor U19622 (N_19622,N_19421,N_19517);
xnor U19623 (N_19623,N_19442,N_19428);
nor U19624 (N_19624,N_19414,N_19389);
xor U19625 (N_19625,N_19393,N_19422);
nor U19626 (N_19626,N_19416,N_19417);
or U19627 (N_19627,N_19388,N_19462);
and U19628 (N_19628,N_19473,N_19382);
nand U19629 (N_19629,N_19444,N_19431);
nand U19630 (N_19630,N_19418,N_19446);
and U19631 (N_19631,N_19517,N_19503);
nor U19632 (N_19632,N_19502,N_19364);
xor U19633 (N_19633,N_19360,N_19441);
or U19634 (N_19634,N_19430,N_19438);
and U19635 (N_19635,N_19454,N_19488);
xnor U19636 (N_19636,N_19415,N_19370);
or U19637 (N_19637,N_19458,N_19476);
and U19638 (N_19638,N_19515,N_19498);
nor U19639 (N_19639,N_19473,N_19416);
or U19640 (N_19640,N_19414,N_19519);
and U19641 (N_19641,N_19424,N_19367);
xnor U19642 (N_19642,N_19444,N_19419);
nor U19643 (N_19643,N_19428,N_19440);
nand U19644 (N_19644,N_19508,N_19452);
nor U19645 (N_19645,N_19469,N_19417);
xor U19646 (N_19646,N_19369,N_19454);
and U19647 (N_19647,N_19462,N_19428);
xor U19648 (N_19648,N_19361,N_19478);
xnor U19649 (N_19649,N_19409,N_19425);
nand U19650 (N_19650,N_19436,N_19453);
nand U19651 (N_19651,N_19415,N_19411);
or U19652 (N_19652,N_19401,N_19444);
xnor U19653 (N_19653,N_19419,N_19367);
nor U19654 (N_19654,N_19380,N_19399);
or U19655 (N_19655,N_19440,N_19431);
or U19656 (N_19656,N_19460,N_19397);
xor U19657 (N_19657,N_19373,N_19504);
or U19658 (N_19658,N_19440,N_19439);
nor U19659 (N_19659,N_19417,N_19387);
nand U19660 (N_19660,N_19497,N_19393);
nor U19661 (N_19661,N_19491,N_19394);
or U19662 (N_19662,N_19435,N_19383);
and U19663 (N_19663,N_19477,N_19426);
nand U19664 (N_19664,N_19496,N_19518);
xor U19665 (N_19665,N_19485,N_19464);
or U19666 (N_19666,N_19483,N_19446);
xor U19667 (N_19667,N_19440,N_19401);
nor U19668 (N_19668,N_19384,N_19401);
nor U19669 (N_19669,N_19394,N_19487);
or U19670 (N_19670,N_19410,N_19491);
nand U19671 (N_19671,N_19459,N_19477);
nor U19672 (N_19672,N_19421,N_19419);
nand U19673 (N_19673,N_19506,N_19500);
and U19674 (N_19674,N_19431,N_19482);
or U19675 (N_19675,N_19476,N_19486);
and U19676 (N_19676,N_19481,N_19487);
or U19677 (N_19677,N_19436,N_19423);
or U19678 (N_19678,N_19488,N_19472);
and U19679 (N_19679,N_19462,N_19506);
nor U19680 (N_19680,N_19607,N_19660);
or U19681 (N_19681,N_19530,N_19652);
or U19682 (N_19682,N_19608,N_19525);
or U19683 (N_19683,N_19570,N_19628);
nand U19684 (N_19684,N_19665,N_19558);
nand U19685 (N_19685,N_19542,N_19595);
or U19686 (N_19686,N_19635,N_19528);
xnor U19687 (N_19687,N_19675,N_19648);
nor U19688 (N_19688,N_19526,N_19537);
or U19689 (N_19689,N_19644,N_19611);
and U19690 (N_19690,N_19671,N_19565);
nand U19691 (N_19691,N_19610,N_19645);
nand U19692 (N_19692,N_19641,N_19549);
nor U19693 (N_19693,N_19605,N_19544);
nand U19694 (N_19694,N_19560,N_19657);
xnor U19695 (N_19695,N_19620,N_19541);
or U19696 (N_19696,N_19543,N_19545);
nand U19697 (N_19697,N_19520,N_19661);
xnor U19698 (N_19698,N_19677,N_19667);
or U19699 (N_19699,N_19574,N_19532);
nor U19700 (N_19700,N_19581,N_19650);
nor U19701 (N_19701,N_19594,N_19668);
nor U19702 (N_19702,N_19552,N_19625);
or U19703 (N_19703,N_19531,N_19533);
and U19704 (N_19704,N_19658,N_19592);
nand U19705 (N_19705,N_19673,N_19632);
nor U19706 (N_19706,N_19554,N_19584);
nor U19707 (N_19707,N_19521,N_19578);
xor U19708 (N_19708,N_19567,N_19550);
xor U19709 (N_19709,N_19599,N_19672);
xor U19710 (N_19710,N_19575,N_19583);
nor U19711 (N_19711,N_19571,N_19534);
nand U19712 (N_19712,N_19585,N_19612);
nand U19713 (N_19713,N_19564,N_19591);
nor U19714 (N_19714,N_19636,N_19539);
xor U19715 (N_19715,N_19676,N_19639);
or U19716 (N_19716,N_19664,N_19629);
nand U19717 (N_19717,N_19559,N_19582);
xnor U19718 (N_19718,N_19656,N_19623);
or U19719 (N_19719,N_19662,N_19535);
or U19720 (N_19720,N_19524,N_19615);
nor U19721 (N_19721,N_19569,N_19654);
xor U19722 (N_19722,N_19630,N_19556);
nor U19723 (N_19723,N_19631,N_19638);
xnor U19724 (N_19724,N_19646,N_19572);
nand U19725 (N_19725,N_19562,N_19555);
nand U19726 (N_19726,N_19557,N_19643);
or U19727 (N_19727,N_19653,N_19568);
nand U19728 (N_19728,N_19566,N_19598);
nand U19729 (N_19729,N_19621,N_19538);
xor U19730 (N_19730,N_19593,N_19600);
nand U19731 (N_19731,N_19602,N_19573);
or U19732 (N_19732,N_19640,N_19655);
or U19733 (N_19733,N_19561,N_19637);
xor U19734 (N_19734,N_19527,N_19576);
xnor U19735 (N_19735,N_19597,N_19669);
xnor U19736 (N_19736,N_19522,N_19619);
nor U19737 (N_19737,N_19553,N_19614);
xnor U19738 (N_19738,N_19586,N_19659);
xnor U19739 (N_19739,N_19551,N_19523);
nand U19740 (N_19740,N_19678,N_19587);
nor U19741 (N_19741,N_19617,N_19589);
and U19742 (N_19742,N_19626,N_19624);
or U19743 (N_19743,N_19546,N_19579);
or U19744 (N_19744,N_19647,N_19601);
xnor U19745 (N_19745,N_19606,N_19577);
nand U19746 (N_19746,N_19588,N_19666);
and U19747 (N_19747,N_19540,N_19649);
and U19748 (N_19748,N_19609,N_19651);
nor U19749 (N_19749,N_19670,N_19618);
nor U19750 (N_19750,N_19679,N_19663);
and U19751 (N_19751,N_19580,N_19674);
and U19752 (N_19752,N_19622,N_19634);
or U19753 (N_19753,N_19590,N_19536);
or U19754 (N_19754,N_19633,N_19596);
nand U19755 (N_19755,N_19613,N_19563);
and U19756 (N_19756,N_19642,N_19548);
or U19757 (N_19757,N_19616,N_19627);
nand U19758 (N_19758,N_19547,N_19603);
or U19759 (N_19759,N_19529,N_19604);
nand U19760 (N_19760,N_19583,N_19663);
nand U19761 (N_19761,N_19539,N_19635);
nor U19762 (N_19762,N_19660,N_19584);
nor U19763 (N_19763,N_19649,N_19663);
nand U19764 (N_19764,N_19567,N_19589);
and U19765 (N_19765,N_19659,N_19656);
nor U19766 (N_19766,N_19663,N_19550);
and U19767 (N_19767,N_19575,N_19660);
or U19768 (N_19768,N_19571,N_19589);
and U19769 (N_19769,N_19559,N_19629);
or U19770 (N_19770,N_19571,N_19537);
xor U19771 (N_19771,N_19577,N_19639);
and U19772 (N_19772,N_19565,N_19676);
nor U19773 (N_19773,N_19597,N_19555);
and U19774 (N_19774,N_19548,N_19619);
nor U19775 (N_19775,N_19580,N_19597);
nand U19776 (N_19776,N_19574,N_19592);
or U19777 (N_19777,N_19557,N_19548);
or U19778 (N_19778,N_19564,N_19629);
xor U19779 (N_19779,N_19565,N_19585);
and U19780 (N_19780,N_19668,N_19522);
and U19781 (N_19781,N_19631,N_19556);
nand U19782 (N_19782,N_19637,N_19668);
nand U19783 (N_19783,N_19631,N_19590);
nor U19784 (N_19784,N_19633,N_19584);
nand U19785 (N_19785,N_19522,N_19664);
xor U19786 (N_19786,N_19640,N_19636);
or U19787 (N_19787,N_19576,N_19594);
or U19788 (N_19788,N_19657,N_19592);
xor U19789 (N_19789,N_19574,N_19593);
or U19790 (N_19790,N_19632,N_19597);
or U19791 (N_19791,N_19641,N_19617);
xnor U19792 (N_19792,N_19590,N_19544);
or U19793 (N_19793,N_19618,N_19608);
nor U19794 (N_19794,N_19546,N_19663);
nor U19795 (N_19795,N_19572,N_19641);
xor U19796 (N_19796,N_19614,N_19670);
nor U19797 (N_19797,N_19523,N_19596);
nand U19798 (N_19798,N_19610,N_19677);
and U19799 (N_19799,N_19651,N_19673);
and U19800 (N_19800,N_19602,N_19619);
nand U19801 (N_19801,N_19628,N_19632);
nor U19802 (N_19802,N_19602,N_19607);
or U19803 (N_19803,N_19539,N_19656);
xnor U19804 (N_19804,N_19667,N_19623);
nor U19805 (N_19805,N_19537,N_19599);
nor U19806 (N_19806,N_19677,N_19617);
nand U19807 (N_19807,N_19625,N_19609);
xnor U19808 (N_19808,N_19604,N_19542);
xor U19809 (N_19809,N_19661,N_19668);
xnor U19810 (N_19810,N_19620,N_19522);
xor U19811 (N_19811,N_19619,N_19577);
xor U19812 (N_19812,N_19578,N_19676);
or U19813 (N_19813,N_19617,N_19660);
and U19814 (N_19814,N_19603,N_19542);
nor U19815 (N_19815,N_19595,N_19523);
and U19816 (N_19816,N_19564,N_19601);
or U19817 (N_19817,N_19644,N_19622);
and U19818 (N_19818,N_19592,N_19537);
xor U19819 (N_19819,N_19626,N_19621);
nand U19820 (N_19820,N_19606,N_19562);
xnor U19821 (N_19821,N_19583,N_19528);
or U19822 (N_19822,N_19642,N_19597);
or U19823 (N_19823,N_19673,N_19659);
or U19824 (N_19824,N_19619,N_19585);
nand U19825 (N_19825,N_19642,N_19591);
nor U19826 (N_19826,N_19637,N_19599);
or U19827 (N_19827,N_19669,N_19585);
nor U19828 (N_19828,N_19594,N_19631);
nand U19829 (N_19829,N_19570,N_19529);
nand U19830 (N_19830,N_19649,N_19608);
nand U19831 (N_19831,N_19564,N_19577);
or U19832 (N_19832,N_19585,N_19529);
nor U19833 (N_19833,N_19651,N_19643);
nor U19834 (N_19834,N_19639,N_19567);
nand U19835 (N_19835,N_19537,N_19521);
or U19836 (N_19836,N_19616,N_19549);
and U19837 (N_19837,N_19544,N_19641);
xnor U19838 (N_19838,N_19589,N_19677);
nand U19839 (N_19839,N_19545,N_19537);
or U19840 (N_19840,N_19832,N_19826);
xnor U19841 (N_19841,N_19717,N_19827);
xnor U19842 (N_19842,N_19810,N_19735);
xnor U19843 (N_19843,N_19798,N_19799);
nor U19844 (N_19844,N_19745,N_19834);
and U19845 (N_19845,N_19707,N_19777);
nand U19846 (N_19846,N_19728,N_19782);
nand U19847 (N_19847,N_19775,N_19738);
xnor U19848 (N_19848,N_19816,N_19751);
xnor U19849 (N_19849,N_19822,N_19756);
nor U19850 (N_19850,N_19807,N_19757);
nor U19851 (N_19851,N_19763,N_19715);
nor U19852 (N_19852,N_19802,N_19733);
or U19853 (N_19853,N_19831,N_19772);
nor U19854 (N_19854,N_19811,N_19731);
nor U19855 (N_19855,N_19712,N_19683);
nor U19856 (N_19856,N_19760,N_19783);
xnor U19857 (N_19857,N_19706,N_19836);
nand U19858 (N_19858,N_19698,N_19781);
and U19859 (N_19859,N_19729,N_19721);
xor U19860 (N_19860,N_19696,N_19752);
and U19861 (N_19861,N_19795,N_19746);
nor U19862 (N_19862,N_19703,N_19797);
nand U19863 (N_19863,N_19766,N_19803);
nand U19864 (N_19864,N_19820,N_19688);
xnor U19865 (N_19865,N_19743,N_19689);
nor U19866 (N_19866,N_19699,N_19747);
xnor U19867 (N_19867,N_19788,N_19771);
and U19868 (N_19868,N_19705,N_19749);
xnor U19869 (N_19869,N_19837,N_19785);
or U19870 (N_19870,N_19690,N_19710);
nor U19871 (N_19871,N_19794,N_19817);
or U19872 (N_19872,N_19693,N_19830);
nand U19873 (N_19873,N_19769,N_19708);
nor U19874 (N_19874,N_19818,N_19790);
nand U19875 (N_19875,N_19814,N_19744);
or U19876 (N_19876,N_19838,N_19704);
nor U19877 (N_19877,N_19724,N_19716);
and U19878 (N_19878,N_19692,N_19714);
or U19879 (N_19879,N_19806,N_19687);
nor U19880 (N_19880,N_19736,N_19718);
and U19881 (N_19881,N_19713,N_19813);
nand U19882 (N_19882,N_19700,N_19789);
and U19883 (N_19883,N_19737,N_19694);
or U19884 (N_19884,N_19739,N_19725);
xnor U19885 (N_19885,N_19800,N_19796);
and U19886 (N_19886,N_19759,N_19768);
or U19887 (N_19887,N_19748,N_19730);
nand U19888 (N_19888,N_19740,N_19770);
xnor U19889 (N_19889,N_19753,N_19819);
nor U19890 (N_19890,N_19758,N_19824);
nor U19891 (N_19891,N_19711,N_19825);
and U19892 (N_19892,N_19821,N_19726);
nand U19893 (N_19893,N_19754,N_19686);
or U19894 (N_19894,N_19742,N_19681);
xor U19895 (N_19895,N_19767,N_19815);
and U19896 (N_19896,N_19808,N_19761);
nor U19897 (N_19897,N_19701,N_19773);
or U19898 (N_19898,N_19829,N_19702);
nand U19899 (N_19899,N_19764,N_19684);
nor U19900 (N_19900,N_19750,N_19695);
xor U19901 (N_19901,N_19709,N_19734);
or U19902 (N_19902,N_19828,N_19755);
xnor U19903 (N_19903,N_19685,N_19787);
nor U19904 (N_19904,N_19723,N_19805);
or U19905 (N_19905,N_19776,N_19780);
nand U19906 (N_19906,N_19697,N_19741);
xor U19907 (N_19907,N_19784,N_19792);
xnor U19908 (N_19908,N_19680,N_19833);
xnor U19909 (N_19909,N_19719,N_19793);
xor U19910 (N_19910,N_19809,N_19812);
xnor U19911 (N_19911,N_19691,N_19722);
nand U19912 (N_19912,N_19804,N_19774);
xnor U19913 (N_19913,N_19778,N_19765);
xnor U19914 (N_19914,N_19839,N_19801);
nor U19915 (N_19915,N_19762,N_19786);
nand U19916 (N_19916,N_19682,N_19727);
xnor U19917 (N_19917,N_19823,N_19720);
and U19918 (N_19918,N_19835,N_19779);
or U19919 (N_19919,N_19732,N_19791);
and U19920 (N_19920,N_19733,N_19747);
and U19921 (N_19921,N_19787,N_19753);
xnor U19922 (N_19922,N_19680,N_19723);
or U19923 (N_19923,N_19778,N_19698);
nand U19924 (N_19924,N_19701,N_19791);
xor U19925 (N_19925,N_19761,N_19697);
or U19926 (N_19926,N_19799,N_19833);
or U19927 (N_19927,N_19697,N_19831);
xor U19928 (N_19928,N_19783,N_19779);
nand U19929 (N_19929,N_19779,N_19706);
and U19930 (N_19930,N_19779,N_19742);
and U19931 (N_19931,N_19735,N_19785);
or U19932 (N_19932,N_19731,N_19807);
xor U19933 (N_19933,N_19705,N_19824);
xnor U19934 (N_19934,N_19720,N_19701);
and U19935 (N_19935,N_19685,N_19698);
or U19936 (N_19936,N_19787,N_19684);
nand U19937 (N_19937,N_19757,N_19768);
xor U19938 (N_19938,N_19766,N_19789);
xor U19939 (N_19939,N_19681,N_19772);
or U19940 (N_19940,N_19754,N_19715);
or U19941 (N_19941,N_19693,N_19776);
nand U19942 (N_19942,N_19733,N_19777);
or U19943 (N_19943,N_19780,N_19812);
xor U19944 (N_19944,N_19700,N_19814);
xor U19945 (N_19945,N_19827,N_19784);
nor U19946 (N_19946,N_19705,N_19683);
and U19947 (N_19947,N_19697,N_19810);
and U19948 (N_19948,N_19793,N_19739);
and U19949 (N_19949,N_19805,N_19834);
xnor U19950 (N_19950,N_19752,N_19749);
nor U19951 (N_19951,N_19732,N_19716);
and U19952 (N_19952,N_19711,N_19788);
nand U19953 (N_19953,N_19833,N_19721);
nand U19954 (N_19954,N_19687,N_19816);
xor U19955 (N_19955,N_19693,N_19821);
nor U19956 (N_19956,N_19765,N_19825);
and U19957 (N_19957,N_19805,N_19687);
xnor U19958 (N_19958,N_19800,N_19695);
or U19959 (N_19959,N_19791,N_19804);
xor U19960 (N_19960,N_19711,N_19757);
and U19961 (N_19961,N_19695,N_19802);
or U19962 (N_19962,N_19776,N_19753);
and U19963 (N_19963,N_19803,N_19741);
or U19964 (N_19964,N_19764,N_19720);
xor U19965 (N_19965,N_19693,N_19777);
or U19966 (N_19966,N_19820,N_19702);
or U19967 (N_19967,N_19725,N_19832);
or U19968 (N_19968,N_19754,N_19832);
xor U19969 (N_19969,N_19714,N_19839);
xnor U19970 (N_19970,N_19835,N_19838);
xor U19971 (N_19971,N_19717,N_19805);
nand U19972 (N_19972,N_19736,N_19814);
and U19973 (N_19973,N_19732,N_19727);
nand U19974 (N_19974,N_19812,N_19726);
or U19975 (N_19975,N_19796,N_19834);
nand U19976 (N_19976,N_19714,N_19732);
nand U19977 (N_19977,N_19806,N_19814);
and U19978 (N_19978,N_19823,N_19824);
and U19979 (N_19979,N_19811,N_19702);
nor U19980 (N_19980,N_19798,N_19808);
xnor U19981 (N_19981,N_19770,N_19788);
and U19982 (N_19982,N_19712,N_19834);
nor U19983 (N_19983,N_19778,N_19732);
nand U19984 (N_19984,N_19750,N_19811);
nor U19985 (N_19985,N_19680,N_19683);
nand U19986 (N_19986,N_19834,N_19765);
nor U19987 (N_19987,N_19824,N_19813);
or U19988 (N_19988,N_19726,N_19746);
nor U19989 (N_19989,N_19732,N_19689);
and U19990 (N_19990,N_19822,N_19798);
nor U19991 (N_19991,N_19744,N_19767);
xnor U19992 (N_19992,N_19791,N_19683);
nor U19993 (N_19993,N_19828,N_19826);
or U19994 (N_19994,N_19729,N_19764);
and U19995 (N_19995,N_19815,N_19818);
and U19996 (N_19996,N_19707,N_19724);
and U19997 (N_19997,N_19691,N_19696);
xnor U19998 (N_19998,N_19796,N_19830);
nor U19999 (N_19999,N_19830,N_19825);
nand UO_0 (O_0,N_19969,N_19928);
nand UO_1 (O_1,N_19985,N_19997);
or UO_2 (O_2,N_19879,N_19858);
or UO_3 (O_3,N_19899,N_19945);
or UO_4 (O_4,N_19937,N_19894);
nand UO_5 (O_5,N_19848,N_19860);
xor UO_6 (O_6,N_19962,N_19992);
xor UO_7 (O_7,N_19942,N_19993);
and UO_8 (O_8,N_19967,N_19966);
and UO_9 (O_9,N_19973,N_19947);
or UO_10 (O_10,N_19949,N_19955);
or UO_11 (O_11,N_19850,N_19878);
or UO_12 (O_12,N_19911,N_19913);
nor UO_13 (O_13,N_19920,N_19882);
nor UO_14 (O_14,N_19953,N_19853);
or UO_15 (O_15,N_19995,N_19988);
nand UO_16 (O_16,N_19972,N_19940);
and UO_17 (O_17,N_19999,N_19975);
and UO_18 (O_18,N_19867,N_19871);
xnor UO_19 (O_19,N_19873,N_19888);
nor UO_20 (O_20,N_19959,N_19932);
xor UO_21 (O_21,N_19880,N_19885);
or UO_22 (O_22,N_19883,N_19840);
or UO_23 (O_23,N_19986,N_19857);
xor UO_24 (O_24,N_19989,N_19896);
nor UO_25 (O_25,N_19842,N_19902);
or UO_26 (O_26,N_19977,N_19892);
or UO_27 (O_27,N_19889,N_19951);
xor UO_28 (O_28,N_19960,N_19968);
nand UO_29 (O_29,N_19930,N_19861);
nand UO_30 (O_30,N_19965,N_19874);
nand UO_31 (O_31,N_19983,N_19907);
or UO_32 (O_32,N_19895,N_19897);
nor UO_33 (O_33,N_19869,N_19927);
xnor UO_34 (O_34,N_19870,N_19944);
or UO_35 (O_35,N_19923,N_19996);
nand UO_36 (O_36,N_19938,N_19991);
nand UO_37 (O_37,N_19964,N_19963);
nand UO_38 (O_38,N_19990,N_19909);
nor UO_39 (O_39,N_19931,N_19979);
nand UO_40 (O_40,N_19906,N_19844);
and UO_41 (O_41,N_19854,N_19961);
xor UO_42 (O_42,N_19987,N_19946);
nand UO_43 (O_43,N_19903,N_19865);
nand UO_44 (O_44,N_19957,N_19912);
and UO_45 (O_45,N_19855,N_19981);
nor UO_46 (O_46,N_19916,N_19877);
xor UO_47 (O_47,N_19971,N_19856);
and UO_48 (O_48,N_19956,N_19875);
and UO_49 (O_49,N_19954,N_19939);
nor UO_50 (O_50,N_19970,N_19925);
xnor UO_51 (O_51,N_19893,N_19978);
or UO_52 (O_52,N_19851,N_19926);
or UO_53 (O_53,N_19864,N_19974);
nor UO_54 (O_54,N_19859,N_19886);
and UO_55 (O_55,N_19845,N_19862);
nor UO_56 (O_56,N_19900,N_19918);
nand UO_57 (O_57,N_19872,N_19982);
nor UO_58 (O_58,N_19922,N_19881);
nand UO_59 (O_59,N_19921,N_19948);
nand UO_60 (O_60,N_19905,N_19976);
xnor UO_61 (O_61,N_19958,N_19950);
and UO_62 (O_62,N_19904,N_19924);
nor UO_63 (O_63,N_19887,N_19915);
nand UO_64 (O_64,N_19941,N_19943);
nor UO_65 (O_65,N_19884,N_19934);
and UO_66 (O_66,N_19852,N_19863);
or UO_67 (O_67,N_19843,N_19917);
nor UO_68 (O_68,N_19846,N_19908);
nand UO_69 (O_69,N_19876,N_19935);
and UO_70 (O_70,N_19933,N_19929);
or UO_71 (O_71,N_19994,N_19984);
xnor UO_72 (O_72,N_19866,N_19952);
xnor UO_73 (O_73,N_19901,N_19980);
or UO_74 (O_74,N_19841,N_19891);
nand UO_75 (O_75,N_19998,N_19847);
and UO_76 (O_76,N_19910,N_19849);
and UO_77 (O_77,N_19890,N_19914);
nand UO_78 (O_78,N_19868,N_19919);
nor UO_79 (O_79,N_19936,N_19898);
or UO_80 (O_80,N_19873,N_19891);
or UO_81 (O_81,N_19993,N_19875);
and UO_82 (O_82,N_19967,N_19979);
nor UO_83 (O_83,N_19845,N_19940);
nand UO_84 (O_84,N_19853,N_19994);
and UO_85 (O_85,N_19845,N_19914);
nor UO_86 (O_86,N_19846,N_19979);
xor UO_87 (O_87,N_19843,N_19912);
nor UO_88 (O_88,N_19957,N_19876);
xnor UO_89 (O_89,N_19999,N_19902);
and UO_90 (O_90,N_19964,N_19865);
and UO_91 (O_91,N_19934,N_19938);
nor UO_92 (O_92,N_19866,N_19916);
and UO_93 (O_93,N_19840,N_19862);
xnor UO_94 (O_94,N_19996,N_19865);
and UO_95 (O_95,N_19860,N_19855);
nand UO_96 (O_96,N_19871,N_19912);
and UO_97 (O_97,N_19918,N_19894);
or UO_98 (O_98,N_19964,N_19993);
and UO_99 (O_99,N_19963,N_19842);
xor UO_100 (O_100,N_19884,N_19885);
or UO_101 (O_101,N_19943,N_19949);
xor UO_102 (O_102,N_19849,N_19992);
nand UO_103 (O_103,N_19905,N_19855);
nor UO_104 (O_104,N_19861,N_19981);
or UO_105 (O_105,N_19883,N_19872);
nand UO_106 (O_106,N_19949,N_19876);
xnor UO_107 (O_107,N_19988,N_19940);
nand UO_108 (O_108,N_19867,N_19977);
or UO_109 (O_109,N_19905,N_19925);
nor UO_110 (O_110,N_19868,N_19996);
nor UO_111 (O_111,N_19885,N_19866);
and UO_112 (O_112,N_19874,N_19883);
nand UO_113 (O_113,N_19951,N_19987);
nand UO_114 (O_114,N_19924,N_19956);
or UO_115 (O_115,N_19964,N_19909);
nor UO_116 (O_116,N_19931,N_19986);
nor UO_117 (O_117,N_19845,N_19962);
and UO_118 (O_118,N_19852,N_19961);
nor UO_119 (O_119,N_19899,N_19886);
nor UO_120 (O_120,N_19956,N_19976);
nand UO_121 (O_121,N_19994,N_19980);
nand UO_122 (O_122,N_19996,N_19903);
xor UO_123 (O_123,N_19927,N_19969);
and UO_124 (O_124,N_19917,N_19887);
nand UO_125 (O_125,N_19985,N_19946);
nand UO_126 (O_126,N_19888,N_19851);
nand UO_127 (O_127,N_19884,N_19978);
xor UO_128 (O_128,N_19934,N_19966);
and UO_129 (O_129,N_19961,N_19934);
or UO_130 (O_130,N_19871,N_19859);
nor UO_131 (O_131,N_19932,N_19843);
xor UO_132 (O_132,N_19950,N_19845);
nor UO_133 (O_133,N_19908,N_19857);
nand UO_134 (O_134,N_19935,N_19860);
xnor UO_135 (O_135,N_19899,N_19936);
xnor UO_136 (O_136,N_19853,N_19979);
xor UO_137 (O_137,N_19889,N_19963);
or UO_138 (O_138,N_19903,N_19986);
xnor UO_139 (O_139,N_19866,N_19951);
nand UO_140 (O_140,N_19964,N_19863);
nand UO_141 (O_141,N_19985,N_19973);
xnor UO_142 (O_142,N_19876,N_19842);
and UO_143 (O_143,N_19983,N_19863);
or UO_144 (O_144,N_19911,N_19925);
nand UO_145 (O_145,N_19863,N_19944);
xor UO_146 (O_146,N_19846,N_19926);
nand UO_147 (O_147,N_19913,N_19984);
xor UO_148 (O_148,N_19889,N_19859);
and UO_149 (O_149,N_19918,N_19965);
xor UO_150 (O_150,N_19929,N_19854);
and UO_151 (O_151,N_19884,N_19962);
or UO_152 (O_152,N_19855,N_19959);
nor UO_153 (O_153,N_19846,N_19929);
and UO_154 (O_154,N_19905,N_19848);
xnor UO_155 (O_155,N_19941,N_19870);
nand UO_156 (O_156,N_19844,N_19941);
xor UO_157 (O_157,N_19921,N_19846);
or UO_158 (O_158,N_19948,N_19856);
nor UO_159 (O_159,N_19847,N_19889);
xnor UO_160 (O_160,N_19929,N_19989);
nor UO_161 (O_161,N_19982,N_19854);
xor UO_162 (O_162,N_19953,N_19954);
nor UO_163 (O_163,N_19983,N_19867);
xor UO_164 (O_164,N_19850,N_19950);
or UO_165 (O_165,N_19904,N_19909);
nor UO_166 (O_166,N_19944,N_19886);
xnor UO_167 (O_167,N_19865,N_19919);
nor UO_168 (O_168,N_19915,N_19922);
nor UO_169 (O_169,N_19951,N_19991);
nor UO_170 (O_170,N_19847,N_19869);
or UO_171 (O_171,N_19856,N_19923);
nor UO_172 (O_172,N_19968,N_19882);
nand UO_173 (O_173,N_19995,N_19985);
nand UO_174 (O_174,N_19868,N_19915);
and UO_175 (O_175,N_19919,N_19876);
nand UO_176 (O_176,N_19971,N_19877);
and UO_177 (O_177,N_19840,N_19869);
or UO_178 (O_178,N_19852,N_19926);
nand UO_179 (O_179,N_19856,N_19913);
or UO_180 (O_180,N_19893,N_19931);
or UO_181 (O_181,N_19849,N_19883);
and UO_182 (O_182,N_19849,N_19892);
nor UO_183 (O_183,N_19954,N_19846);
xor UO_184 (O_184,N_19855,N_19849);
xnor UO_185 (O_185,N_19906,N_19864);
nand UO_186 (O_186,N_19969,N_19995);
nand UO_187 (O_187,N_19973,N_19962);
nor UO_188 (O_188,N_19929,N_19922);
nand UO_189 (O_189,N_19871,N_19895);
xnor UO_190 (O_190,N_19902,N_19847);
nor UO_191 (O_191,N_19932,N_19926);
and UO_192 (O_192,N_19891,N_19865);
and UO_193 (O_193,N_19962,N_19891);
nor UO_194 (O_194,N_19860,N_19842);
nand UO_195 (O_195,N_19862,N_19934);
nand UO_196 (O_196,N_19912,N_19964);
and UO_197 (O_197,N_19875,N_19997);
nand UO_198 (O_198,N_19941,N_19891);
xnor UO_199 (O_199,N_19918,N_19966);
or UO_200 (O_200,N_19959,N_19878);
or UO_201 (O_201,N_19911,N_19975);
xnor UO_202 (O_202,N_19901,N_19912);
and UO_203 (O_203,N_19919,N_19877);
or UO_204 (O_204,N_19955,N_19994);
nand UO_205 (O_205,N_19959,N_19996);
and UO_206 (O_206,N_19994,N_19986);
xor UO_207 (O_207,N_19974,N_19920);
or UO_208 (O_208,N_19854,N_19927);
nand UO_209 (O_209,N_19907,N_19865);
or UO_210 (O_210,N_19872,N_19975);
and UO_211 (O_211,N_19932,N_19994);
nor UO_212 (O_212,N_19914,N_19895);
or UO_213 (O_213,N_19920,N_19923);
nand UO_214 (O_214,N_19934,N_19947);
nor UO_215 (O_215,N_19949,N_19975);
or UO_216 (O_216,N_19889,N_19923);
and UO_217 (O_217,N_19893,N_19872);
or UO_218 (O_218,N_19852,N_19910);
nor UO_219 (O_219,N_19977,N_19936);
or UO_220 (O_220,N_19927,N_19910);
nand UO_221 (O_221,N_19894,N_19975);
or UO_222 (O_222,N_19975,N_19992);
and UO_223 (O_223,N_19971,N_19908);
and UO_224 (O_224,N_19934,N_19911);
and UO_225 (O_225,N_19975,N_19997);
nor UO_226 (O_226,N_19945,N_19846);
nor UO_227 (O_227,N_19861,N_19935);
and UO_228 (O_228,N_19875,N_19939);
and UO_229 (O_229,N_19924,N_19870);
xor UO_230 (O_230,N_19988,N_19966);
xor UO_231 (O_231,N_19975,N_19959);
and UO_232 (O_232,N_19905,N_19900);
xor UO_233 (O_233,N_19983,N_19916);
nor UO_234 (O_234,N_19923,N_19932);
xor UO_235 (O_235,N_19899,N_19859);
nor UO_236 (O_236,N_19856,N_19915);
xor UO_237 (O_237,N_19893,N_19948);
xnor UO_238 (O_238,N_19925,N_19941);
or UO_239 (O_239,N_19990,N_19892);
or UO_240 (O_240,N_19877,N_19890);
or UO_241 (O_241,N_19941,N_19942);
or UO_242 (O_242,N_19989,N_19917);
nor UO_243 (O_243,N_19879,N_19938);
xor UO_244 (O_244,N_19958,N_19867);
xnor UO_245 (O_245,N_19934,N_19856);
nor UO_246 (O_246,N_19976,N_19922);
and UO_247 (O_247,N_19963,N_19953);
nand UO_248 (O_248,N_19957,N_19971);
nand UO_249 (O_249,N_19931,N_19847);
xor UO_250 (O_250,N_19888,N_19881);
or UO_251 (O_251,N_19986,N_19874);
xnor UO_252 (O_252,N_19927,N_19944);
and UO_253 (O_253,N_19863,N_19860);
xor UO_254 (O_254,N_19963,N_19906);
and UO_255 (O_255,N_19912,N_19851);
nand UO_256 (O_256,N_19965,N_19990);
and UO_257 (O_257,N_19928,N_19917);
nor UO_258 (O_258,N_19940,N_19881);
nand UO_259 (O_259,N_19976,N_19915);
and UO_260 (O_260,N_19988,N_19893);
and UO_261 (O_261,N_19888,N_19857);
and UO_262 (O_262,N_19888,N_19981);
or UO_263 (O_263,N_19890,N_19944);
xor UO_264 (O_264,N_19944,N_19906);
nand UO_265 (O_265,N_19857,N_19860);
and UO_266 (O_266,N_19872,N_19969);
nand UO_267 (O_267,N_19856,N_19960);
or UO_268 (O_268,N_19886,N_19909);
and UO_269 (O_269,N_19936,N_19949);
or UO_270 (O_270,N_19903,N_19889);
nor UO_271 (O_271,N_19959,N_19945);
or UO_272 (O_272,N_19968,N_19852);
xnor UO_273 (O_273,N_19855,N_19867);
and UO_274 (O_274,N_19912,N_19988);
nand UO_275 (O_275,N_19891,N_19930);
and UO_276 (O_276,N_19949,N_19989);
xor UO_277 (O_277,N_19928,N_19978);
nor UO_278 (O_278,N_19943,N_19992);
xor UO_279 (O_279,N_19895,N_19841);
nor UO_280 (O_280,N_19909,N_19845);
xor UO_281 (O_281,N_19968,N_19972);
nor UO_282 (O_282,N_19974,N_19841);
and UO_283 (O_283,N_19853,N_19965);
nor UO_284 (O_284,N_19861,N_19896);
and UO_285 (O_285,N_19996,N_19891);
nor UO_286 (O_286,N_19934,N_19920);
nand UO_287 (O_287,N_19974,N_19871);
or UO_288 (O_288,N_19854,N_19926);
xor UO_289 (O_289,N_19892,N_19942);
xor UO_290 (O_290,N_19897,N_19953);
xnor UO_291 (O_291,N_19965,N_19912);
nor UO_292 (O_292,N_19935,N_19847);
nand UO_293 (O_293,N_19856,N_19975);
nor UO_294 (O_294,N_19889,N_19991);
nand UO_295 (O_295,N_19920,N_19848);
nor UO_296 (O_296,N_19883,N_19892);
and UO_297 (O_297,N_19931,N_19876);
xnor UO_298 (O_298,N_19961,N_19954);
and UO_299 (O_299,N_19981,N_19971);
or UO_300 (O_300,N_19954,N_19986);
xor UO_301 (O_301,N_19936,N_19978);
nand UO_302 (O_302,N_19886,N_19875);
nor UO_303 (O_303,N_19927,N_19980);
nor UO_304 (O_304,N_19967,N_19928);
or UO_305 (O_305,N_19876,N_19970);
xnor UO_306 (O_306,N_19976,N_19926);
or UO_307 (O_307,N_19954,N_19902);
or UO_308 (O_308,N_19989,N_19928);
and UO_309 (O_309,N_19914,N_19851);
nor UO_310 (O_310,N_19881,N_19902);
or UO_311 (O_311,N_19888,N_19897);
nand UO_312 (O_312,N_19845,N_19854);
xor UO_313 (O_313,N_19931,N_19897);
nor UO_314 (O_314,N_19919,N_19941);
xor UO_315 (O_315,N_19946,N_19896);
nor UO_316 (O_316,N_19983,N_19997);
nor UO_317 (O_317,N_19921,N_19922);
nor UO_318 (O_318,N_19988,N_19954);
nor UO_319 (O_319,N_19977,N_19864);
xor UO_320 (O_320,N_19846,N_19897);
xor UO_321 (O_321,N_19847,N_19936);
xnor UO_322 (O_322,N_19842,N_19911);
nand UO_323 (O_323,N_19968,N_19858);
xnor UO_324 (O_324,N_19879,N_19976);
nand UO_325 (O_325,N_19860,N_19950);
nand UO_326 (O_326,N_19926,N_19943);
xnor UO_327 (O_327,N_19925,N_19878);
xnor UO_328 (O_328,N_19886,N_19989);
and UO_329 (O_329,N_19989,N_19905);
or UO_330 (O_330,N_19993,N_19904);
and UO_331 (O_331,N_19920,N_19988);
or UO_332 (O_332,N_19931,N_19875);
nor UO_333 (O_333,N_19844,N_19982);
xnor UO_334 (O_334,N_19923,N_19947);
xor UO_335 (O_335,N_19843,N_19846);
nand UO_336 (O_336,N_19856,N_19843);
nor UO_337 (O_337,N_19936,N_19997);
nand UO_338 (O_338,N_19973,N_19860);
xnor UO_339 (O_339,N_19946,N_19876);
and UO_340 (O_340,N_19967,N_19941);
xnor UO_341 (O_341,N_19926,N_19965);
and UO_342 (O_342,N_19902,N_19998);
or UO_343 (O_343,N_19860,N_19890);
or UO_344 (O_344,N_19859,N_19888);
nor UO_345 (O_345,N_19951,N_19858);
nand UO_346 (O_346,N_19890,N_19874);
nand UO_347 (O_347,N_19856,N_19985);
or UO_348 (O_348,N_19854,N_19899);
nor UO_349 (O_349,N_19908,N_19909);
and UO_350 (O_350,N_19976,N_19914);
and UO_351 (O_351,N_19876,N_19894);
nand UO_352 (O_352,N_19909,N_19953);
or UO_353 (O_353,N_19844,N_19938);
nand UO_354 (O_354,N_19957,N_19906);
or UO_355 (O_355,N_19938,N_19936);
or UO_356 (O_356,N_19989,N_19892);
or UO_357 (O_357,N_19922,N_19935);
xnor UO_358 (O_358,N_19875,N_19887);
and UO_359 (O_359,N_19855,N_19858);
nand UO_360 (O_360,N_19951,N_19878);
and UO_361 (O_361,N_19845,N_19877);
xor UO_362 (O_362,N_19933,N_19915);
and UO_363 (O_363,N_19842,N_19878);
nor UO_364 (O_364,N_19944,N_19980);
nor UO_365 (O_365,N_19870,N_19890);
or UO_366 (O_366,N_19975,N_19899);
or UO_367 (O_367,N_19857,N_19913);
nor UO_368 (O_368,N_19923,N_19875);
nand UO_369 (O_369,N_19883,N_19930);
nand UO_370 (O_370,N_19866,N_19892);
and UO_371 (O_371,N_19879,N_19981);
nor UO_372 (O_372,N_19930,N_19885);
nor UO_373 (O_373,N_19882,N_19876);
xor UO_374 (O_374,N_19987,N_19998);
or UO_375 (O_375,N_19850,N_19976);
or UO_376 (O_376,N_19902,N_19858);
and UO_377 (O_377,N_19926,N_19842);
nor UO_378 (O_378,N_19990,N_19982);
nor UO_379 (O_379,N_19914,N_19977);
or UO_380 (O_380,N_19985,N_19858);
nor UO_381 (O_381,N_19965,N_19919);
or UO_382 (O_382,N_19851,N_19871);
nor UO_383 (O_383,N_19919,N_19898);
nand UO_384 (O_384,N_19888,N_19848);
or UO_385 (O_385,N_19928,N_19921);
or UO_386 (O_386,N_19931,N_19862);
xnor UO_387 (O_387,N_19980,N_19849);
or UO_388 (O_388,N_19982,N_19963);
and UO_389 (O_389,N_19991,N_19882);
nand UO_390 (O_390,N_19853,N_19887);
or UO_391 (O_391,N_19871,N_19978);
nand UO_392 (O_392,N_19915,N_19934);
nor UO_393 (O_393,N_19923,N_19931);
nor UO_394 (O_394,N_19924,N_19926);
or UO_395 (O_395,N_19980,N_19920);
nand UO_396 (O_396,N_19961,N_19981);
xnor UO_397 (O_397,N_19959,N_19892);
xnor UO_398 (O_398,N_19864,N_19924);
xnor UO_399 (O_399,N_19911,N_19974);
xnor UO_400 (O_400,N_19996,N_19984);
nand UO_401 (O_401,N_19931,N_19991);
and UO_402 (O_402,N_19896,N_19957);
and UO_403 (O_403,N_19958,N_19880);
xor UO_404 (O_404,N_19987,N_19960);
xnor UO_405 (O_405,N_19932,N_19976);
nand UO_406 (O_406,N_19870,N_19878);
or UO_407 (O_407,N_19979,N_19915);
and UO_408 (O_408,N_19969,N_19967);
nand UO_409 (O_409,N_19906,N_19940);
and UO_410 (O_410,N_19853,N_19926);
or UO_411 (O_411,N_19960,N_19851);
and UO_412 (O_412,N_19973,N_19954);
nand UO_413 (O_413,N_19875,N_19911);
nand UO_414 (O_414,N_19908,N_19933);
or UO_415 (O_415,N_19993,N_19892);
or UO_416 (O_416,N_19848,N_19929);
and UO_417 (O_417,N_19840,N_19863);
and UO_418 (O_418,N_19996,N_19949);
or UO_419 (O_419,N_19863,N_19958);
xor UO_420 (O_420,N_19938,N_19976);
xor UO_421 (O_421,N_19905,N_19997);
nand UO_422 (O_422,N_19936,N_19942);
and UO_423 (O_423,N_19926,N_19923);
nand UO_424 (O_424,N_19922,N_19864);
or UO_425 (O_425,N_19900,N_19997);
xnor UO_426 (O_426,N_19852,N_19953);
xor UO_427 (O_427,N_19937,N_19884);
or UO_428 (O_428,N_19875,N_19965);
and UO_429 (O_429,N_19884,N_19996);
or UO_430 (O_430,N_19987,N_19986);
nand UO_431 (O_431,N_19951,N_19975);
and UO_432 (O_432,N_19961,N_19918);
nor UO_433 (O_433,N_19841,N_19993);
nand UO_434 (O_434,N_19910,N_19998);
nor UO_435 (O_435,N_19993,N_19972);
nor UO_436 (O_436,N_19856,N_19957);
and UO_437 (O_437,N_19879,N_19965);
xnor UO_438 (O_438,N_19851,N_19884);
and UO_439 (O_439,N_19852,N_19908);
xor UO_440 (O_440,N_19916,N_19862);
and UO_441 (O_441,N_19845,N_19976);
and UO_442 (O_442,N_19856,N_19855);
and UO_443 (O_443,N_19964,N_19926);
and UO_444 (O_444,N_19931,N_19973);
and UO_445 (O_445,N_19842,N_19922);
or UO_446 (O_446,N_19928,N_19954);
nand UO_447 (O_447,N_19862,N_19881);
nor UO_448 (O_448,N_19899,N_19979);
nand UO_449 (O_449,N_19903,N_19968);
xor UO_450 (O_450,N_19965,N_19868);
nand UO_451 (O_451,N_19914,N_19978);
or UO_452 (O_452,N_19887,N_19981);
nor UO_453 (O_453,N_19953,N_19955);
and UO_454 (O_454,N_19944,N_19952);
nand UO_455 (O_455,N_19897,N_19993);
xor UO_456 (O_456,N_19915,N_19997);
nor UO_457 (O_457,N_19926,N_19949);
or UO_458 (O_458,N_19889,N_19973);
or UO_459 (O_459,N_19872,N_19964);
nor UO_460 (O_460,N_19943,N_19852);
xnor UO_461 (O_461,N_19948,N_19851);
nor UO_462 (O_462,N_19896,N_19948);
and UO_463 (O_463,N_19951,N_19977);
xnor UO_464 (O_464,N_19942,N_19900);
xor UO_465 (O_465,N_19956,N_19860);
or UO_466 (O_466,N_19939,N_19879);
xnor UO_467 (O_467,N_19926,N_19909);
or UO_468 (O_468,N_19869,N_19970);
and UO_469 (O_469,N_19959,N_19901);
nand UO_470 (O_470,N_19840,N_19907);
and UO_471 (O_471,N_19931,N_19902);
nand UO_472 (O_472,N_19860,N_19968);
xor UO_473 (O_473,N_19843,N_19980);
nor UO_474 (O_474,N_19992,N_19852);
xor UO_475 (O_475,N_19894,N_19860);
or UO_476 (O_476,N_19924,N_19900);
xnor UO_477 (O_477,N_19972,N_19912);
or UO_478 (O_478,N_19859,N_19840);
and UO_479 (O_479,N_19848,N_19935);
nand UO_480 (O_480,N_19860,N_19959);
xnor UO_481 (O_481,N_19880,N_19875);
nand UO_482 (O_482,N_19973,N_19981);
xor UO_483 (O_483,N_19940,N_19937);
or UO_484 (O_484,N_19977,N_19863);
nor UO_485 (O_485,N_19930,N_19860);
nand UO_486 (O_486,N_19987,N_19956);
nand UO_487 (O_487,N_19909,N_19916);
or UO_488 (O_488,N_19953,N_19947);
xnor UO_489 (O_489,N_19992,N_19870);
xnor UO_490 (O_490,N_19892,N_19937);
or UO_491 (O_491,N_19867,N_19961);
and UO_492 (O_492,N_19904,N_19925);
nand UO_493 (O_493,N_19906,N_19934);
nor UO_494 (O_494,N_19934,N_19921);
nor UO_495 (O_495,N_19921,N_19858);
nor UO_496 (O_496,N_19916,N_19861);
xnor UO_497 (O_497,N_19984,N_19900);
or UO_498 (O_498,N_19890,N_19861);
xnor UO_499 (O_499,N_19842,N_19875);
and UO_500 (O_500,N_19987,N_19959);
nor UO_501 (O_501,N_19860,N_19958);
or UO_502 (O_502,N_19884,N_19899);
nand UO_503 (O_503,N_19933,N_19918);
or UO_504 (O_504,N_19948,N_19994);
nor UO_505 (O_505,N_19947,N_19916);
and UO_506 (O_506,N_19847,N_19903);
and UO_507 (O_507,N_19842,N_19916);
nand UO_508 (O_508,N_19948,N_19876);
nand UO_509 (O_509,N_19971,N_19876);
nor UO_510 (O_510,N_19918,N_19872);
nand UO_511 (O_511,N_19960,N_19929);
or UO_512 (O_512,N_19865,N_19979);
nand UO_513 (O_513,N_19907,N_19970);
or UO_514 (O_514,N_19921,N_19894);
nor UO_515 (O_515,N_19986,N_19946);
nor UO_516 (O_516,N_19885,N_19959);
or UO_517 (O_517,N_19903,N_19899);
nor UO_518 (O_518,N_19913,N_19883);
xor UO_519 (O_519,N_19885,N_19982);
nand UO_520 (O_520,N_19957,N_19840);
nor UO_521 (O_521,N_19864,N_19887);
xor UO_522 (O_522,N_19853,N_19987);
nor UO_523 (O_523,N_19845,N_19896);
nor UO_524 (O_524,N_19951,N_19910);
nand UO_525 (O_525,N_19955,N_19866);
xor UO_526 (O_526,N_19960,N_19939);
xor UO_527 (O_527,N_19964,N_19984);
nor UO_528 (O_528,N_19925,N_19906);
nand UO_529 (O_529,N_19863,N_19845);
xor UO_530 (O_530,N_19994,N_19859);
nor UO_531 (O_531,N_19974,N_19847);
xnor UO_532 (O_532,N_19879,N_19842);
xor UO_533 (O_533,N_19948,N_19881);
nor UO_534 (O_534,N_19970,N_19911);
or UO_535 (O_535,N_19963,N_19862);
nand UO_536 (O_536,N_19843,N_19940);
nor UO_537 (O_537,N_19870,N_19873);
and UO_538 (O_538,N_19920,N_19856);
or UO_539 (O_539,N_19980,N_19975);
nor UO_540 (O_540,N_19883,N_19976);
or UO_541 (O_541,N_19951,N_19929);
xnor UO_542 (O_542,N_19882,N_19969);
or UO_543 (O_543,N_19993,N_19903);
nand UO_544 (O_544,N_19913,N_19841);
and UO_545 (O_545,N_19951,N_19985);
nor UO_546 (O_546,N_19877,N_19855);
or UO_547 (O_547,N_19907,N_19902);
or UO_548 (O_548,N_19849,N_19905);
nand UO_549 (O_549,N_19881,N_19864);
nand UO_550 (O_550,N_19984,N_19883);
nand UO_551 (O_551,N_19939,N_19950);
or UO_552 (O_552,N_19957,N_19955);
nor UO_553 (O_553,N_19896,N_19904);
nor UO_554 (O_554,N_19926,N_19942);
nand UO_555 (O_555,N_19998,N_19945);
xnor UO_556 (O_556,N_19961,N_19968);
nand UO_557 (O_557,N_19882,N_19905);
xor UO_558 (O_558,N_19950,N_19843);
or UO_559 (O_559,N_19997,N_19842);
or UO_560 (O_560,N_19930,N_19961);
or UO_561 (O_561,N_19872,N_19890);
xor UO_562 (O_562,N_19980,N_19961);
and UO_563 (O_563,N_19855,N_19955);
nand UO_564 (O_564,N_19886,N_19910);
nand UO_565 (O_565,N_19939,N_19889);
and UO_566 (O_566,N_19880,N_19865);
nor UO_567 (O_567,N_19913,N_19967);
or UO_568 (O_568,N_19921,N_19920);
or UO_569 (O_569,N_19978,N_19960);
nand UO_570 (O_570,N_19881,N_19966);
xor UO_571 (O_571,N_19993,N_19901);
xor UO_572 (O_572,N_19918,N_19913);
xnor UO_573 (O_573,N_19911,N_19919);
nand UO_574 (O_574,N_19858,N_19986);
nand UO_575 (O_575,N_19969,N_19860);
nor UO_576 (O_576,N_19872,N_19877);
xnor UO_577 (O_577,N_19897,N_19876);
nand UO_578 (O_578,N_19862,N_19941);
nor UO_579 (O_579,N_19908,N_19904);
nand UO_580 (O_580,N_19859,N_19950);
nand UO_581 (O_581,N_19859,N_19929);
xor UO_582 (O_582,N_19913,N_19848);
and UO_583 (O_583,N_19888,N_19964);
nand UO_584 (O_584,N_19948,N_19981);
or UO_585 (O_585,N_19986,N_19991);
xnor UO_586 (O_586,N_19856,N_19893);
nand UO_587 (O_587,N_19981,N_19847);
nor UO_588 (O_588,N_19999,N_19944);
nand UO_589 (O_589,N_19970,N_19969);
xor UO_590 (O_590,N_19860,N_19856);
and UO_591 (O_591,N_19866,N_19964);
nor UO_592 (O_592,N_19945,N_19888);
xnor UO_593 (O_593,N_19999,N_19917);
xor UO_594 (O_594,N_19907,N_19984);
and UO_595 (O_595,N_19881,N_19893);
nor UO_596 (O_596,N_19907,N_19845);
nor UO_597 (O_597,N_19980,N_19865);
nand UO_598 (O_598,N_19879,N_19882);
and UO_599 (O_599,N_19959,N_19943);
nand UO_600 (O_600,N_19997,N_19887);
nand UO_601 (O_601,N_19861,N_19860);
nor UO_602 (O_602,N_19843,N_19840);
and UO_603 (O_603,N_19863,N_19933);
xnor UO_604 (O_604,N_19994,N_19916);
and UO_605 (O_605,N_19892,N_19921);
xnor UO_606 (O_606,N_19885,N_19944);
and UO_607 (O_607,N_19842,N_19859);
nand UO_608 (O_608,N_19849,N_19891);
nor UO_609 (O_609,N_19856,N_19914);
nor UO_610 (O_610,N_19898,N_19870);
nand UO_611 (O_611,N_19980,N_19883);
nand UO_612 (O_612,N_19843,N_19849);
or UO_613 (O_613,N_19983,N_19915);
nand UO_614 (O_614,N_19902,N_19868);
nand UO_615 (O_615,N_19911,N_19954);
nand UO_616 (O_616,N_19928,N_19960);
and UO_617 (O_617,N_19911,N_19985);
and UO_618 (O_618,N_19871,N_19855);
nor UO_619 (O_619,N_19871,N_19841);
nor UO_620 (O_620,N_19988,N_19857);
nand UO_621 (O_621,N_19954,N_19847);
xor UO_622 (O_622,N_19963,N_19928);
and UO_623 (O_623,N_19976,N_19983);
or UO_624 (O_624,N_19919,N_19924);
nand UO_625 (O_625,N_19945,N_19995);
or UO_626 (O_626,N_19960,N_19841);
nor UO_627 (O_627,N_19872,N_19981);
xnor UO_628 (O_628,N_19864,N_19932);
and UO_629 (O_629,N_19970,N_19965);
or UO_630 (O_630,N_19906,N_19958);
xor UO_631 (O_631,N_19943,N_19924);
nor UO_632 (O_632,N_19974,N_19959);
and UO_633 (O_633,N_19999,N_19983);
nand UO_634 (O_634,N_19867,N_19869);
nand UO_635 (O_635,N_19889,N_19968);
nor UO_636 (O_636,N_19866,N_19886);
or UO_637 (O_637,N_19987,N_19900);
and UO_638 (O_638,N_19888,N_19874);
or UO_639 (O_639,N_19840,N_19999);
and UO_640 (O_640,N_19931,N_19858);
and UO_641 (O_641,N_19978,N_19933);
xnor UO_642 (O_642,N_19874,N_19904);
nand UO_643 (O_643,N_19947,N_19970);
and UO_644 (O_644,N_19960,N_19950);
nand UO_645 (O_645,N_19889,N_19947);
nand UO_646 (O_646,N_19875,N_19990);
nand UO_647 (O_647,N_19902,N_19993);
nor UO_648 (O_648,N_19923,N_19887);
nor UO_649 (O_649,N_19969,N_19915);
nand UO_650 (O_650,N_19996,N_19945);
or UO_651 (O_651,N_19915,N_19902);
or UO_652 (O_652,N_19920,N_19861);
and UO_653 (O_653,N_19871,N_19940);
nand UO_654 (O_654,N_19984,N_19867);
xnor UO_655 (O_655,N_19917,N_19853);
nand UO_656 (O_656,N_19869,N_19929);
and UO_657 (O_657,N_19992,N_19931);
or UO_658 (O_658,N_19998,N_19879);
and UO_659 (O_659,N_19854,N_19985);
nor UO_660 (O_660,N_19926,N_19960);
nand UO_661 (O_661,N_19953,N_19925);
nand UO_662 (O_662,N_19840,N_19866);
and UO_663 (O_663,N_19844,N_19855);
nor UO_664 (O_664,N_19908,N_19974);
nand UO_665 (O_665,N_19887,N_19849);
nor UO_666 (O_666,N_19892,N_19857);
nand UO_667 (O_667,N_19935,N_19853);
nor UO_668 (O_668,N_19886,N_19925);
xor UO_669 (O_669,N_19922,N_19875);
nand UO_670 (O_670,N_19977,N_19954);
nor UO_671 (O_671,N_19913,N_19999);
nand UO_672 (O_672,N_19960,N_19965);
and UO_673 (O_673,N_19910,N_19930);
and UO_674 (O_674,N_19937,N_19928);
nand UO_675 (O_675,N_19948,N_19995);
or UO_676 (O_676,N_19888,N_19908);
xnor UO_677 (O_677,N_19930,N_19950);
xnor UO_678 (O_678,N_19931,N_19939);
nor UO_679 (O_679,N_19842,N_19914);
or UO_680 (O_680,N_19896,N_19966);
nor UO_681 (O_681,N_19977,N_19969);
nor UO_682 (O_682,N_19884,N_19964);
and UO_683 (O_683,N_19893,N_19889);
nor UO_684 (O_684,N_19995,N_19923);
nand UO_685 (O_685,N_19929,N_19979);
xnor UO_686 (O_686,N_19865,N_19871);
xnor UO_687 (O_687,N_19923,N_19912);
xnor UO_688 (O_688,N_19991,N_19911);
nor UO_689 (O_689,N_19956,N_19843);
nor UO_690 (O_690,N_19938,N_19914);
nor UO_691 (O_691,N_19844,N_19887);
or UO_692 (O_692,N_19883,N_19842);
xor UO_693 (O_693,N_19881,N_19870);
or UO_694 (O_694,N_19950,N_19968);
or UO_695 (O_695,N_19851,N_19971);
xnor UO_696 (O_696,N_19953,N_19988);
xnor UO_697 (O_697,N_19993,N_19866);
nor UO_698 (O_698,N_19923,N_19914);
nand UO_699 (O_699,N_19874,N_19998);
xnor UO_700 (O_700,N_19904,N_19996);
xnor UO_701 (O_701,N_19980,N_19971);
nor UO_702 (O_702,N_19901,N_19937);
nor UO_703 (O_703,N_19854,N_19840);
nor UO_704 (O_704,N_19850,N_19959);
nand UO_705 (O_705,N_19963,N_19843);
and UO_706 (O_706,N_19879,N_19997);
nand UO_707 (O_707,N_19871,N_19847);
nand UO_708 (O_708,N_19848,N_19958);
xnor UO_709 (O_709,N_19951,N_19905);
nand UO_710 (O_710,N_19844,N_19868);
and UO_711 (O_711,N_19967,N_19992);
or UO_712 (O_712,N_19931,N_19859);
xnor UO_713 (O_713,N_19919,N_19847);
or UO_714 (O_714,N_19888,N_19895);
nor UO_715 (O_715,N_19900,N_19986);
nand UO_716 (O_716,N_19956,N_19906);
xor UO_717 (O_717,N_19904,N_19910);
xnor UO_718 (O_718,N_19903,N_19908);
or UO_719 (O_719,N_19960,N_19843);
or UO_720 (O_720,N_19902,N_19941);
or UO_721 (O_721,N_19860,N_19892);
and UO_722 (O_722,N_19857,N_19871);
nand UO_723 (O_723,N_19919,N_19912);
xnor UO_724 (O_724,N_19878,N_19896);
and UO_725 (O_725,N_19989,N_19969);
or UO_726 (O_726,N_19880,N_19960);
or UO_727 (O_727,N_19877,N_19880);
or UO_728 (O_728,N_19954,N_19982);
nor UO_729 (O_729,N_19889,N_19961);
nor UO_730 (O_730,N_19928,N_19905);
and UO_731 (O_731,N_19891,N_19972);
nand UO_732 (O_732,N_19955,N_19999);
xor UO_733 (O_733,N_19901,N_19893);
and UO_734 (O_734,N_19886,N_19853);
or UO_735 (O_735,N_19909,N_19971);
or UO_736 (O_736,N_19901,N_19891);
and UO_737 (O_737,N_19923,N_19901);
xnor UO_738 (O_738,N_19965,N_19867);
and UO_739 (O_739,N_19913,N_19937);
xor UO_740 (O_740,N_19887,N_19880);
or UO_741 (O_741,N_19911,N_19854);
nor UO_742 (O_742,N_19927,N_19923);
nand UO_743 (O_743,N_19905,N_19970);
nand UO_744 (O_744,N_19869,N_19999);
or UO_745 (O_745,N_19928,N_19903);
or UO_746 (O_746,N_19930,N_19863);
or UO_747 (O_747,N_19869,N_19996);
and UO_748 (O_748,N_19930,N_19858);
xor UO_749 (O_749,N_19898,N_19941);
and UO_750 (O_750,N_19920,N_19863);
xnor UO_751 (O_751,N_19868,N_19913);
or UO_752 (O_752,N_19882,N_19862);
nand UO_753 (O_753,N_19933,N_19984);
or UO_754 (O_754,N_19977,N_19990);
or UO_755 (O_755,N_19917,N_19966);
and UO_756 (O_756,N_19845,N_19915);
and UO_757 (O_757,N_19886,N_19956);
xor UO_758 (O_758,N_19845,N_19971);
nand UO_759 (O_759,N_19881,N_19894);
or UO_760 (O_760,N_19965,N_19941);
or UO_761 (O_761,N_19887,N_19952);
nor UO_762 (O_762,N_19919,N_19922);
nor UO_763 (O_763,N_19874,N_19988);
and UO_764 (O_764,N_19960,N_19936);
and UO_765 (O_765,N_19987,N_19908);
xnor UO_766 (O_766,N_19937,N_19946);
nand UO_767 (O_767,N_19977,N_19962);
nand UO_768 (O_768,N_19937,N_19895);
or UO_769 (O_769,N_19936,N_19940);
and UO_770 (O_770,N_19985,N_19981);
and UO_771 (O_771,N_19858,N_19874);
nor UO_772 (O_772,N_19945,N_19984);
and UO_773 (O_773,N_19874,N_19975);
or UO_774 (O_774,N_19950,N_19913);
nand UO_775 (O_775,N_19920,N_19841);
nor UO_776 (O_776,N_19899,N_19983);
xnor UO_777 (O_777,N_19912,N_19898);
or UO_778 (O_778,N_19973,N_19845);
or UO_779 (O_779,N_19909,N_19984);
and UO_780 (O_780,N_19968,N_19988);
or UO_781 (O_781,N_19982,N_19901);
xor UO_782 (O_782,N_19976,N_19991);
xor UO_783 (O_783,N_19896,N_19859);
nand UO_784 (O_784,N_19947,N_19968);
and UO_785 (O_785,N_19985,N_19938);
nand UO_786 (O_786,N_19972,N_19885);
nand UO_787 (O_787,N_19990,N_19950);
xnor UO_788 (O_788,N_19983,N_19892);
xor UO_789 (O_789,N_19924,N_19845);
xnor UO_790 (O_790,N_19894,N_19960);
xnor UO_791 (O_791,N_19887,N_19945);
nand UO_792 (O_792,N_19943,N_19883);
nand UO_793 (O_793,N_19974,N_19906);
nand UO_794 (O_794,N_19973,N_19858);
and UO_795 (O_795,N_19895,N_19933);
nor UO_796 (O_796,N_19965,N_19967);
xor UO_797 (O_797,N_19880,N_19987);
or UO_798 (O_798,N_19903,N_19943);
and UO_799 (O_799,N_19919,N_19870);
xnor UO_800 (O_800,N_19850,N_19881);
or UO_801 (O_801,N_19985,N_19924);
xnor UO_802 (O_802,N_19978,N_19887);
nand UO_803 (O_803,N_19946,N_19884);
nor UO_804 (O_804,N_19924,N_19967);
or UO_805 (O_805,N_19942,N_19946);
xnor UO_806 (O_806,N_19969,N_19876);
or UO_807 (O_807,N_19844,N_19926);
or UO_808 (O_808,N_19868,N_19978);
xnor UO_809 (O_809,N_19962,N_19934);
nand UO_810 (O_810,N_19939,N_19885);
nand UO_811 (O_811,N_19964,N_19907);
xnor UO_812 (O_812,N_19958,N_19857);
nand UO_813 (O_813,N_19905,N_19846);
and UO_814 (O_814,N_19865,N_19931);
or UO_815 (O_815,N_19918,N_19922);
or UO_816 (O_816,N_19918,N_19856);
or UO_817 (O_817,N_19853,N_19913);
and UO_818 (O_818,N_19932,N_19974);
nand UO_819 (O_819,N_19962,N_19982);
and UO_820 (O_820,N_19955,N_19950);
nand UO_821 (O_821,N_19929,N_19865);
nand UO_822 (O_822,N_19974,N_19894);
xnor UO_823 (O_823,N_19846,N_19906);
xor UO_824 (O_824,N_19912,N_19942);
nor UO_825 (O_825,N_19872,N_19867);
or UO_826 (O_826,N_19978,N_19859);
or UO_827 (O_827,N_19986,N_19878);
nor UO_828 (O_828,N_19910,N_19943);
xnor UO_829 (O_829,N_19841,N_19992);
nor UO_830 (O_830,N_19959,N_19953);
nand UO_831 (O_831,N_19940,N_19925);
or UO_832 (O_832,N_19931,N_19906);
or UO_833 (O_833,N_19946,N_19895);
and UO_834 (O_834,N_19888,N_19917);
xor UO_835 (O_835,N_19907,N_19941);
or UO_836 (O_836,N_19983,N_19935);
or UO_837 (O_837,N_19881,N_19843);
xor UO_838 (O_838,N_19913,N_19939);
xnor UO_839 (O_839,N_19996,N_19879);
xor UO_840 (O_840,N_19944,N_19912);
xor UO_841 (O_841,N_19930,N_19945);
and UO_842 (O_842,N_19945,N_19980);
and UO_843 (O_843,N_19973,N_19847);
and UO_844 (O_844,N_19891,N_19932);
nor UO_845 (O_845,N_19915,N_19861);
xnor UO_846 (O_846,N_19850,N_19871);
xor UO_847 (O_847,N_19985,N_19869);
nor UO_848 (O_848,N_19866,N_19872);
nor UO_849 (O_849,N_19877,N_19928);
and UO_850 (O_850,N_19852,N_19931);
nor UO_851 (O_851,N_19840,N_19846);
nand UO_852 (O_852,N_19898,N_19984);
and UO_853 (O_853,N_19855,N_19882);
xnor UO_854 (O_854,N_19948,N_19933);
or UO_855 (O_855,N_19997,N_19857);
nor UO_856 (O_856,N_19926,N_19874);
nand UO_857 (O_857,N_19927,N_19992);
or UO_858 (O_858,N_19849,N_19899);
and UO_859 (O_859,N_19852,N_19854);
nand UO_860 (O_860,N_19883,N_19985);
or UO_861 (O_861,N_19867,N_19995);
and UO_862 (O_862,N_19928,N_19986);
xor UO_863 (O_863,N_19908,N_19853);
nor UO_864 (O_864,N_19999,N_19851);
nor UO_865 (O_865,N_19982,N_19866);
xor UO_866 (O_866,N_19952,N_19864);
xor UO_867 (O_867,N_19891,N_19904);
nor UO_868 (O_868,N_19935,N_19949);
nand UO_869 (O_869,N_19879,N_19878);
nor UO_870 (O_870,N_19978,N_19891);
nor UO_871 (O_871,N_19920,N_19862);
xnor UO_872 (O_872,N_19920,N_19967);
or UO_873 (O_873,N_19979,N_19859);
or UO_874 (O_874,N_19980,N_19907);
nand UO_875 (O_875,N_19869,N_19948);
or UO_876 (O_876,N_19925,N_19873);
and UO_877 (O_877,N_19971,N_19844);
xnor UO_878 (O_878,N_19937,N_19987);
nand UO_879 (O_879,N_19964,N_19856);
nor UO_880 (O_880,N_19917,N_19976);
xor UO_881 (O_881,N_19962,N_19840);
or UO_882 (O_882,N_19917,N_19867);
or UO_883 (O_883,N_19893,N_19958);
nand UO_884 (O_884,N_19903,N_19983);
or UO_885 (O_885,N_19966,N_19886);
and UO_886 (O_886,N_19905,N_19964);
and UO_887 (O_887,N_19989,N_19898);
nor UO_888 (O_888,N_19840,N_19929);
or UO_889 (O_889,N_19920,N_19910);
nand UO_890 (O_890,N_19917,N_19873);
xnor UO_891 (O_891,N_19918,N_19932);
nor UO_892 (O_892,N_19975,N_19966);
nor UO_893 (O_893,N_19927,N_19931);
nand UO_894 (O_894,N_19955,N_19973);
or UO_895 (O_895,N_19884,N_19973);
and UO_896 (O_896,N_19919,N_19983);
nor UO_897 (O_897,N_19851,N_19962);
nand UO_898 (O_898,N_19860,N_19884);
nand UO_899 (O_899,N_19848,N_19991);
and UO_900 (O_900,N_19885,N_19855);
xnor UO_901 (O_901,N_19933,N_19959);
or UO_902 (O_902,N_19960,N_19904);
or UO_903 (O_903,N_19964,N_19871);
or UO_904 (O_904,N_19919,N_19878);
and UO_905 (O_905,N_19895,N_19944);
or UO_906 (O_906,N_19914,N_19901);
nor UO_907 (O_907,N_19996,N_19858);
or UO_908 (O_908,N_19860,N_19859);
or UO_909 (O_909,N_19901,N_19847);
nor UO_910 (O_910,N_19984,N_19989);
xor UO_911 (O_911,N_19972,N_19868);
nand UO_912 (O_912,N_19975,N_19851);
or UO_913 (O_913,N_19881,N_19951);
and UO_914 (O_914,N_19889,N_19984);
nand UO_915 (O_915,N_19931,N_19879);
and UO_916 (O_916,N_19959,N_19877);
xnor UO_917 (O_917,N_19904,N_19888);
nor UO_918 (O_918,N_19951,N_19915);
xnor UO_919 (O_919,N_19889,N_19860);
nand UO_920 (O_920,N_19902,N_19949);
and UO_921 (O_921,N_19909,N_19864);
nand UO_922 (O_922,N_19967,N_19871);
or UO_923 (O_923,N_19934,N_19888);
and UO_924 (O_924,N_19998,N_19954);
xor UO_925 (O_925,N_19969,N_19843);
and UO_926 (O_926,N_19842,N_19918);
or UO_927 (O_927,N_19859,N_19942);
and UO_928 (O_928,N_19983,N_19868);
and UO_929 (O_929,N_19959,N_19916);
and UO_930 (O_930,N_19905,N_19910);
nand UO_931 (O_931,N_19892,N_19944);
nand UO_932 (O_932,N_19934,N_19942);
nand UO_933 (O_933,N_19984,N_19969);
or UO_934 (O_934,N_19967,N_19898);
nor UO_935 (O_935,N_19897,N_19945);
nand UO_936 (O_936,N_19921,N_19900);
nand UO_937 (O_937,N_19916,N_19964);
nand UO_938 (O_938,N_19904,N_19873);
nand UO_939 (O_939,N_19844,N_19977);
or UO_940 (O_940,N_19963,N_19975);
nand UO_941 (O_941,N_19853,N_19918);
nand UO_942 (O_942,N_19909,N_19941);
and UO_943 (O_943,N_19868,N_19883);
xnor UO_944 (O_944,N_19988,N_19894);
nor UO_945 (O_945,N_19916,N_19917);
nor UO_946 (O_946,N_19872,N_19854);
or UO_947 (O_947,N_19908,N_19872);
nor UO_948 (O_948,N_19927,N_19877);
and UO_949 (O_949,N_19868,N_19975);
or UO_950 (O_950,N_19948,N_19942);
nor UO_951 (O_951,N_19844,N_19996);
nand UO_952 (O_952,N_19973,N_19922);
and UO_953 (O_953,N_19996,N_19913);
nor UO_954 (O_954,N_19841,N_19966);
nand UO_955 (O_955,N_19950,N_19897);
nand UO_956 (O_956,N_19980,N_19987);
xnor UO_957 (O_957,N_19916,N_19918);
xor UO_958 (O_958,N_19937,N_19891);
nor UO_959 (O_959,N_19956,N_19898);
nand UO_960 (O_960,N_19928,N_19919);
and UO_961 (O_961,N_19909,N_19980);
or UO_962 (O_962,N_19840,N_19856);
xor UO_963 (O_963,N_19854,N_19998);
nand UO_964 (O_964,N_19948,N_19949);
and UO_965 (O_965,N_19937,N_19898);
xnor UO_966 (O_966,N_19879,N_19911);
and UO_967 (O_967,N_19900,N_19844);
nor UO_968 (O_968,N_19841,N_19943);
nand UO_969 (O_969,N_19865,N_19909);
or UO_970 (O_970,N_19888,N_19847);
nor UO_971 (O_971,N_19964,N_19969);
nand UO_972 (O_972,N_19919,N_19994);
and UO_973 (O_973,N_19903,N_19982);
nor UO_974 (O_974,N_19982,N_19907);
or UO_975 (O_975,N_19922,N_19873);
nand UO_976 (O_976,N_19953,N_19842);
xor UO_977 (O_977,N_19963,N_19970);
nor UO_978 (O_978,N_19935,N_19958);
xor UO_979 (O_979,N_19897,N_19966);
and UO_980 (O_980,N_19876,N_19896);
and UO_981 (O_981,N_19874,N_19927);
nand UO_982 (O_982,N_19868,N_19921);
or UO_983 (O_983,N_19976,N_19856);
xor UO_984 (O_984,N_19943,N_19871);
or UO_985 (O_985,N_19974,N_19926);
nor UO_986 (O_986,N_19880,N_19985);
and UO_987 (O_987,N_19842,N_19987);
xor UO_988 (O_988,N_19904,N_19900);
nand UO_989 (O_989,N_19974,N_19943);
nor UO_990 (O_990,N_19884,N_19912);
nor UO_991 (O_991,N_19995,N_19939);
nand UO_992 (O_992,N_19940,N_19899);
nor UO_993 (O_993,N_19855,N_19899);
xor UO_994 (O_994,N_19881,N_19979);
nand UO_995 (O_995,N_19866,N_19844);
and UO_996 (O_996,N_19897,N_19856);
nor UO_997 (O_997,N_19842,N_19912);
nand UO_998 (O_998,N_19928,N_19953);
and UO_999 (O_999,N_19848,N_19868);
nor UO_1000 (O_1000,N_19903,N_19932);
and UO_1001 (O_1001,N_19866,N_19959);
nand UO_1002 (O_1002,N_19912,N_19900);
nand UO_1003 (O_1003,N_19939,N_19863);
xnor UO_1004 (O_1004,N_19916,N_19850);
or UO_1005 (O_1005,N_19951,N_19911);
xor UO_1006 (O_1006,N_19857,N_19926);
or UO_1007 (O_1007,N_19933,N_19882);
xor UO_1008 (O_1008,N_19878,N_19955);
nand UO_1009 (O_1009,N_19916,N_19886);
or UO_1010 (O_1010,N_19940,N_19859);
nor UO_1011 (O_1011,N_19925,N_19889);
xor UO_1012 (O_1012,N_19913,N_19945);
nor UO_1013 (O_1013,N_19921,N_19867);
nor UO_1014 (O_1014,N_19924,N_19993);
xor UO_1015 (O_1015,N_19974,N_19953);
nand UO_1016 (O_1016,N_19937,N_19879);
and UO_1017 (O_1017,N_19917,N_19980);
nor UO_1018 (O_1018,N_19946,N_19870);
and UO_1019 (O_1019,N_19845,N_19988);
xor UO_1020 (O_1020,N_19973,N_19876);
and UO_1021 (O_1021,N_19994,N_19974);
xnor UO_1022 (O_1022,N_19863,N_19867);
and UO_1023 (O_1023,N_19975,N_19958);
and UO_1024 (O_1024,N_19932,N_19915);
nor UO_1025 (O_1025,N_19863,N_19966);
xnor UO_1026 (O_1026,N_19986,N_19893);
or UO_1027 (O_1027,N_19952,N_19996);
nor UO_1028 (O_1028,N_19953,N_19886);
nor UO_1029 (O_1029,N_19981,N_19979);
or UO_1030 (O_1030,N_19915,N_19912);
xnor UO_1031 (O_1031,N_19906,N_19996);
nand UO_1032 (O_1032,N_19980,N_19959);
nor UO_1033 (O_1033,N_19948,N_19974);
or UO_1034 (O_1034,N_19864,N_19890);
or UO_1035 (O_1035,N_19903,N_19912);
and UO_1036 (O_1036,N_19951,N_19989);
xnor UO_1037 (O_1037,N_19883,N_19919);
nand UO_1038 (O_1038,N_19850,N_19920);
xnor UO_1039 (O_1039,N_19999,N_19961);
nor UO_1040 (O_1040,N_19969,N_19846);
nand UO_1041 (O_1041,N_19970,N_19847);
nor UO_1042 (O_1042,N_19984,N_19920);
nand UO_1043 (O_1043,N_19957,N_19908);
nand UO_1044 (O_1044,N_19937,N_19943);
nor UO_1045 (O_1045,N_19957,N_19996);
nor UO_1046 (O_1046,N_19981,N_19893);
nor UO_1047 (O_1047,N_19969,N_19879);
nor UO_1048 (O_1048,N_19865,N_19957);
and UO_1049 (O_1049,N_19968,N_19842);
xor UO_1050 (O_1050,N_19969,N_19900);
or UO_1051 (O_1051,N_19908,N_19964);
nor UO_1052 (O_1052,N_19864,N_19851);
xnor UO_1053 (O_1053,N_19890,N_19980);
and UO_1054 (O_1054,N_19859,N_19918);
and UO_1055 (O_1055,N_19933,N_19965);
nand UO_1056 (O_1056,N_19966,N_19919);
or UO_1057 (O_1057,N_19926,N_19919);
and UO_1058 (O_1058,N_19982,N_19883);
xnor UO_1059 (O_1059,N_19880,N_19912);
or UO_1060 (O_1060,N_19954,N_19936);
nor UO_1061 (O_1061,N_19943,N_19895);
nand UO_1062 (O_1062,N_19866,N_19968);
xnor UO_1063 (O_1063,N_19882,N_19967);
nor UO_1064 (O_1064,N_19973,N_19846);
or UO_1065 (O_1065,N_19935,N_19916);
nand UO_1066 (O_1066,N_19902,N_19850);
xor UO_1067 (O_1067,N_19977,N_19855);
xor UO_1068 (O_1068,N_19913,N_19891);
or UO_1069 (O_1069,N_19972,N_19906);
or UO_1070 (O_1070,N_19907,N_19972);
nand UO_1071 (O_1071,N_19909,N_19851);
xor UO_1072 (O_1072,N_19921,N_19955);
or UO_1073 (O_1073,N_19924,N_19997);
and UO_1074 (O_1074,N_19858,N_19903);
nor UO_1075 (O_1075,N_19847,N_19999);
or UO_1076 (O_1076,N_19967,N_19911);
nor UO_1077 (O_1077,N_19996,N_19910);
and UO_1078 (O_1078,N_19866,N_19948);
xnor UO_1079 (O_1079,N_19895,N_19857);
or UO_1080 (O_1080,N_19901,N_19984);
or UO_1081 (O_1081,N_19921,N_19880);
xnor UO_1082 (O_1082,N_19961,N_19872);
or UO_1083 (O_1083,N_19921,N_19910);
xor UO_1084 (O_1084,N_19975,N_19875);
or UO_1085 (O_1085,N_19968,N_19985);
and UO_1086 (O_1086,N_19959,N_19888);
nand UO_1087 (O_1087,N_19956,N_19927);
xor UO_1088 (O_1088,N_19990,N_19922);
xor UO_1089 (O_1089,N_19920,N_19877);
xnor UO_1090 (O_1090,N_19871,N_19962);
xor UO_1091 (O_1091,N_19973,N_19926);
nand UO_1092 (O_1092,N_19951,N_19902);
or UO_1093 (O_1093,N_19931,N_19869);
nand UO_1094 (O_1094,N_19869,N_19862);
and UO_1095 (O_1095,N_19869,N_19846);
xor UO_1096 (O_1096,N_19965,N_19934);
or UO_1097 (O_1097,N_19909,N_19981);
and UO_1098 (O_1098,N_19995,N_19887);
nand UO_1099 (O_1099,N_19939,N_19934);
nand UO_1100 (O_1100,N_19926,N_19848);
or UO_1101 (O_1101,N_19956,N_19917);
or UO_1102 (O_1102,N_19908,N_19890);
nand UO_1103 (O_1103,N_19861,N_19945);
nor UO_1104 (O_1104,N_19870,N_19949);
or UO_1105 (O_1105,N_19975,N_19991);
xnor UO_1106 (O_1106,N_19853,N_19962);
or UO_1107 (O_1107,N_19865,N_19918);
nand UO_1108 (O_1108,N_19886,N_19852);
or UO_1109 (O_1109,N_19897,N_19951);
nor UO_1110 (O_1110,N_19880,N_19924);
xnor UO_1111 (O_1111,N_19936,N_19916);
nand UO_1112 (O_1112,N_19969,N_19898);
xnor UO_1113 (O_1113,N_19877,N_19848);
xor UO_1114 (O_1114,N_19962,N_19997);
nand UO_1115 (O_1115,N_19894,N_19900);
and UO_1116 (O_1116,N_19899,N_19927);
nand UO_1117 (O_1117,N_19922,N_19897);
nand UO_1118 (O_1118,N_19897,N_19955);
nor UO_1119 (O_1119,N_19900,N_19898);
nor UO_1120 (O_1120,N_19889,N_19901);
xor UO_1121 (O_1121,N_19969,N_19980);
or UO_1122 (O_1122,N_19889,N_19851);
and UO_1123 (O_1123,N_19965,N_19956);
and UO_1124 (O_1124,N_19901,N_19971);
nor UO_1125 (O_1125,N_19906,N_19921);
nand UO_1126 (O_1126,N_19962,N_19927);
xor UO_1127 (O_1127,N_19902,N_19978);
and UO_1128 (O_1128,N_19841,N_19965);
nand UO_1129 (O_1129,N_19978,N_19981);
and UO_1130 (O_1130,N_19930,N_19929);
nor UO_1131 (O_1131,N_19973,N_19977);
nand UO_1132 (O_1132,N_19947,N_19978);
nor UO_1133 (O_1133,N_19903,N_19873);
or UO_1134 (O_1134,N_19986,N_19964);
or UO_1135 (O_1135,N_19985,N_19888);
nand UO_1136 (O_1136,N_19898,N_19955);
xor UO_1137 (O_1137,N_19973,N_19904);
and UO_1138 (O_1138,N_19866,N_19943);
nor UO_1139 (O_1139,N_19870,N_19877);
or UO_1140 (O_1140,N_19922,N_19982);
or UO_1141 (O_1141,N_19929,N_19910);
xor UO_1142 (O_1142,N_19887,N_19986);
and UO_1143 (O_1143,N_19887,N_19999);
and UO_1144 (O_1144,N_19943,N_19961);
nor UO_1145 (O_1145,N_19974,N_19937);
nand UO_1146 (O_1146,N_19987,N_19864);
and UO_1147 (O_1147,N_19985,N_19984);
and UO_1148 (O_1148,N_19861,N_19975);
nor UO_1149 (O_1149,N_19989,N_19942);
nand UO_1150 (O_1150,N_19918,N_19941);
nand UO_1151 (O_1151,N_19916,N_19855);
xnor UO_1152 (O_1152,N_19880,N_19859);
or UO_1153 (O_1153,N_19945,N_19933);
xor UO_1154 (O_1154,N_19975,N_19906);
nand UO_1155 (O_1155,N_19991,N_19977);
and UO_1156 (O_1156,N_19921,N_19938);
nor UO_1157 (O_1157,N_19868,N_19872);
nor UO_1158 (O_1158,N_19850,N_19843);
nor UO_1159 (O_1159,N_19938,N_19863);
or UO_1160 (O_1160,N_19944,N_19878);
and UO_1161 (O_1161,N_19846,N_19853);
nor UO_1162 (O_1162,N_19999,N_19884);
and UO_1163 (O_1163,N_19880,N_19996);
or UO_1164 (O_1164,N_19995,N_19931);
nand UO_1165 (O_1165,N_19951,N_19844);
xnor UO_1166 (O_1166,N_19999,N_19984);
nor UO_1167 (O_1167,N_19873,N_19938);
xnor UO_1168 (O_1168,N_19847,N_19875);
nand UO_1169 (O_1169,N_19946,N_19944);
xnor UO_1170 (O_1170,N_19904,N_19862);
and UO_1171 (O_1171,N_19932,N_19922);
or UO_1172 (O_1172,N_19963,N_19947);
nand UO_1173 (O_1173,N_19962,N_19970);
nand UO_1174 (O_1174,N_19873,N_19881);
or UO_1175 (O_1175,N_19906,N_19987);
or UO_1176 (O_1176,N_19904,N_19931);
nor UO_1177 (O_1177,N_19993,N_19997);
and UO_1178 (O_1178,N_19988,N_19855);
nand UO_1179 (O_1179,N_19918,N_19946);
nand UO_1180 (O_1180,N_19983,N_19898);
nor UO_1181 (O_1181,N_19924,N_19920);
or UO_1182 (O_1182,N_19892,N_19879);
and UO_1183 (O_1183,N_19921,N_19999);
or UO_1184 (O_1184,N_19894,N_19952);
or UO_1185 (O_1185,N_19976,N_19870);
nand UO_1186 (O_1186,N_19889,N_19866);
and UO_1187 (O_1187,N_19845,N_19968);
nand UO_1188 (O_1188,N_19889,N_19985);
or UO_1189 (O_1189,N_19992,N_19953);
or UO_1190 (O_1190,N_19937,N_19851);
xor UO_1191 (O_1191,N_19971,N_19939);
nor UO_1192 (O_1192,N_19925,N_19977);
or UO_1193 (O_1193,N_19880,N_19884);
xnor UO_1194 (O_1194,N_19962,N_19957);
xor UO_1195 (O_1195,N_19929,N_19992);
nand UO_1196 (O_1196,N_19889,N_19909);
and UO_1197 (O_1197,N_19884,N_19870);
or UO_1198 (O_1198,N_19918,N_19958);
nor UO_1199 (O_1199,N_19986,N_19943);
nor UO_1200 (O_1200,N_19960,N_19876);
nand UO_1201 (O_1201,N_19920,N_19883);
nand UO_1202 (O_1202,N_19910,N_19863);
xor UO_1203 (O_1203,N_19962,N_19858);
or UO_1204 (O_1204,N_19888,N_19911);
nor UO_1205 (O_1205,N_19932,N_19860);
or UO_1206 (O_1206,N_19851,N_19846);
and UO_1207 (O_1207,N_19956,N_19899);
nor UO_1208 (O_1208,N_19988,N_19992);
xor UO_1209 (O_1209,N_19843,N_19947);
xor UO_1210 (O_1210,N_19967,N_19868);
xor UO_1211 (O_1211,N_19902,N_19899);
nor UO_1212 (O_1212,N_19976,N_19854);
nor UO_1213 (O_1213,N_19849,N_19954);
and UO_1214 (O_1214,N_19950,N_19895);
nor UO_1215 (O_1215,N_19871,N_19935);
nor UO_1216 (O_1216,N_19906,N_19882);
nor UO_1217 (O_1217,N_19909,N_19957);
xnor UO_1218 (O_1218,N_19883,N_19889);
nor UO_1219 (O_1219,N_19857,N_19948);
or UO_1220 (O_1220,N_19981,N_19929);
nand UO_1221 (O_1221,N_19938,N_19854);
nand UO_1222 (O_1222,N_19977,N_19994);
nand UO_1223 (O_1223,N_19883,N_19940);
and UO_1224 (O_1224,N_19986,N_19984);
nand UO_1225 (O_1225,N_19905,N_19935);
nor UO_1226 (O_1226,N_19961,N_19949);
nor UO_1227 (O_1227,N_19869,N_19890);
nand UO_1228 (O_1228,N_19948,N_19943);
nor UO_1229 (O_1229,N_19889,N_19919);
nand UO_1230 (O_1230,N_19935,N_19868);
nor UO_1231 (O_1231,N_19916,N_19982);
nor UO_1232 (O_1232,N_19956,N_19885);
xor UO_1233 (O_1233,N_19936,N_19865);
and UO_1234 (O_1234,N_19874,N_19993);
or UO_1235 (O_1235,N_19899,N_19890);
or UO_1236 (O_1236,N_19957,N_19858);
xor UO_1237 (O_1237,N_19851,N_19921);
nor UO_1238 (O_1238,N_19999,N_19925);
xor UO_1239 (O_1239,N_19887,N_19956);
nor UO_1240 (O_1240,N_19873,N_19926);
and UO_1241 (O_1241,N_19881,N_19866);
or UO_1242 (O_1242,N_19959,N_19997);
xnor UO_1243 (O_1243,N_19858,N_19899);
xnor UO_1244 (O_1244,N_19957,N_19843);
and UO_1245 (O_1245,N_19969,N_19999);
nand UO_1246 (O_1246,N_19906,N_19945);
xnor UO_1247 (O_1247,N_19998,N_19916);
or UO_1248 (O_1248,N_19976,N_19840);
and UO_1249 (O_1249,N_19996,N_19854);
nor UO_1250 (O_1250,N_19853,N_19934);
xnor UO_1251 (O_1251,N_19928,N_19914);
or UO_1252 (O_1252,N_19913,N_19877);
and UO_1253 (O_1253,N_19957,N_19985);
or UO_1254 (O_1254,N_19879,N_19923);
or UO_1255 (O_1255,N_19850,N_19854);
nand UO_1256 (O_1256,N_19916,N_19905);
xor UO_1257 (O_1257,N_19947,N_19943);
nand UO_1258 (O_1258,N_19939,N_19949);
or UO_1259 (O_1259,N_19845,N_19908);
nor UO_1260 (O_1260,N_19855,N_19998);
and UO_1261 (O_1261,N_19871,N_19942);
nand UO_1262 (O_1262,N_19928,N_19860);
or UO_1263 (O_1263,N_19988,N_19901);
and UO_1264 (O_1264,N_19919,N_19849);
xnor UO_1265 (O_1265,N_19886,N_19911);
and UO_1266 (O_1266,N_19996,N_19915);
xor UO_1267 (O_1267,N_19886,N_19951);
nand UO_1268 (O_1268,N_19895,N_19911);
nand UO_1269 (O_1269,N_19938,N_19945);
or UO_1270 (O_1270,N_19978,N_19962);
nor UO_1271 (O_1271,N_19982,N_19924);
nand UO_1272 (O_1272,N_19901,N_19888);
nand UO_1273 (O_1273,N_19990,N_19841);
nor UO_1274 (O_1274,N_19920,N_19943);
and UO_1275 (O_1275,N_19891,N_19944);
xor UO_1276 (O_1276,N_19965,N_19860);
nand UO_1277 (O_1277,N_19991,N_19843);
and UO_1278 (O_1278,N_19984,N_19967);
nand UO_1279 (O_1279,N_19982,N_19846);
and UO_1280 (O_1280,N_19970,N_19865);
nand UO_1281 (O_1281,N_19845,N_19890);
xnor UO_1282 (O_1282,N_19995,N_19951);
or UO_1283 (O_1283,N_19907,N_19842);
nor UO_1284 (O_1284,N_19855,N_19927);
or UO_1285 (O_1285,N_19926,N_19876);
nand UO_1286 (O_1286,N_19983,N_19991);
and UO_1287 (O_1287,N_19967,N_19843);
nor UO_1288 (O_1288,N_19889,N_19884);
nand UO_1289 (O_1289,N_19978,N_19927);
nand UO_1290 (O_1290,N_19972,N_19961);
xor UO_1291 (O_1291,N_19875,N_19980);
and UO_1292 (O_1292,N_19952,N_19884);
xnor UO_1293 (O_1293,N_19933,N_19979);
xor UO_1294 (O_1294,N_19921,N_19914);
and UO_1295 (O_1295,N_19974,N_19876);
and UO_1296 (O_1296,N_19890,N_19956);
nor UO_1297 (O_1297,N_19848,N_19934);
xnor UO_1298 (O_1298,N_19937,N_19893);
nor UO_1299 (O_1299,N_19876,N_19976);
xnor UO_1300 (O_1300,N_19950,N_19942);
nand UO_1301 (O_1301,N_19883,N_19959);
nand UO_1302 (O_1302,N_19997,N_19914);
nand UO_1303 (O_1303,N_19991,N_19902);
xnor UO_1304 (O_1304,N_19929,N_19918);
or UO_1305 (O_1305,N_19929,N_19968);
and UO_1306 (O_1306,N_19852,N_19875);
and UO_1307 (O_1307,N_19914,N_19973);
or UO_1308 (O_1308,N_19920,N_19976);
xnor UO_1309 (O_1309,N_19941,N_19860);
nand UO_1310 (O_1310,N_19992,N_19983);
or UO_1311 (O_1311,N_19898,N_19883);
nand UO_1312 (O_1312,N_19937,N_19964);
and UO_1313 (O_1313,N_19955,N_19961);
xnor UO_1314 (O_1314,N_19994,N_19876);
nor UO_1315 (O_1315,N_19932,N_19892);
or UO_1316 (O_1316,N_19916,N_19897);
nand UO_1317 (O_1317,N_19869,N_19912);
and UO_1318 (O_1318,N_19924,N_19869);
nand UO_1319 (O_1319,N_19968,N_19850);
xor UO_1320 (O_1320,N_19852,N_19980);
xnor UO_1321 (O_1321,N_19871,N_19861);
nor UO_1322 (O_1322,N_19950,N_19893);
nand UO_1323 (O_1323,N_19841,N_19937);
and UO_1324 (O_1324,N_19876,N_19922);
nor UO_1325 (O_1325,N_19916,N_19938);
and UO_1326 (O_1326,N_19967,N_19985);
or UO_1327 (O_1327,N_19952,N_19914);
nand UO_1328 (O_1328,N_19981,N_19885);
and UO_1329 (O_1329,N_19866,N_19869);
and UO_1330 (O_1330,N_19982,N_19840);
nor UO_1331 (O_1331,N_19988,N_19923);
nor UO_1332 (O_1332,N_19989,N_19855);
nand UO_1333 (O_1333,N_19978,N_19921);
xor UO_1334 (O_1334,N_19933,N_19944);
or UO_1335 (O_1335,N_19995,N_19963);
or UO_1336 (O_1336,N_19950,N_19863);
nand UO_1337 (O_1337,N_19992,N_19856);
xnor UO_1338 (O_1338,N_19894,N_19979);
or UO_1339 (O_1339,N_19853,N_19877);
nand UO_1340 (O_1340,N_19934,N_19979);
nand UO_1341 (O_1341,N_19995,N_19912);
xnor UO_1342 (O_1342,N_19869,N_19983);
nand UO_1343 (O_1343,N_19916,N_19868);
nor UO_1344 (O_1344,N_19860,N_19937);
nand UO_1345 (O_1345,N_19890,N_19942);
nand UO_1346 (O_1346,N_19992,N_19980);
xor UO_1347 (O_1347,N_19928,N_19904);
or UO_1348 (O_1348,N_19990,N_19870);
nor UO_1349 (O_1349,N_19866,N_19851);
nor UO_1350 (O_1350,N_19958,N_19977);
nand UO_1351 (O_1351,N_19892,N_19968);
nand UO_1352 (O_1352,N_19965,N_19909);
xnor UO_1353 (O_1353,N_19935,N_19882);
nor UO_1354 (O_1354,N_19918,N_19931);
nand UO_1355 (O_1355,N_19878,N_19962);
or UO_1356 (O_1356,N_19906,N_19893);
or UO_1357 (O_1357,N_19986,N_19944);
xnor UO_1358 (O_1358,N_19952,N_19926);
xnor UO_1359 (O_1359,N_19974,N_19870);
and UO_1360 (O_1360,N_19910,N_19870);
or UO_1361 (O_1361,N_19862,N_19929);
nor UO_1362 (O_1362,N_19941,N_19972);
and UO_1363 (O_1363,N_19930,N_19972);
and UO_1364 (O_1364,N_19986,N_19843);
nor UO_1365 (O_1365,N_19869,N_19902);
or UO_1366 (O_1366,N_19913,N_19921);
nand UO_1367 (O_1367,N_19950,N_19854);
nand UO_1368 (O_1368,N_19955,N_19890);
nand UO_1369 (O_1369,N_19843,N_19941);
or UO_1370 (O_1370,N_19995,N_19920);
nand UO_1371 (O_1371,N_19895,N_19954);
and UO_1372 (O_1372,N_19908,N_19961);
nand UO_1373 (O_1373,N_19946,N_19892);
xor UO_1374 (O_1374,N_19932,N_19845);
nor UO_1375 (O_1375,N_19894,N_19983);
or UO_1376 (O_1376,N_19851,N_19967);
nor UO_1377 (O_1377,N_19871,N_19845);
nor UO_1378 (O_1378,N_19989,N_19860);
nor UO_1379 (O_1379,N_19969,N_19848);
or UO_1380 (O_1380,N_19895,N_19840);
xnor UO_1381 (O_1381,N_19966,N_19901);
xnor UO_1382 (O_1382,N_19965,N_19940);
nor UO_1383 (O_1383,N_19842,N_19903);
nand UO_1384 (O_1384,N_19973,N_19938);
xor UO_1385 (O_1385,N_19846,N_19988);
nor UO_1386 (O_1386,N_19934,N_19878);
nor UO_1387 (O_1387,N_19887,N_19868);
nand UO_1388 (O_1388,N_19996,N_19960);
xnor UO_1389 (O_1389,N_19981,N_19965);
nor UO_1390 (O_1390,N_19949,N_19956);
xor UO_1391 (O_1391,N_19848,N_19876);
nor UO_1392 (O_1392,N_19924,N_19865);
or UO_1393 (O_1393,N_19978,N_19923);
xnor UO_1394 (O_1394,N_19933,N_19881);
nand UO_1395 (O_1395,N_19842,N_19935);
xnor UO_1396 (O_1396,N_19875,N_19890);
and UO_1397 (O_1397,N_19854,N_19913);
xor UO_1398 (O_1398,N_19965,N_19858);
nand UO_1399 (O_1399,N_19954,N_19883);
or UO_1400 (O_1400,N_19904,N_19880);
and UO_1401 (O_1401,N_19888,N_19977);
nand UO_1402 (O_1402,N_19922,N_19882);
nand UO_1403 (O_1403,N_19951,N_19964);
xnor UO_1404 (O_1404,N_19870,N_19859);
nor UO_1405 (O_1405,N_19880,N_19911);
and UO_1406 (O_1406,N_19919,N_19866);
nand UO_1407 (O_1407,N_19981,N_19928);
xor UO_1408 (O_1408,N_19924,N_19891);
nand UO_1409 (O_1409,N_19869,N_19955);
or UO_1410 (O_1410,N_19840,N_19847);
or UO_1411 (O_1411,N_19994,N_19862);
nor UO_1412 (O_1412,N_19888,N_19899);
xnor UO_1413 (O_1413,N_19942,N_19953);
nand UO_1414 (O_1414,N_19903,N_19924);
nand UO_1415 (O_1415,N_19893,N_19863);
or UO_1416 (O_1416,N_19964,N_19990);
or UO_1417 (O_1417,N_19843,N_19865);
or UO_1418 (O_1418,N_19941,N_19954);
or UO_1419 (O_1419,N_19951,N_19927);
xnor UO_1420 (O_1420,N_19913,N_19840);
or UO_1421 (O_1421,N_19956,N_19928);
and UO_1422 (O_1422,N_19918,N_19948);
xnor UO_1423 (O_1423,N_19966,N_19880);
nand UO_1424 (O_1424,N_19911,N_19987);
nand UO_1425 (O_1425,N_19850,N_19899);
and UO_1426 (O_1426,N_19887,N_19854);
nand UO_1427 (O_1427,N_19867,N_19954);
xor UO_1428 (O_1428,N_19993,N_19856);
xor UO_1429 (O_1429,N_19893,N_19905);
xor UO_1430 (O_1430,N_19955,N_19883);
xor UO_1431 (O_1431,N_19919,N_19934);
xor UO_1432 (O_1432,N_19887,N_19850);
or UO_1433 (O_1433,N_19989,N_19932);
and UO_1434 (O_1434,N_19905,N_19930);
and UO_1435 (O_1435,N_19994,N_19868);
nand UO_1436 (O_1436,N_19870,N_19867);
and UO_1437 (O_1437,N_19896,N_19898);
nand UO_1438 (O_1438,N_19891,N_19906);
or UO_1439 (O_1439,N_19921,N_19904);
xnor UO_1440 (O_1440,N_19869,N_19876);
or UO_1441 (O_1441,N_19872,N_19875);
nor UO_1442 (O_1442,N_19880,N_19933);
nand UO_1443 (O_1443,N_19849,N_19893);
or UO_1444 (O_1444,N_19959,N_19847);
nand UO_1445 (O_1445,N_19863,N_19891);
and UO_1446 (O_1446,N_19851,N_19931);
nor UO_1447 (O_1447,N_19953,N_19907);
nor UO_1448 (O_1448,N_19925,N_19966);
nand UO_1449 (O_1449,N_19990,N_19877);
nor UO_1450 (O_1450,N_19895,N_19861);
or UO_1451 (O_1451,N_19912,N_19934);
xor UO_1452 (O_1452,N_19895,N_19903);
and UO_1453 (O_1453,N_19944,N_19963);
xnor UO_1454 (O_1454,N_19918,N_19989);
xnor UO_1455 (O_1455,N_19975,N_19986);
nor UO_1456 (O_1456,N_19914,N_19991);
or UO_1457 (O_1457,N_19907,N_19886);
xnor UO_1458 (O_1458,N_19874,N_19923);
nand UO_1459 (O_1459,N_19911,N_19916);
xnor UO_1460 (O_1460,N_19892,N_19882);
xor UO_1461 (O_1461,N_19852,N_19898);
nor UO_1462 (O_1462,N_19859,N_19879);
xor UO_1463 (O_1463,N_19904,N_19898);
and UO_1464 (O_1464,N_19955,N_19899);
nand UO_1465 (O_1465,N_19906,N_19970);
or UO_1466 (O_1466,N_19865,N_19982);
or UO_1467 (O_1467,N_19912,N_19940);
nor UO_1468 (O_1468,N_19956,N_19966);
xor UO_1469 (O_1469,N_19864,N_19921);
or UO_1470 (O_1470,N_19853,N_19907);
and UO_1471 (O_1471,N_19921,N_19844);
nand UO_1472 (O_1472,N_19896,N_19920);
and UO_1473 (O_1473,N_19898,N_19921);
nor UO_1474 (O_1474,N_19979,N_19995);
xnor UO_1475 (O_1475,N_19856,N_19944);
nand UO_1476 (O_1476,N_19863,N_19869);
nand UO_1477 (O_1477,N_19976,N_19852);
and UO_1478 (O_1478,N_19926,N_19951);
and UO_1479 (O_1479,N_19918,N_19858);
and UO_1480 (O_1480,N_19941,N_19966);
nand UO_1481 (O_1481,N_19891,N_19946);
or UO_1482 (O_1482,N_19924,N_19937);
nor UO_1483 (O_1483,N_19964,N_19982);
xor UO_1484 (O_1484,N_19990,N_19908);
nand UO_1485 (O_1485,N_19995,N_19895);
and UO_1486 (O_1486,N_19861,N_19907);
or UO_1487 (O_1487,N_19964,N_19965);
xor UO_1488 (O_1488,N_19874,N_19958);
and UO_1489 (O_1489,N_19914,N_19913);
nor UO_1490 (O_1490,N_19871,N_19846);
xnor UO_1491 (O_1491,N_19879,N_19944);
nor UO_1492 (O_1492,N_19906,N_19969);
and UO_1493 (O_1493,N_19920,N_19847);
or UO_1494 (O_1494,N_19884,N_19871);
nand UO_1495 (O_1495,N_19941,N_19956);
nor UO_1496 (O_1496,N_19942,N_19972);
nand UO_1497 (O_1497,N_19853,N_19952);
and UO_1498 (O_1498,N_19958,N_19855);
and UO_1499 (O_1499,N_19929,N_19983);
nor UO_1500 (O_1500,N_19962,N_19906);
and UO_1501 (O_1501,N_19888,N_19896);
nand UO_1502 (O_1502,N_19987,N_19888);
nor UO_1503 (O_1503,N_19906,N_19901);
and UO_1504 (O_1504,N_19870,N_19942);
xnor UO_1505 (O_1505,N_19940,N_19856);
and UO_1506 (O_1506,N_19970,N_19928);
nand UO_1507 (O_1507,N_19864,N_19876);
nor UO_1508 (O_1508,N_19851,N_19951);
xnor UO_1509 (O_1509,N_19934,N_19937);
nand UO_1510 (O_1510,N_19888,N_19846);
xor UO_1511 (O_1511,N_19845,N_19923);
nand UO_1512 (O_1512,N_19913,N_19865);
xor UO_1513 (O_1513,N_19890,N_19928);
xnor UO_1514 (O_1514,N_19876,N_19988);
and UO_1515 (O_1515,N_19857,N_19981);
or UO_1516 (O_1516,N_19995,N_19964);
xnor UO_1517 (O_1517,N_19977,N_19841);
and UO_1518 (O_1518,N_19851,N_19932);
nor UO_1519 (O_1519,N_19947,N_19966);
nand UO_1520 (O_1520,N_19894,N_19965);
nor UO_1521 (O_1521,N_19844,N_19913);
nor UO_1522 (O_1522,N_19873,N_19861);
xnor UO_1523 (O_1523,N_19927,N_19922);
or UO_1524 (O_1524,N_19990,N_19861);
or UO_1525 (O_1525,N_19985,N_19972);
xnor UO_1526 (O_1526,N_19879,N_19898);
xor UO_1527 (O_1527,N_19966,N_19962);
or UO_1528 (O_1528,N_19868,N_19856);
xor UO_1529 (O_1529,N_19963,N_19846);
and UO_1530 (O_1530,N_19919,N_19967);
and UO_1531 (O_1531,N_19899,N_19874);
xnor UO_1532 (O_1532,N_19939,N_19991);
nand UO_1533 (O_1533,N_19923,N_19900);
or UO_1534 (O_1534,N_19867,N_19967);
nor UO_1535 (O_1535,N_19848,N_19890);
nor UO_1536 (O_1536,N_19957,N_19910);
nand UO_1537 (O_1537,N_19920,N_19922);
nand UO_1538 (O_1538,N_19847,N_19975);
nand UO_1539 (O_1539,N_19927,N_19903);
or UO_1540 (O_1540,N_19862,N_19866);
and UO_1541 (O_1541,N_19936,N_19855);
and UO_1542 (O_1542,N_19952,N_19971);
nand UO_1543 (O_1543,N_19975,N_19962);
and UO_1544 (O_1544,N_19991,N_19943);
nor UO_1545 (O_1545,N_19968,N_19908);
nor UO_1546 (O_1546,N_19848,N_19881);
or UO_1547 (O_1547,N_19920,N_19969);
nand UO_1548 (O_1548,N_19977,N_19873);
xnor UO_1549 (O_1549,N_19939,N_19897);
xor UO_1550 (O_1550,N_19929,N_19944);
or UO_1551 (O_1551,N_19900,N_19872);
xor UO_1552 (O_1552,N_19874,N_19871);
nand UO_1553 (O_1553,N_19842,N_19871);
xnor UO_1554 (O_1554,N_19908,N_19953);
and UO_1555 (O_1555,N_19951,N_19907);
xor UO_1556 (O_1556,N_19848,N_19856);
or UO_1557 (O_1557,N_19928,N_19979);
nor UO_1558 (O_1558,N_19958,N_19944);
or UO_1559 (O_1559,N_19974,N_19882);
nand UO_1560 (O_1560,N_19950,N_19867);
or UO_1561 (O_1561,N_19986,N_19897);
nor UO_1562 (O_1562,N_19843,N_19983);
nor UO_1563 (O_1563,N_19843,N_19958);
or UO_1564 (O_1564,N_19894,N_19855);
and UO_1565 (O_1565,N_19954,N_19990);
nand UO_1566 (O_1566,N_19896,N_19988);
xor UO_1567 (O_1567,N_19882,N_19970);
nor UO_1568 (O_1568,N_19921,N_19957);
and UO_1569 (O_1569,N_19952,N_19925);
nor UO_1570 (O_1570,N_19983,N_19922);
or UO_1571 (O_1571,N_19895,N_19962);
nand UO_1572 (O_1572,N_19999,N_19867);
nor UO_1573 (O_1573,N_19865,N_19915);
and UO_1574 (O_1574,N_19924,N_19998);
or UO_1575 (O_1575,N_19934,N_19945);
xor UO_1576 (O_1576,N_19990,N_19958);
or UO_1577 (O_1577,N_19919,N_19908);
nor UO_1578 (O_1578,N_19997,N_19998);
nor UO_1579 (O_1579,N_19917,N_19981);
nor UO_1580 (O_1580,N_19978,N_19956);
nor UO_1581 (O_1581,N_19886,N_19964);
and UO_1582 (O_1582,N_19862,N_19991);
nand UO_1583 (O_1583,N_19934,N_19953);
nand UO_1584 (O_1584,N_19891,N_19848);
xnor UO_1585 (O_1585,N_19856,N_19890);
xor UO_1586 (O_1586,N_19976,N_19948);
xor UO_1587 (O_1587,N_19931,N_19936);
nand UO_1588 (O_1588,N_19933,N_19923);
or UO_1589 (O_1589,N_19857,N_19929);
and UO_1590 (O_1590,N_19862,N_19969);
and UO_1591 (O_1591,N_19916,N_19847);
nand UO_1592 (O_1592,N_19997,N_19849);
nor UO_1593 (O_1593,N_19909,N_19931);
nand UO_1594 (O_1594,N_19981,N_19951);
nor UO_1595 (O_1595,N_19882,N_19963);
nor UO_1596 (O_1596,N_19987,N_19981);
nor UO_1597 (O_1597,N_19973,N_19992);
and UO_1598 (O_1598,N_19951,N_19979);
xnor UO_1599 (O_1599,N_19940,N_19967);
and UO_1600 (O_1600,N_19928,N_19966);
nand UO_1601 (O_1601,N_19962,N_19946);
or UO_1602 (O_1602,N_19987,N_19977);
nand UO_1603 (O_1603,N_19862,N_19895);
nor UO_1604 (O_1604,N_19926,N_19967);
nand UO_1605 (O_1605,N_19970,N_19955);
xnor UO_1606 (O_1606,N_19917,N_19970);
xor UO_1607 (O_1607,N_19969,N_19905);
and UO_1608 (O_1608,N_19948,N_19916);
and UO_1609 (O_1609,N_19857,N_19882);
and UO_1610 (O_1610,N_19899,N_19910);
nor UO_1611 (O_1611,N_19872,N_19902);
xnor UO_1612 (O_1612,N_19909,N_19843);
xor UO_1613 (O_1613,N_19938,N_19850);
nand UO_1614 (O_1614,N_19994,N_19917);
or UO_1615 (O_1615,N_19923,N_19877);
or UO_1616 (O_1616,N_19856,N_19970);
xnor UO_1617 (O_1617,N_19934,N_19843);
nand UO_1618 (O_1618,N_19933,N_19942);
xor UO_1619 (O_1619,N_19989,N_19912);
or UO_1620 (O_1620,N_19966,N_19957);
nor UO_1621 (O_1621,N_19852,N_19997);
xor UO_1622 (O_1622,N_19860,N_19867);
xnor UO_1623 (O_1623,N_19921,N_19932);
xor UO_1624 (O_1624,N_19887,N_19876);
or UO_1625 (O_1625,N_19960,N_19884);
or UO_1626 (O_1626,N_19906,N_19926);
and UO_1627 (O_1627,N_19858,N_19945);
nor UO_1628 (O_1628,N_19853,N_19925);
or UO_1629 (O_1629,N_19845,N_19880);
nand UO_1630 (O_1630,N_19930,N_19841);
nand UO_1631 (O_1631,N_19900,N_19993);
or UO_1632 (O_1632,N_19877,N_19925);
nor UO_1633 (O_1633,N_19932,N_19952);
or UO_1634 (O_1634,N_19919,N_19935);
xor UO_1635 (O_1635,N_19948,N_19889);
nand UO_1636 (O_1636,N_19984,N_19843);
nor UO_1637 (O_1637,N_19964,N_19943);
and UO_1638 (O_1638,N_19900,N_19842);
and UO_1639 (O_1639,N_19999,N_19862);
xor UO_1640 (O_1640,N_19912,N_19953);
nor UO_1641 (O_1641,N_19892,N_19954);
nand UO_1642 (O_1642,N_19859,N_19989);
and UO_1643 (O_1643,N_19956,N_19995);
and UO_1644 (O_1644,N_19944,N_19981);
and UO_1645 (O_1645,N_19904,N_19842);
nor UO_1646 (O_1646,N_19919,N_19850);
nand UO_1647 (O_1647,N_19974,N_19966);
xnor UO_1648 (O_1648,N_19954,N_19840);
and UO_1649 (O_1649,N_19960,N_19903);
nand UO_1650 (O_1650,N_19853,N_19884);
or UO_1651 (O_1651,N_19948,N_19878);
nor UO_1652 (O_1652,N_19953,N_19939);
or UO_1653 (O_1653,N_19988,N_19885);
nor UO_1654 (O_1654,N_19935,N_19844);
or UO_1655 (O_1655,N_19973,N_19854);
xor UO_1656 (O_1656,N_19881,N_19944);
and UO_1657 (O_1657,N_19891,N_19981);
nand UO_1658 (O_1658,N_19964,N_19972);
xor UO_1659 (O_1659,N_19920,N_19931);
and UO_1660 (O_1660,N_19891,N_19846);
nor UO_1661 (O_1661,N_19968,N_19867);
or UO_1662 (O_1662,N_19910,N_19909);
nand UO_1663 (O_1663,N_19911,N_19977);
xnor UO_1664 (O_1664,N_19914,N_19850);
and UO_1665 (O_1665,N_19846,N_19976);
nand UO_1666 (O_1666,N_19849,N_19924);
and UO_1667 (O_1667,N_19848,N_19970);
and UO_1668 (O_1668,N_19899,N_19954);
or UO_1669 (O_1669,N_19945,N_19855);
nand UO_1670 (O_1670,N_19846,N_19967);
xor UO_1671 (O_1671,N_19971,N_19906);
or UO_1672 (O_1672,N_19909,N_19868);
nor UO_1673 (O_1673,N_19921,N_19845);
xnor UO_1674 (O_1674,N_19982,N_19971);
or UO_1675 (O_1675,N_19844,N_19936);
nand UO_1676 (O_1676,N_19943,N_19967);
or UO_1677 (O_1677,N_19917,N_19937);
nor UO_1678 (O_1678,N_19970,N_19931);
or UO_1679 (O_1679,N_19848,N_19864);
xnor UO_1680 (O_1680,N_19841,N_19981);
xnor UO_1681 (O_1681,N_19894,N_19953);
xnor UO_1682 (O_1682,N_19905,N_19854);
xnor UO_1683 (O_1683,N_19946,N_19956);
nand UO_1684 (O_1684,N_19844,N_19983);
and UO_1685 (O_1685,N_19966,N_19895);
nand UO_1686 (O_1686,N_19933,N_19873);
or UO_1687 (O_1687,N_19888,N_19882);
nand UO_1688 (O_1688,N_19853,N_19980);
or UO_1689 (O_1689,N_19903,N_19871);
and UO_1690 (O_1690,N_19953,N_19916);
nand UO_1691 (O_1691,N_19856,N_19875);
or UO_1692 (O_1692,N_19930,N_19996);
nor UO_1693 (O_1693,N_19869,N_19977);
nor UO_1694 (O_1694,N_19848,N_19962);
xor UO_1695 (O_1695,N_19926,N_19860);
and UO_1696 (O_1696,N_19881,N_19867);
and UO_1697 (O_1697,N_19982,N_19958);
xnor UO_1698 (O_1698,N_19929,N_19878);
nor UO_1699 (O_1699,N_19953,N_19989);
xnor UO_1700 (O_1700,N_19971,N_19860);
and UO_1701 (O_1701,N_19961,N_19988);
nor UO_1702 (O_1702,N_19972,N_19975);
nand UO_1703 (O_1703,N_19954,N_19993);
and UO_1704 (O_1704,N_19915,N_19967);
or UO_1705 (O_1705,N_19993,N_19908);
and UO_1706 (O_1706,N_19875,N_19891);
and UO_1707 (O_1707,N_19853,N_19966);
nand UO_1708 (O_1708,N_19972,N_19957);
xnor UO_1709 (O_1709,N_19977,N_19865);
or UO_1710 (O_1710,N_19956,N_19930);
nand UO_1711 (O_1711,N_19997,N_19881);
xnor UO_1712 (O_1712,N_19938,N_19881);
or UO_1713 (O_1713,N_19865,N_19969);
xor UO_1714 (O_1714,N_19911,N_19847);
nand UO_1715 (O_1715,N_19907,N_19858);
nand UO_1716 (O_1716,N_19909,N_19930);
or UO_1717 (O_1717,N_19965,N_19848);
or UO_1718 (O_1718,N_19963,N_19891);
and UO_1719 (O_1719,N_19996,N_19863);
nand UO_1720 (O_1720,N_19993,N_19907);
nand UO_1721 (O_1721,N_19997,N_19874);
xnor UO_1722 (O_1722,N_19898,N_19991);
xnor UO_1723 (O_1723,N_19856,N_19939);
nor UO_1724 (O_1724,N_19866,N_19913);
or UO_1725 (O_1725,N_19860,N_19993);
and UO_1726 (O_1726,N_19998,N_19961);
nand UO_1727 (O_1727,N_19974,N_19923);
nor UO_1728 (O_1728,N_19961,N_19859);
and UO_1729 (O_1729,N_19938,N_19930);
or UO_1730 (O_1730,N_19868,N_19922);
nor UO_1731 (O_1731,N_19970,N_19995);
nand UO_1732 (O_1732,N_19914,N_19950);
and UO_1733 (O_1733,N_19852,N_19951);
and UO_1734 (O_1734,N_19994,N_19844);
or UO_1735 (O_1735,N_19918,N_19969);
nor UO_1736 (O_1736,N_19878,N_19947);
nor UO_1737 (O_1737,N_19945,N_19852);
or UO_1738 (O_1738,N_19961,N_19941);
xnor UO_1739 (O_1739,N_19984,N_19860);
and UO_1740 (O_1740,N_19895,N_19931);
xor UO_1741 (O_1741,N_19988,N_19888);
xnor UO_1742 (O_1742,N_19998,N_19860);
and UO_1743 (O_1743,N_19854,N_19869);
nand UO_1744 (O_1744,N_19886,N_19954);
nand UO_1745 (O_1745,N_19926,N_19858);
or UO_1746 (O_1746,N_19952,N_19974);
or UO_1747 (O_1747,N_19960,N_19875);
or UO_1748 (O_1748,N_19914,N_19911);
nand UO_1749 (O_1749,N_19958,N_19943);
xor UO_1750 (O_1750,N_19950,N_19884);
or UO_1751 (O_1751,N_19861,N_19949);
or UO_1752 (O_1752,N_19991,N_19960);
xnor UO_1753 (O_1753,N_19865,N_19987);
nand UO_1754 (O_1754,N_19977,N_19924);
nor UO_1755 (O_1755,N_19842,N_19992);
nand UO_1756 (O_1756,N_19850,N_19894);
nand UO_1757 (O_1757,N_19878,N_19961);
nand UO_1758 (O_1758,N_19850,N_19877);
xnor UO_1759 (O_1759,N_19841,N_19906);
xor UO_1760 (O_1760,N_19878,N_19960);
nor UO_1761 (O_1761,N_19977,N_19916);
or UO_1762 (O_1762,N_19901,N_19903);
xnor UO_1763 (O_1763,N_19944,N_19900);
or UO_1764 (O_1764,N_19951,N_19937);
xor UO_1765 (O_1765,N_19939,N_19849);
nand UO_1766 (O_1766,N_19974,N_19924);
xnor UO_1767 (O_1767,N_19867,N_19902);
xnor UO_1768 (O_1768,N_19950,N_19998);
and UO_1769 (O_1769,N_19895,N_19981);
nand UO_1770 (O_1770,N_19990,N_19946);
and UO_1771 (O_1771,N_19985,N_19841);
and UO_1772 (O_1772,N_19941,N_19890);
xor UO_1773 (O_1773,N_19851,N_19940);
xor UO_1774 (O_1774,N_19930,N_19949);
and UO_1775 (O_1775,N_19928,N_19874);
and UO_1776 (O_1776,N_19847,N_19863);
nand UO_1777 (O_1777,N_19954,N_19868);
and UO_1778 (O_1778,N_19934,N_19950);
xnor UO_1779 (O_1779,N_19874,N_19900);
nand UO_1780 (O_1780,N_19851,N_19973);
or UO_1781 (O_1781,N_19968,N_19924);
or UO_1782 (O_1782,N_19968,N_19921);
nor UO_1783 (O_1783,N_19849,N_19987);
xnor UO_1784 (O_1784,N_19882,N_19895);
and UO_1785 (O_1785,N_19915,N_19977);
or UO_1786 (O_1786,N_19911,N_19857);
xor UO_1787 (O_1787,N_19985,N_19953);
or UO_1788 (O_1788,N_19861,N_19962);
xnor UO_1789 (O_1789,N_19904,N_19980);
nand UO_1790 (O_1790,N_19842,N_19920);
xnor UO_1791 (O_1791,N_19930,N_19989);
nand UO_1792 (O_1792,N_19903,N_19967);
nor UO_1793 (O_1793,N_19999,N_19929);
xnor UO_1794 (O_1794,N_19979,N_19954);
nor UO_1795 (O_1795,N_19984,N_19844);
and UO_1796 (O_1796,N_19967,N_19879);
and UO_1797 (O_1797,N_19986,N_19909);
and UO_1798 (O_1798,N_19890,N_19994);
nor UO_1799 (O_1799,N_19988,N_19993);
xor UO_1800 (O_1800,N_19904,N_19994);
nor UO_1801 (O_1801,N_19993,N_19938);
nor UO_1802 (O_1802,N_19913,N_19976);
nand UO_1803 (O_1803,N_19979,N_19862);
or UO_1804 (O_1804,N_19993,N_19926);
xor UO_1805 (O_1805,N_19970,N_19959);
or UO_1806 (O_1806,N_19995,N_19986);
xnor UO_1807 (O_1807,N_19997,N_19973);
or UO_1808 (O_1808,N_19852,N_19870);
and UO_1809 (O_1809,N_19959,N_19900);
nor UO_1810 (O_1810,N_19853,N_19923);
nor UO_1811 (O_1811,N_19940,N_19918);
xnor UO_1812 (O_1812,N_19958,N_19889);
or UO_1813 (O_1813,N_19880,N_19843);
and UO_1814 (O_1814,N_19991,N_19966);
and UO_1815 (O_1815,N_19862,N_19967);
nand UO_1816 (O_1816,N_19874,N_19935);
xnor UO_1817 (O_1817,N_19977,N_19910);
nand UO_1818 (O_1818,N_19879,N_19852);
and UO_1819 (O_1819,N_19986,N_19849);
and UO_1820 (O_1820,N_19964,N_19988);
nor UO_1821 (O_1821,N_19981,N_19844);
nand UO_1822 (O_1822,N_19959,N_19873);
xnor UO_1823 (O_1823,N_19955,N_19934);
and UO_1824 (O_1824,N_19884,N_19971);
nor UO_1825 (O_1825,N_19963,N_19961);
or UO_1826 (O_1826,N_19915,N_19854);
and UO_1827 (O_1827,N_19882,N_19869);
nand UO_1828 (O_1828,N_19931,N_19891);
nor UO_1829 (O_1829,N_19947,N_19995);
nand UO_1830 (O_1830,N_19984,N_19926);
and UO_1831 (O_1831,N_19981,N_19894);
nor UO_1832 (O_1832,N_19938,N_19913);
nor UO_1833 (O_1833,N_19847,N_19982);
or UO_1834 (O_1834,N_19962,N_19999);
nor UO_1835 (O_1835,N_19955,N_19982);
xnor UO_1836 (O_1836,N_19858,N_19843);
xnor UO_1837 (O_1837,N_19982,N_19859);
and UO_1838 (O_1838,N_19997,N_19982);
nand UO_1839 (O_1839,N_19982,N_19858);
xnor UO_1840 (O_1840,N_19861,N_19936);
or UO_1841 (O_1841,N_19851,N_19872);
and UO_1842 (O_1842,N_19983,N_19979);
xor UO_1843 (O_1843,N_19918,N_19944);
nor UO_1844 (O_1844,N_19975,N_19974);
nor UO_1845 (O_1845,N_19984,N_19873);
nand UO_1846 (O_1846,N_19867,N_19953);
nor UO_1847 (O_1847,N_19965,N_19903);
and UO_1848 (O_1848,N_19937,N_19973);
or UO_1849 (O_1849,N_19981,N_19930);
nand UO_1850 (O_1850,N_19983,N_19857);
or UO_1851 (O_1851,N_19888,N_19919);
nor UO_1852 (O_1852,N_19893,N_19858);
nand UO_1853 (O_1853,N_19924,N_19860);
and UO_1854 (O_1854,N_19936,N_19856);
or UO_1855 (O_1855,N_19906,N_19854);
or UO_1856 (O_1856,N_19890,N_19894);
nand UO_1857 (O_1857,N_19990,N_19996);
nor UO_1858 (O_1858,N_19932,N_19999);
xor UO_1859 (O_1859,N_19937,N_19864);
nor UO_1860 (O_1860,N_19947,N_19917);
or UO_1861 (O_1861,N_19888,N_19864);
nand UO_1862 (O_1862,N_19920,N_19939);
xnor UO_1863 (O_1863,N_19909,N_19841);
nor UO_1864 (O_1864,N_19973,N_19958);
nand UO_1865 (O_1865,N_19874,N_19945);
or UO_1866 (O_1866,N_19882,N_19870);
and UO_1867 (O_1867,N_19856,N_19901);
nor UO_1868 (O_1868,N_19982,N_19931);
nor UO_1869 (O_1869,N_19859,N_19919);
or UO_1870 (O_1870,N_19848,N_19999);
or UO_1871 (O_1871,N_19958,N_19938);
nor UO_1872 (O_1872,N_19983,N_19874);
or UO_1873 (O_1873,N_19949,N_19976);
or UO_1874 (O_1874,N_19862,N_19972);
nor UO_1875 (O_1875,N_19965,N_19904);
or UO_1876 (O_1876,N_19962,N_19944);
nand UO_1877 (O_1877,N_19982,N_19942);
nor UO_1878 (O_1878,N_19930,N_19985);
or UO_1879 (O_1879,N_19842,N_19966);
xnor UO_1880 (O_1880,N_19867,N_19970);
and UO_1881 (O_1881,N_19870,N_19936);
nand UO_1882 (O_1882,N_19897,N_19924);
nor UO_1883 (O_1883,N_19860,N_19917);
xor UO_1884 (O_1884,N_19977,N_19938);
nand UO_1885 (O_1885,N_19891,N_19973);
nor UO_1886 (O_1886,N_19908,N_19912);
xnor UO_1887 (O_1887,N_19899,N_19998);
and UO_1888 (O_1888,N_19907,N_19999);
nand UO_1889 (O_1889,N_19983,N_19978);
nor UO_1890 (O_1890,N_19840,N_19878);
and UO_1891 (O_1891,N_19891,N_19976);
or UO_1892 (O_1892,N_19943,N_19939);
nor UO_1893 (O_1893,N_19878,N_19875);
or UO_1894 (O_1894,N_19875,N_19994);
or UO_1895 (O_1895,N_19933,N_19964);
and UO_1896 (O_1896,N_19841,N_19857);
or UO_1897 (O_1897,N_19881,N_19913);
and UO_1898 (O_1898,N_19959,N_19913);
and UO_1899 (O_1899,N_19971,N_19977);
and UO_1900 (O_1900,N_19945,N_19925);
nor UO_1901 (O_1901,N_19975,N_19846);
and UO_1902 (O_1902,N_19997,N_19911);
or UO_1903 (O_1903,N_19910,N_19974);
and UO_1904 (O_1904,N_19892,N_19984);
nor UO_1905 (O_1905,N_19956,N_19959);
nor UO_1906 (O_1906,N_19892,N_19867);
or UO_1907 (O_1907,N_19844,N_19877);
nor UO_1908 (O_1908,N_19912,N_19948);
or UO_1909 (O_1909,N_19909,N_19970);
nand UO_1910 (O_1910,N_19926,N_19936);
nor UO_1911 (O_1911,N_19845,N_19884);
xnor UO_1912 (O_1912,N_19930,N_19875);
or UO_1913 (O_1913,N_19896,N_19976);
xor UO_1914 (O_1914,N_19977,N_19983);
nor UO_1915 (O_1915,N_19917,N_19944);
nand UO_1916 (O_1916,N_19855,N_19852);
or UO_1917 (O_1917,N_19939,N_19959);
and UO_1918 (O_1918,N_19972,N_19899);
and UO_1919 (O_1919,N_19907,N_19896);
and UO_1920 (O_1920,N_19897,N_19926);
nor UO_1921 (O_1921,N_19920,N_19961);
and UO_1922 (O_1922,N_19927,N_19898);
xnor UO_1923 (O_1923,N_19955,N_19996);
nand UO_1924 (O_1924,N_19952,N_19840);
and UO_1925 (O_1925,N_19933,N_19962);
nand UO_1926 (O_1926,N_19859,N_19992);
xor UO_1927 (O_1927,N_19981,N_19984);
nor UO_1928 (O_1928,N_19860,N_19864);
xor UO_1929 (O_1929,N_19947,N_19931);
and UO_1930 (O_1930,N_19968,N_19897);
and UO_1931 (O_1931,N_19895,N_19901);
xor UO_1932 (O_1932,N_19913,N_19861);
and UO_1933 (O_1933,N_19944,N_19921);
or UO_1934 (O_1934,N_19865,N_19941);
nor UO_1935 (O_1935,N_19913,N_19962);
nand UO_1936 (O_1936,N_19993,N_19974);
or UO_1937 (O_1937,N_19922,N_19992);
nor UO_1938 (O_1938,N_19957,N_19848);
xnor UO_1939 (O_1939,N_19948,N_19985);
and UO_1940 (O_1940,N_19942,N_19910);
or UO_1941 (O_1941,N_19887,N_19885);
nand UO_1942 (O_1942,N_19869,N_19853);
nand UO_1943 (O_1943,N_19950,N_19994);
nor UO_1944 (O_1944,N_19932,N_19867);
or UO_1945 (O_1945,N_19865,N_19947);
or UO_1946 (O_1946,N_19890,N_19876);
nor UO_1947 (O_1947,N_19995,N_19990);
xor UO_1948 (O_1948,N_19968,N_19873);
nand UO_1949 (O_1949,N_19900,N_19840);
nor UO_1950 (O_1950,N_19865,N_19951);
or UO_1951 (O_1951,N_19855,N_19961);
or UO_1952 (O_1952,N_19929,N_19945);
nor UO_1953 (O_1953,N_19841,N_19860);
and UO_1954 (O_1954,N_19849,N_19850);
xnor UO_1955 (O_1955,N_19946,N_19882);
or UO_1956 (O_1956,N_19900,N_19957);
nor UO_1957 (O_1957,N_19961,N_19901);
nand UO_1958 (O_1958,N_19887,N_19857);
nor UO_1959 (O_1959,N_19966,N_19997);
nor UO_1960 (O_1960,N_19877,N_19994);
and UO_1961 (O_1961,N_19988,N_19999);
or UO_1962 (O_1962,N_19965,N_19930);
and UO_1963 (O_1963,N_19857,N_19920);
nand UO_1964 (O_1964,N_19960,N_19908);
xnor UO_1965 (O_1965,N_19970,N_19984);
nor UO_1966 (O_1966,N_19978,N_19934);
or UO_1967 (O_1967,N_19979,N_19912);
xor UO_1968 (O_1968,N_19997,N_19956);
xor UO_1969 (O_1969,N_19987,N_19858);
and UO_1970 (O_1970,N_19873,N_19902);
or UO_1971 (O_1971,N_19963,N_19957);
nor UO_1972 (O_1972,N_19928,N_19972);
xor UO_1973 (O_1973,N_19965,N_19962);
xnor UO_1974 (O_1974,N_19973,N_19843);
xor UO_1975 (O_1975,N_19927,N_19861);
or UO_1976 (O_1976,N_19874,N_19880);
and UO_1977 (O_1977,N_19988,N_19976);
or UO_1978 (O_1978,N_19936,N_19853);
or UO_1979 (O_1979,N_19924,N_19936);
or UO_1980 (O_1980,N_19935,N_19934);
and UO_1981 (O_1981,N_19847,N_19842);
or UO_1982 (O_1982,N_19862,N_19984);
xnor UO_1983 (O_1983,N_19911,N_19866);
or UO_1984 (O_1984,N_19970,N_19966);
nor UO_1985 (O_1985,N_19993,N_19932);
nand UO_1986 (O_1986,N_19882,N_19964);
or UO_1987 (O_1987,N_19933,N_19939);
and UO_1988 (O_1988,N_19948,N_19953);
and UO_1989 (O_1989,N_19981,N_19905);
nand UO_1990 (O_1990,N_19859,N_19984);
or UO_1991 (O_1991,N_19856,N_19977);
nor UO_1992 (O_1992,N_19858,N_19943);
and UO_1993 (O_1993,N_19852,N_19932);
and UO_1994 (O_1994,N_19928,N_19859);
and UO_1995 (O_1995,N_19896,N_19991);
xor UO_1996 (O_1996,N_19883,N_19960);
xnor UO_1997 (O_1997,N_19999,N_19850);
and UO_1998 (O_1998,N_19932,N_19910);
and UO_1999 (O_1999,N_19994,N_19936);
nor UO_2000 (O_2000,N_19879,N_19854);
xor UO_2001 (O_2001,N_19846,N_19930);
or UO_2002 (O_2002,N_19935,N_19900);
and UO_2003 (O_2003,N_19852,N_19927);
nor UO_2004 (O_2004,N_19939,N_19870);
xor UO_2005 (O_2005,N_19945,N_19865);
nand UO_2006 (O_2006,N_19883,N_19853);
nor UO_2007 (O_2007,N_19909,N_19911);
and UO_2008 (O_2008,N_19927,N_19997);
nand UO_2009 (O_2009,N_19963,N_19915);
xor UO_2010 (O_2010,N_19990,N_19910);
or UO_2011 (O_2011,N_19858,N_19872);
nand UO_2012 (O_2012,N_19868,N_19881);
nor UO_2013 (O_2013,N_19916,N_19864);
xor UO_2014 (O_2014,N_19975,N_19885);
nor UO_2015 (O_2015,N_19935,N_19948);
nand UO_2016 (O_2016,N_19921,N_19875);
xor UO_2017 (O_2017,N_19922,N_19953);
nor UO_2018 (O_2018,N_19859,N_19926);
or UO_2019 (O_2019,N_19902,N_19897);
and UO_2020 (O_2020,N_19863,N_19932);
or UO_2021 (O_2021,N_19932,N_19978);
nor UO_2022 (O_2022,N_19880,N_19925);
xnor UO_2023 (O_2023,N_19976,N_19842);
and UO_2024 (O_2024,N_19858,N_19974);
or UO_2025 (O_2025,N_19877,N_19860);
and UO_2026 (O_2026,N_19952,N_19980);
and UO_2027 (O_2027,N_19914,N_19992);
and UO_2028 (O_2028,N_19950,N_19943);
nand UO_2029 (O_2029,N_19933,N_19904);
or UO_2030 (O_2030,N_19852,N_19876);
nor UO_2031 (O_2031,N_19848,N_19842);
and UO_2032 (O_2032,N_19853,N_19968);
xnor UO_2033 (O_2033,N_19873,N_19971);
or UO_2034 (O_2034,N_19847,N_19992);
xnor UO_2035 (O_2035,N_19870,N_19909);
nand UO_2036 (O_2036,N_19997,N_19919);
nor UO_2037 (O_2037,N_19962,N_19989);
and UO_2038 (O_2038,N_19969,N_19855);
nor UO_2039 (O_2039,N_19964,N_19851);
nand UO_2040 (O_2040,N_19862,N_19898);
or UO_2041 (O_2041,N_19862,N_19860);
nand UO_2042 (O_2042,N_19963,N_19876);
nor UO_2043 (O_2043,N_19924,N_19941);
and UO_2044 (O_2044,N_19856,N_19945);
xnor UO_2045 (O_2045,N_19899,N_19916);
nand UO_2046 (O_2046,N_19992,N_19866);
or UO_2047 (O_2047,N_19849,N_19925);
or UO_2048 (O_2048,N_19879,N_19993);
xor UO_2049 (O_2049,N_19956,N_19937);
xnor UO_2050 (O_2050,N_19991,N_19933);
xnor UO_2051 (O_2051,N_19986,N_19996);
or UO_2052 (O_2052,N_19954,N_19932);
nand UO_2053 (O_2053,N_19987,N_19890);
or UO_2054 (O_2054,N_19988,N_19851);
nand UO_2055 (O_2055,N_19922,N_19989);
nand UO_2056 (O_2056,N_19934,N_19889);
nor UO_2057 (O_2057,N_19976,N_19877);
nor UO_2058 (O_2058,N_19924,N_19960);
and UO_2059 (O_2059,N_19847,N_19894);
xnor UO_2060 (O_2060,N_19901,N_19885);
xnor UO_2061 (O_2061,N_19968,N_19975);
or UO_2062 (O_2062,N_19928,N_19924);
nand UO_2063 (O_2063,N_19864,N_19934);
or UO_2064 (O_2064,N_19887,N_19918);
nand UO_2065 (O_2065,N_19856,N_19929);
or UO_2066 (O_2066,N_19877,N_19961);
nand UO_2067 (O_2067,N_19851,N_19934);
xor UO_2068 (O_2068,N_19847,N_19941);
nor UO_2069 (O_2069,N_19846,N_19842);
xor UO_2070 (O_2070,N_19998,N_19941);
and UO_2071 (O_2071,N_19889,N_19869);
and UO_2072 (O_2072,N_19914,N_19951);
and UO_2073 (O_2073,N_19849,N_19865);
nor UO_2074 (O_2074,N_19898,N_19986);
xor UO_2075 (O_2075,N_19870,N_19887);
and UO_2076 (O_2076,N_19908,N_19975);
and UO_2077 (O_2077,N_19906,N_19995);
xor UO_2078 (O_2078,N_19915,N_19971);
or UO_2079 (O_2079,N_19978,N_19925);
xor UO_2080 (O_2080,N_19893,N_19932);
nor UO_2081 (O_2081,N_19867,N_19896);
xnor UO_2082 (O_2082,N_19964,N_19941);
xnor UO_2083 (O_2083,N_19976,N_19868);
xor UO_2084 (O_2084,N_19907,N_19969);
or UO_2085 (O_2085,N_19971,N_19907);
and UO_2086 (O_2086,N_19999,N_19992);
nand UO_2087 (O_2087,N_19982,N_19863);
and UO_2088 (O_2088,N_19840,N_19877);
or UO_2089 (O_2089,N_19942,N_19898);
xor UO_2090 (O_2090,N_19888,N_19999);
and UO_2091 (O_2091,N_19889,N_19918);
nand UO_2092 (O_2092,N_19935,N_19967);
nand UO_2093 (O_2093,N_19853,N_19930);
and UO_2094 (O_2094,N_19866,N_19983);
xor UO_2095 (O_2095,N_19847,N_19858);
nand UO_2096 (O_2096,N_19851,N_19949);
and UO_2097 (O_2097,N_19967,N_19870);
and UO_2098 (O_2098,N_19939,N_19848);
nand UO_2099 (O_2099,N_19848,N_19956);
and UO_2100 (O_2100,N_19925,N_19961);
or UO_2101 (O_2101,N_19931,N_19914);
nand UO_2102 (O_2102,N_19985,N_19902);
and UO_2103 (O_2103,N_19888,N_19878);
or UO_2104 (O_2104,N_19924,N_19886);
and UO_2105 (O_2105,N_19865,N_19988);
xnor UO_2106 (O_2106,N_19884,N_19930);
nor UO_2107 (O_2107,N_19887,N_19897);
and UO_2108 (O_2108,N_19914,N_19939);
or UO_2109 (O_2109,N_19945,N_19975);
nor UO_2110 (O_2110,N_19855,N_19943);
nor UO_2111 (O_2111,N_19842,N_19913);
nor UO_2112 (O_2112,N_19927,N_19949);
xor UO_2113 (O_2113,N_19904,N_19847);
or UO_2114 (O_2114,N_19986,N_19992);
or UO_2115 (O_2115,N_19971,N_19975);
or UO_2116 (O_2116,N_19986,N_19885);
nor UO_2117 (O_2117,N_19918,N_19998);
nor UO_2118 (O_2118,N_19963,N_19857);
or UO_2119 (O_2119,N_19945,N_19843);
nand UO_2120 (O_2120,N_19874,N_19882);
or UO_2121 (O_2121,N_19881,N_19970);
and UO_2122 (O_2122,N_19896,N_19912);
and UO_2123 (O_2123,N_19951,N_19840);
xnor UO_2124 (O_2124,N_19943,N_19982);
nor UO_2125 (O_2125,N_19904,N_19982);
xnor UO_2126 (O_2126,N_19956,N_19943);
and UO_2127 (O_2127,N_19955,N_19888);
and UO_2128 (O_2128,N_19863,N_19953);
nand UO_2129 (O_2129,N_19950,N_19909);
and UO_2130 (O_2130,N_19925,N_19934);
nand UO_2131 (O_2131,N_19934,N_19860);
or UO_2132 (O_2132,N_19853,N_19959);
xor UO_2133 (O_2133,N_19910,N_19856);
or UO_2134 (O_2134,N_19971,N_19927);
nand UO_2135 (O_2135,N_19958,N_19890);
xnor UO_2136 (O_2136,N_19931,N_19971);
nor UO_2137 (O_2137,N_19885,N_19946);
and UO_2138 (O_2138,N_19963,N_19919);
or UO_2139 (O_2139,N_19855,N_19934);
nand UO_2140 (O_2140,N_19842,N_19940);
nand UO_2141 (O_2141,N_19870,N_19869);
or UO_2142 (O_2142,N_19895,N_19891);
nand UO_2143 (O_2143,N_19876,N_19886);
or UO_2144 (O_2144,N_19901,N_19894);
nor UO_2145 (O_2145,N_19879,N_19864);
or UO_2146 (O_2146,N_19978,N_19856);
and UO_2147 (O_2147,N_19857,N_19921);
and UO_2148 (O_2148,N_19943,N_19874);
nand UO_2149 (O_2149,N_19870,N_19979);
xor UO_2150 (O_2150,N_19860,N_19945);
nand UO_2151 (O_2151,N_19872,N_19924);
nand UO_2152 (O_2152,N_19909,N_19961);
nor UO_2153 (O_2153,N_19968,N_19949);
nand UO_2154 (O_2154,N_19998,N_19862);
and UO_2155 (O_2155,N_19914,N_19909);
or UO_2156 (O_2156,N_19869,N_19982);
nor UO_2157 (O_2157,N_19848,N_19961);
or UO_2158 (O_2158,N_19924,N_19889);
nor UO_2159 (O_2159,N_19852,N_19995);
nand UO_2160 (O_2160,N_19984,N_19869);
or UO_2161 (O_2161,N_19934,N_19847);
nor UO_2162 (O_2162,N_19910,N_19948);
nand UO_2163 (O_2163,N_19855,N_19987);
xor UO_2164 (O_2164,N_19973,N_19967);
and UO_2165 (O_2165,N_19883,N_19906);
xor UO_2166 (O_2166,N_19963,N_19850);
nand UO_2167 (O_2167,N_19893,N_19926);
and UO_2168 (O_2168,N_19910,N_19995);
nor UO_2169 (O_2169,N_19966,N_19898);
nand UO_2170 (O_2170,N_19879,N_19867);
and UO_2171 (O_2171,N_19850,N_19993);
or UO_2172 (O_2172,N_19920,N_19846);
or UO_2173 (O_2173,N_19905,N_19952);
nand UO_2174 (O_2174,N_19931,N_19899);
nand UO_2175 (O_2175,N_19995,N_19849);
nand UO_2176 (O_2176,N_19898,N_19867);
xor UO_2177 (O_2177,N_19979,N_19927);
nor UO_2178 (O_2178,N_19877,N_19986);
and UO_2179 (O_2179,N_19859,N_19951);
and UO_2180 (O_2180,N_19960,N_19858);
and UO_2181 (O_2181,N_19852,N_19959);
nand UO_2182 (O_2182,N_19887,N_19928);
and UO_2183 (O_2183,N_19969,N_19947);
nand UO_2184 (O_2184,N_19916,N_19929);
xnor UO_2185 (O_2185,N_19990,N_19844);
nand UO_2186 (O_2186,N_19868,N_19953);
xnor UO_2187 (O_2187,N_19928,N_19933);
nand UO_2188 (O_2188,N_19982,N_19888);
and UO_2189 (O_2189,N_19963,N_19884);
and UO_2190 (O_2190,N_19919,N_19940);
nor UO_2191 (O_2191,N_19990,N_19923);
nor UO_2192 (O_2192,N_19901,N_19995);
nor UO_2193 (O_2193,N_19955,N_19845);
or UO_2194 (O_2194,N_19964,N_19881);
nor UO_2195 (O_2195,N_19989,N_19857);
or UO_2196 (O_2196,N_19928,N_19906);
nand UO_2197 (O_2197,N_19957,N_19953);
nor UO_2198 (O_2198,N_19996,N_19907);
nand UO_2199 (O_2199,N_19868,N_19854);
or UO_2200 (O_2200,N_19896,N_19959);
or UO_2201 (O_2201,N_19875,N_19951);
nand UO_2202 (O_2202,N_19850,N_19954);
or UO_2203 (O_2203,N_19963,N_19902);
nor UO_2204 (O_2204,N_19846,N_19991);
xor UO_2205 (O_2205,N_19884,N_19886);
xor UO_2206 (O_2206,N_19935,N_19992);
xor UO_2207 (O_2207,N_19919,N_19972);
and UO_2208 (O_2208,N_19855,N_19887);
nor UO_2209 (O_2209,N_19907,N_19931);
nand UO_2210 (O_2210,N_19979,N_19945);
nor UO_2211 (O_2211,N_19938,N_19925);
xnor UO_2212 (O_2212,N_19966,N_19848);
nand UO_2213 (O_2213,N_19875,N_19915);
or UO_2214 (O_2214,N_19871,N_19998);
and UO_2215 (O_2215,N_19855,N_19917);
or UO_2216 (O_2216,N_19989,N_19993);
nor UO_2217 (O_2217,N_19956,N_19847);
nor UO_2218 (O_2218,N_19995,N_19937);
and UO_2219 (O_2219,N_19980,N_19910);
xor UO_2220 (O_2220,N_19898,N_19960);
and UO_2221 (O_2221,N_19995,N_19929);
xnor UO_2222 (O_2222,N_19885,N_19951);
or UO_2223 (O_2223,N_19846,N_19876);
xor UO_2224 (O_2224,N_19982,N_19953);
nand UO_2225 (O_2225,N_19954,N_19910);
nor UO_2226 (O_2226,N_19954,N_19912);
and UO_2227 (O_2227,N_19886,N_19921);
xnor UO_2228 (O_2228,N_19941,N_19985);
nor UO_2229 (O_2229,N_19841,N_19900);
or UO_2230 (O_2230,N_19872,N_19860);
or UO_2231 (O_2231,N_19948,N_19905);
nand UO_2232 (O_2232,N_19978,N_19920);
or UO_2233 (O_2233,N_19992,N_19893);
and UO_2234 (O_2234,N_19858,N_19940);
nor UO_2235 (O_2235,N_19984,N_19930);
xnor UO_2236 (O_2236,N_19870,N_19841);
nand UO_2237 (O_2237,N_19843,N_19879);
xnor UO_2238 (O_2238,N_19885,N_19962);
or UO_2239 (O_2239,N_19959,N_19978);
xnor UO_2240 (O_2240,N_19886,N_19933);
or UO_2241 (O_2241,N_19877,N_19903);
and UO_2242 (O_2242,N_19900,N_19922);
nand UO_2243 (O_2243,N_19929,N_19931);
nor UO_2244 (O_2244,N_19892,N_19979);
xor UO_2245 (O_2245,N_19953,N_19855);
nand UO_2246 (O_2246,N_19869,N_19952);
and UO_2247 (O_2247,N_19882,N_19900);
nor UO_2248 (O_2248,N_19863,N_19918);
xor UO_2249 (O_2249,N_19952,N_19897);
and UO_2250 (O_2250,N_19840,N_19844);
nor UO_2251 (O_2251,N_19878,N_19963);
nor UO_2252 (O_2252,N_19923,N_19904);
or UO_2253 (O_2253,N_19895,N_19899);
xnor UO_2254 (O_2254,N_19893,N_19944);
nand UO_2255 (O_2255,N_19987,N_19921);
xor UO_2256 (O_2256,N_19990,N_19975);
xor UO_2257 (O_2257,N_19993,N_19884);
xor UO_2258 (O_2258,N_19845,N_19857);
and UO_2259 (O_2259,N_19877,N_19943);
or UO_2260 (O_2260,N_19852,N_19942);
xor UO_2261 (O_2261,N_19853,N_19874);
xor UO_2262 (O_2262,N_19904,N_19916);
and UO_2263 (O_2263,N_19880,N_19976);
xor UO_2264 (O_2264,N_19941,N_19975);
nand UO_2265 (O_2265,N_19972,N_19901);
and UO_2266 (O_2266,N_19883,N_19953);
or UO_2267 (O_2267,N_19924,N_19988);
or UO_2268 (O_2268,N_19872,N_19932);
nand UO_2269 (O_2269,N_19889,N_19902);
and UO_2270 (O_2270,N_19968,N_19888);
and UO_2271 (O_2271,N_19912,N_19960);
or UO_2272 (O_2272,N_19901,N_19863);
and UO_2273 (O_2273,N_19947,N_19951);
or UO_2274 (O_2274,N_19945,N_19955);
xnor UO_2275 (O_2275,N_19928,N_19998);
nand UO_2276 (O_2276,N_19932,N_19958);
xnor UO_2277 (O_2277,N_19889,N_19950);
nand UO_2278 (O_2278,N_19863,N_19879);
nor UO_2279 (O_2279,N_19963,N_19980);
nor UO_2280 (O_2280,N_19853,N_19937);
nor UO_2281 (O_2281,N_19886,N_19971);
and UO_2282 (O_2282,N_19998,N_19974);
or UO_2283 (O_2283,N_19993,N_19961);
xnor UO_2284 (O_2284,N_19995,N_19936);
nand UO_2285 (O_2285,N_19874,N_19994);
nor UO_2286 (O_2286,N_19959,N_19936);
or UO_2287 (O_2287,N_19890,N_19926);
and UO_2288 (O_2288,N_19991,N_19928);
and UO_2289 (O_2289,N_19997,N_19955);
nor UO_2290 (O_2290,N_19884,N_19953);
and UO_2291 (O_2291,N_19897,N_19877);
nor UO_2292 (O_2292,N_19941,N_19842);
or UO_2293 (O_2293,N_19980,N_19997);
nor UO_2294 (O_2294,N_19848,N_19950);
nand UO_2295 (O_2295,N_19921,N_19995);
or UO_2296 (O_2296,N_19958,N_19905);
nor UO_2297 (O_2297,N_19844,N_19875);
nor UO_2298 (O_2298,N_19992,N_19875);
nor UO_2299 (O_2299,N_19911,N_19966);
and UO_2300 (O_2300,N_19880,N_19940);
nor UO_2301 (O_2301,N_19947,N_19856);
and UO_2302 (O_2302,N_19931,N_19960);
or UO_2303 (O_2303,N_19972,N_19864);
nand UO_2304 (O_2304,N_19945,N_19868);
xor UO_2305 (O_2305,N_19840,N_19909);
and UO_2306 (O_2306,N_19860,N_19844);
and UO_2307 (O_2307,N_19919,N_19945);
xnor UO_2308 (O_2308,N_19876,N_19992);
or UO_2309 (O_2309,N_19847,N_19948);
nor UO_2310 (O_2310,N_19841,N_19961);
and UO_2311 (O_2311,N_19905,N_19974);
xnor UO_2312 (O_2312,N_19915,N_19982);
nor UO_2313 (O_2313,N_19879,N_19940);
and UO_2314 (O_2314,N_19915,N_19882);
or UO_2315 (O_2315,N_19889,N_19891);
or UO_2316 (O_2316,N_19915,N_19862);
nand UO_2317 (O_2317,N_19980,N_19899);
and UO_2318 (O_2318,N_19942,N_19863);
nor UO_2319 (O_2319,N_19857,N_19998);
nor UO_2320 (O_2320,N_19863,N_19955);
nor UO_2321 (O_2321,N_19924,N_19934);
or UO_2322 (O_2322,N_19841,N_19946);
nor UO_2323 (O_2323,N_19854,N_19883);
xnor UO_2324 (O_2324,N_19863,N_19949);
nand UO_2325 (O_2325,N_19862,N_19854);
and UO_2326 (O_2326,N_19912,N_19971);
or UO_2327 (O_2327,N_19879,N_19891);
nor UO_2328 (O_2328,N_19955,N_19941);
nor UO_2329 (O_2329,N_19856,N_19999);
nor UO_2330 (O_2330,N_19994,N_19907);
nor UO_2331 (O_2331,N_19993,N_19970);
and UO_2332 (O_2332,N_19881,N_19995);
nor UO_2333 (O_2333,N_19908,N_19849);
nand UO_2334 (O_2334,N_19998,N_19984);
nand UO_2335 (O_2335,N_19899,N_19915);
nor UO_2336 (O_2336,N_19884,N_19947);
nor UO_2337 (O_2337,N_19842,N_19844);
or UO_2338 (O_2338,N_19889,N_19979);
xor UO_2339 (O_2339,N_19951,N_19934);
nor UO_2340 (O_2340,N_19850,N_19862);
and UO_2341 (O_2341,N_19861,N_19979);
and UO_2342 (O_2342,N_19936,N_19906);
nor UO_2343 (O_2343,N_19960,N_19971);
and UO_2344 (O_2344,N_19953,N_19981);
nor UO_2345 (O_2345,N_19846,N_19959);
xnor UO_2346 (O_2346,N_19844,N_19879);
xor UO_2347 (O_2347,N_19983,N_19865);
and UO_2348 (O_2348,N_19940,N_19973);
and UO_2349 (O_2349,N_19913,N_19928);
xor UO_2350 (O_2350,N_19859,N_19884);
or UO_2351 (O_2351,N_19931,N_19900);
nand UO_2352 (O_2352,N_19856,N_19883);
or UO_2353 (O_2353,N_19919,N_19953);
xnor UO_2354 (O_2354,N_19993,N_19889);
or UO_2355 (O_2355,N_19868,N_19932);
nor UO_2356 (O_2356,N_19942,N_19952);
nand UO_2357 (O_2357,N_19853,N_19982);
xor UO_2358 (O_2358,N_19937,N_19967);
nand UO_2359 (O_2359,N_19998,N_19841);
xnor UO_2360 (O_2360,N_19958,N_19852);
nand UO_2361 (O_2361,N_19856,N_19861);
or UO_2362 (O_2362,N_19937,N_19919);
xnor UO_2363 (O_2363,N_19979,N_19883);
and UO_2364 (O_2364,N_19973,N_19946);
nand UO_2365 (O_2365,N_19966,N_19914);
nor UO_2366 (O_2366,N_19984,N_19951);
xnor UO_2367 (O_2367,N_19925,N_19898);
nor UO_2368 (O_2368,N_19999,N_19989);
and UO_2369 (O_2369,N_19856,N_19857);
nand UO_2370 (O_2370,N_19898,N_19995);
nor UO_2371 (O_2371,N_19920,N_19994);
nand UO_2372 (O_2372,N_19908,N_19878);
or UO_2373 (O_2373,N_19933,N_19875);
and UO_2374 (O_2374,N_19950,N_19842);
and UO_2375 (O_2375,N_19874,N_19846);
or UO_2376 (O_2376,N_19861,N_19911);
or UO_2377 (O_2377,N_19853,N_19973);
and UO_2378 (O_2378,N_19941,N_19866);
or UO_2379 (O_2379,N_19986,N_19899);
or UO_2380 (O_2380,N_19898,N_19985);
nor UO_2381 (O_2381,N_19901,N_19957);
nand UO_2382 (O_2382,N_19883,N_19932);
and UO_2383 (O_2383,N_19917,N_19979);
and UO_2384 (O_2384,N_19984,N_19936);
or UO_2385 (O_2385,N_19970,N_19903);
and UO_2386 (O_2386,N_19958,N_19896);
or UO_2387 (O_2387,N_19850,N_19948);
nand UO_2388 (O_2388,N_19967,N_19991);
nor UO_2389 (O_2389,N_19946,N_19845);
or UO_2390 (O_2390,N_19937,N_19915);
nand UO_2391 (O_2391,N_19964,N_19945);
or UO_2392 (O_2392,N_19958,N_19872);
and UO_2393 (O_2393,N_19904,N_19966);
or UO_2394 (O_2394,N_19943,N_19868);
or UO_2395 (O_2395,N_19903,N_19933);
xor UO_2396 (O_2396,N_19981,N_19977);
nor UO_2397 (O_2397,N_19961,N_19935);
xor UO_2398 (O_2398,N_19972,N_19842);
nand UO_2399 (O_2399,N_19896,N_19954);
nand UO_2400 (O_2400,N_19966,N_19915);
and UO_2401 (O_2401,N_19840,N_19941);
nand UO_2402 (O_2402,N_19938,N_19984);
nor UO_2403 (O_2403,N_19959,N_19972);
or UO_2404 (O_2404,N_19860,N_19847);
or UO_2405 (O_2405,N_19912,N_19985);
and UO_2406 (O_2406,N_19917,N_19971);
nand UO_2407 (O_2407,N_19878,N_19943);
or UO_2408 (O_2408,N_19944,N_19867);
nor UO_2409 (O_2409,N_19856,N_19919);
or UO_2410 (O_2410,N_19950,N_19882);
and UO_2411 (O_2411,N_19876,N_19953);
nor UO_2412 (O_2412,N_19902,N_19857);
xnor UO_2413 (O_2413,N_19909,N_19999);
or UO_2414 (O_2414,N_19968,N_19967);
nor UO_2415 (O_2415,N_19875,N_19982);
or UO_2416 (O_2416,N_19897,N_19879);
xnor UO_2417 (O_2417,N_19875,N_19973);
nand UO_2418 (O_2418,N_19932,N_19986);
or UO_2419 (O_2419,N_19983,N_19940);
nand UO_2420 (O_2420,N_19883,N_19841);
or UO_2421 (O_2421,N_19871,N_19917);
xor UO_2422 (O_2422,N_19978,N_19965);
xnor UO_2423 (O_2423,N_19855,N_19861);
nor UO_2424 (O_2424,N_19843,N_19874);
xnor UO_2425 (O_2425,N_19901,N_19886);
and UO_2426 (O_2426,N_19984,N_19864);
nand UO_2427 (O_2427,N_19859,N_19901);
and UO_2428 (O_2428,N_19949,N_19988);
or UO_2429 (O_2429,N_19873,N_19943);
nand UO_2430 (O_2430,N_19988,N_19960);
or UO_2431 (O_2431,N_19875,N_19928);
or UO_2432 (O_2432,N_19948,N_19877);
nand UO_2433 (O_2433,N_19913,N_19879);
xor UO_2434 (O_2434,N_19925,N_19841);
nand UO_2435 (O_2435,N_19873,N_19878);
nand UO_2436 (O_2436,N_19858,N_19862);
or UO_2437 (O_2437,N_19922,N_19892);
or UO_2438 (O_2438,N_19892,N_19957);
nor UO_2439 (O_2439,N_19855,N_19964);
and UO_2440 (O_2440,N_19987,N_19866);
or UO_2441 (O_2441,N_19952,N_19857);
xnor UO_2442 (O_2442,N_19880,N_19946);
nand UO_2443 (O_2443,N_19879,N_19855);
nor UO_2444 (O_2444,N_19924,N_19885);
nand UO_2445 (O_2445,N_19877,N_19847);
or UO_2446 (O_2446,N_19847,N_19991);
xor UO_2447 (O_2447,N_19921,N_19895);
and UO_2448 (O_2448,N_19891,N_19871);
nor UO_2449 (O_2449,N_19942,N_19897);
nor UO_2450 (O_2450,N_19954,N_19937);
nand UO_2451 (O_2451,N_19869,N_19935);
nor UO_2452 (O_2452,N_19935,N_19946);
and UO_2453 (O_2453,N_19994,N_19959);
xnor UO_2454 (O_2454,N_19970,N_19888);
nor UO_2455 (O_2455,N_19993,N_19950);
and UO_2456 (O_2456,N_19944,N_19961);
and UO_2457 (O_2457,N_19980,N_19911);
nand UO_2458 (O_2458,N_19861,N_19854);
or UO_2459 (O_2459,N_19968,N_19974);
xor UO_2460 (O_2460,N_19935,N_19901);
nor UO_2461 (O_2461,N_19898,N_19957);
nand UO_2462 (O_2462,N_19929,N_19913);
nor UO_2463 (O_2463,N_19901,N_19915);
nor UO_2464 (O_2464,N_19959,N_19960);
nor UO_2465 (O_2465,N_19984,N_19903);
and UO_2466 (O_2466,N_19847,N_19983);
nor UO_2467 (O_2467,N_19937,N_19840);
nor UO_2468 (O_2468,N_19980,N_19870);
or UO_2469 (O_2469,N_19900,N_19846);
nand UO_2470 (O_2470,N_19894,N_19910);
xor UO_2471 (O_2471,N_19849,N_19989);
xor UO_2472 (O_2472,N_19909,N_19857);
xnor UO_2473 (O_2473,N_19929,N_19860);
nand UO_2474 (O_2474,N_19840,N_19918);
or UO_2475 (O_2475,N_19999,N_19875);
nor UO_2476 (O_2476,N_19845,N_19998);
or UO_2477 (O_2477,N_19864,N_19896);
and UO_2478 (O_2478,N_19987,N_19845);
nand UO_2479 (O_2479,N_19953,N_19927);
or UO_2480 (O_2480,N_19940,N_19841);
and UO_2481 (O_2481,N_19878,N_19976);
or UO_2482 (O_2482,N_19934,N_19971);
or UO_2483 (O_2483,N_19977,N_19887);
or UO_2484 (O_2484,N_19856,N_19968);
and UO_2485 (O_2485,N_19967,N_19976);
and UO_2486 (O_2486,N_19942,N_19841);
xor UO_2487 (O_2487,N_19918,N_19846);
and UO_2488 (O_2488,N_19867,N_19976);
or UO_2489 (O_2489,N_19917,N_19939);
nand UO_2490 (O_2490,N_19951,N_19860);
nand UO_2491 (O_2491,N_19976,N_19997);
nand UO_2492 (O_2492,N_19888,N_19952);
and UO_2493 (O_2493,N_19958,N_19959);
or UO_2494 (O_2494,N_19884,N_19919);
or UO_2495 (O_2495,N_19949,N_19921);
nand UO_2496 (O_2496,N_19973,N_19972);
nand UO_2497 (O_2497,N_19853,N_19983);
xor UO_2498 (O_2498,N_19896,N_19887);
xnor UO_2499 (O_2499,N_19928,N_19968);
endmodule