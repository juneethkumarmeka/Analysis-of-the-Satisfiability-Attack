module basic_2500_25000_3000_40_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_132,In_2167);
nor U1 (N_1,In_1108,In_541);
or U2 (N_2,In_1533,In_148);
nand U3 (N_3,In_842,In_1520);
and U4 (N_4,In_1237,In_884);
nor U5 (N_5,In_445,In_304);
xnor U6 (N_6,In_1889,In_612);
nor U7 (N_7,In_264,In_1503);
nand U8 (N_8,In_1893,In_2438);
or U9 (N_9,In_1225,In_378);
and U10 (N_10,In_1834,In_2051);
nor U11 (N_11,In_620,In_1591);
nand U12 (N_12,In_1551,In_1512);
or U13 (N_13,In_24,In_2221);
and U14 (N_14,In_166,In_513);
xor U15 (N_15,In_2363,In_740);
nor U16 (N_16,In_982,In_1907);
xor U17 (N_17,In_979,In_184);
xor U18 (N_18,In_370,In_2120);
and U19 (N_19,In_2003,In_1660);
nand U20 (N_20,In_593,In_2431);
nand U21 (N_21,In_556,In_443);
xor U22 (N_22,In_806,In_1358);
or U23 (N_23,In_160,In_1273);
and U24 (N_24,In_2397,In_1214);
xor U25 (N_25,In_867,In_1943);
nand U26 (N_26,In_2483,In_877);
and U27 (N_27,In_1836,In_1364);
or U28 (N_28,In_907,In_38);
or U29 (N_29,In_377,In_1190);
nor U30 (N_30,In_2097,In_138);
xnor U31 (N_31,In_1601,In_983);
and U32 (N_32,In_727,In_2172);
nor U33 (N_33,In_515,In_2420);
and U34 (N_34,In_2157,In_150);
nor U35 (N_35,In_274,In_1752);
or U36 (N_36,In_1861,In_598);
nor U37 (N_37,In_1789,In_2008);
and U38 (N_38,In_1847,In_911);
nor U39 (N_39,In_1179,In_2432);
nor U40 (N_40,In_316,In_2465);
and U41 (N_41,In_469,In_2240);
xor U42 (N_42,In_195,In_2133);
nand U43 (N_43,In_325,In_411);
nor U44 (N_44,In_2115,In_668);
or U45 (N_45,In_540,In_1234);
nand U46 (N_46,In_1445,In_2122);
nand U47 (N_47,In_1478,In_1295);
xnor U48 (N_48,In_2213,In_500);
or U49 (N_49,In_152,In_1121);
and U50 (N_50,In_2031,In_348);
nand U51 (N_51,In_2391,In_714);
xnor U52 (N_52,In_1022,In_199);
or U53 (N_53,In_584,In_1288);
xnor U54 (N_54,In_1598,In_2169);
or U55 (N_55,In_203,In_1620);
and U56 (N_56,In_653,In_1914);
or U57 (N_57,In_454,In_8);
nor U58 (N_58,In_1542,In_2360);
xor U59 (N_59,In_2373,In_1338);
or U60 (N_60,In_2000,In_876);
nor U61 (N_61,In_788,In_86);
nand U62 (N_62,In_2152,In_497);
or U63 (N_63,In_546,In_1916);
and U64 (N_64,In_64,In_1386);
xor U65 (N_65,In_1350,In_209);
or U66 (N_66,In_338,In_1267);
or U67 (N_67,In_333,In_1536);
nand U68 (N_68,In_1672,In_1159);
or U69 (N_69,In_853,In_2139);
nand U70 (N_70,In_262,In_1546);
nand U71 (N_71,In_2155,In_2472);
and U72 (N_72,In_2100,In_1053);
nor U73 (N_73,In_2018,In_303);
nor U74 (N_74,In_1815,In_1284);
nand U75 (N_75,In_1770,In_2324);
or U76 (N_76,In_2093,In_782);
nand U77 (N_77,In_1744,In_1149);
nand U78 (N_78,In_464,In_2477);
and U79 (N_79,In_75,In_90);
nor U80 (N_80,In_1946,In_435);
nand U81 (N_81,In_2065,In_349);
nor U82 (N_82,In_1649,In_1263);
or U83 (N_83,In_2058,In_2118);
nor U84 (N_84,In_2022,In_574);
xor U85 (N_85,In_1575,In_1679);
and U86 (N_86,In_923,In_421);
nand U87 (N_87,In_1795,In_226);
nor U88 (N_88,In_1927,In_939);
nand U89 (N_89,In_1710,In_906);
nand U90 (N_90,In_1125,In_1348);
nor U91 (N_91,In_2439,In_1768);
or U92 (N_92,In_1439,In_1504);
xnor U93 (N_93,In_858,In_278);
or U94 (N_94,In_2125,In_1540);
nor U95 (N_95,In_623,In_2173);
xor U96 (N_96,In_1527,In_1655);
nand U97 (N_97,In_1928,In_1608);
nand U98 (N_98,In_1743,In_1972);
and U99 (N_99,In_337,In_1217);
or U100 (N_100,In_1563,In_429);
and U101 (N_101,In_47,In_403);
and U102 (N_102,In_1991,In_996);
or U103 (N_103,In_936,In_2250);
or U104 (N_104,In_1537,In_2239);
and U105 (N_105,In_1185,In_530);
and U106 (N_106,In_1509,In_1457);
and U107 (N_107,In_213,In_775);
nor U108 (N_108,In_2321,In_830);
and U109 (N_109,In_857,In_1957);
nor U110 (N_110,In_657,In_753);
xor U111 (N_111,In_122,In_2182);
xor U112 (N_112,In_467,In_843);
nor U113 (N_113,In_1857,In_1923);
and U114 (N_114,In_1229,In_803);
and U115 (N_115,In_0,In_1161);
and U116 (N_116,In_1039,In_892);
or U117 (N_117,In_124,In_2194);
xnor U118 (N_118,In_528,In_1623);
nand U119 (N_119,In_1393,In_521);
nand U120 (N_120,In_994,In_1290);
or U121 (N_121,In_1103,In_280);
and U122 (N_122,In_297,In_1902);
xor U123 (N_123,In_279,In_437);
xnor U124 (N_124,In_1994,In_660);
nand U125 (N_125,In_1312,In_872);
or U126 (N_126,In_783,In_1633);
or U127 (N_127,In_1055,In_182);
xor U128 (N_128,In_36,In_256);
nor U129 (N_129,In_1280,In_2482);
or U130 (N_130,In_424,In_551);
xnor U131 (N_131,In_1488,In_746);
nor U132 (N_132,In_2,In_1981);
nor U133 (N_133,In_1337,In_2143);
xor U134 (N_134,In_1345,In_960);
or U135 (N_135,In_1332,In_2076);
nand U136 (N_136,In_2318,In_395);
xor U137 (N_137,In_1707,In_1115);
and U138 (N_138,In_733,In_2338);
nand U139 (N_139,In_719,In_1172);
xor U140 (N_140,In_2231,In_1024);
nor U141 (N_141,In_575,In_1549);
nand U142 (N_142,In_364,In_210);
xnor U143 (N_143,In_328,In_96);
nand U144 (N_144,In_852,In_2333);
or U145 (N_145,In_2440,In_1791);
or U146 (N_146,In_1778,In_1316);
and U147 (N_147,In_434,In_807);
xor U148 (N_148,In_369,In_652);
or U149 (N_149,In_120,In_2346);
xnor U150 (N_150,In_1343,In_1147);
and U151 (N_151,In_2303,In_1662);
xnor U152 (N_152,In_933,In_1865);
nand U153 (N_153,In_1557,In_1081);
xnor U154 (N_154,In_975,In_550);
or U155 (N_155,In_1731,In_88);
xor U156 (N_156,In_2208,In_499);
nor U157 (N_157,In_102,In_1614);
and U158 (N_158,In_26,In_2461);
and U159 (N_159,In_760,In_3);
nand U160 (N_160,In_687,In_323);
nand U161 (N_161,In_1028,In_1772);
nor U162 (N_162,In_539,In_365);
or U163 (N_163,In_743,In_744);
xnor U164 (N_164,In_2108,In_2015);
nand U165 (N_165,In_1278,In_2136);
or U166 (N_166,In_1939,In_1429);
and U167 (N_167,In_1440,In_12);
or U168 (N_168,In_1102,In_2343);
nor U169 (N_169,In_1719,In_394);
xor U170 (N_170,In_1049,In_1820);
nor U171 (N_171,In_965,In_1494);
nor U172 (N_172,In_931,In_110);
and U173 (N_173,In_1265,In_2047);
and U174 (N_174,In_1210,In_255);
or U175 (N_175,In_277,In_848);
or U176 (N_176,In_2080,In_1398);
nand U177 (N_177,In_1133,In_639);
nand U178 (N_178,In_180,In_1112);
nor U179 (N_179,In_2301,In_1418);
nor U180 (N_180,In_610,In_17);
and U181 (N_181,In_2029,In_2110);
and U182 (N_182,In_399,In_1019);
nor U183 (N_183,In_1838,In_1286);
xor U184 (N_184,In_459,In_2489);
xor U185 (N_185,In_1687,In_494);
nand U186 (N_186,In_367,In_70);
and U187 (N_187,In_1974,In_1846);
nor U188 (N_188,In_410,In_736);
nand U189 (N_189,In_1232,In_758);
or U190 (N_190,In_1754,In_1841);
and U191 (N_191,In_1835,In_2428);
xor U192 (N_192,In_417,In_1068);
and U193 (N_193,In_2066,In_393);
and U194 (N_194,In_1023,In_1733);
and U195 (N_195,In_973,In_1248);
or U196 (N_196,In_2014,In_1640);
and U197 (N_197,In_1031,In_2473);
or U198 (N_198,In_1944,In_1352);
or U199 (N_199,In_413,In_1901);
nand U200 (N_200,In_1645,In_267);
xnor U201 (N_201,In_531,In_863);
nand U202 (N_202,In_1244,In_181);
nor U203 (N_203,In_913,In_1532);
nor U204 (N_204,In_1766,In_813);
nand U205 (N_205,In_1682,In_1326);
and U206 (N_206,In_1075,In_2445);
xor U207 (N_207,In_480,In_966);
nor U208 (N_208,In_1956,In_969);
nand U209 (N_209,In_1716,In_589);
or U210 (N_210,In_2415,In_817);
or U211 (N_211,In_2130,In_1309);
nor U212 (N_212,In_1750,In_2222);
and U213 (N_213,In_1658,In_441);
or U214 (N_214,In_32,In_880);
nand U215 (N_215,In_371,In_1335);
xor U216 (N_216,In_648,In_1208);
or U217 (N_217,In_2450,In_1178);
or U218 (N_218,In_914,In_1524);
and U219 (N_219,In_777,In_1048);
or U220 (N_220,In_2279,In_1490);
nor U221 (N_221,In_331,In_402);
or U222 (N_222,In_2209,In_873);
nor U223 (N_223,In_1665,In_103);
nand U224 (N_224,In_2429,In_289);
or U225 (N_225,In_1452,In_2200);
and U226 (N_226,In_2087,In_1813);
nand U227 (N_227,In_583,In_709);
and U228 (N_228,In_1405,In_2496);
and U229 (N_229,In_1152,In_761);
xnor U230 (N_230,In_2305,In_1430);
and U231 (N_231,In_832,In_140);
nand U232 (N_232,In_2012,In_189);
or U233 (N_233,In_2214,In_961);
and U234 (N_234,In_694,In_868);
nand U235 (N_235,In_169,In_1450);
or U236 (N_236,In_2228,In_2290);
or U237 (N_237,In_1381,In_1775);
nor U238 (N_238,In_60,In_1144);
nand U239 (N_239,In_1628,In_161);
xor U240 (N_240,In_95,In_1058);
nor U241 (N_241,In_1460,In_1711);
and U242 (N_242,In_1955,In_1489);
nand U243 (N_243,In_2463,In_2426);
or U244 (N_244,In_1362,In_239);
nor U245 (N_245,In_2412,In_340);
nand U246 (N_246,In_801,In_241);
or U247 (N_247,In_1817,In_1207);
nor U248 (N_248,In_2163,In_1126);
nor U249 (N_249,In_1980,In_1032);
or U250 (N_250,In_1869,In_2225);
or U251 (N_251,In_1414,In_2366);
or U252 (N_252,In_354,In_2236);
nand U253 (N_253,In_2005,In_2356);
nand U254 (N_254,In_444,In_1762);
and U255 (N_255,In_1463,In_2096);
and U256 (N_256,In_578,In_1123);
and U257 (N_257,In_387,In_456);
and U258 (N_258,In_1759,In_1359);
nor U259 (N_259,In_1093,In_1571);
and U260 (N_260,In_208,In_251);
or U261 (N_261,In_998,In_27);
nand U262 (N_262,In_959,In_1874);
xnor U263 (N_263,In_609,In_2336);
nor U264 (N_264,In_2424,In_31);
xnor U265 (N_265,In_948,In_909);
and U266 (N_266,In_670,In_2331);
or U267 (N_267,In_2437,In_861);
nand U268 (N_268,In_748,In_2191);
nor U269 (N_269,In_1690,In_361);
or U270 (N_270,In_2410,In_614);
nor U271 (N_271,In_1993,In_1127);
nor U272 (N_272,In_1281,In_2430);
or U273 (N_273,In_854,In_926);
and U274 (N_274,In_1468,In_272);
xor U275 (N_275,In_636,In_1885);
and U276 (N_276,In_1084,In_2091);
nor U277 (N_277,In_952,In_860);
or U278 (N_278,In_353,In_193);
and U279 (N_279,In_1043,In_2238);
xnor U280 (N_280,In_118,In_1180);
and U281 (N_281,In_1124,In_1798);
nor U282 (N_282,In_1168,In_233);
and U283 (N_283,In_475,In_127);
nand U284 (N_284,In_1970,In_1844);
nand U285 (N_285,In_2009,In_1498);
or U286 (N_286,In_696,In_811);
xor U287 (N_287,In_1984,In_1819);
nand U288 (N_288,In_1243,In_2416);
and U289 (N_289,In_1186,In_1958);
xnor U290 (N_290,In_776,In_1580);
or U291 (N_291,In_537,In_1877);
or U292 (N_292,In_642,In_1277);
and U293 (N_293,In_572,In_2007);
nand U294 (N_294,In_2421,In_186);
and U295 (N_295,In_43,In_54);
and U296 (N_296,In_146,In_1007);
or U297 (N_297,In_2184,In_119);
nand U298 (N_298,In_1008,In_894);
xnor U299 (N_299,In_2105,In_1931);
and U300 (N_300,In_2006,In_1654);
or U301 (N_301,In_1245,In_1631);
and U302 (N_302,In_997,In_1171);
nand U303 (N_303,In_1014,In_577);
xnor U304 (N_304,In_1275,In_1936);
nor U305 (N_305,In_1330,In_1822);
or U306 (N_306,In_1044,In_579);
nand U307 (N_307,In_1569,In_1246);
xnor U308 (N_308,In_2109,In_764);
xnor U309 (N_309,In_170,In_1270);
or U310 (N_310,In_1903,In_1856);
xor U311 (N_311,In_2380,In_56);
and U312 (N_312,In_2081,In_827);
xnor U313 (N_313,In_1385,In_123);
or U314 (N_314,In_631,In_91);
xor U315 (N_315,In_1333,In_2187);
and U316 (N_316,In_755,In_1);
nor U317 (N_317,In_314,In_177);
and U318 (N_318,In_1590,In_1354);
xnor U319 (N_319,In_1453,In_2234);
or U320 (N_320,In_388,In_918);
xor U321 (N_321,In_763,In_2446);
xnor U322 (N_322,In_1866,In_2486);
xor U323 (N_323,In_1680,In_1505);
nand U324 (N_324,In_2306,In_1585);
and U325 (N_325,In_766,In_870);
and U326 (N_326,In_1197,In_597);
and U327 (N_327,In_1547,In_2113);
nor U328 (N_328,In_240,In_2059);
or U329 (N_329,In_1369,In_1948);
or U330 (N_330,In_493,In_1810);
nand U331 (N_331,In_2223,In_1389);
xor U332 (N_332,In_1455,In_554);
xor U333 (N_333,In_1691,In_198);
nor U334 (N_334,In_1285,In_1896);
xnor U335 (N_335,In_1131,In_608);
and U336 (N_336,In_33,In_223);
or U337 (N_337,In_157,In_1804);
or U338 (N_338,In_2335,In_134);
xor U339 (N_339,In_2341,In_2253);
xor U340 (N_340,In_1971,In_2131);
and U341 (N_341,In_729,In_749);
xor U342 (N_342,In_908,In_185);
and U343 (N_343,In_963,In_2064);
and U344 (N_344,In_473,In_617);
and U345 (N_345,In_1926,In_780);
xor U346 (N_346,In_1739,In_1458);
xor U347 (N_347,In_1106,In_347);
xnor U348 (N_348,In_1771,In_732);
or U349 (N_349,In_1289,In_1477);
xnor U350 (N_350,In_1891,In_40);
and U351 (N_351,In_2114,In_1787);
or U352 (N_352,In_978,In_1515);
and U353 (N_353,In_1483,In_871);
xor U354 (N_354,In_265,In_2146);
or U355 (N_355,In_1561,In_1807);
or U356 (N_356,In_168,In_1182);
and U357 (N_357,In_2078,In_1424);
or U358 (N_358,In_1924,In_634);
nor U359 (N_359,In_1009,In_2203);
and U360 (N_360,In_1443,In_2362);
or U361 (N_361,In_1906,In_432);
and U362 (N_362,In_2442,In_1796);
and U363 (N_363,In_1525,In_1293);
or U364 (N_364,In_1037,In_350);
nor U365 (N_365,In_1388,In_1833);
xnor U366 (N_366,In_1878,In_243);
and U367 (N_367,In_2045,In_2375);
or U368 (N_368,In_1090,In_980);
nand U369 (N_369,In_615,In_1809);
and U370 (N_370,In_2095,In_2037);
nor U371 (N_371,In_519,In_1411);
or U372 (N_372,In_1274,In_534);
or U373 (N_373,In_1346,In_1578);
nor U374 (N_374,In_2206,In_599);
nor U375 (N_375,In_1670,In_153);
and U376 (N_376,In_2403,In_94);
nand U377 (N_377,In_1753,In_2049);
or U378 (N_378,In_2141,In_856);
nand U379 (N_379,In_920,In_1915);
nor U380 (N_380,In_1556,In_61);
and U381 (N_381,In_665,In_1220);
xor U382 (N_382,In_1935,In_569);
nand U383 (N_383,In_2205,In_404);
xor U384 (N_384,In_1749,In_2170);
xnor U385 (N_385,In_1447,In_896);
or U386 (N_386,In_522,In_1307);
or U387 (N_387,In_2308,In_1908);
nor U388 (N_388,In_1545,In_1203);
nor U389 (N_389,In_1918,In_326);
nand U390 (N_390,In_400,In_1269);
xnor U391 (N_391,In_1045,In_942);
xor U392 (N_392,In_318,In_1164);
xor U393 (N_393,In_1712,In_69);
or U394 (N_394,In_2270,In_1806);
and U395 (N_395,In_677,In_478);
xor U396 (N_396,In_334,In_2409);
xnor U397 (N_397,In_2088,In_159);
and U398 (N_398,In_487,In_2418);
nand U399 (N_399,In_362,In_1384);
and U400 (N_400,In_1999,In_1110);
nand U401 (N_401,In_205,In_1060);
nand U402 (N_402,In_1464,In_2354);
and U403 (N_403,In_1723,In_673);
and U404 (N_404,In_2471,In_2298);
or U405 (N_405,In_1538,In_1738);
or U406 (N_406,In_1859,In_692);
nor U407 (N_407,In_372,In_1195);
and U408 (N_408,In_1621,In_1882);
or U409 (N_409,In_845,In_716);
nor U410 (N_410,In_1607,In_335);
xnor U411 (N_411,In_1374,In_483);
xnor U412 (N_412,In_29,In_2148);
nor U413 (N_413,In_812,In_1165);
nand U414 (N_414,In_1715,In_254);
nor U415 (N_415,In_2385,In_2199);
xnor U416 (N_416,In_286,In_618);
or U417 (N_417,In_675,In_526);
xor U418 (N_418,In_2106,In_1085);
xor U419 (N_419,In_1432,In_1784);
xnor U420 (N_420,In_283,In_1884);
xor U421 (N_421,In_1412,In_1259);
nand U422 (N_422,In_2307,In_971);
xnor U423 (N_423,In_795,In_1261);
xor U424 (N_424,In_1327,In_1426);
nand U425 (N_425,In_671,In_1684);
and U426 (N_426,In_2462,In_1818);
nor U427 (N_427,In_1572,In_34);
and U428 (N_428,In_1905,In_1839);
xnor U429 (N_429,In_1298,In_436);
xor U430 (N_430,In_2372,In_1850);
nor U431 (N_431,In_790,In_560);
xor U432 (N_432,In_2179,In_2123);
xnor U433 (N_433,In_1721,In_2368);
nand U434 (N_434,In_23,In_1666);
nor U435 (N_435,In_2476,In_2323);
xor U436 (N_436,In_2396,In_10);
and U437 (N_437,In_1100,In_953);
nand U438 (N_438,In_28,In_2475);
and U439 (N_439,In_1036,In_533);
and U440 (N_440,In_1170,In_580);
or U441 (N_441,In_310,In_1848);
nand U442 (N_442,In_1191,In_207);
xor U443 (N_443,In_904,In_1247);
xnor U444 (N_444,In_222,In_2484);
and U445 (N_445,In_2399,In_2258);
nand U446 (N_446,In_1500,In_1729);
xnor U447 (N_447,In_1392,In_887);
nand U448 (N_448,In_2264,In_1786);
and U449 (N_449,In_1173,In_151);
or U450 (N_450,In_1674,In_1592);
and U451 (N_451,In_52,In_767);
xor U452 (N_452,In_2400,In_25);
or U453 (N_453,In_419,In_2293);
xor U454 (N_454,In_2406,In_452);
nor U455 (N_455,In_373,In_358);
nand U456 (N_456,In_1317,In_275);
xnor U457 (N_457,In_288,In_2315);
and U458 (N_458,In_1158,In_1154);
or U459 (N_459,In_910,In_1587);
and U460 (N_460,In_885,In_641);
nand U461 (N_461,In_895,In_351);
or U462 (N_462,In_1624,In_1748);
nand U463 (N_463,In_805,In_772);
nand U464 (N_464,In_2077,In_1376);
nand U465 (N_465,In_2312,In_2337);
nand U466 (N_466,In_477,In_2243);
xor U467 (N_467,In_2302,In_1522);
or U468 (N_468,In_602,In_244);
nand U469 (N_469,In_149,In_2075);
nor U470 (N_470,In_506,In_1417);
nand U471 (N_471,In_555,In_1011);
nor U472 (N_472,In_2061,In_527);
nand U473 (N_473,In_1199,In_1648);
nand U474 (N_474,In_558,In_1669);
xnor U475 (N_475,In_2386,In_839);
and U476 (N_476,In_2299,In_266);
nand U477 (N_477,In_703,In_2153);
nand U478 (N_478,In_988,In_1605);
and U479 (N_479,In_1995,In_601);
and U480 (N_480,In_1700,In_1616);
xor U481 (N_481,In_1013,In_955);
and U482 (N_482,In_831,In_2073);
and U483 (N_483,In_1613,In_355);
nor U484 (N_484,In_603,In_1831);
nand U485 (N_485,In_1967,In_81);
xor U486 (N_486,In_287,In_1029);
and U487 (N_487,In_232,In_1484);
nand U488 (N_488,In_1436,In_202);
nand U489 (N_489,In_2070,In_479);
nor U490 (N_490,In_734,In_2292);
and U491 (N_491,In_238,In_320);
nand U492 (N_492,In_462,In_2089);
or U493 (N_493,In_862,In_750);
nor U494 (N_494,In_1399,In_1073);
xnor U495 (N_495,In_225,In_1644);
or U496 (N_496,In_2069,In_268);
nor U497 (N_497,In_449,In_2453);
and U498 (N_498,In_512,In_927);
nor U499 (N_499,In_834,In_65);
nor U500 (N_500,In_1162,In_1686);
nand U501 (N_501,In_2408,In_944);
and U502 (N_502,In_1097,In_1198);
xor U503 (N_503,In_882,In_1105);
nor U504 (N_504,In_1975,In_423);
nor U505 (N_505,In_74,In_2092);
nand U506 (N_506,In_2224,In_128);
or U507 (N_507,In_2013,In_139);
or U508 (N_508,In_1310,In_1034);
nor U509 (N_509,In_1637,In_792);
nand U510 (N_510,In_2028,In_2062);
nand U511 (N_511,In_967,In_1074);
and U512 (N_512,In_1832,In_903);
xnor U513 (N_513,In_765,In_735);
nand U514 (N_514,In_290,In_2371);
xor U515 (N_515,In_536,In_1650);
nor U516 (N_516,In_1952,In_379);
or U517 (N_517,In_2459,In_155);
or U518 (N_518,In_142,In_1740);
xor U519 (N_519,In_1929,In_2230);
nand U520 (N_520,In_212,In_178);
nor U521 (N_521,In_1438,In_2435);
xor U522 (N_522,In_2344,In_154);
and U523 (N_523,In_689,In_1705);
nand U524 (N_524,In_1151,In_680);
and U525 (N_525,In_131,In_42);
and U526 (N_526,In_2150,In_396);
and U527 (N_527,In_1276,In_455);
nand U528 (N_528,In_2288,In_2149);
and U529 (N_529,In_1095,In_276);
or U530 (N_530,In_586,In_1146);
and U531 (N_531,In_99,In_701);
and U532 (N_532,In_1027,In_1925);
and U533 (N_533,In_1420,In_376);
or U534 (N_534,In_1415,In_787);
or U535 (N_535,In_2499,In_1258);
nand U536 (N_536,In_428,In_1745);
nand U537 (N_537,In_1018,In_1402);
and U538 (N_538,In_282,In_327);
and U539 (N_539,In_2126,In_2322);
or U540 (N_540,In_2124,In_1437);
nor U541 (N_541,In_2478,In_1219);
or U542 (N_542,In_1855,In_1982);
or U543 (N_543,In_581,In_2481);
or U544 (N_544,In_1382,In_562);
and U545 (N_545,In_756,In_1224);
nand U546 (N_546,In_2389,In_2458);
nand U547 (N_547,In_1435,In_1720);
or U548 (N_548,In_401,In_190);
and U549 (N_549,In_2068,In_1132);
nand U550 (N_550,In_20,In_63);
and U551 (N_551,In_1004,In_2246);
and U552 (N_552,In_68,In_1603);
nand U553 (N_553,In_2056,In_1187);
nand U554 (N_554,In_1619,In_2355);
or U555 (N_555,In_804,In_2378);
and U556 (N_556,In_446,In_1260);
or U557 (N_557,In_2168,In_1779);
nor U558 (N_558,In_2116,In_616);
nand U559 (N_559,In_1883,In_345);
and U560 (N_560,In_1356,In_1881);
or U561 (N_561,In_649,In_1202);
and U562 (N_562,In_1065,In_1747);
xnor U563 (N_563,In_1709,In_1837);
nor U564 (N_564,In_1442,In_438);
or U565 (N_565,In_624,In_167);
xor U566 (N_566,In_1797,In_564);
nor U567 (N_567,In_79,In_458);
nor U568 (N_568,In_2281,In_809);
nand U569 (N_569,In_1609,In_829);
nand U570 (N_570,In_828,In_1803);
nand U571 (N_571,In_818,In_62);
and U572 (N_572,In_2485,In_228);
or U573 (N_573,In_993,In_1030);
xnor U574 (N_574,In_2151,In_794);
xnor U575 (N_575,In_1104,In_1635);
xor U576 (N_576,In_1727,In_1653);
nor U577 (N_577,In_925,In_1718);
xor U578 (N_578,In_1871,In_201);
or U579 (N_579,In_1911,In_1063);
and U580 (N_580,In_2487,In_1782);
xnor U581 (N_581,In_1968,In_2217);
or U582 (N_582,In_2449,In_1947);
or U583 (N_583,In_802,In_715);
xnor U584 (N_584,In_1175,In_2404);
and U585 (N_585,In_1553,In_1769);
nand U586 (N_586,In_330,In_2142);
and U587 (N_587,In_1618,In_1067);
or U588 (N_588,In_1373,In_2198);
nor U589 (N_589,In_1552,In_570);
nor U590 (N_590,In_977,In_485);
xor U591 (N_591,In_1143,In_1454);
nor U592 (N_592,In_723,In_784);
nor U593 (N_593,In_346,In_269);
or U594 (N_594,In_1047,In_1502);
nor U595 (N_595,In_1940,In_622);
nor U596 (N_596,In_543,In_491);
nor U597 (N_597,In_1689,In_1138);
and U598 (N_598,In_1978,In_1814);
xor U599 (N_599,In_1942,In_791);
xor U600 (N_600,In_650,In_1529);
and U601 (N_601,In_633,In_1713);
xnor U602 (N_602,In_1148,In_1543);
nand U603 (N_603,In_2491,In_2137);
xnor U604 (N_604,In_107,In_1308);
or U605 (N_605,In_18,In_1560);
and U606 (N_606,In_1419,In_313);
or U607 (N_607,In_188,In_1963);
nand U608 (N_608,In_1015,In_661);
or U609 (N_609,In_1919,In_2320);
nor U610 (N_610,In_84,In_964);
nor U611 (N_611,In_2024,In_799);
or U612 (N_612,In_221,In_2176);
nor U613 (N_613,In_1567,In_2433);
nand U614 (N_614,In_415,In_1630);
nand U615 (N_615,In_1272,In_669);
nor U616 (N_616,In_2101,In_2017);
or U617 (N_617,In_707,In_2313);
nand U618 (N_618,In_2218,In_2189);
or U619 (N_619,In_2180,In_2370);
nand U620 (N_620,In_720,In_1643);
nand U621 (N_621,In_638,In_1909);
xor U622 (N_622,In_1794,In_1586);
nand U623 (N_623,In_2495,In_1268);
or U624 (N_624,In_1890,In_561);
and U625 (N_625,N_205,N_283);
and U626 (N_626,In_105,In_611);
and U627 (N_627,N_115,In_344);
nand U628 (N_628,In_2016,In_2351);
or U629 (N_629,In_2464,In_2226);
nand U630 (N_630,N_162,In_1087);
or U631 (N_631,N_475,In_1678);
nand U632 (N_632,In_999,In_1755);
nor U633 (N_633,In_2229,In_711);
xnor U634 (N_634,In_1262,In_1231);
and U635 (N_635,In_1328,N_354);
xnor U636 (N_636,In_1035,In_300);
nand U637 (N_637,N_418,In_15);
or U638 (N_638,In_143,In_662);
nor U639 (N_639,N_190,N_353);
and U640 (N_640,N_368,N_208);
nor U641 (N_641,In_1843,N_174);
and U642 (N_642,In_591,In_2285);
xor U643 (N_643,In_947,N_466);
nor U644 (N_644,In_1101,In_1657);
or U645 (N_645,N_32,In_1378);
and U646 (N_646,N_377,N_603);
and U647 (N_647,In_563,N_94);
or U648 (N_648,In_943,In_1499);
and U649 (N_649,N_599,In_898);
xnor U650 (N_650,In_9,In_643);
or U651 (N_651,In_1150,N_580);
xnor U652 (N_652,In_191,In_2252);
nor U653 (N_653,In_2383,In_2283);
nor U654 (N_654,In_2268,In_628);
and U655 (N_655,In_2135,In_58);
nand U656 (N_656,In_135,N_317);
nor U657 (N_657,In_1236,In_592);
and U658 (N_658,In_1910,N_201);
nand U659 (N_659,N_457,N_610);
or U660 (N_660,N_181,N_93);
nand U661 (N_661,In_2492,N_72);
xnor U662 (N_662,In_76,In_1223);
xor U663 (N_663,N_114,In_147);
nor U664 (N_664,In_1823,In_2393);
or U665 (N_665,In_2291,N_171);
and U666 (N_666,In_405,N_122);
and U667 (N_667,In_496,N_524);
xor U668 (N_668,N_41,N_503);
nand U669 (N_669,N_566,In_751);
or U670 (N_670,N_58,N_428);
nand U671 (N_671,In_1615,In_2103);
and U672 (N_672,In_114,In_2296);
nor U673 (N_673,In_798,In_1589);
nand U674 (N_674,In_2402,N_95);
and U675 (N_675,In_1530,In_2019);
and U676 (N_676,In_793,N_460);
nand U677 (N_677,In_1681,N_28);
or U678 (N_678,N_5,In_250);
and U679 (N_679,In_2490,N_382);
nand U680 (N_680,In_1706,N_425);
and U681 (N_681,N_62,In_710);
and U682 (N_682,N_336,In_2183);
nand U683 (N_683,N_472,In_1465);
or U684 (N_684,In_214,In_1677);
nand U685 (N_685,In_1544,N_40);
and U686 (N_686,In_1344,In_2147);
and U687 (N_687,In_1339,N_213);
and U688 (N_688,In_468,In_89);
xor U689 (N_689,In_1826,N_442);
or U690 (N_690,In_950,In_949);
nand U691 (N_691,In_2035,N_441);
or U692 (N_692,In_585,In_2247);
and U693 (N_693,In_2441,N_31);
and U694 (N_694,N_493,N_361);
xnor U695 (N_695,In_137,N_454);
nor U696 (N_696,In_4,N_611);
and U697 (N_697,In_45,In_1256);
or U698 (N_698,N_204,In_1042);
or U699 (N_699,In_745,In_463);
xor U700 (N_700,In_1760,In_1020);
and U701 (N_701,In_1266,In_545);
nor U702 (N_702,In_890,In_1319);
nand U703 (N_703,In_1579,In_1122);
or U704 (N_704,N_84,N_197);
nor U705 (N_705,N_411,In_846);
and U706 (N_706,N_65,In_1306);
xnor U707 (N_707,In_768,In_1086);
or U708 (N_708,In_1213,In_2259);
nor U709 (N_709,N_343,N_146);
xor U710 (N_710,N_104,N_46);
xor U711 (N_711,N_274,In_879);
and U712 (N_712,In_1325,In_2055);
nor U713 (N_713,N_562,In_1360);
nand U714 (N_714,N_4,In_2251);
nand U715 (N_715,N_557,In_1765);
and U716 (N_716,In_1699,In_2325);
or U717 (N_717,N_79,N_167);
nand U718 (N_718,N_291,N_431);
nand U719 (N_719,In_1107,In_810);
and U720 (N_720,N_360,In_718);
nor U721 (N_721,In_218,In_433);
and U722 (N_722,N_262,In_14);
and U723 (N_723,In_984,N_138);
and U724 (N_724,In_229,N_150);
nand U725 (N_725,In_1583,In_2232);
and U726 (N_726,N_199,N_71);
nor U727 (N_727,In_2041,In_1862);
and U728 (N_728,In_2210,In_426);
nor U729 (N_729,N_281,N_469);
nand U730 (N_730,In_1938,In_235);
and U731 (N_731,In_1239,In_954);
xor U732 (N_732,N_455,In_263);
xnor U733 (N_733,N_364,In_565);
nor U734 (N_734,In_1964,In_1329);
and U735 (N_735,In_2423,In_1238);
xor U736 (N_736,N_82,N_59);
xor U737 (N_737,In_1998,N_438);
nand U738 (N_738,In_2392,In_738);
nor U739 (N_739,In_1200,N_192);
nor U740 (N_740,N_594,In_2367);
xor U741 (N_741,In_1296,In_247);
nor U742 (N_742,N_482,In_1320);
xor U743 (N_743,In_2384,In_1401);
nor U744 (N_744,In_1612,In_1830);
and U745 (N_745,In_1781,In_2162);
nand U746 (N_746,In_2140,N_595);
xnor U747 (N_747,In_940,In_215);
or U748 (N_748,In_951,In_1922);
nand U749 (N_749,In_881,In_1698);
nand U750 (N_750,In_1230,In_2479);
or U751 (N_751,In_2090,In_2039);
or U752 (N_752,In_1257,N_381);
xor U753 (N_753,N_49,In_1471);
nor U754 (N_754,In_2286,N_390);
nor U755 (N_755,In_1304,In_1730);
or U756 (N_756,In_2265,In_1912);
or U757 (N_757,In_1156,N_11);
or U758 (N_758,In_724,N_556);
or U759 (N_759,In_2339,In_666);
or U760 (N_760,In_835,In_1516);
or U761 (N_761,In_1321,N_25);
nand U762 (N_762,In_220,N_301);
xor U763 (N_763,N_144,In_204);
and U764 (N_764,In_606,N_80);
xnor U765 (N_765,In_406,In_1076);
or U766 (N_766,In_1704,In_1361);
xor U767 (N_767,N_156,In_2020);
nor U768 (N_768,In_1194,In_1641);
nand U769 (N_769,In_1900,In_1961);
or U770 (N_770,In_385,N_277);
nand U771 (N_771,In_886,In_366);
xor U772 (N_772,In_2452,N_177);
and U773 (N_773,N_429,In_1174);
xnor U774 (N_774,N_543,In_605);
nand U775 (N_775,N_452,N_1);
nor U776 (N_776,N_315,N_226);
xor U777 (N_777,In_1145,In_1751);
nor U778 (N_778,In_231,In_548);
nand U779 (N_779,N_507,N_123);
and U780 (N_780,N_598,N_124);
or U781 (N_781,In_595,N_279);
and U782 (N_782,In_1921,N_0);
nand U783 (N_783,In_97,N_483);
or U784 (N_784,In_246,In_109);
nand U785 (N_785,N_568,In_739);
xor U786 (N_786,In_1240,In_1774);
nor U787 (N_787,N_165,In_663);
nor U788 (N_788,N_394,In_2289);
or U789 (N_789,N_103,N_545);
nor U790 (N_790,In_1593,In_2361);
and U791 (N_791,N_619,In_1867);
nor U792 (N_792,In_1780,N_558);
nor U793 (N_793,In_1334,In_2190);
nor U794 (N_794,In_98,In_1080);
xor U795 (N_795,N_539,N_335);
or U796 (N_796,In_1582,In_1279);
nand U797 (N_797,N_397,N_613);
nor U798 (N_798,In_2197,N_30);
or U799 (N_799,N_501,N_334);
and U800 (N_800,N_17,In_418);
and U801 (N_801,In_1722,In_1486);
nor U802 (N_802,In_1851,N_67);
and U803 (N_803,N_447,In_2036);
nor U804 (N_804,In_1167,In_1064);
and U805 (N_805,N_518,N_561);
nand U806 (N_806,In_2161,In_2414);
or U807 (N_807,In_1470,N_129);
nand U808 (N_808,N_366,N_609);
xor U809 (N_809,In_2233,N_304);
and U810 (N_810,In_1254,In_431);
nand U811 (N_811,N_66,N_575);
or U812 (N_812,In_1390,N_222);
and U813 (N_813,In_1314,In_568);
or U814 (N_814,N_232,N_554);
xnor U815 (N_815,N_107,N_513);
or U816 (N_816,N_355,In_1089);
and U817 (N_817,In_664,In_2004);
nand U818 (N_818,N_464,In_566);
or U819 (N_819,In_390,N_384);
nor U820 (N_820,In_1870,In_206);
xnor U821 (N_821,In_1735,In_1479);
xor U822 (N_822,N_374,In_2417);
nor U823 (N_823,N_591,In_2001);
and U824 (N_824,In_427,N_285);
or U825 (N_825,In_1685,N_231);
xnor U826 (N_826,In_2177,N_272);
nor U827 (N_827,In_1659,In_826);
xnor U828 (N_828,N_597,In_630);
xnor U829 (N_829,In_175,N_166);
or U830 (N_830,In_824,In_712);
xor U831 (N_831,In_2498,In_416);
xnor U832 (N_832,N_365,N_321);
and U833 (N_833,N_579,In_517);
and U834 (N_834,N_169,N_37);
nand U835 (N_835,N_461,N_616);
nor U836 (N_836,N_376,In_271);
nand U837 (N_837,N_424,N_39);
or U838 (N_838,In_488,In_1375);
nor U839 (N_839,In_117,N_111);
nor U840 (N_840,In_1221,In_1573);
nor U841 (N_841,In_1577,In_781);
or U842 (N_842,In_5,In_1444);
and U843 (N_843,N_326,In_514);
nor U844 (N_844,In_2304,In_2309);
nand U845 (N_845,N_253,In_1434);
xor U846 (N_846,In_1611,In_1886);
nand U847 (N_847,N_38,In_111);
and U848 (N_848,N_12,In_359);
nor U849 (N_849,In_259,N_21);
and U850 (N_850,In_307,N_221);
nor U851 (N_851,N_587,In_2054);
nor U852 (N_852,N_540,In_679);
or U853 (N_853,In_921,N_548);
xor U854 (N_854,N_305,In_332);
nand U855 (N_855,N_478,In_476);
or U856 (N_856,In_1079,In_1351);
nor U857 (N_857,In_771,In_683);
and U858 (N_858,N_409,In_1576);
xor U859 (N_859,N_242,In_7);
or U860 (N_860,In_389,In_71);
nand U861 (N_861,N_266,In_1888);
and U862 (N_862,N_560,In_2027);
nor U863 (N_863,N_333,In_1741);
nor U864 (N_864,In_2044,In_398);
xor U865 (N_865,N_399,N_371);
or U866 (N_866,In_956,In_2407);
or U867 (N_867,N_276,N_207);
nor U868 (N_868,In_1466,In_295);
nand U869 (N_869,In_825,In_1676);
nand U870 (N_870,In_133,In_1783);
or U871 (N_871,In_6,N_314);
or U872 (N_872,N_142,In_121);
and U873 (N_873,N_102,N_584);
and U874 (N_874,In_2271,In_46);
nor U875 (N_875,In_557,In_2212);
and U876 (N_876,In_2138,N_259);
nand U877 (N_877,In_21,In_1355);
nand U878 (N_878,N_459,N_18);
or U879 (N_879,N_170,In_2310);
xnor U880 (N_880,In_1449,N_10);
xnor U881 (N_881,In_1930,In_44);
and U882 (N_882,In_635,N_517);
nor U883 (N_883,N_81,N_588);
nand U884 (N_884,N_55,In_1188);
and U885 (N_885,In_237,In_2493);
nand U886 (N_886,N_617,N_362);
nand U887 (N_887,N_306,In_1973);
nor U888 (N_888,N_396,In_640);
nand U889 (N_889,In_1427,N_43);
nand U890 (N_890,In_2350,In_1997);
or U891 (N_891,In_1983,N_63);
nor U892 (N_892,In_73,In_2365);
nor U893 (N_893,In_883,In_1255);
or U894 (N_894,N_295,N_578);
nand U895 (N_895,In_1383,In_900);
and U896 (N_896,In_922,In_1550);
nor U897 (N_897,In_2357,In_875);
and U898 (N_898,In_1094,N_357);
xor U899 (N_899,In_343,N_458);
or U900 (N_900,In_106,In_1863);
nor U901 (N_901,In_2099,In_850);
and U902 (N_902,In_1302,In_2317);
and U903 (N_903,In_291,In_524);
or U904 (N_904,In_457,N_329);
nand U905 (N_905,In_484,N_99);
and U906 (N_906,N_48,N_297);
nand U907 (N_907,N_87,In_646);
xor U908 (N_908,In_888,In_2447);
or U909 (N_909,In_1555,In_1109);
xor U910 (N_910,In_2079,N_209);
nor U911 (N_911,In_708,In_1136);
or U912 (N_912,N_338,In_1128);
nor U913 (N_913,In_645,In_507);
and U914 (N_914,In_1380,In_1481);
or U915 (N_915,In_1507,In_2112);
and U916 (N_916,N_504,In_741);
or U917 (N_917,In_2353,In_1693);
and U918 (N_918,N_56,N_350);
and U919 (N_919,N_569,N_367);
xor U920 (N_920,N_271,N_14);
or U921 (N_921,In_2457,In_1410);
or U922 (N_922,In_2166,In_1895);
or U923 (N_923,N_433,In_2023);
xnor U924 (N_924,N_252,N_515);
nand U925 (N_925,N_551,N_16);
or U926 (N_926,In_249,N_511);
nand U927 (N_927,In_752,N_330);
nor U928 (N_928,In_747,In_183);
xor U929 (N_929,N_522,In_136);
xnor U930 (N_930,In_1370,In_2220);
and U931 (N_931,In_2181,N_110);
xnor U932 (N_932,In_596,N_92);
and U933 (N_933,In_471,N_117);
nand U934 (N_934,N_509,In_1606);
and U935 (N_935,N_20,In_619);
or U936 (N_936,In_2158,N_140);
and U937 (N_937,In_1407,In_690);
nand U938 (N_938,In_869,In_1318);
xor U939 (N_939,In_1461,N_563);
nor U940 (N_940,In_625,N_553);
and U941 (N_941,N_173,In_2379);
xor U942 (N_942,In_1026,N_555);
and U943 (N_943,In_392,In_2348);
and U944 (N_944,In_1467,In_80);
or U945 (N_945,In_1459,N_303);
and U946 (N_946,N_331,In_1596);
nor U947 (N_947,In_442,In_2256);
xnor U948 (N_948,In_1005,In_686);
or U949 (N_949,In_878,In_2276);
and U950 (N_950,N_574,In_2072);
and U951 (N_951,In_261,N_249);
nor U952 (N_952,In_1253,In_571);
nand U953 (N_953,In_447,In_2010);
or U954 (N_954,N_161,In_995);
nor U955 (N_955,In_713,In_1664);
or U956 (N_956,In_851,In_637);
nand U957 (N_957,In_1756,In_481);
and U958 (N_958,In_200,N_289);
nand U959 (N_959,In_1409,N_141);
or U960 (N_960,In_2382,In_1431);
nand U961 (N_961,N_370,In_1875);
xor U962 (N_962,In_104,In_1242);
and U963 (N_963,In_1315,In_194);
or U964 (N_964,N_131,N_526);
xnor U965 (N_965,In_2332,N_119);
nand U966 (N_966,In_1416,N_340);
xor U967 (N_967,In_1340,N_529);
and U968 (N_968,In_66,In_2002);
nor U969 (N_969,In_1297,In_651);
nand U970 (N_970,In_1189,N_78);
and U971 (N_971,In_108,N_258);
xor U972 (N_972,N_541,In_164);
xnor U973 (N_973,In_1737,In_2395);
or U974 (N_974,In_1012,In_83);
xor U975 (N_975,In_1282,In_1292);
and U976 (N_976,In_217,In_1140);
xor U977 (N_977,N_327,In_306);
nor U978 (N_978,In_549,N_550);
xnor U979 (N_979,N_133,In_1696);
and U980 (N_980,N_521,In_1379);
nor U981 (N_981,N_440,N_83);
nand U982 (N_982,N_163,In_864);
nor U983 (N_983,In_1366,In_2328);
and U984 (N_984,In_567,In_1116);
and U985 (N_985,N_348,In_2171);
and U986 (N_986,N_359,In_1986);
nor U987 (N_987,In_1827,In_1157);
nand U988 (N_988,N_311,N_246);
nand U989 (N_989,In_270,N_332);
nand U990 (N_990,N_488,In_672);
and U991 (N_991,In_1038,In_731);
xor U992 (N_992,In_1732,In_2129);
or U993 (N_993,In_1941,N_615);
nor U994 (N_994,In_704,In_284);
xor U995 (N_995,In_1617,N_270);
xor U996 (N_996,In_1724,In_2497);
and U997 (N_997,N_101,In_1568);
and U998 (N_998,In_1228,In_1887);
and U999 (N_999,N_175,N_497);
nand U1000 (N_1000,In_654,In_211);
nand U1001 (N_1001,In_688,N_113);
nor U1002 (N_1002,In_440,N_51);
nor U1003 (N_1003,In_1675,In_981);
xor U1004 (N_1004,In_1323,N_230);
and U1005 (N_1005,In_1990,In_1066);
nor U1006 (N_1006,In_1176,In_789);
or U1007 (N_1007,In_257,N_347);
or U1008 (N_1008,In_1668,In_472);
nor U1009 (N_1009,In_382,In_1462);
xor U1010 (N_1010,N_136,N_76);
and U1011 (N_1011,N_415,N_600);
xor U1012 (N_1012,In_2201,N_407);
or U1013 (N_1013,In_439,In_1801);
nor U1014 (N_1014,N_320,In_1311);
nor U1015 (N_1015,In_498,In_1003);
and U1016 (N_1016,N_22,N_116);
nand U1017 (N_1017,N_189,In_2398);
nor U1018 (N_1018,In_1010,In_451);
nor U1019 (N_1019,In_1757,N_484);
nand U1020 (N_1020,In_2063,In_242);
nand U1021 (N_1021,N_534,N_538);
nor U1022 (N_1022,N_261,In_778);
nand U1023 (N_1023,In_1584,In_2207);
or U1024 (N_1024,N_430,In_1651);
nand U1025 (N_1025,In_1853,In_523);
nand U1026 (N_1026,N_153,In_1283);
or U1027 (N_1027,N_468,In_916);
and U1028 (N_1028,In_2278,In_450);
nand U1029 (N_1029,In_700,In_30);
xnor U1030 (N_1030,N_180,In_1192);
or U1031 (N_1031,N_307,In_691);
xor U1032 (N_1032,In_2330,In_409);
xnor U1033 (N_1033,In_1371,N_393);
nor U1034 (N_1034,In_1849,N_477);
nor U1035 (N_1035,In_1433,In_889);
xor U1036 (N_1036,In_1142,In_2052);
nand U1037 (N_1037,In_1209,In_958);
or U1038 (N_1038,In_2083,In_2467);
nand U1039 (N_1039,In_1493,N_589);
xor U1040 (N_1040,In_693,N_128);
or U1041 (N_1041,N_145,In_656);
xnor U1042 (N_1042,In_397,In_1932);
nand U1043 (N_1043,N_528,N_451);
nand U1044 (N_1044,In_2144,In_1714);
nor U1045 (N_1045,N_624,In_360);
nand U1046 (N_1046,In_305,N_446);
nor U1047 (N_1047,In_779,N_256);
and U1048 (N_1048,N_322,N_255);
xor U1049 (N_1049,N_436,In_2434);
nor U1050 (N_1050,In_2195,N_198);
and U1051 (N_1051,In_1353,In_1510);
nor U1052 (N_1052,N_248,In_647);
and U1053 (N_1053,In_2377,In_934);
nand U1054 (N_1054,N_251,In_698);
nor U1055 (N_1055,In_2451,In_1241);
nand U1056 (N_1056,N_176,In_1496);
or U1057 (N_1057,In_836,N_533);
nand U1058 (N_1058,In_2127,In_928);
and U1059 (N_1059,N_215,In_363);
nor U1060 (N_1060,N_24,N_217);
and U1061 (N_1061,In_785,N_622);
or U1062 (N_1062,In_1250,N_224);
xnor U1063 (N_1063,N_422,In_901);
nand U1064 (N_1064,In_2107,In_930);
nor U1065 (N_1065,In_2050,In_722);
nor U1066 (N_1066,In_2134,In_1497);
xor U1067 (N_1067,In_1372,In_1341);
nor U1068 (N_1068,N_109,In_1959);
xor U1069 (N_1069,In_1078,In_1021);
xor U1070 (N_1070,In_1052,In_759);
or U1071 (N_1071,N_218,In_1717);
or U1072 (N_1072,In_559,N_178);
nor U1073 (N_1073,N_316,N_449);
and U1074 (N_1074,In_1858,N_465);
xnor U1075 (N_1075,N_349,In_281);
nor U1076 (N_1076,N_586,In_2266);
nand U1077 (N_1077,In_2419,In_1083);
and U1078 (N_1078,In_2164,In_2074);
nor U1079 (N_1079,In_2319,N_308);
nor U1080 (N_1080,N_200,N_86);
nor U1081 (N_1081,In_219,In_1033);
nor U1082 (N_1082,N_35,In_1950);
and U1083 (N_1083,N_342,In_1777);
or U1084 (N_1084,N_375,N_378);
nand U1085 (N_1085,In_972,In_695);
nor U1086 (N_1086,N_490,N_416);
nand U1087 (N_1087,In_1072,In_976);
xor U1088 (N_1088,N_188,In_607);
nand U1089 (N_1089,In_1876,In_1917);
nand U1090 (N_1090,In_2038,In_1040);
and U1091 (N_1091,In_816,In_2267);
nand U1092 (N_1092,In_224,N_42);
and U1093 (N_1093,In_460,In_1904);
xor U1094 (N_1094,N_453,In_1291);
and U1095 (N_1095,In_1130,N_505);
or U1096 (N_1096,In_2011,In_1016);
nand U1097 (N_1097,In_1701,N_294);
and U1098 (N_1098,N_489,In_129);
or U1099 (N_1099,In_1595,In_465);
and U1100 (N_1100,In_2128,In_520);
xor U1101 (N_1101,In_2117,In_590);
nand U1102 (N_1102,In_2216,In_1742);
and U1103 (N_1103,In_357,In_1120);
and U1104 (N_1104,N_318,In_962);
and U1105 (N_1105,In_1322,In_932);
xor U1106 (N_1106,In_1091,N_388);
and U1107 (N_1107,In_859,In_2260);
xnor U1108 (N_1108,N_75,In_2154);
nor U1109 (N_1109,N_168,N_582);
xnor U1110 (N_1110,N_450,In_547);
and U1111 (N_1111,In_1534,In_2394);
nor U1112 (N_1112,N_275,N_263);
nor U1113 (N_1113,In_820,In_1056);
nand U1114 (N_1114,N_293,In_987);
nand U1115 (N_1115,In_2043,In_1523);
xor U1116 (N_1116,In_1894,N_552);
nand U1117 (N_1117,In_1137,N_34);
nor U1118 (N_1118,In_1646,N_137);
nand U1119 (N_1119,In_116,In_1632);
nand U1120 (N_1120,N_403,In_893);
xnor U1121 (N_1121,In_1129,N_618);
xnor U1122 (N_1122,In_2263,In_1949);
xnor U1123 (N_1123,In_505,In_1491);
nand U1124 (N_1124,N_212,In_2192);
or U1125 (N_1125,N_426,In_502);
xor U1126 (N_1126,In_726,N_462);
nand U1127 (N_1127,N_612,In_1726);
nor U1128 (N_1128,In_1271,In_2327);
and U1129 (N_1129,N_583,N_604);
xnor U1130 (N_1130,N_50,N_269);
or U1131 (N_1131,In_294,N_96);
nor U1132 (N_1132,N_471,In_172);
nand U1133 (N_1133,In_2425,N_427);
xnor U1134 (N_1134,N_54,In_41);
nor U1135 (N_1135,N_596,In_1597);
nand U1136 (N_1136,N_273,In_1599);
nand U1137 (N_1137,In_1528,In_2174);
nor U1138 (N_1138,In_774,N_476);
nand U1139 (N_1139,In_1446,In_1495);
and U1140 (N_1140,In_917,In_823);
or U1141 (N_1141,N_351,N_395);
nand U1142 (N_1142,In_1331,N_398);
nor U1143 (N_1143,In_762,In_1204);
or U1144 (N_1144,In_2053,In_1626);
or U1145 (N_1145,In_302,In_1099);
nand U1146 (N_1146,In_2443,In_1057);
xor U1147 (N_1147,N_214,In_992);
or U1148 (N_1148,In_1736,N_147);
and U1149 (N_1149,In_1508,In_13);
nor U1150 (N_1150,In_19,N_267);
nand U1151 (N_1151,In_717,In_1694);
xor U1152 (N_1152,N_499,In_2244);
or U1153 (N_1153,In_2294,In_2086);
nor U1154 (N_1154,In_489,In_1811);
nor U1155 (N_1155,In_2269,In_115);
nor U1156 (N_1156,In_525,In_1349);
nand U1157 (N_1157,N_445,N_479);
or U1158 (N_1158,In_1487,In_518);
nor U1159 (N_1159,In_1965,N_444);
xor U1160 (N_1160,In_1294,In_706);
and U1161 (N_1161,N_184,N_29);
or U1162 (N_1162,In_1824,N_203);
nand U1163 (N_1163,In_101,N_268);
xnor U1164 (N_1164,N_565,In_352);
nor U1165 (N_1165,In_613,In_39);
nor U1166 (N_1166,In_1868,In_2277);
or U1167 (N_1167,In_1792,In_833);
and U1168 (N_1168,In_2282,In_538);
or U1169 (N_1169,In_1647,In_1472);
and U1170 (N_1170,In_412,In_1184);
xnor U1171 (N_1171,In_1396,In_800);
nand U1172 (N_1172,N_9,In_173);
xor U1173 (N_1173,N_481,N_206);
nand U1174 (N_1174,In_510,N_149);
xor U1175 (N_1175,In_702,In_298);
and U1176 (N_1176,In_2427,In_420);
nand U1177 (N_1177,In_1475,In_1492);
or U1178 (N_1178,In_658,In_912);
xor U1179 (N_1179,In_466,In_2436);
and U1180 (N_1180,N_53,In_2242);
xor U1181 (N_1181,In_1703,In_1996);
and U1182 (N_1182,In_1873,In_2480);
xnor U1183 (N_1183,N_97,In_705);
or U1184 (N_1184,In_380,In_1249);
xor U1185 (N_1185,In_1945,In_604);
nor U1186 (N_1186,In_171,In_990);
and U1187 (N_1187,In_1061,N_410);
nor U1188 (N_1188,In_655,In_573);
nand U1189 (N_1189,N_401,N_216);
xnor U1190 (N_1190,In_486,N_510);
nand U1191 (N_1191,In_855,In_1363);
and U1192 (N_1192,In_319,In_384);
nor U1193 (N_1193,In_1287,In_582);
nor U1194 (N_1194,In_2468,N_19);
xor U1195 (N_1195,In_919,In_1139);
nand U1196 (N_1196,N_121,In_1365);
nor U1197 (N_1197,N_309,N_514);
nand U1198 (N_1198,In_356,In_1548);
or U1199 (N_1199,In_2098,In_797);
and U1200 (N_1200,In_492,In_1667);
nor U1201 (N_1201,In_1793,N_155);
nor U1202 (N_1202,In_197,N_531);
nand U1203 (N_1203,N_234,In_1788);
nand U1204 (N_1204,In_2295,In_1299);
nand U1205 (N_1205,In_721,N_157);
xor U1206 (N_1206,N_434,In_594);
xnor U1207 (N_1207,In_2042,N_152);
and U1208 (N_1208,N_379,In_1166);
xor U1209 (N_1209,In_1695,N_404);
and U1210 (N_1210,In_158,In_632);
or U1211 (N_1211,In_2121,N_494);
and U1212 (N_1212,N_33,In_1933);
nor U1213 (N_1213,In_1169,In_1357);
xnor U1214 (N_1214,N_135,In_341);
and U1215 (N_1215,In_2193,In_1473);
nor U1216 (N_1216,N_187,In_82);
and U1217 (N_1217,N_239,In_2413);
nor U1218 (N_1218,N_225,In_407);
nand U1219 (N_1219,N_470,In_408);
xnor U1220 (N_1220,In_844,N_100);
nor U1221 (N_1221,In_374,In_1050);
nand U1222 (N_1222,In_1469,N_202);
nand U1223 (N_1223,N_417,N_546);
nor U1224 (N_1224,N_564,In_838);
and U1225 (N_1225,In_2494,In_1135);
nand U1226 (N_1226,In_1776,N_130);
nand U1227 (N_1227,In_1828,In_725);
xnor U1228 (N_1228,In_1521,In_2272);
nand U1229 (N_1229,In_968,N_535);
and U1230 (N_1230,In_769,In_1554);
nor U1231 (N_1231,N_238,N_341);
xor U1232 (N_1232,In_299,In_227);
or U1233 (N_1233,N_284,In_667);
and U1234 (N_1234,N_508,N_77);
xnor U1235 (N_1235,In_1233,In_1539);
and U1236 (N_1236,N_573,N_486);
xor U1237 (N_1237,In_1117,In_1802);
and U1238 (N_1238,In_1181,N_312);
and U1239 (N_1239,In_974,In_1702);
nor U1240 (N_1240,N_391,In_929);
or U1241 (N_1241,In_1092,N_61);
or U1242 (N_1242,N_15,In_1134);
and U1243 (N_1243,N_323,In_1852);
and U1244 (N_1244,N_120,N_369);
or U1245 (N_1245,In_2025,In_1183);
and U1246 (N_1246,In_1559,In_386);
xor U1247 (N_1247,In_2376,In_1800);
or U1248 (N_1248,In_1441,In_1088);
or U1249 (N_1249,In_544,In_1480);
nand U1250 (N_1250,In_1966,N_1025);
and U1251 (N_1251,In_85,N_1136);
and U1252 (N_1252,In_1531,N_940);
nor U1253 (N_1253,N_975,In_1193);
nor U1254 (N_1254,N_795,In_629);
nor U1255 (N_1255,In_48,N_1239);
nor U1256 (N_1256,In_627,N_862);
and U1257 (N_1257,In_2102,N_815);
nand U1258 (N_1258,N_210,N_1068);
xnor U1259 (N_1259,In_2314,N_664);
and U1260 (N_1260,N_44,N_1199);
nand U1261 (N_1261,N_643,N_1005);
or U1262 (N_1262,N_480,N_1009);
nand U1263 (N_1263,N_770,In_1368);
and U1264 (N_1264,In_1977,N_666);
nand U1265 (N_1265,In_1062,N_1177);
nor U1266 (N_1266,In_324,N_194);
nor U1267 (N_1267,N_1028,In_1638);
xor U1268 (N_1268,In_1842,N_894);
nand U1269 (N_1269,In_383,N_768);
nor U1270 (N_1270,N_1030,N_960);
nand U1271 (N_1271,N_682,N_910);
nand U1272 (N_1272,In_2460,N_991);
nor U1273 (N_1273,In_542,In_448);
nand U1274 (N_1274,N_776,N_738);
nand U1275 (N_1275,N_1017,In_1000);
nor U1276 (N_1276,N_694,N_873);
xor U1277 (N_1277,In_141,In_684);
xnor U1278 (N_1278,In_1511,N_858);
xnor U1279 (N_1279,In_1324,N_423);
or U1280 (N_1280,In_2145,N_125);
xor U1281 (N_1281,N_319,In_1118);
xor U1282 (N_1282,In_470,N_1127);
xor U1283 (N_1283,N_1007,In_1934);
nor U1284 (N_1284,In_126,N_665);
nor U1285 (N_1285,N_774,N_85);
xor U1286 (N_1286,N_983,N_930);
and U1287 (N_1287,In_1216,In_1602);
xnor U1288 (N_1288,N_673,N_608);
xnor U1289 (N_1289,N_1131,In_125);
nor U1290 (N_1290,N_1162,In_1394);
nor U1291 (N_1291,N_134,N_658);
nand U1292 (N_1292,N_985,N_1070);
or U1293 (N_1293,N_993,N_799);
nand U1294 (N_1294,N_1145,N_1058);
nor U1295 (N_1295,N_925,N_976);
nand U1296 (N_1296,N_1212,In_678);
nor U1297 (N_1297,N_663,In_2159);
nand U1298 (N_1298,In_1177,In_1692);
xor U1299 (N_1299,N_106,In_1954);
xor U1300 (N_1300,N_869,N_899);
nand U1301 (N_1301,N_547,In_2235);
or U1302 (N_1302,N_832,N_1148);
nor U1303 (N_1303,N_1107,N_825);
nor U1304 (N_1304,N_819,N_620);
or U1305 (N_1305,In_273,In_659);
nand U1306 (N_1306,N_626,N_1167);
xor U1307 (N_1307,N_1076,N_952);
and U1308 (N_1308,In_1300,In_2359);
or U1309 (N_1309,In_1017,N_753);
nor U1310 (N_1310,In_2033,In_2032);
or U1311 (N_1311,N_747,In_1474);
and U1312 (N_1312,In_1077,N_929);
nor U1313 (N_1313,N_953,In_1953);
nand U1314 (N_1314,In_1111,In_309);
or U1315 (N_1315,In_2257,N_1186);
xor U1316 (N_1316,In_145,N_857);
nor U1317 (N_1317,N_808,N_196);
nor U1318 (N_1318,In_1625,In_474);
or U1319 (N_1319,In_1812,In_1519);
xnor U1320 (N_1320,N_1066,N_741);
xor U1321 (N_1321,N_1151,N_567);
nor U1322 (N_1322,In_1758,N_1140);
or U1323 (N_1323,N_678,In_2474);
or U1324 (N_1324,In_1211,N_581);
nor U1325 (N_1325,In_92,In_1406);
nor U1326 (N_1326,N_127,N_1115);
nand U1327 (N_1327,N_851,In_315);
or U1328 (N_1328,N_860,N_1072);
xnor U1329 (N_1329,N_831,N_720);
nor U1330 (N_1330,N_651,N_845);
or U1331 (N_1331,N_628,N_967);
nor U1332 (N_1332,N_1051,N_1243);
nand U1333 (N_1333,N_804,N_1108);
nor U1334 (N_1334,N_1088,In_1119);
nand U1335 (N_1335,In_1400,In_588);
nand U1336 (N_1336,N_244,In_2211);
and U1337 (N_1337,N_1218,N_1132);
or U1338 (N_1338,N_264,N_840);
xnor U1339 (N_1339,N_220,In_529);
or U1340 (N_1340,N_160,In_179);
nand U1341 (N_1341,N_1056,N_1112);
xor U1342 (N_1342,N_344,N_674);
nand U1343 (N_1343,In_1845,In_849);
xor U1344 (N_1344,N_52,In_57);
nor U1345 (N_1345,N_1096,In_2334);
xnor U1346 (N_1346,N_653,N_926);
nor U1347 (N_1347,In_2030,N_310);
and U1348 (N_1348,In_100,N_1159);
nor U1349 (N_1349,N_773,N_1079);
or U1350 (N_1350,In_535,N_638);
or U1351 (N_1351,N_1143,N_820);
nor U1352 (N_1352,N_601,N_1024);
nand U1353 (N_1353,In_1059,N_704);
xnor U1354 (N_1354,N_532,N_1094);
or U1355 (N_1355,In_1513,N_542);
nand U1356 (N_1356,In_786,N_1073);
or U1357 (N_1357,N_70,In_322);
xnor U1358 (N_1358,In_1141,N_1090);
nand U1359 (N_1359,N_633,In_1336);
nor U1360 (N_1360,In_2160,N_516);
xor U1361 (N_1361,N_1099,In_1391);
or U1362 (N_1362,N_1205,N_386);
and U1363 (N_1363,N_1008,N_769);
xor U1364 (N_1364,N_1166,N_1211);
nand U1365 (N_1365,In_1201,In_508);
xnor U1366 (N_1366,In_2364,N_383);
and U1367 (N_1367,In_1448,N_108);
xnor U1368 (N_1368,In_1763,In_2401);
nand U1369 (N_1369,N_324,In_1879);
and U1370 (N_1370,N_413,N_1045);
and U1371 (N_1371,N_287,In_516);
and U1372 (N_1372,In_1205,N_726);
nor U1373 (N_1373,In_2390,N_408);
and U1374 (N_1374,In_1864,N_576);
nand U1375 (N_1375,N_235,N_435);
xnor U1376 (N_1376,N_570,N_211);
or U1377 (N_1377,N_1237,In_2248);
and U1378 (N_1378,N_105,In_511);
or U1379 (N_1379,N_265,N_699);
and U1380 (N_1380,In_453,N_996);
xor U1381 (N_1381,N_406,N_158);
or U1382 (N_1382,In_1988,N_1035);
and U1383 (N_1383,N_903,N_1144);
and U1384 (N_1384,N_977,N_1175);
nor U1385 (N_1385,In_899,N_495);
or U1386 (N_1386,N_856,N_1055);
nand U1387 (N_1387,In_22,N_1187);
nand U1388 (N_1388,In_2300,N_683);
nand U1389 (N_1389,N_648,N_727);
and U1390 (N_1390,In_2466,In_1854);
nor U1391 (N_1391,N_1161,N_760);
nand U1392 (N_1392,N_280,N_1149);
or U1393 (N_1393,N_792,N_743);
xor U1394 (N_1394,In_2352,In_482);
and U1395 (N_1395,N_1133,N_1246);
or U1396 (N_1396,N_1019,N_672);
xor U1397 (N_1397,N_865,N_419);
xnor U1398 (N_1398,N_463,N_904);
xnor U1399 (N_1399,In_2329,In_165);
or U1400 (N_1400,In_49,In_587);
nand U1401 (N_1401,In_260,N_988);
nand U1402 (N_1402,N_736,In_248);
xnor U1403 (N_1403,In_1002,N_402);
xor U1404 (N_1404,N_842,N_380);
nor U1405 (N_1405,In_682,N_1016);
xor U1406 (N_1406,N_1021,N_1113);
or U1407 (N_1407,In_2165,In_339);
and U1408 (N_1408,N_732,N_346);
nor U1409 (N_1409,In_1155,N_650);
and U1410 (N_1410,In_296,N_1157);
nand U1411 (N_1411,N_838,N_237);
nand U1412 (N_1412,In_1840,N_723);
xor U1413 (N_1413,In_685,N_1209);
and U1414 (N_1414,N_686,N_872);
and U1415 (N_1415,In_1960,In_1041);
or U1416 (N_1416,N_502,In_2456);
nor U1417 (N_1417,N_1014,In_2411);
and U1418 (N_1418,N_1047,In_1196);
or U1419 (N_1419,N_183,N_778);
nor U1420 (N_1420,N_998,In_1212);
xor U1421 (N_1421,N_126,N_939);
nand U1422 (N_1422,N_765,N_762);
nand U1423 (N_1423,N_182,N_313);
nand U1424 (N_1424,In_87,In_681);
nand U1425 (N_1425,N_864,N_949);
or U1426 (N_1426,N_966,N_836);
nand U1427 (N_1427,N_392,N_1208);
nand U1428 (N_1428,N_729,N_725);
or U1429 (N_1429,In_1913,N_1114);
or U1430 (N_1430,N_636,N_1207);
or U1431 (N_1431,N_1103,N_846);
nand U1432 (N_1432,N_866,N_448);
and U1433 (N_1433,N_1137,N_630);
nor U1434 (N_1434,N_922,In_2111);
and U1435 (N_1435,N_657,N_195);
and U1436 (N_1436,N_1223,N_861);
xor U1437 (N_1437,N_757,N_979);
nor U1438 (N_1438,N_1204,N_523);
xor U1439 (N_1439,N_875,N_965);
xor U1440 (N_1440,In_253,N_236);
or U1441 (N_1441,N_1213,In_1898);
xor U1442 (N_1442,N_572,N_414);
or U1443 (N_1443,N_668,N_1128);
and U1444 (N_1444,N_730,N_676);
xor U1445 (N_1445,In_1451,N_809);
or U1446 (N_1446,N_372,In_55);
nor U1447 (N_1447,N_1098,N_811);
and U1448 (N_1448,N_837,In_1728);
nand U1449 (N_1449,N_1180,N_1033);
xnor U1450 (N_1450,In_945,N_299);
xor U1451 (N_1451,N_750,N_512);
nor U1452 (N_1452,In_837,N_296);
and U1453 (N_1453,N_537,In_1562);
nand U1454 (N_1454,In_329,In_311);
xor U1455 (N_1455,N_530,N_695);
nor U1456 (N_1456,N_1078,N_1083);
nor U1457 (N_1457,N_764,In_2488);
nor U1458 (N_1458,N_789,N_1238);
and U1459 (N_1459,In_2448,In_1303);
xor U1460 (N_1460,N_853,N_854);
nor U1461 (N_1461,N_1210,N_585);
nand U1462 (N_1462,N_886,N_571);
nor U1463 (N_1463,N_937,N_1013);
xor U1464 (N_1464,In_891,In_1683);
nand U1465 (N_1465,N_1053,In_730);
nand U1466 (N_1466,N_739,N_1102);
nor U1467 (N_1467,In_1153,N_942);
nand U1468 (N_1468,N_1003,N_644);
and U1469 (N_1469,N_759,In_1594);
xnor U1470 (N_1470,N_824,N_345);
nand U1471 (N_1471,In_292,N_662);
or U1472 (N_1472,In_1421,In_1218);
and U1473 (N_1473,N_742,N_1119);
nand U1474 (N_1474,In_1098,N_1052);
xor U1475 (N_1475,N_954,In_293);
and U1476 (N_1476,N_1117,N_980);
or U1477 (N_1477,In_2094,N_1069);
nor U1478 (N_1478,N_680,N_1020);
xnor U1479 (N_1479,N_485,N_621);
and U1480 (N_1480,In_742,N_1062);
nand U1481 (N_1481,N_944,N_763);
or U1482 (N_1482,N_919,In_1629);
nor U1483 (N_1483,N_1121,In_1251);
and U1484 (N_1484,In_368,N_797);
xnor U1485 (N_1485,N_1054,In_1816);
nand U1486 (N_1486,N_1084,N_1106);
and U1487 (N_1487,In_2227,N_716);
xnor U1488 (N_1488,N_761,In_1872);
nand U1489 (N_1489,N_1123,N_1206);
and U1490 (N_1490,In_2347,N_913);
or U1491 (N_1491,N_1184,N_647);
and U1492 (N_1492,N_1022,N_1118);
or U1493 (N_1493,In_1114,In_1082);
nand U1494 (N_1494,N_286,In_342);
nand U1495 (N_1495,N_219,N_328);
or U1496 (N_1496,N_1242,N_946);
nor U1497 (N_1497,In_1604,N_1043);
nand U1498 (N_1498,N_1183,N_822);
nor U1499 (N_1499,In_1821,In_754);
or U1500 (N_1500,N_655,N_1129);
or U1501 (N_1501,N_1219,In_2349);
nor U1502 (N_1502,In_11,N_1227);
nor U1503 (N_1503,N_772,N_498);
nor U1504 (N_1504,In_2241,In_1535);
nand U1505 (N_1505,N_519,In_532);
xnor U1506 (N_1506,N_844,In_59);
or U1507 (N_1507,In_1992,N_923);
or U1508 (N_1508,N_1093,N_1160);
and U1509 (N_1509,In_1526,N_839);
or U1510 (N_1510,N_1067,In_915);
nor U1511 (N_1511,N_250,N_740);
nand U1512 (N_1512,In_1785,In_902);
nand U1513 (N_1513,N_544,N_834);
xnor U1514 (N_1514,In_2326,In_422);
nor U1515 (N_1515,In_1558,In_50);
nand U1516 (N_1516,N_290,In_847);
xor U1517 (N_1517,N_1126,N_506);
xor U1518 (N_1518,In_2297,N_766);
and U1519 (N_1519,N_389,N_1075);
nor U1520 (N_1520,In_1570,N_240);
nand U1521 (N_1521,In_1387,N_916);
and U1522 (N_1522,In_1226,In_2255);
nor U1523 (N_1523,N_652,N_1232);
and U1524 (N_1524,N_669,N_800);
nor U1525 (N_1525,N_520,N_1109);
xnor U1526 (N_1526,N_719,N_642);
and U1527 (N_1527,N_1059,N_936);
and U1528 (N_1528,In_1403,N_876);
nor U1529 (N_1529,N_1015,N_6);
nand U1530 (N_1530,N_635,N_292);
or U1531 (N_1531,N_902,In_2204);
and U1532 (N_1532,N_994,N_639);
nand U1533 (N_1533,N_358,In_991);
nor U1534 (N_1534,N_577,In_321);
and U1535 (N_1535,N_385,N_1225);
nor U1536 (N_1536,N_68,N_1231);
nor U1537 (N_1537,In_1673,N_900);
or U1538 (N_1538,N_847,N_715);
nand U1539 (N_1539,N_1170,N_829);
xor U1540 (N_1540,N_1203,N_785);
or U1541 (N_1541,N_614,N_1018);
xor U1542 (N_1542,In_576,N_487);
or U1543 (N_1543,N_257,In_2261);
or U1544 (N_1544,N_995,N_57);
nand U1545 (N_1545,N_1116,N_1189);
or U1546 (N_1546,N_684,N_660);
xnor U1547 (N_1547,N_631,N_914);
nor U1548 (N_1548,In_626,N_833);
or U1549 (N_1549,In_1627,In_336);
and U1550 (N_1550,In_1808,In_495);
and U1551 (N_1551,N_1217,N_1200);
nor U1552 (N_1552,N_637,N_951);
or U1553 (N_1553,N_755,In_1588);
or U1554 (N_1554,N_828,N_112);
or U1555 (N_1555,N_895,In_2274);
or U1556 (N_1556,N_645,N_1027);
nand U1557 (N_1557,N_387,N_897);
and U1558 (N_1558,N_737,N_1006);
nor U1559 (N_1559,In_2342,N_654);
xnor U1560 (N_1560,N_432,N_179);
or U1561 (N_1561,In_2469,N_1176);
xor U1562 (N_1562,In_2284,N_1074);
and U1563 (N_1563,N_1138,N_909);
xor U1564 (N_1564,In_2104,In_1518);
or U1565 (N_1565,N_1233,In_130);
nand U1566 (N_1566,N_3,N_756);
nand U1567 (N_1567,N_987,N_992);
nor U1568 (N_1568,N_981,In_174);
nand U1569 (N_1569,N_911,N_982);
nand U1570 (N_1570,In_1773,N_978);
and U1571 (N_1571,N_972,In_1051);
nor U1572 (N_1572,N_891,In_938);
nand U1573 (N_1573,N_661,N_927);
and U1574 (N_1574,In_1096,N_933);
nand U1575 (N_1575,N_1010,In_821);
nand U1576 (N_1576,N_714,N_1039);
and U1577 (N_1577,N_356,In_1252);
nor U1578 (N_1578,N_649,In_970);
xor U1579 (N_1579,N_1004,N_1125);
and U1580 (N_1580,N_1150,N_782);
and U1581 (N_1581,N_692,N_288);
or U1582 (N_1582,N_689,N_412);
xor U1583 (N_1583,In_1163,N_969);
and U1584 (N_1584,In_1610,N_841);
nor U1585 (N_1585,N_1048,In_2470);
or U1586 (N_1586,In_1227,In_317);
nor U1587 (N_1587,N_1046,In_1404);
and U1588 (N_1588,N_708,N_1156);
nand U1589 (N_1589,N_606,N_827);
nand U1590 (N_1590,N_787,N_790);
and U1591 (N_1591,N_1182,N_300);
nand U1592 (N_1592,N_1248,N_997);
nand U1593 (N_1593,N_859,N_947);
nand U1594 (N_1594,N_705,N_1241);
and U1595 (N_1595,In_1514,N_1092);
xnor U1596 (N_1596,N_2,In_234);
xnor U1597 (N_1597,N_1195,N_26);
or U1598 (N_1598,N_883,In_552);
and U1599 (N_1599,N_7,N_1071);
nor U1600 (N_1600,N_1050,N_687);
nand U1601 (N_1601,N_802,N_807);
and U1602 (N_1602,N_420,In_1825);
nor U1603 (N_1603,N_971,In_1301);
or U1604 (N_1604,N_1080,In_37);
xor U1605 (N_1605,In_874,N_701);
nand U1606 (N_1606,In_2156,In_216);
xor U1607 (N_1607,In_1235,In_1206);
xor U1608 (N_1608,In_509,N_777);
nand U1609 (N_1609,N_803,In_1541);
and U1610 (N_1610,N_118,N_1141);
nand U1611 (N_1611,N_905,In_381);
nor U1612 (N_1612,In_815,In_67);
or U1613 (N_1613,N_989,In_1054);
and U1614 (N_1614,In_1880,N_1222);
xnor U1615 (N_1615,N_898,N_711);
and U1616 (N_1616,N_794,In_1564);
and U1617 (N_1617,N_691,In_2455);
nor U1618 (N_1618,In_2132,N_89);
nor U1619 (N_1619,In_2381,N_1041);
xnor U1620 (N_1620,N_151,N_1155);
xor U1621 (N_1621,N_670,In_1969);
nand U1622 (N_1622,In_1656,N_813);
nand U1623 (N_1623,N_702,In_985);
nand U1624 (N_1624,In_644,N_912);
and U1625 (N_1625,In_1661,N_1110);
and U1626 (N_1626,N_559,N_849);
or U1627 (N_1627,N_986,N_634);
xor U1628 (N_1628,N_1192,N_1057);
or U1629 (N_1629,N_1245,N_625);
nor U1630 (N_1630,N_1142,N_1026);
nand U1631 (N_1631,In_1395,N_1089);
and U1632 (N_1632,N_806,N_921);
nor U1633 (N_1633,N_1174,In_156);
nand U1634 (N_1634,N_801,In_676);
nand U1635 (N_1635,In_2422,N_685);
or U1636 (N_1636,N_302,N_627);
xor U1637 (N_1637,In_2196,In_490);
and U1638 (N_1638,In_245,N_781);
and U1639 (N_1639,N_974,N_964);
or U1640 (N_1640,N_1168,In_2185);
and U1641 (N_1641,In_2202,N_920);
and U1642 (N_1642,N_1224,N_896);
xor U1643 (N_1643,In_986,N_1165);
or U1644 (N_1644,N_700,N_492);
nor U1645 (N_1645,In_2316,In_163);
or U1646 (N_1646,In_2186,In_78);
nand U1647 (N_1647,N_735,N_1169);
nor U1648 (N_1648,N_901,N_363);
nand U1649 (N_1649,In_819,In_2405);
nor U1650 (N_1650,N_746,In_196);
and U1651 (N_1651,In_935,In_72);
nand U1652 (N_1652,In_946,N_1135);
nor U1653 (N_1653,N_632,N_1023);
xnor U1654 (N_1654,In_2046,In_1517);
and U1655 (N_1655,In_2071,In_93);
and U1656 (N_1656,N_90,N_439);
or U1657 (N_1657,In_1829,N_775);
xor U1658 (N_1658,In_1397,In_1799);
and U1659 (N_1659,In_1113,N_1139);
or U1660 (N_1660,In_1069,N_999);
and U1661 (N_1661,N_881,In_2219);
and U1662 (N_1662,In_2034,N_1158);
nand U1663 (N_1663,N_1172,In_503);
xnor U1664 (N_1664,N_870,N_1001);
nand U1665 (N_1665,N_880,N_751);
nor U1666 (N_1666,N_882,N_1100);
and U1667 (N_1667,N_721,N_805);
or U1668 (N_1668,N_1122,N_867);
or U1669 (N_1669,N_758,In_1423);
or U1670 (N_1670,N_843,In_2082);
nand U1671 (N_1671,N_1095,In_2021);
and U1672 (N_1672,N_784,In_1725);
or U1673 (N_1673,In_2358,N_848);
xnor U1674 (N_1674,N_1012,In_1962);
nor U1675 (N_1675,In_2454,N_1034);
or U1676 (N_1676,N_679,N_1193);
nor U1677 (N_1677,N_852,N_1124);
and U1678 (N_1678,In_2287,In_144);
nand U1679 (N_1679,In_1790,In_1600);
nor U1680 (N_1680,In_1897,N_879);
xnor U1681 (N_1681,In_1001,N_823);
xnor U1682 (N_1682,In_425,N_863);
or U1683 (N_1683,In_112,N_928);
xnor U1684 (N_1684,In_2369,N_1134);
xor U1685 (N_1685,In_728,In_897);
and U1686 (N_1686,N_973,In_162);
nor U1687 (N_1687,In_1367,N_1229);
or U1688 (N_1688,N_592,In_1006);
or U1689 (N_1689,In_1663,N_443);
nor U1690 (N_1690,N_1228,N_47);
and U1691 (N_1691,In_1987,N_185);
nor U1692 (N_1692,In_822,N_228);
and U1693 (N_1693,N_45,N_703);
nand U1694 (N_1694,N_278,In_1708);
nand U1695 (N_1695,N_1152,N_1236);
xnor U1696 (N_1696,N_659,N_500);
nor U1697 (N_1697,N_1235,N_60);
and U1698 (N_1698,N_796,N_821);
xor U1699 (N_1699,In_1805,In_757);
xor U1700 (N_1700,N_1037,In_1565);
or U1701 (N_1701,In_236,N_607);
or U1702 (N_1702,In_1215,N_64);
and U1703 (N_1703,N_1190,N_1040);
nor U1704 (N_1704,N_893,N_698);
nand U1705 (N_1705,In_1639,In_814);
or U1706 (N_1706,N_955,N_1154);
and U1707 (N_1707,In_1485,In_600);
xnor U1708 (N_1708,N_473,In_16);
nand U1709 (N_1709,N_817,N_906);
and U1710 (N_1710,N_73,N_1036);
nor U1711 (N_1711,In_1264,N_1105);
and U1712 (N_1712,In_1976,N_990);
nand U1713 (N_1713,N_941,In_2085);
or U1714 (N_1714,N_1179,N_437);
nor U1715 (N_1715,In_1652,N_223);
xnor U1716 (N_1716,N_888,N_1042);
nand U1717 (N_1717,N_677,N_260);
nand U1718 (N_1718,N_850,In_2444);
nand U1719 (N_1719,N_728,N_688);
nand U1720 (N_1720,In_2048,N_889);
and U1721 (N_1721,N_1215,N_496);
and U1722 (N_1722,In_1951,N_935);
or U1723 (N_1723,In_77,In_1734);
or U1724 (N_1724,N_1230,N_908);
xnor U1725 (N_1725,In_1476,In_2254);
xnor U1726 (N_1726,In_2060,In_841);
and U1727 (N_1727,N_884,In_957);
nor U1728 (N_1728,N_767,N_247);
xor U1729 (N_1729,N_1031,In_1746);
and U1730 (N_1730,N_325,In_1671);
or U1731 (N_1731,In_1408,N_1044);
and U1732 (N_1732,N_706,N_826);
and U1733 (N_1733,N_132,N_1077);
and U1734 (N_1734,N_298,N_1086);
or U1735 (N_1735,N_885,N_887);
and U1736 (N_1736,N_172,N_812);
and U1737 (N_1737,N_754,In_1697);
and U1738 (N_1738,In_1764,N_1153);
and U1739 (N_1739,N_1185,N_233);
nand U1740 (N_1740,N_1147,N_1104);
nor U1741 (N_1741,In_1899,In_2345);
nor U1742 (N_1742,In_1634,In_301);
or U1743 (N_1743,In_697,N_918);
and U1744 (N_1744,In_1892,N_1221);
nand U1745 (N_1745,N_1063,N_1201);
xnor U1746 (N_1746,In_2311,In_113);
and U1747 (N_1747,N_734,N_791);
xor U1748 (N_1748,N_962,N_143);
nor U1749 (N_1749,In_1425,N_629);
nand U1750 (N_1750,N_984,N_1064);
nand U1751 (N_1751,N_675,In_1071);
nand U1752 (N_1752,In_375,In_1482);
or U1753 (N_1753,N_713,N_722);
nand U1754 (N_1754,N_1146,N_788);
nand U1755 (N_1755,In_2275,N_186);
nand U1756 (N_1756,N_241,N_1234);
and U1757 (N_1757,In_1761,N_602);
nand U1758 (N_1758,N_786,In_1642);
nand U1759 (N_1759,In_1305,N_779);
and U1760 (N_1760,In_461,N_970);
nor U1761 (N_1761,N_23,In_1566);
and U1762 (N_1762,N_798,N_710);
nor U1763 (N_1763,N_1011,In_230);
and U1764 (N_1764,In_924,In_989);
nor U1765 (N_1765,N_1247,In_51);
nand U1766 (N_1766,N_1197,In_1622);
nor U1767 (N_1767,N_924,N_352);
nor U1768 (N_1768,In_1422,In_1574);
nand U1769 (N_1769,N_605,N_697);
nand U1770 (N_1770,N_1244,N_1216);
nand U1771 (N_1771,N_1061,N_623);
xnor U1772 (N_1772,N_139,N_1188);
or U1773 (N_1773,In_35,In_2057);
nor U1774 (N_1774,N_948,N_878);
or U1775 (N_1775,N_931,N_793);
xnor U1776 (N_1776,N_400,N_525);
and U1777 (N_1777,N_724,In_2388);
nor U1778 (N_1778,In_1501,N_771);
or U1779 (N_1779,N_871,N_945);
xor U1780 (N_1780,In_2178,N_957);
xor U1781 (N_1781,In_2188,N_1181);
and U1782 (N_1782,N_830,In_1313);
nand U1783 (N_1783,N_1032,N_943);
nor U1784 (N_1784,In_1937,In_192);
nand U1785 (N_1785,N_491,N_1101);
xnor U1786 (N_1786,N_814,N_748);
xnor U1787 (N_1787,In_770,In_2119);
nand U1788 (N_1788,N_456,N_818);
and U1789 (N_1789,N_749,N_593);
nor U1790 (N_1790,In_176,N_1120);
nor U1791 (N_1791,In_2237,N_1164);
nand U1792 (N_1792,N_373,In_796);
or U1793 (N_1793,N_733,N_810);
nor U1794 (N_1794,N_74,N_907);
nand U1795 (N_1795,N_707,N_1065);
or U1796 (N_1796,N_229,N_671);
nand U1797 (N_1797,In_2374,N_917);
xnor U1798 (N_1798,N_681,N_227);
nand U1799 (N_1799,N_855,In_1347);
nor U1800 (N_1800,N_1091,N_963);
nor U1801 (N_1801,In_1222,N_339);
and U1802 (N_1802,N_1196,In_187);
xor U1803 (N_1803,N_1097,In_1636);
xnor U1804 (N_1804,In_1985,N_1082);
nor U1805 (N_1805,N_474,In_501);
xor U1806 (N_1806,N_1029,N_958);
xor U1807 (N_1807,N_709,N_950);
nand U1808 (N_1808,N_1087,In_308);
or U1809 (N_1809,N_1060,N_717);
xnor U1810 (N_1810,N_1085,In_1342);
nand U1811 (N_1811,N_245,N_731);
or U1812 (N_1812,N_590,In_737);
nand U1813 (N_1813,In_1070,In_1581);
xnor U1814 (N_1814,In_252,In_1860);
xor U1815 (N_1815,In_1920,N_1191);
xnor U1816 (N_1816,N_1163,In_1046);
nor U1817 (N_1817,N_783,In_2280);
and U1818 (N_1818,In_1688,N_243);
and U1819 (N_1819,N_934,N_1249);
nand U1820 (N_1820,N_536,In_285);
xnor U1821 (N_1821,N_646,N_191);
nand U1822 (N_1822,In_1456,In_2387);
or U1823 (N_1823,N_148,In_1160);
or U1824 (N_1824,N_656,N_956);
xor U1825 (N_1825,N_405,N_159);
nand U1826 (N_1826,In_941,In_621);
nand U1827 (N_1827,In_1979,N_1002);
nor U1828 (N_1828,N_337,N_961);
nand U1829 (N_1829,In_2273,N_27);
nand U1830 (N_1830,N_1049,In_865);
nand U1831 (N_1831,N_1194,In_391);
and U1832 (N_1832,N_91,N_282);
nor U1833 (N_1833,In_1428,In_2175);
nor U1834 (N_1834,N_932,N_892);
nand U1835 (N_1835,In_937,N_890);
and U1836 (N_1836,In_773,In_2245);
nand U1837 (N_1837,N_36,In_1989);
xor U1838 (N_1838,N_874,N_88);
and U1839 (N_1839,N_1240,N_193);
nand U1840 (N_1840,N_744,In_258);
or U1841 (N_1841,N_1226,In_312);
nor U1842 (N_1842,In_2026,N_712);
and U1843 (N_1843,N_1000,N_527);
or U1844 (N_1844,N_780,N_1198);
xor U1845 (N_1845,N_745,N_968);
nand U1846 (N_1846,In_808,N_816);
and U1847 (N_1847,N_693,In_1506);
xor U1848 (N_1848,In_504,N_1171);
xor U1849 (N_1849,In_699,N_667);
nor U1850 (N_1850,N_1214,N_13);
nand U1851 (N_1851,In_2262,N_696);
nor U1852 (N_1852,In_1413,N_1220);
nor U1853 (N_1853,N_98,N_877);
or U1854 (N_1854,In_2084,N_718);
nor U1855 (N_1855,In_2215,N_915);
xor U1856 (N_1856,N_421,In_430);
and U1857 (N_1857,N_69,In_1025);
and U1858 (N_1858,N_1038,N_254);
or U1859 (N_1859,N_868,N_1178);
xnor U1860 (N_1860,N_835,In_840);
xnor U1861 (N_1861,N_1111,In_674);
nor U1862 (N_1862,In_1377,N_1173);
xor U1863 (N_1863,In_1767,N_467);
xor U1864 (N_1864,In_2340,N_752);
xor U1865 (N_1865,In_905,N_959);
or U1866 (N_1866,In_2040,In_553);
nand U1867 (N_1867,In_2067,N_690);
nor U1868 (N_1868,In_866,N_1130);
or U1869 (N_1869,N_8,N_154);
or U1870 (N_1870,N_938,N_164);
nand U1871 (N_1871,N_640,In_414);
nor U1872 (N_1872,In_53,In_2249);
nand U1873 (N_1873,N_1202,N_641);
nand U1874 (N_1874,N_549,N_1081);
nor U1875 (N_1875,N_1787,N_1360);
xnor U1876 (N_1876,N_1683,N_1761);
and U1877 (N_1877,N_1476,N_1505);
and U1878 (N_1878,N_1276,N_1722);
and U1879 (N_1879,N_1731,N_1517);
and U1880 (N_1880,N_1661,N_1638);
or U1881 (N_1881,N_1350,N_1671);
or U1882 (N_1882,N_1569,N_1481);
nand U1883 (N_1883,N_1670,N_1837);
nand U1884 (N_1884,N_1448,N_1408);
or U1885 (N_1885,N_1327,N_1858);
nand U1886 (N_1886,N_1834,N_1654);
xnor U1887 (N_1887,N_1778,N_1462);
xor U1888 (N_1888,N_1873,N_1449);
or U1889 (N_1889,N_1277,N_1690);
or U1890 (N_1890,N_1788,N_1428);
nor U1891 (N_1891,N_1635,N_1626);
and U1892 (N_1892,N_1715,N_1378);
and U1893 (N_1893,N_1496,N_1744);
xnor U1894 (N_1894,N_1805,N_1599);
nand U1895 (N_1895,N_1550,N_1803);
nand U1896 (N_1896,N_1824,N_1321);
nor U1897 (N_1897,N_1614,N_1820);
nand U1898 (N_1898,N_1611,N_1868);
or U1899 (N_1899,N_1621,N_1774);
nor U1900 (N_1900,N_1827,N_1594);
xor U1901 (N_1901,N_1632,N_1431);
or U1902 (N_1902,N_1850,N_1831);
xor U1903 (N_1903,N_1395,N_1317);
or U1904 (N_1904,N_1328,N_1301);
and U1905 (N_1905,N_1846,N_1510);
nand U1906 (N_1906,N_1374,N_1392);
nor U1907 (N_1907,N_1798,N_1503);
nor U1908 (N_1908,N_1602,N_1736);
nor U1909 (N_1909,N_1261,N_1279);
nand U1910 (N_1910,N_1764,N_1393);
nor U1911 (N_1911,N_1734,N_1274);
xnor U1912 (N_1912,N_1582,N_1718);
or U1913 (N_1913,N_1482,N_1367);
xor U1914 (N_1914,N_1862,N_1593);
nand U1915 (N_1915,N_1441,N_1511);
or U1916 (N_1916,N_1800,N_1600);
xnor U1917 (N_1917,N_1664,N_1813);
nand U1918 (N_1918,N_1839,N_1304);
nor U1919 (N_1919,N_1291,N_1863);
xor U1920 (N_1920,N_1762,N_1561);
and U1921 (N_1921,N_1598,N_1270);
or U1922 (N_1922,N_1533,N_1292);
nor U1923 (N_1923,N_1495,N_1275);
xor U1924 (N_1924,N_1676,N_1865);
xor U1925 (N_1925,N_1283,N_1498);
nand U1926 (N_1926,N_1713,N_1405);
nor U1927 (N_1927,N_1775,N_1726);
or U1928 (N_1928,N_1413,N_1695);
nor U1929 (N_1929,N_1337,N_1456);
and U1930 (N_1930,N_1454,N_1287);
nor U1931 (N_1931,N_1361,N_1332);
nor U1932 (N_1932,N_1771,N_1544);
nand U1933 (N_1933,N_1346,N_1570);
xor U1934 (N_1934,N_1564,N_1601);
xor U1935 (N_1935,N_1860,N_1869);
and U1936 (N_1936,N_1574,N_1555);
nor U1937 (N_1937,N_1535,N_1520);
nor U1938 (N_1938,N_1766,N_1375);
and U1939 (N_1939,N_1747,N_1484);
nor U1940 (N_1940,N_1595,N_1382);
xnor U1941 (N_1941,N_1351,N_1666);
or U1942 (N_1942,N_1607,N_1492);
and U1943 (N_1943,N_1323,N_1272);
xnor U1944 (N_1944,N_1667,N_1857);
or U1945 (N_1945,N_1723,N_1658);
and U1946 (N_1946,N_1606,N_1821);
nand U1947 (N_1947,N_1825,N_1490);
nand U1948 (N_1948,N_1310,N_1547);
or U1949 (N_1949,N_1467,N_1325);
xor U1950 (N_1950,N_1864,N_1721);
xor U1951 (N_1951,N_1472,N_1515);
or U1952 (N_1952,N_1725,N_1802);
or U1953 (N_1953,N_1478,N_1406);
xor U1954 (N_1954,N_1691,N_1302);
nand U1955 (N_1955,N_1712,N_1772);
and U1956 (N_1956,N_1866,N_1296);
nor U1957 (N_1957,N_1369,N_1501);
and U1958 (N_1958,N_1315,N_1700);
nor U1959 (N_1959,N_1568,N_1603);
xor U1960 (N_1960,N_1388,N_1326);
xnor U1961 (N_1961,N_1684,N_1765);
nand U1962 (N_1962,N_1580,N_1330);
nand U1963 (N_1963,N_1256,N_1319);
nor U1964 (N_1964,N_1612,N_1303);
and U1965 (N_1965,N_1266,N_1867);
xnor U1966 (N_1966,N_1417,N_1453);
nand U1967 (N_1967,N_1280,N_1767);
and U1968 (N_1968,N_1814,N_1504);
and U1969 (N_1969,N_1331,N_1259);
nor U1970 (N_1970,N_1418,N_1724);
nand U1971 (N_1971,N_1752,N_1347);
nor U1972 (N_1972,N_1450,N_1500);
nand U1973 (N_1973,N_1349,N_1760);
or U1974 (N_1974,N_1634,N_1565);
xnor U1975 (N_1975,N_1637,N_1556);
nor U1976 (N_1976,N_1459,N_1297);
nand U1977 (N_1977,N_1733,N_1542);
or U1978 (N_1978,N_1491,N_1642);
nor U1979 (N_1979,N_1541,N_1719);
and U1980 (N_1980,N_1681,N_1262);
nor U1981 (N_1981,N_1659,N_1352);
or U1982 (N_1982,N_1548,N_1845);
and U1983 (N_1983,N_1797,N_1464);
nand U1984 (N_1984,N_1759,N_1358);
nor U1985 (N_1985,N_1372,N_1306);
and U1986 (N_1986,N_1288,N_1414);
and U1987 (N_1987,N_1750,N_1465);
nand U1988 (N_1988,N_1420,N_1438);
nor U1989 (N_1989,N_1596,N_1651);
xor U1990 (N_1990,N_1730,N_1540);
xor U1991 (N_1991,N_1254,N_1429);
xor U1992 (N_1992,N_1471,N_1436);
xor U1993 (N_1993,N_1625,N_1604);
nor U1994 (N_1994,N_1322,N_1313);
nand U1995 (N_1995,N_1631,N_1257);
and U1996 (N_1996,N_1353,N_1575);
xnor U1997 (N_1997,N_1644,N_1793);
nor U1998 (N_1998,N_1763,N_1697);
xor U1999 (N_1999,N_1253,N_1649);
xor U2000 (N_2000,N_1679,N_1529);
xnor U2001 (N_2001,N_1663,N_1460);
or U2002 (N_2002,N_1271,N_1410);
nor U2003 (N_2003,N_1320,N_1615);
or U2004 (N_2004,N_1545,N_1657);
or U2005 (N_2005,N_1693,N_1300);
nor U2006 (N_2006,N_1643,N_1489);
nand U2007 (N_2007,N_1707,N_1412);
xor U2008 (N_2008,N_1610,N_1789);
and U2009 (N_2009,N_1356,N_1342);
xor U2010 (N_2010,N_1870,N_1442);
or U2011 (N_2011,N_1250,N_1399);
xor U2012 (N_2012,N_1488,N_1840);
nand U2013 (N_2013,N_1779,N_1776);
nor U2014 (N_2014,N_1251,N_1578);
nand U2015 (N_2015,N_1738,N_1385);
and U2016 (N_2016,N_1507,N_1685);
or U2017 (N_2017,N_1512,N_1377);
or U2018 (N_2018,N_1808,N_1758);
nor U2019 (N_2019,N_1427,N_1841);
nand U2020 (N_2020,N_1397,N_1407);
xnor U2021 (N_2021,N_1656,N_1794);
nor U2022 (N_2022,N_1273,N_1451);
nand U2023 (N_2023,N_1403,N_1588);
or U2024 (N_2024,N_1745,N_1716);
nand U2025 (N_2025,N_1314,N_1849);
nor U2026 (N_2026,N_1391,N_1786);
nor U2027 (N_2027,N_1648,N_1720);
or U2028 (N_2028,N_1608,N_1781);
nor U2029 (N_2029,N_1305,N_1461);
xor U2030 (N_2030,N_1286,N_1483);
xnor U2031 (N_2031,N_1526,N_1368);
nand U2032 (N_2032,N_1636,N_1829);
xnor U2033 (N_2033,N_1267,N_1335);
and U2034 (N_2034,N_1307,N_1737);
nand U2035 (N_2035,N_1662,N_1514);
xnor U2036 (N_2036,N_1705,N_1255);
xor U2037 (N_2037,N_1530,N_1572);
or U2038 (N_2038,N_1424,N_1379);
nand U2039 (N_2039,N_1795,N_1422);
nor U2040 (N_2040,N_1586,N_1702);
and U2041 (N_2041,N_1278,N_1419);
or U2042 (N_2042,N_1289,N_1842);
nand U2043 (N_2043,N_1861,N_1401);
nand U2044 (N_2044,N_1852,N_1411);
nor U2045 (N_2045,N_1345,N_1708);
nor U2046 (N_2046,N_1282,N_1365);
or U2047 (N_2047,N_1680,N_1381);
nand U2048 (N_2048,N_1640,N_1576);
xnor U2049 (N_2049,N_1329,N_1415);
nand U2050 (N_2050,N_1284,N_1872);
xor U2051 (N_2051,N_1728,N_1435);
nor U2052 (N_2052,N_1742,N_1366);
nor U2053 (N_2053,N_1669,N_1573);
nor U2054 (N_2054,N_1689,N_1692);
xor U2055 (N_2055,N_1686,N_1466);
nor U2056 (N_2056,N_1694,N_1710);
and U2057 (N_2057,N_1709,N_1387);
nor U2058 (N_2058,N_1566,N_1613);
xor U2059 (N_2059,N_1359,N_1678);
nand U2060 (N_2060,N_1717,N_1318);
nor U2061 (N_2061,N_1749,N_1784);
nor U2062 (N_2062,N_1714,N_1704);
nor U2063 (N_2063,N_1457,N_1502);
or U2064 (N_2064,N_1609,N_1258);
nand U2065 (N_2065,N_1735,N_1437);
xor U2066 (N_2066,N_1687,N_1620);
or U2067 (N_2067,N_1826,N_1477);
or U2068 (N_2068,N_1660,N_1338);
nor U2069 (N_2069,N_1421,N_1818);
nor U2070 (N_2070,N_1536,N_1316);
and U2071 (N_2071,N_1344,N_1809);
and U2072 (N_2072,N_1398,N_1558);
nor U2073 (N_2073,N_1592,N_1295);
or U2074 (N_2074,N_1812,N_1706);
and U2075 (N_2075,N_1519,N_1807);
or U2076 (N_2076,N_1581,N_1518);
nor U2077 (N_2077,N_1817,N_1384);
and U2078 (N_2078,N_1754,N_1383);
xnor U2079 (N_2079,N_1843,N_1585);
xor U2080 (N_2080,N_1755,N_1551);
xor U2081 (N_2081,N_1538,N_1583);
or U2082 (N_2082,N_1554,N_1757);
or U2083 (N_2083,N_1783,N_1339);
xnor U2084 (N_2084,N_1348,N_1523);
nand U2085 (N_2085,N_1486,N_1796);
nor U2086 (N_2086,N_1298,N_1263);
and U2087 (N_2087,N_1838,N_1311);
nand U2088 (N_2088,N_1493,N_1739);
xor U2089 (N_2089,N_1562,N_1380);
nor U2090 (N_2090,N_1853,N_1455);
nand U2091 (N_2091,N_1357,N_1816);
or U2092 (N_2092,N_1355,N_1376);
and U2093 (N_2093,N_1688,N_1790);
xnor U2094 (N_2094,N_1506,N_1281);
nor U2095 (N_2095,N_1285,N_1268);
or U2096 (N_2096,N_1452,N_1597);
nand U2097 (N_2097,N_1830,N_1605);
nand U2098 (N_2098,N_1426,N_1549);
nor U2099 (N_2099,N_1468,N_1386);
or U2100 (N_2100,N_1823,N_1703);
xor U2101 (N_2101,N_1537,N_1434);
nor U2102 (N_2102,N_1782,N_1701);
xor U2103 (N_2103,N_1336,N_1856);
or U2104 (N_2104,N_1364,N_1832);
or U2105 (N_2105,N_1851,N_1645);
and U2106 (N_2106,N_1447,N_1470);
or U2107 (N_2107,N_1354,N_1362);
nand U2108 (N_2108,N_1810,N_1390);
xor U2109 (N_2109,N_1508,N_1652);
and U2110 (N_2110,N_1756,N_1539);
nor U2111 (N_2111,N_1532,N_1463);
nand U2112 (N_2112,N_1524,N_1633);
or U2113 (N_2113,N_1743,N_1469);
or U2114 (N_2114,N_1650,N_1698);
nand U2115 (N_2115,N_1553,N_1741);
nand U2116 (N_2116,N_1677,N_1416);
nand U2117 (N_2117,N_1711,N_1836);
xor U2118 (N_2118,N_1647,N_1260);
nand U2119 (N_2119,N_1509,N_1440);
nor U2120 (N_2120,N_1293,N_1567);
nand U2121 (N_2121,N_1806,N_1312);
nor U2122 (N_2122,N_1859,N_1373);
and U2123 (N_2123,N_1791,N_1815);
and U2124 (N_2124,N_1389,N_1425);
nand U2125 (N_2125,N_1430,N_1522);
xor U2126 (N_2126,N_1521,N_1753);
xor U2127 (N_2127,N_1871,N_1400);
nand U2128 (N_2128,N_1746,N_1579);
nor U2129 (N_2129,N_1528,N_1627);
nor U2130 (N_2130,N_1363,N_1732);
xnor U2131 (N_2131,N_1748,N_1264);
or U2132 (N_2132,N_1404,N_1497);
nor U2133 (N_2133,N_1773,N_1458);
nor U2134 (N_2134,N_1584,N_1444);
or U2135 (N_2135,N_1785,N_1623);
or U2136 (N_2136,N_1780,N_1587);
or U2137 (N_2137,N_1769,N_1480);
nand U2138 (N_2138,N_1618,N_1443);
or U2139 (N_2139,N_1801,N_1409);
and U2140 (N_2140,N_1655,N_1252);
nor U2141 (N_2141,N_1591,N_1619);
and U2142 (N_2142,N_1616,N_1854);
xnor U2143 (N_2143,N_1396,N_1751);
nand U2144 (N_2144,N_1699,N_1768);
or U2145 (N_2145,N_1835,N_1475);
nand U2146 (N_2146,N_1589,N_1848);
nand U2147 (N_2147,N_1527,N_1792);
or U2148 (N_2148,N_1729,N_1653);
nor U2149 (N_2149,N_1543,N_1639);
or U2150 (N_2150,N_1665,N_1622);
or U2151 (N_2151,N_1674,N_1646);
nor U2152 (N_2152,N_1308,N_1499);
nor U2153 (N_2153,N_1534,N_1474);
and U2154 (N_2154,N_1855,N_1770);
or U2155 (N_2155,N_1672,N_1727);
nor U2156 (N_2156,N_1552,N_1560);
nand U2157 (N_2157,N_1847,N_1571);
nand U2158 (N_2158,N_1673,N_1269);
nor U2159 (N_2159,N_1628,N_1516);
nor U2160 (N_2160,N_1682,N_1402);
nand U2161 (N_2161,N_1844,N_1371);
or U2162 (N_2162,N_1799,N_1370);
or U2163 (N_2163,N_1333,N_1828);
nor U2164 (N_2164,N_1324,N_1675);
nor U2165 (N_2165,N_1341,N_1433);
nor U2166 (N_2166,N_1513,N_1432);
xor U2167 (N_2167,N_1479,N_1696);
nor U2168 (N_2168,N_1577,N_1531);
nand U2169 (N_2169,N_1343,N_1439);
nand U2170 (N_2170,N_1874,N_1334);
or U2171 (N_2171,N_1777,N_1309);
nor U2172 (N_2172,N_1819,N_1546);
and U2173 (N_2173,N_1423,N_1446);
or U2174 (N_2174,N_1294,N_1559);
or U2175 (N_2175,N_1485,N_1822);
or U2176 (N_2176,N_1629,N_1590);
nor U2177 (N_2177,N_1804,N_1487);
nor U2178 (N_2178,N_1624,N_1265);
nor U2179 (N_2179,N_1494,N_1668);
or U2180 (N_2180,N_1630,N_1340);
nand U2181 (N_2181,N_1740,N_1525);
and U2182 (N_2182,N_1473,N_1557);
and U2183 (N_2183,N_1290,N_1811);
nand U2184 (N_2184,N_1641,N_1445);
or U2185 (N_2185,N_1299,N_1563);
and U2186 (N_2186,N_1617,N_1394);
and U2187 (N_2187,N_1833,N_1358);
nor U2188 (N_2188,N_1450,N_1463);
nand U2189 (N_2189,N_1367,N_1437);
xnor U2190 (N_2190,N_1813,N_1289);
xnor U2191 (N_2191,N_1806,N_1560);
nand U2192 (N_2192,N_1838,N_1732);
or U2193 (N_2193,N_1751,N_1448);
xor U2194 (N_2194,N_1257,N_1861);
or U2195 (N_2195,N_1745,N_1277);
xor U2196 (N_2196,N_1386,N_1463);
xnor U2197 (N_2197,N_1380,N_1743);
and U2198 (N_2198,N_1282,N_1777);
nor U2199 (N_2199,N_1250,N_1619);
and U2200 (N_2200,N_1312,N_1531);
and U2201 (N_2201,N_1549,N_1828);
xnor U2202 (N_2202,N_1486,N_1778);
or U2203 (N_2203,N_1742,N_1447);
xor U2204 (N_2204,N_1329,N_1670);
and U2205 (N_2205,N_1670,N_1510);
nor U2206 (N_2206,N_1825,N_1851);
nor U2207 (N_2207,N_1479,N_1395);
or U2208 (N_2208,N_1325,N_1716);
nand U2209 (N_2209,N_1403,N_1639);
or U2210 (N_2210,N_1863,N_1678);
nand U2211 (N_2211,N_1403,N_1830);
nand U2212 (N_2212,N_1834,N_1755);
xor U2213 (N_2213,N_1576,N_1547);
and U2214 (N_2214,N_1720,N_1553);
nor U2215 (N_2215,N_1769,N_1753);
or U2216 (N_2216,N_1547,N_1299);
xnor U2217 (N_2217,N_1259,N_1743);
and U2218 (N_2218,N_1504,N_1372);
xor U2219 (N_2219,N_1535,N_1707);
nand U2220 (N_2220,N_1411,N_1737);
or U2221 (N_2221,N_1390,N_1421);
nand U2222 (N_2222,N_1779,N_1812);
and U2223 (N_2223,N_1406,N_1402);
or U2224 (N_2224,N_1869,N_1854);
nor U2225 (N_2225,N_1495,N_1724);
or U2226 (N_2226,N_1406,N_1491);
xor U2227 (N_2227,N_1499,N_1855);
or U2228 (N_2228,N_1806,N_1327);
nor U2229 (N_2229,N_1563,N_1475);
nand U2230 (N_2230,N_1835,N_1364);
and U2231 (N_2231,N_1632,N_1866);
nor U2232 (N_2232,N_1551,N_1509);
nand U2233 (N_2233,N_1653,N_1322);
xor U2234 (N_2234,N_1577,N_1399);
nand U2235 (N_2235,N_1807,N_1300);
nor U2236 (N_2236,N_1480,N_1333);
and U2237 (N_2237,N_1657,N_1612);
nand U2238 (N_2238,N_1551,N_1474);
and U2239 (N_2239,N_1346,N_1751);
or U2240 (N_2240,N_1641,N_1380);
or U2241 (N_2241,N_1532,N_1768);
and U2242 (N_2242,N_1716,N_1595);
nor U2243 (N_2243,N_1722,N_1455);
nand U2244 (N_2244,N_1589,N_1594);
xor U2245 (N_2245,N_1574,N_1556);
nand U2246 (N_2246,N_1718,N_1792);
and U2247 (N_2247,N_1444,N_1554);
nand U2248 (N_2248,N_1725,N_1615);
nand U2249 (N_2249,N_1690,N_1568);
xnor U2250 (N_2250,N_1441,N_1855);
xor U2251 (N_2251,N_1773,N_1313);
nand U2252 (N_2252,N_1450,N_1526);
nor U2253 (N_2253,N_1693,N_1597);
xnor U2254 (N_2254,N_1250,N_1761);
or U2255 (N_2255,N_1287,N_1532);
xnor U2256 (N_2256,N_1637,N_1291);
and U2257 (N_2257,N_1748,N_1425);
xor U2258 (N_2258,N_1834,N_1362);
and U2259 (N_2259,N_1633,N_1579);
and U2260 (N_2260,N_1325,N_1418);
nand U2261 (N_2261,N_1768,N_1849);
or U2262 (N_2262,N_1364,N_1713);
nor U2263 (N_2263,N_1742,N_1275);
nand U2264 (N_2264,N_1687,N_1780);
nor U2265 (N_2265,N_1297,N_1618);
and U2266 (N_2266,N_1262,N_1538);
or U2267 (N_2267,N_1784,N_1868);
nand U2268 (N_2268,N_1418,N_1574);
or U2269 (N_2269,N_1710,N_1386);
xor U2270 (N_2270,N_1842,N_1632);
nor U2271 (N_2271,N_1429,N_1826);
nand U2272 (N_2272,N_1296,N_1315);
and U2273 (N_2273,N_1413,N_1381);
nor U2274 (N_2274,N_1554,N_1502);
and U2275 (N_2275,N_1504,N_1714);
or U2276 (N_2276,N_1417,N_1797);
or U2277 (N_2277,N_1717,N_1378);
nor U2278 (N_2278,N_1518,N_1285);
nor U2279 (N_2279,N_1638,N_1843);
or U2280 (N_2280,N_1338,N_1839);
or U2281 (N_2281,N_1866,N_1307);
nor U2282 (N_2282,N_1451,N_1862);
and U2283 (N_2283,N_1403,N_1406);
or U2284 (N_2284,N_1417,N_1265);
nand U2285 (N_2285,N_1768,N_1639);
nor U2286 (N_2286,N_1255,N_1582);
nand U2287 (N_2287,N_1310,N_1278);
and U2288 (N_2288,N_1804,N_1604);
nor U2289 (N_2289,N_1691,N_1495);
or U2290 (N_2290,N_1819,N_1668);
xor U2291 (N_2291,N_1424,N_1335);
nor U2292 (N_2292,N_1270,N_1569);
and U2293 (N_2293,N_1304,N_1408);
or U2294 (N_2294,N_1469,N_1385);
or U2295 (N_2295,N_1632,N_1843);
and U2296 (N_2296,N_1634,N_1599);
nand U2297 (N_2297,N_1855,N_1598);
and U2298 (N_2298,N_1609,N_1379);
nand U2299 (N_2299,N_1763,N_1557);
or U2300 (N_2300,N_1873,N_1814);
nor U2301 (N_2301,N_1710,N_1785);
nand U2302 (N_2302,N_1686,N_1449);
or U2303 (N_2303,N_1497,N_1659);
xor U2304 (N_2304,N_1781,N_1405);
or U2305 (N_2305,N_1575,N_1352);
or U2306 (N_2306,N_1328,N_1807);
or U2307 (N_2307,N_1741,N_1719);
nor U2308 (N_2308,N_1859,N_1595);
xnor U2309 (N_2309,N_1643,N_1727);
or U2310 (N_2310,N_1278,N_1640);
nand U2311 (N_2311,N_1819,N_1284);
xor U2312 (N_2312,N_1570,N_1716);
xor U2313 (N_2313,N_1500,N_1663);
and U2314 (N_2314,N_1347,N_1299);
or U2315 (N_2315,N_1380,N_1596);
and U2316 (N_2316,N_1370,N_1874);
nand U2317 (N_2317,N_1600,N_1415);
nand U2318 (N_2318,N_1708,N_1709);
or U2319 (N_2319,N_1503,N_1822);
xor U2320 (N_2320,N_1326,N_1741);
or U2321 (N_2321,N_1452,N_1725);
nand U2322 (N_2322,N_1611,N_1508);
nand U2323 (N_2323,N_1389,N_1531);
and U2324 (N_2324,N_1526,N_1464);
nand U2325 (N_2325,N_1786,N_1728);
or U2326 (N_2326,N_1852,N_1686);
xor U2327 (N_2327,N_1419,N_1535);
nand U2328 (N_2328,N_1605,N_1395);
nand U2329 (N_2329,N_1473,N_1736);
and U2330 (N_2330,N_1289,N_1547);
nor U2331 (N_2331,N_1285,N_1864);
nand U2332 (N_2332,N_1339,N_1295);
or U2333 (N_2333,N_1586,N_1818);
nor U2334 (N_2334,N_1435,N_1334);
or U2335 (N_2335,N_1450,N_1786);
nand U2336 (N_2336,N_1502,N_1768);
or U2337 (N_2337,N_1288,N_1650);
and U2338 (N_2338,N_1455,N_1348);
or U2339 (N_2339,N_1326,N_1424);
xor U2340 (N_2340,N_1548,N_1777);
and U2341 (N_2341,N_1579,N_1465);
nor U2342 (N_2342,N_1676,N_1488);
nor U2343 (N_2343,N_1709,N_1376);
nand U2344 (N_2344,N_1672,N_1614);
nor U2345 (N_2345,N_1354,N_1459);
and U2346 (N_2346,N_1691,N_1305);
nand U2347 (N_2347,N_1689,N_1501);
nor U2348 (N_2348,N_1618,N_1853);
xor U2349 (N_2349,N_1296,N_1570);
or U2350 (N_2350,N_1700,N_1584);
xor U2351 (N_2351,N_1752,N_1468);
xnor U2352 (N_2352,N_1751,N_1416);
and U2353 (N_2353,N_1686,N_1513);
xnor U2354 (N_2354,N_1679,N_1655);
xnor U2355 (N_2355,N_1595,N_1755);
nor U2356 (N_2356,N_1775,N_1719);
and U2357 (N_2357,N_1633,N_1391);
and U2358 (N_2358,N_1599,N_1661);
nor U2359 (N_2359,N_1520,N_1677);
xnor U2360 (N_2360,N_1301,N_1645);
xor U2361 (N_2361,N_1282,N_1369);
nor U2362 (N_2362,N_1629,N_1528);
nor U2363 (N_2363,N_1631,N_1835);
nand U2364 (N_2364,N_1442,N_1854);
xor U2365 (N_2365,N_1323,N_1683);
or U2366 (N_2366,N_1779,N_1284);
nand U2367 (N_2367,N_1506,N_1497);
nand U2368 (N_2368,N_1460,N_1271);
xnor U2369 (N_2369,N_1648,N_1404);
or U2370 (N_2370,N_1519,N_1861);
nand U2371 (N_2371,N_1521,N_1297);
or U2372 (N_2372,N_1404,N_1672);
xor U2373 (N_2373,N_1701,N_1870);
nand U2374 (N_2374,N_1683,N_1288);
and U2375 (N_2375,N_1582,N_1326);
nand U2376 (N_2376,N_1473,N_1790);
nand U2377 (N_2377,N_1862,N_1314);
and U2378 (N_2378,N_1772,N_1465);
xnor U2379 (N_2379,N_1726,N_1698);
or U2380 (N_2380,N_1535,N_1544);
or U2381 (N_2381,N_1295,N_1279);
nand U2382 (N_2382,N_1457,N_1542);
nor U2383 (N_2383,N_1666,N_1548);
or U2384 (N_2384,N_1266,N_1777);
or U2385 (N_2385,N_1265,N_1266);
xor U2386 (N_2386,N_1514,N_1546);
nand U2387 (N_2387,N_1455,N_1381);
xnor U2388 (N_2388,N_1335,N_1466);
nor U2389 (N_2389,N_1540,N_1529);
nand U2390 (N_2390,N_1397,N_1674);
xnor U2391 (N_2391,N_1437,N_1365);
nand U2392 (N_2392,N_1281,N_1326);
nand U2393 (N_2393,N_1443,N_1778);
or U2394 (N_2394,N_1664,N_1842);
nor U2395 (N_2395,N_1865,N_1352);
or U2396 (N_2396,N_1683,N_1426);
xnor U2397 (N_2397,N_1403,N_1382);
and U2398 (N_2398,N_1322,N_1450);
nor U2399 (N_2399,N_1729,N_1841);
nor U2400 (N_2400,N_1386,N_1788);
nand U2401 (N_2401,N_1796,N_1735);
and U2402 (N_2402,N_1821,N_1868);
nor U2403 (N_2403,N_1486,N_1272);
xnor U2404 (N_2404,N_1462,N_1569);
nor U2405 (N_2405,N_1574,N_1280);
nand U2406 (N_2406,N_1716,N_1486);
xor U2407 (N_2407,N_1660,N_1445);
or U2408 (N_2408,N_1828,N_1820);
nand U2409 (N_2409,N_1659,N_1627);
nor U2410 (N_2410,N_1254,N_1859);
xor U2411 (N_2411,N_1410,N_1346);
xnor U2412 (N_2412,N_1510,N_1286);
and U2413 (N_2413,N_1376,N_1691);
xor U2414 (N_2414,N_1329,N_1324);
nor U2415 (N_2415,N_1354,N_1843);
xnor U2416 (N_2416,N_1347,N_1840);
nand U2417 (N_2417,N_1478,N_1449);
nor U2418 (N_2418,N_1622,N_1628);
xor U2419 (N_2419,N_1337,N_1681);
nand U2420 (N_2420,N_1799,N_1697);
or U2421 (N_2421,N_1715,N_1627);
nor U2422 (N_2422,N_1763,N_1475);
and U2423 (N_2423,N_1524,N_1508);
nand U2424 (N_2424,N_1405,N_1634);
or U2425 (N_2425,N_1791,N_1794);
nand U2426 (N_2426,N_1600,N_1699);
nand U2427 (N_2427,N_1556,N_1800);
nand U2428 (N_2428,N_1684,N_1285);
nor U2429 (N_2429,N_1471,N_1279);
nor U2430 (N_2430,N_1486,N_1654);
nor U2431 (N_2431,N_1856,N_1456);
nand U2432 (N_2432,N_1774,N_1666);
nor U2433 (N_2433,N_1312,N_1518);
nor U2434 (N_2434,N_1719,N_1265);
xor U2435 (N_2435,N_1414,N_1616);
xor U2436 (N_2436,N_1479,N_1506);
xnor U2437 (N_2437,N_1839,N_1366);
xnor U2438 (N_2438,N_1580,N_1797);
or U2439 (N_2439,N_1820,N_1494);
xnor U2440 (N_2440,N_1585,N_1848);
nand U2441 (N_2441,N_1688,N_1669);
nor U2442 (N_2442,N_1642,N_1594);
xnor U2443 (N_2443,N_1593,N_1420);
nand U2444 (N_2444,N_1269,N_1371);
xor U2445 (N_2445,N_1315,N_1498);
nand U2446 (N_2446,N_1403,N_1496);
nor U2447 (N_2447,N_1429,N_1852);
or U2448 (N_2448,N_1657,N_1536);
nor U2449 (N_2449,N_1515,N_1251);
and U2450 (N_2450,N_1493,N_1793);
or U2451 (N_2451,N_1755,N_1325);
nor U2452 (N_2452,N_1795,N_1386);
nor U2453 (N_2453,N_1761,N_1491);
and U2454 (N_2454,N_1872,N_1746);
and U2455 (N_2455,N_1668,N_1816);
nor U2456 (N_2456,N_1864,N_1261);
nand U2457 (N_2457,N_1873,N_1850);
and U2458 (N_2458,N_1368,N_1319);
and U2459 (N_2459,N_1577,N_1665);
nor U2460 (N_2460,N_1319,N_1417);
nor U2461 (N_2461,N_1366,N_1338);
and U2462 (N_2462,N_1443,N_1848);
and U2463 (N_2463,N_1795,N_1686);
or U2464 (N_2464,N_1264,N_1374);
nor U2465 (N_2465,N_1255,N_1755);
nand U2466 (N_2466,N_1810,N_1535);
and U2467 (N_2467,N_1290,N_1481);
nor U2468 (N_2468,N_1443,N_1373);
or U2469 (N_2469,N_1803,N_1709);
nor U2470 (N_2470,N_1443,N_1423);
nor U2471 (N_2471,N_1723,N_1304);
nand U2472 (N_2472,N_1267,N_1847);
and U2473 (N_2473,N_1585,N_1770);
nor U2474 (N_2474,N_1459,N_1253);
nand U2475 (N_2475,N_1491,N_1862);
nor U2476 (N_2476,N_1792,N_1254);
nor U2477 (N_2477,N_1759,N_1781);
and U2478 (N_2478,N_1701,N_1412);
or U2479 (N_2479,N_1722,N_1849);
nor U2480 (N_2480,N_1793,N_1414);
nor U2481 (N_2481,N_1457,N_1454);
or U2482 (N_2482,N_1450,N_1525);
and U2483 (N_2483,N_1524,N_1574);
xor U2484 (N_2484,N_1502,N_1347);
nor U2485 (N_2485,N_1485,N_1609);
xor U2486 (N_2486,N_1776,N_1375);
nor U2487 (N_2487,N_1336,N_1863);
xnor U2488 (N_2488,N_1762,N_1788);
xor U2489 (N_2489,N_1378,N_1285);
or U2490 (N_2490,N_1820,N_1794);
or U2491 (N_2491,N_1293,N_1476);
nor U2492 (N_2492,N_1801,N_1355);
and U2493 (N_2493,N_1673,N_1466);
and U2494 (N_2494,N_1817,N_1582);
xor U2495 (N_2495,N_1729,N_1805);
and U2496 (N_2496,N_1608,N_1533);
nor U2497 (N_2497,N_1500,N_1744);
nand U2498 (N_2498,N_1432,N_1816);
nand U2499 (N_2499,N_1577,N_1520);
nor U2500 (N_2500,N_1931,N_2392);
xor U2501 (N_2501,N_2039,N_2383);
and U2502 (N_2502,N_1907,N_2380);
and U2503 (N_2503,N_2201,N_2299);
or U2504 (N_2504,N_2087,N_2347);
or U2505 (N_2505,N_2377,N_1972);
nand U2506 (N_2506,N_1883,N_2181);
and U2507 (N_2507,N_2387,N_1993);
xor U2508 (N_2508,N_2165,N_2052);
nand U2509 (N_2509,N_2437,N_2375);
and U2510 (N_2510,N_2022,N_2268);
and U2511 (N_2511,N_1937,N_2461);
nand U2512 (N_2512,N_2424,N_2139);
or U2513 (N_2513,N_2489,N_2302);
nand U2514 (N_2514,N_2381,N_2356);
nand U2515 (N_2515,N_2178,N_2338);
or U2516 (N_2516,N_1939,N_1948);
nand U2517 (N_2517,N_2083,N_1949);
xor U2518 (N_2518,N_2072,N_2259);
xnor U2519 (N_2519,N_2099,N_2045);
and U2520 (N_2520,N_2197,N_2007);
or U2521 (N_2521,N_2283,N_2055);
or U2522 (N_2522,N_2315,N_1946);
and U2523 (N_2523,N_2412,N_2333);
or U2524 (N_2524,N_2255,N_2172);
nand U2525 (N_2525,N_1894,N_1991);
xor U2526 (N_2526,N_2361,N_2258);
nand U2527 (N_2527,N_2440,N_2218);
nand U2528 (N_2528,N_2325,N_2360);
nor U2529 (N_2529,N_2161,N_2293);
nor U2530 (N_2530,N_2321,N_1927);
xor U2531 (N_2531,N_1904,N_2390);
nand U2532 (N_2532,N_2183,N_2146);
and U2533 (N_2533,N_2341,N_2442);
and U2534 (N_2534,N_2038,N_1975);
xor U2535 (N_2535,N_2117,N_2213);
or U2536 (N_2536,N_2116,N_1977);
xnor U2537 (N_2537,N_2254,N_2065);
and U2538 (N_2538,N_1965,N_2068);
nand U2539 (N_2539,N_2294,N_2422);
or U2540 (N_2540,N_2173,N_1926);
nor U2541 (N_2541,N_2300,N_1910);
or U2542 (N_2542,N_2168,N_2182);
or U2543 (N_2543,N_2003,N_1921);
or U2544 (N_2544,N_2257,N_2460);
or U2545 (N_2545,N_2133,N_2014);
xor U2546 (N_2546,N_2027,N_2049);
and U2547 (N_2547,N_2285,N_1989);
nor U2548 (N_2548,N_2307,N_2247);
and U2549 (N_2549,N_2203,N_2229);
or U2550 (N_2550,N_2286,N_2102);
or U2551 (N_2551,N_2018,N_2295);
nand U2552 (N_2552,N_2042,N_2110);
xor U2553 (N_2553,N_1885,N_2048);
nor U2554 (N_2554,N_2405,N_2438);
nand U2555 (N_2555,N_1888,N_2417);
or U2556 (N_2556,N_2008,N_2323);
nor U2557 (N_2557,N_2378,N_2297);
xnor U2558 (N_2558,N_2098,N_2451);
xor U2559 (N_2559,N_2089,N_2143);
nand U2560 (N_2560,N_2249,N_1887);
and U2561 (N_2561,N_2135,N_2114);
xnor U2562 (N_2562,N_2407,N_2211);
or U2563 (N_2563,N_1982,N_2267);
xor U2564 (N_2564,N_2043,N_1919);
nand U2565 (N_2565,N_2093,N_2499);
xnor U2566 (N_2566,N_1994,N_1974);
or U2567 (N_2567,N_2192,N_2107);
nor U2568 (N_2568,N_2496,N_2482);
xnor U2569 (N_2569,N_2317,N_2382);
nand U2570 (N_2570,N_2078,N_1950);
nor U2571 (N_2571,N_1914,N_2251);
nand U2572 (N_2572,N_2147,N_2015);
nand U2573 (N_2573,N_2056,N_2033);
and U2574 (N_2574,N_2459,N_2073);
or U2575 (N_2575,N_1953,N_1979);
nor U2576 (N_2576,N_2123,N_2314);
and U2577 (N_2577,N_2063,N_2205);
and U2578 (N_2578,N_2092,N_2242);
and U2579 (N_2579,N_2413,N_2311);
nor U2580 (N_2580,N_1955,N_1875);
and U2581 (N_2581,N_2054,N_2418);
nor U2582 (N_2582,N_2406,N_2270);
and U2583 (N_2583,N_2214,N_1957);
nor U2584 (N_2584,N_2425,N_2059);
or U2585 (N_2585,N_2243,N_1902);
xor U2586 (N_2586,N_2037,N_2432);
and U2587 (N_2587,N_2219,N_2483);
xnor U2588 (N_2588,N_2106,N_2265);
nor U2589 (N_2589,N_2128,N_2109);
nor U2590 (N_2590,N_1981,N_2111);
nand U2591 (N_2591,N_2167,N_2009);
nor U2592 (N_2592,N_2274,N_1898);
nand U2593 (N_2593,N_1942,N_1878);
and U2594 (N_2594,N_2328,N_2041);
and U2595 (N_2595,N_2204,N_2455);
nand U2596 (N_2596,N_2170,N_2053);
nor U2597 (N_2597,N_2449,N_2276);
xnor U2598 (N_2598,N_2101,N_1881);
xnor U2599 (N_2599,N_2095,N_2253);
xor U2600 (N_2600,N_2391,N_2466);
nand U2601 (N_2601,N_1944,N_1935);
and U2602 (N_2602,N_2291,N_1960);
xnor U2603 (N_2603,N_1973,N_2400);
nor U2604 (N_2604,N_2031,N_2200);
and U2605 (N_2605,N_2207,N_2002);
xnor U2606 (N_2606,N_1922,N_1958);
nand U2607 (N_2607,N_2313,N_2290);
nand U2608 (N_2608,N_2419,N_2240);
and U2609 (N_2609,N_2131,N_1938);
nor U2610 (N_2610,N_1951,N_2339);
nor U2611 (N_2611,N_2184,N_2235);
or U2612 (N_2612,N_2004,N_2212);
and U2613 (N_2613,N_2248,N_2058);
xnor U2614 (N_2614,N_2061,N_2318);
xnor U2615 (N_2615,N_2046,N_2138);
or U2616 (N_2616,N_2444,N_1996);
nor U2617 (N_2617,N_1947,N_2281);
and U2618 (N_2618,N_2032,N_2084);
nor U2619 (N_2619,N_1967,N_1889);
and U2620 (N_2620,N_2086,N_2498);
or U2621 (N_2621,N_2067,N_2487);
nand U2622 (N_2622,N_1934,N_1940);
nand U2623 (N_2623,N_2233,N_2337);
and U2624 (N_2624,N_2399,N_2169);
nand U2625 (N_2625,N_2215,N_2224);
or U2626 (N_2626,N_2475,N_2241);
xor U2627 (N_2627,N_2490,N_2209);
or U2628 (N_2628,N_1968,N_2469);
or U2629 (N_2629,N_2234,N_2034);
nand U2630 (N_2630,N_2393,N_2144);
nor U2631 (N_2631,N_2222,N_2385);
xnor U2632 (N_2632,N_2485,N_2113);
and U2633 (N_2633,N_1918,N_1890);
nand U2634 (N_2634,N_2350,N_2456);
nor U2635 (N_2635,N_2035,N_2344);
and U2636 (N_2636,N_2079,N_2225);
or U2637 (N_2637,N_1984,N_1886);
or U2638 (N_2638,N_2326,N_2239);
nor U2639 (N_2639,N_1997,N_2141);
xor U2640 (N_2640,N_1908,N_2404);
and U2641 (N_2641,N_2231,N_2471);
and U2642 (N_2642,N_2023,N_2226);
xor U2643 (N_2643,N_2190,N_1998);
nand U2644 (N_2644,N_1901,N_2436);
nand U2645 (N_2645,N_2386,N_2269);
xor U2646 (N_2646,N_2127,N_2280);
and U2647 (N_2647,N_1945,N_2198);
xor U2648 (N_2648,N_2262,N_1985);
and U2649 (N_2649,N_2175,N_2358);
xor U2650 (N_2650,N_2366,N_2196);
or U2651 (N_2651,N_1900,N_2156);
nor U2652 (N_2652,N_2272,N_2051);
and U2653 (N_2653,N_2151,N_2369);
nor U2654 (N_2654,N_2408,N_2429);
or U2655 (N_2655,N_2335,N_2273);
nor U2656 (N_2656,N_2029,N_1928);
nand U2657 (N_2657,N_2473,N_2357);
nor U2658 (N_2658,N_2388,N_2077);
xnor U2659 (N_2659,N_2125,N_2316);
nand U2660 (N_2660,N_2013,N_1952);
nor U2661 (N_2661,N_2006,N_2091);
xnor U2662 (N_2662,N_1976,N_2071);
nand U2663 (N_2663,N_2403,N_2075);
nand U2664 (N_2664,N_2236,N_2080);
and U2665 (N_2665,N_2005,N_2100);
nand U2666 (N_2666,N_1983,N_2379);
nor U2667 (N_2667,N_2069,N_2465);
nand U2668 (N_2668,N_2130,N_2343);
and U2669 (N_2669,N_2480,N_2044);
and U2670 (N_2670,N_2244,N_2365);
xnor U2671 (N_2671,N_2479,N_2368);
nand U2672 (N_2672,N_2462,N_2463);
nand U2673 (N_2673,N_1970,N_2250);
xor U2674 (N_2674,N_1999,N_2433);
nand U2675 (N_2675,N_2394,N_2028);
or U2676 (N_2676,N_2266,N_2304);
xor U2677 (N_2677,N_2416,N_2186);
or U2678 (N_2678,N_2457,N_2470);
nor U2679 (N_2679,N_2486,N_2327);
nand U2680 (N_2680,N_2352,N_2137);
xnor U2681 (N_2681,N_1992,N_2142);
nor U2682 (N_2682,N_2308,N_2194);
nor U2683 (N_2683,N_2324,N_1980);
and U2684 (N_2684,N_1925,N_2047);
or U2685 (N_2685,N_1963,N_2411);
nand U2686 (N_2686,N_1879,N_2012);
nor U2687 (N_2687,N_2414,N_2094);
nor U2688 (N_2688,N_2070,N_2119);
xor U2689 (N_2689,N_1912,N_2227);
or U2690 (N_2690,N_2309,N_2264);
and U2691 (N_2691,N_2312,N_2491);
and U2692 (N_2692,N_2329,N_2342);
and U2693 (N_2693,N_2148,N_2472);
or U2694 (N_2694,N_2090,N_2395);
or U2695 (N_2695,N_2155,N_2081);
or U2696 (N_2696,N_2359,N_2149);
nand U2697 (N_2697,N_2336,N_2445);
xnor U2698 (N_2698,N_2415,N_2132);
nand U2699 (N_2699,N_2426,N_1932);
nor U2700 (N_2700,N_2064,N_2420);
xnor U2701 (N_2701,N_1961,N_2085);
nand U2702 (N_2702,N_2296,N_2275);
and U2703 (N_2703,N_2252,N_2353);
nand U2704 (N_2704,N_2376,N_2154);
nand U2705 (N_2705,N_1893,N_2474);
nor U2706 (N_2706,N_1954,N_2493);
xnor U2707 (N_2707,N_1913,N_2104);
nand U2708 (N_2708,N_2322,N_2195);
nand U2709 (N_2709,N_2026,N_1905);
xnor U2710 (N_2710,N_2289,N_2367);
nand U2711 (N_2711,N_2096,N_2246);
xnor U2712 (N_2712,N_2040,N_2024);
nand U2713 (N_2713,N_2153,N_1884);
nand U2714 (N_2714,N_2176,N_1971);
xnor U2715 (N_2715,N_2066,N_1995);
nand U2716 (N_2716,N_1987,N_2282);
nand U2717 (N_2717,N_2467,N_2431);
xor U2718 (N_2718,N_2488,N_2410);
or U2719 (N_2719,N_1930,N_2260);
or U2720 (N_2720,N_2331,N_2129);
nor U2721 (N_2721,N_1923,N_1916);
or U2722 (N_2722,N_2163,N_2363);
nor U2723 (N_2723,N_2001,N_2016);
nor U2724 (N_2724,N_2495,N_2428);
nand U2725 (N_2725,N_2208,N_1978);
nor U2726 (N_2726,N_2453,N_1936);
xor U2727 (N_2727,N_1986,N_2171);
or U2728 (N_2728,N_2216,N_2057);
or U2729 (N_2729,N_2370,N_1906);
nor U2730 (N_2730,N_2103,N_2263);
xnor U2731 (N_2731,N_2384,N_2494);
or U2732 (N_2732,N_2020,N_1903);
and U2733 (N_2733,N_2124,N_2036);
xnor U2734 (N_2734,N_2261,N_2217);
xor U2735 (N_2735,N_2160,N_2157);
xor U2736 (N_2736,N_1933,N_2450);
or U2737 (N_2737,N_2292,N_2447);
or U2738 (N_2738,N_1964,N_2346);
and U2739 (N_2739,N_2271,N_1962);
xnor U2740 (N_2740,N_2021,N_2484);
and U2741 (N_2741,N_2373,N_2188);
and U2742 (N_2742,N_2221,N_2468);
nor U2743 (N_2743,N_2189,N_2330);
or U2744 (N_2744,N_2278,N_2166);
nand U2745 (N_2745,N_2332,N_2303);
nor U2746 (N_2746,N_2441,N_2097);
nor U2747 (N_2747,N_2158,N_2396);
xnor U2748 (N_2748,N_2389,N_2134);
nor U2749 (N_2749,N_2019,N_1882);
nor U2750 (N_2750,N_2140,N_1880);
or U2751 (N_2751,N_2232,N_1911);
nor U2752 (N_2752,N_2434,N_2025);
or U2753 (N_2753,N_2464,N_2108);
nor U2754 (N_2754,N_2000,N_2206);
nor U2755 (N_2755,N_2284,N_2398);
or U2756 (N_2756,N_2187,N_2349);
nor U2757 (N_2757,N_2162,N_2372);
xnor U2758 (N_2758,N_2164,N_2310);
and U2759 (N_2759,N_2220,N_1892);
or U2760 (N_2760,N_2062,N_2112);
nand U2761 (N_2761,N_2121,N_1909);
or U2762 (N_2762,N_2237,N_2477);
xor U2763 (N_2763,N_2011,N_2401);
xnor U2764 (N_2764,N_2458,N_1929);
xor U2765 (N_2765,N_2374,N_2319);
nand U2766 (N_2766,N_2118,N_2402);
or U2767 (N_2767,N_2287,N_2288);
xor U2768 (N_2768,N_1943,N_2174);
or U2769 (N_2769,N_2305,N_1966);
or U2770 (N_2770,N_2060,N_2481);
nand U2771 (N_2771,N_2364,N_2421);
or U2772 (N_2772,N_1896,N_2435);
and U2773 (N_2773,N_1877,N_2423);
and U2774 (N_2774,N_2348,N_2152);
nor U2775 (N_2775,N_2448,N_2082);
and U2776 (N_2776,N_2105,N_2202);
xor U2777 (N_2777,N_1891,N_1956);
nor U2778 (N_2778,N_1897,N_2076);
and U2779 (N_2779,N_2088,N_2476);
xor U2780 (N_2780,N_2430,N_2439);
nand U2781 (N_2781,N_2351,N_2030);
and U2782 (N_2782,N_2017,N_2122);
xnor U2783 (N_2783,N_2074,N_1876);
nor U2784 (N_2784,N_2245,N_2159);
or U2785 (N_2785,N_1915,N_2115);
nand U2786 (N_2786,N_2397,N_1990);
and U2787 (N_2787,N_2177,N_2355);
nand U2788 (N_2788,N_2126,N_2256);
and U2789 (N_2789,N_2210,N_2454);
or U2790 (N_2790,N_2345,N_2306);
nand U2791 (N_2791,N_1895,N_2362);
nor U2792 (N_2792,N_2443,N_1988);
nor U2793 (N_2793,N_2446,N_2145);
or U2794 (N_2794,N_2180,N_2120);
nor U2795 (N_2795,N_1924,N_2185);
and U2796 (N_2796,N_2050,N_2409);
nand U2797 (N_2797,N_2193,N_2230);
or U2798 (N_2798,N_2354,N_2228);
nand U2799 (N_2799,N_2334,N_1941);
nor U2800 (N_2800,N_2478,N_2492);
nand U2801 (N_2801,N_1920,N_2301);
nor U2802 (N_2802,N_2320,N_2497);
or U2803 (N_2803,N_2136,N_2191);
or U2804 (N_2804,N_1959,N_2179);
nor U2805 (N_2805,N_2279,N_2340);
xnor U2806 (N_2806,N_2238,N_2199);
or U2807 (N_2807,N_2150,N_1969);
or U2808 (N_2808,N_1917,N_2371);
and U2809 (N_2809,N_2452,N_2298);
and U2810 (N_2810,N_2427,N_2223);
nand U2811 (N_2811,N_2277,N_1899);
nand U2812 (N_2812,N_2010,N_2249);
nor U2813 (N_2813,N_2248,N_2440);
nor U2814 (N_2814,N_2436,N_1957);
nor U2815 (N_2815,N_1972,N_2149);
or U2816 (N_2816,N_2364,N_2212);
and U2817 (N_2817,N_2332,N_1899);
nand U2818 (N_2818,N_2481,N_2378);
nor U2819 (N_2819,N_2381,N_2283);
nor U2820 (N_2820,N_2185,N_2149);
nand U2821 (N_2821,N_2260,N_1994);
and U2822 (N_2822,N_2377,N_2154);
nor U2823 (N_2823,N_2460,N_1941);
nand U2824 (N_2824,N_2297,N_2353);
or U2825 (N_2825,N_2152,N_2186);
or U2826 (N_2826,N_2111,N_2320);
and U2827 (N_2827,N_2390,N_2113);
and U2828 (N_2828,N_2467,N_2052);
nand U2829 (N_2829,N_2241,N_2481);
nor U2830 (N_2830,N_1954,N_2370);
and U2831 (N_2831,N_2000,N_1973);
or U2832 (N_2832,N_2038,N_2157);
xor U2833 (N_2833,N_2209,N_2496);
and U2834 (N_2834,N_2018,N_2197);
or U2835 (N_2835,N_1979,N_2122);
nor U2836 (N_2836,N_2037,N_2431);
or U2837 (N_2837,N_2144,N_1916);
nand U2838 (N_2838,N_2076,N_2380);
xnor U2839 (N_2839,N_2415,N_1971);
xor U2840 (N_2840,N_2497,N_2063);
nand U2841 (N_2841,N_2214,N_1933);
nor U2842 (N_2842,N_2263,N_2295);
xor U2843 (N_2843,N_1877,N_1964);
nor U2844 (N_2844,N_2099,N_2489);
nor U2845 (N_2845,N_2025,N_2384);
nor U2846 (N_2846,N_2230,N_2034);
nor U2847 (N_2847,N_2083,N_1884);
nor U2848 (N_2848,N_1901,N_2388);
nor U2849 (N_2849,N_2079,N_2351);
nor U2850 (N_2850,N_1985,N_2361);
nor U2851 (N_2851,N_2119,N_2387);
xor U2852 (N_2852,N_2345,N_2219);
xor U2853 (N_2853,N_2084,N_2367);
nor U2854 (N_2854,N_2335,N_2079);
or U2855 (N_2855,N_2218,N_1888);
nand U2856 (N_2856,N_2143,N_2014);
nand U2857 (N_2857,N_2074,N_2234);
or U2858 (N_2858,N_1896,N_2474);
and U2859 (N_2859,N_2039,N_1955);
xor U2860 (N_2860,N_2326,N_2367);
nor U2861 (N_2861,N_1977,N_2259);
and U2862 (N_2862,N_2327,N_1971);
nor U2863 (N_2863,N_2323,N_1963);
and U2864 (N_2864,N_2491,N_1886);
nor U2865 (N_2865,N_2055,N_2237);
nor U2866 (N_2866,N_1972,N_2029);
nor U2867 (N_2867,N_1989,N_1884);
and U2868 (N_2868,N_1907,N_2220);
or U2869 (N_2869,N_1887,N_2075);
and U2870 (N_2870,N_2045,N_1984);
xor U2871 (N_2871,N_2499,N_2164);
and U2872 (N_2872,N_1880,N_1991);
and U2873 (N_2873,N_2107,N_1983);
or U2874 (N_2874,N_2466,N_2467);
xnor U2875 (N_2875,N_2304,N_2302);
nor U2876 (N_2876,N_1927,N_2338);
nor U2877 (N_2877,N_2172,N_2446);
or U2878 (N_2878,N_2359,N_2059);
and U2879 (N_2879,N_2498,N_2111);
nand U2880 (N_2880,N_1917,N_2313);
and U2881 (N_2881,N_2268,N_2284);
nand U2882 (N_2882,N_2418,N_2438);
nor U2883 (N_2883,N_2422,N_2372);
or U2884 (N_2884,N_2464,N_1955);
xor U2885 (N_2885,N_2444,N_1912);
nor U2886 (N_2886,N_2292,N_2082);
xor U2887 (N_2887,N_2199,N_2119);
or U2888 (N_2888,N_2377,N_2018);
and U2889 (N_2889,N_2124,N_2127);
nand U2890 (N_2890,N_2304,N_2357);
nand U2891 (N_2891,N_1875,N_2036);
nor U2892 (N_2892,N_2434,N_2216);
and U2893 (N_2893,N_2002,N_2031);
xor U2894 (N_2894,N_2482,N_2052);
nand U2895 (N_2895,N_2272,N_1936);
xnor U2896 (N_2896,N_2088,N_2251);
nand U2897 (N_2897,N_2033,N_2477);
nand U2898 (N_2898,N_1875,N_1998);
and U2899 (N_2899,N_2251,N_2265);
and U2900 (N_2900,N_1894,N_2347);
xnor U2901 (N_2901,N_1891,N_2144);
or U2902 (N_2902,N_2008,N_2356);
xor U2903 (N_2903,N_2480,N_2023);
nand U2904 (N_2904,N_1978,N_1900);
or U2905 (N_2905,N_2168,N_2422);
or U2906 (N_2906,N_2303,N_2065);
or U2907 (N_2907,N_2280,N_2304);
or U2908 (N_2908,N_2023,N_2106);
nand U2909 (N_2909,N_2117,N_2424);
nor U2910 (N_2910,N_2026,N_2053);
and U2911 (N_2911,N_2264,N_1895);
xor U2912 (N_2912,N_2189,N_2029);
nor U2913 (N_2913,N_2492,N_2224);
and U2914 (N_2914,N_2124,N_2141);
and U2915 (N_2915,N_1906,N_2007);
and U2916 (N_2916,N_2103,N_2373);
or U2917 (N_2917,N_2110,N_2262);
nand U2918 (N_2918,N_2258,N_1979);
or U2919 (N_2919,N_1960,N_1986);
or U2920 (N_2920,N_2348,N_1894);
or U2921 (N_2921,N_2243,N_2216);
nor U2922 (N_2922,N_2197,N_2067);
xnor U2923 (N_2923,N_1963,N_2364);
xnor U2924 (N_2924,N_2451,N_1941);
and U2925 (N_2925,N_2056,N_2366);
nor U2926 (N_2926,N_2332,N_2218);
and U2927 (N_2927,N_1902,N_2321);
and U2928 (N_2928,N_2092,N_2437);
xor U2929 (N_2929,N_2363,N_2100);
and U2930 (N_2930,N_2176,N_2047);
nor U2931 (N_2931,N_2471,N_2172);
nand U2932 (N_2932,N_1945,N_1973);
or U2933 (N_2933,N_2167,N_2203);
xnor U2934 (N_2934,N_2483,N_2223);
or U2935 (N_2935,N_2468,N_2268);
and U2936 (N_2936,N_1966,N_1929);
xor U2937 (N_2937,N_2403,N_2259);
xnor U2938 (N_2938,N_2448,N_2486);
nor U2939 (N_2939,N_1984,N_2160);
xor U2940 (N_2940,N_2251,N_2178);
nor U2941 (N_2941,N_2415,N_2059);
or U2942 (N_2942,N_2484,N_2260);
xnor U2943 (N_2943,N_2443,N_2260);
xor U2944 (N_2944,N_2117,N_2163);
nand U2945 (N_2945,N_2347,N_1877);
or U2946 (N_2946,N_2441,N_2126);
or U2947 (N_2947,N_2276,N_2336);
or U2948 (N_2948,N_2430,N_2319);
and U2949 (N_2949,N_2137,N_2069);
nor U2950 (N_2950,N_2332,N_1975);
and U2951 (N_2951,N_2191,N_2433);
or U2952 (N_2952,N_2226,N_1929);
nor U2953 (N_2953,N_2179,N_2135);
xnor U2954 (N_2954,N_2465,N_1878);
xnor U2955 (N_2955,N_1987,N_2130);
xor U2956 (N_2956,N_2119,N_2099);
and U2957 (N_2957,N_1942,N_1889);
xnor U2958 (N_2958,N_2142,N_2025);
and U2959 (N_2959,N_2050,N_2084);
or U2960 (N_2960,N_1901,N_2384);
and U2961 (N_2961,N_2149,N_1884);
or U2962 (N_2962,N_1972,N_2380);
nor U2963 (N_2963,N_2329,N_2219);
nand U2964 (N_2964,N_1967,N_2385);
xnor U2965 (N_2965,N_1960,N_1954);
nand U2966 (N_2966,N_1967,N_2425);
nand U2967 (N_2967,N_1928,N_2305);
or U2968 (N_2968,N_2321,N_2246);
nor U2969 (N_2969,N_2392,N_2275);
nor U2970 (N_2970,N_2022,N_1949);
xnor U2971 (N_2971,N_1913,N_1950);
xor U2972 (N_2972,N_2191,N_1943);
or U2973 (N_2973,N_2083,N_2364);
xor U2974 (N_2974,N_1907,N_1968);
nand U2975 (N_2975,N_2195,N_1924);
xnor U2976 (N_2976,N_2216,N_1875);
nor U2977 (N_2977,N_2240,N_2078);
nand U2978 (N_2978,N_2219,N_1895);
nand U2979 (N_2979,N_1907,N_2462);
nand U2980 (N_2980,N_2229,N_2226);
and U2981 (N_2981,N_2150,N_2063);
nand U2982 (N_2982,N_2469,N_1965);
or U2983 (N_2983,N_2477,N_2096);
or U2984 (N_2984,N_2226,N_1907);
or U2985 (N_2985,N_2087,N_2277);
xnor U2986 (N_2986,N_2009,N_2067);
and U2987 (N_2987,N_2276,N_2003);
nand U2988 (N_2988,N_2401,N_1924);
nand U2989 (N_2989,N_2098,N_2090);
or U2990 (N_2990,N_1903,N_2246);
and U2991 (N_2991,N_2094,N_2276);
nor U2992 (N_2992,N_2455,N_2005);
xor U2993 (N_2993,N_2447,N_2478);
xnor U2994 (N_2994,N_2428,N_2320);
or U2995 (N_2995,N_2118,N_2048);
nand U2996 (N_2996,N_2296,N_1935);
and U2997 (N_2997,N_2341,N_2257);
and U2998 (N_2998,N_1974,N_2363);
and U2999 (N_2999,N_2141,N_2389);
or U3000 (N_3000,N_2465,N_2481);
or U3001 (N_3001,N_2210,N_2005);
or U3002 (N_3002,N_2484,N_1965);
or U3003 (N_3003,N_2024,N_2226);
nor U3004 (N_3004,N_1901,N_2182);
and U3005 (N_3005,N_2366,N_1935);
nand U3006 (N_3006,N_2400,N_1899);
nor U3007 (N_3007,N_2159,N_2071);
nor U3008 (N_3008,N_2484,N_2108);
xnor U3009 (N_3009,N_2101,N_2464);
nand U3010 (N_3010,N_1913,N_2216);
nand U3011 (N_3011,N_1915,N_2255);
xnor U3012 (N_3012,N_2094,N_2247);
xnor U3013 (N_3013,N_2018,N_2276);
xor U3014 (N_3014,N_2440,N_2391);
nor U3015 (N_3015,N_1984,N_2371);
and U3016 (N_3016,N_2335,N_1920);
xnor U3017 (N_3017,N_2282,N_2131);
nand U3018 (N_3018,N_2008,N_2112);
xnor U3019 (N_3019,N_2422,N_2165);
and U3020 (N_3020,N_1984,N_2305);
or U3021 (N_3021,N_1955,N_2181);
xor U3022 (N_3022,N_2156,N_2187);
nand U3023 (N_3023,N_2086,N_2372);
nor U3024 (N_3024,N_2274,N_2219);
nor U3025 (N_3025,N_2385,N_2236);
nand U3026 (N_3026,N_2090,N_2264);
nand U3027 (N_3027,N_2170,N_1894);
or U3028 (N_3028,N_1994,N_2121);
and U3029 (N_3029,N_1977,N_2362);
and U3030 (N_3030,N_2476,N_2474);
and U3031 (N_3031,N_1993,N_2322);
and U3032 (N_3032,N_2295,N_2262);
nor U3033 (N_3033,N_2181,N_2231);
nand U3034 (N_3034,N_1930,N_2359);
nand U3035 (N_3035,N_2054,N_2063);
and U3036 (N_3036,N_2300,N_2262);
nor U3037 (N_3037,N_1996,N_2387);
xnor U3038 (N_3038,N_2365,N_1918);
and U3039 (N_3039,N_1878,N_2060);
nor U3040 (N_3040,N_2364,N_2006);
or U3041 (N_3041,N_2352,N_2446);
nor U3042 (N_3042,N_2214,N_2303);
and U3043 (N_3043,N_2437,N_2038);
or U3044 (N_3044,N_2434,N_2421);
nor U3045 (N_3045,N_2358,N_2284);
nand U3046 (N_3046,N_2288,N_1930);
xnor U3047 (N_3047,N_2164,N_1880);
xor U3048 (N_3048,N_1929,N_1883);
or U3049 (N_3049,N_2181,N_2218);
nand U3050 (N_3050,N_2260,N_2143);
xnor U3051 (N_3051,N_2363,N_2153);
or U3052 (N_3052,N_2076,N_2110);
and U3053 (N_3053,N_2268,N_2190);
and U3054 (N_3054,N_2317,N_1994);
or U3055 (N_3055,N_1970,N_2379);
xor U3056 (N_3056,N_1943,N_2213);
nor U3057 (N_3057,N_1994,N_2294);
nor U3058 (N_3058,N_1964,N_2493);
and U3059 (N_3059,N_2047,N_2440);
xnor U3060 (N_3060,N_2173,N_2414);
and U3061 (N_3061,N_2198,N_2123);
nand U3062 (N_3062,N_1959,N_2471);
or U3063 (N_3063,N_2052,N_2474);
nand U3064 (N_3064,N_1982,N_2236);
xnor U3065 (N_3065,N_2307,N_2265);
nand U3066 (N_3066,N_1986,N_2095);
nor U3067 (N_3067,N_2291,N_2477);
xor U3068 (N_3068,N_2361,N_2175);
xor U3069 (N_3069,N_2460,N_2465);
and U3070 (N_3070,N_2437,N_2164);
nand U3071 (N_3071,N_1929,N_2368);
nand U3072 (N_3072,N_2401,N_2232);
and U3073 (N_3073,N_2360,N_1876);
nor U3074 (N_3074,N_2274,N_1904);
nor U3075 (N_3075,N_2237,N_1896);
xor U3076 (N_3076,N_2306,N_2186);
or U3077 (N_3077,N_2057,N_2046);
xnor U3078 (N_3078,N_2131,N_2098);
nor U3079 (N_3079,N_2469,N_2461);
nand U3080 (N_3080,N_2014,N_2151);
or U3081 (N_3081,N_1936,N_2390);
and U3082 (N_3082,N_2177,N_2009);
and U3083 (N_3083,N_2156,N_1904);
xnor U3084 (N_3084,N_2025,N_2462);
nand U3085 (N_3085,N_1922,N_2382);
or U3086 (N_3086,N_1878,N_2386);
and U3087 (N_3087,N_2155,N_2036);
and U3088 (N_3088,N_2198,N_2311);
xor U3089 (N_3089,N_2011,N_2246);
or U3090 (N_3090,N_1974,N_2484);
or U3091 (N_3091,N_1945,N_2459);
nor U3092 (N_3092,N_2338,N_2441);
or U3093 (N_3093,N_2153,N_1905);
nand U3094 (N_3094,N_2371,N_2052);
nand U3095 (N_3095,N_2190,N_2000);
or U3096 (N_3096,N_2199,N_2274);
xor U3097 (N_3097,N_1965,N_1887);
and U3098 (N_3098,N_2032,N_2265);
nand U3099 (N_3099,N_2156,N_2294);
or U3100 (N_3100,N_1978,N_2216);
xor U3101 (N_3101,N_1886,N_2332);
and U3102 (N_3102,N_2263,N_2432);
nor U3103 (N_3103,N_2167,N_1913);
nand U3104 (N_3104,N_2093,N_2270);
and U3105 (N_3105,N_1917,N_2138);
or U3106 (N_3106,N_2167,N_2461);
or U3107 (N_3107,N_2033,N_2331);
nor U3108 (N_3108,N_2071,N_2425);
or U3109 (N_3109,N_2211,N_1894);
nor U3110 (N_3110,N_2346,N_1933);
xor U3111 (N_3111,N_1876,N_1966);
nor U3112 (N_3112,N_2318,N_2464);
nor U3113 (N_3113,N_1950,N_2408);
or U3114 (N_3114,N_1952,N_2015);
xor U3115 (N_3115,N_2312,N_2091);
or U3116 (N_3116,N_2396,N_2464);
or U3117 (N_3117,N_2143,N_2485);
nand U3118 (N_3118,N_2451,N_2103);
nor U3119 (N_3119,N_1999,N_2161);
nor U3120 (N_3120,N_2308,N_2345);
nor U3121 (N_3121,N_2460,N_2033);
xor U3122 (N_3122,N_2106,N_2365);
nand U3123 (N_3123,N_2083,N_2186);
nor U3124 (N_3124,N_2357,N_1981);
or U3125 (N_3125,N_3008,N_2813);
nor U3126 (N_3126,N_2866,N_2693);
and U3127 (N_3127,N_2911,N_2996);
and U3128 (N_3128,N_2987,N_2915);
nor U3129 (N_3129,N_2835,N_2700);
xnor U3130 (N_3130,N_3103,N_2758);
nand U3131 (N_3131,N_2861,N_2778);
xnor U3132 (N_3132,N_2878,N_2559);
nand U3133 (N_3133,N_2775,N_2762);
and U3134 (N_3134,N_2501,N_3023);
or U3135 (N_3135,N_2964,N_2578);
nor U3136 (N_3136,N_3026,N_2672);
or U3137 (N_3137,N_2746,N_2570);
xor U3138 (N_3138,N_2873,N_2849);
and U3139 (N_3139,N_2920,N_2753);
or U3140 (N_3140,N_2895,N_2634);
nor U3141 (N_3141,N_2612,N_2949);
and U3142 (N_3142,N_2818,N_3096);
xnor U3143 (N_3143,N_2887,N_2825);
xnor U3144 (N_3144,N_2973,N_2549);
xor U3145 (N_3145,N_2514,N_2936);
nand U3146 (N_3146,N_2704,N_2780);
xnor U3147 (N_3147,N_2604,N_2609);
or U3148 (N_3148,N_2536,N_2785);
or U3149 (N_3149,N_2796,N_2982);
or U3150 (N_3150,N_3047,N_2793);
nor U3151 (N_3151,N_2523,N_2884);
nor U3152 (N_3152,N_2644,N_2801);
nor U3153 (N_3153,N_2872,N_2591);
nand U3154 (N_3154,N_3118,N_2614);
xor U3155 (N_3155,N_2730,N_2662);
xnor U3156 (N_3156,N_2642,N_2682);
and U3157 (N_3157,N_2544,N_2513);
nor U3158 (N_3158,N_2891,N_2763);
nand U3159 (N_3159,N_2711,N_2510);
nand U3160 (N_3160,N_3073,N_2940);
or U3161 (N_3161,N_2622,N_2565);
and U3162 (N_3162,N_2894,N_2717);
nor U3163 (N_3163,N_2515,N_2984);
or U3164 (N_3164,N_2649,N_2581);
xor U3165 (N_3165,N_2930,N_2550);
nand U3166 (N_3166,N_2990,N_2674);
nor U3167 (N_3167,N_3031,N_2502);
xnor U3168 (N_3168,N_3074,N_2923);
nand U3169 (N_3169,N_2820,N_2542);
and U3170 (N_3170,N_2545,N_3033);
and U3171 (N_3171,N_3038,N_2563);
nor U3172 (N_3172,N_2522,N_2955);
xor U3173 (N_3173,N_3095,N_3042);
nor U3174 (N_3174,N_2684,N_3001);
nor U3175 (N_3175,N_2774,N_2781);
and U3176 (N_3176,N_2899,N_2689);
and U3177 (N_3177,N_2760,N_2532);
nor U3178 (N_3178,N_2766,N_2875);
nor U3179 (N_3179,N_2991,N_3088);
nand U3180 (N_3180,N_2713,N_2521);
and U3181 (N_3181,N_2588,N_2543);
or U3182 (N_3182,N_2924,N_2858);
nor U3183 (N_3183,N_2828,N_3029);
xor U3184 (N_3184,N_2986,N_2770);
xor U3185 (N_3185,N_2592,N_2902);
or U3186 (N_3186,N_2843,N_2837);
or U3187 (N_3187,N_2716,N_3089);
or U3188 (N_3188,N_2666,N_2686);
nand U3189 (N_3189,N_2978,N_3082);
xnor U3190 (N_3190,N_2508,N_2822);
xor U3191 (N_3191,N_2919,N_2962);
nor U3192 (N_3192,N_2896,N_2597);
or U3193 (N_3193,N_2690,N_2506);
nor U3194 (N_3194,N_2747,N_3013);
and U3195 (N_3195,N_2665,N_2657);
and U3196 (N_3196,N_2658,N_2772);
or U3197 (N_3197,N_3065,N_2643);
xnor U3198 (N_3198,N_2699,N_3079);
and U3199 (N_3199,N_3071,N_2957);
and U3200 (N_3200,N_2958,N_2767);
and U3201 (N_3201,N_2553,N_2632);
nor U3202 (N_3202,N_2997,N_2739);
or U3203 (N_3203,N_3107,N_2918);
or U3204 (N_3204,N_2733,N_2925);
xnor U3205 (N_3205,N_3122,N_2668);
and U3206 (N_3206,N_2616,N_2719);
and U3207 (N_3207,N_2939,N_3045);
xnor U3208 (N_3208,N_3116,N_3025);
or U3209 (N_3209,N_2909,N_2963);
nand U3210 (N_3210,N_2571,N_2976);
nand U3211 (N_3211,N_2580,N_2710);
and U3212 (N_3212,N_3120,N_2970);
nor U3213 (N_3213,N_3087,N_3044);
and U3214 (N_3214,N_3027,N_2630);
nor U3215 (N_3215,N_3022,N_2562);
or U3216 (N_3216,N_2722,N_2914);
or U3217 (N_3217,N_2901,N_2737);
and U3218 (N_3218,N_2855,N_2783);
and U3219 (N_3219,N_3017,N_2846);
and U3220 (N_3220,N_3014,N_3059);
nor U3221 (N_3221,N_2922,N_2735);
nor U3222 (N_3222,N_3024,N_2708);
and U3223 (N_3223,N_3068,N_2596);
nand U3224 (N_3224,N_2535,N_2589);
xor U3225 (N_3225,N_3086,N_2933);
nand U3226 (N_3226,N_2777,N_2965);
xnor U3227 (N_3227,N_2981,N_2720);
xor U3228 (N_3228,N_2511,N_2627);
nor U3229 (N_3229,N_2824,N_2790);
xnor U3230 (N_3230,N_2905,N_3021);
nand U3231 (N_3231,N_2754,N_2947);
xor U3232 (N_3232,N_2800,N_2631);
or U3233 (N_3233,N_2787,N_2723);
and U3234 (N_3234,N_2811,N_2756);
xnor U3235 (N_3235,N_2829,N_2539);
and U3236 (N_3236,N_2845,N_2966);
and U3237 (N_3237,N_2857,N_2847);
or U3238 (N_3238,N_3077,N_2583);
and U3239 (N_3239,N_2650,N_3046);
or U3240 (N_3240,N_2879,N_2712);
or U3241 (N_3241,N_3063,N_2529);
and U3242 (N_3242,N_2664,N_2572);
or U3243 (N_3243,N_2505,N_2653);
xnor U3244 (N_3244,N_2607,N_2641);
or U3245 (N_3245,N_2838,N_2624);
nor U3246 (N_3246,N_2740,N_2590);
nand U3247 (N_3247,N_2679,N_2751);
or U3248 (N_3248,N_2500,N_2728);
or U3249 (N_3249,N_2725,N_2874);
or U3250 (N_3250,N_3050,N_2692);
and U3251 (N_3251,N_2937,N_3111);
nor U3252 (N_3252,N_2629,N_3006);
nand U3253 (N_3253,N_2890,N_2582);
nand U3254 (N_3254,N_2912,N_2640);
nor U3255 (N_3255,N_2533,N_2577);
and U3256 (N_3256,N_2906,N_2794);
nand U3257 (N_3257,N_2921,N_2576);
xor U3258 (N_3258,N_2574,N_2842);
nor U3259 (N_3259,N_3119,N_2695);
nand U3260 (N_3260,N_2537,N_2615);
nand U3261 (N_3261,N_2669,N_2795);
xor U3262 (N_3262,N_2637,N_2897);
nand U3263 (N_3263,N_2769,N_3012);
xor U3264 (N_3264,N_3099,N_3002);
xnor U3265 (N_3265,N_2859,N_2967);
nor U3266 (N_3266,N_2706,N_2531);
or U3267 (N_3267,N_3035,N_2876);
and U3268 (N_3268,N_2786,N_2864);
and U3269 (N_3269,N_2619,N_2675);
and U3270 (N_3270,N_2618,N_2677);
xnor U3271 (N_3271,N_3080,N_2603);
and U3272 (N_3272,N_2517,N_3067);
xor U3273 (N_3273,N_2673,N_2871);
nor U3274 (N_3274,N_2600,N_2881);
nor U3275 (N_3275,N_3060,N_3019);
or U3276 (N_3276,N_3034,N_2865);
nand U3277 (N_3277,N_2752,N_2839);
or U3278 (N_3278,N_2598,N_2900);
and U3279 (N_3279,N_2636,N_2652);
nand U3280 (N_3280,N_2848,N_3062);
xnor U3281 (N_3281,N_2678,N_3090);
xor U3282 (N_3282,N_2687,N_2748);
nor U3283 (N_3283,N_2782,N_3100);
nand U3284 (N_3284,N_2681,N_3084);
or U3285 (N_3285,N_3115,N_3083);
nor U3286 (N_3286,N_2701,N_2821);
and U3287 (N_3287,N_2744,N_2798);
or U3288 (N_3288,N_2860,N_3085);
or U3289 (N_3289,N_2908,N_2663);
nand U3290 (N_3290,N_2883,N_2819);
nor U3291 (N_3291,N_2509,N_2646);
xor U3292 (N_3292,N_2983,N_2836);
or U3293 (N_3293,N_2812,N_2602);
xor U3294 (N_3294,N_2575,N_3092);
or U3295 (N_3295,N_2558,N_2703);
or U3296 (N_3296,N_2810,N_2952);
or U3297 (N_3297,N_2755,N_2888);
nor U3298 (N_3298,N_2799,N_2610);
or U3299 (N_3299,N_2994,N_2776);
and U3300 (N_3300,N_2613,N_2867);
and U3301 (N_3301,N_2546,N_3010);
and U3302 (N_3302,N_2525,N_2750);
and U3303 (N_3303,N_2738,N_2954);
nor U3304 (N_3304,N_2512,N_2948);
xor U3305 (N_3305,N_2826,N_2992);
xor U3306 (N_3306,N_2568,N_2547);
or U3307 (N_3307,N_2691,N_3066);
nand U3308 (N_3308,N_3104,N_2953);
nor U3309 (N_3309,N_2726,N_2606);
nand U3310 (N_3310,N_2654,N_2893);
xnor U3311 (N_3311,N_2683,N_2540);
nand U3312 (N_3312,N_2870,N_2913);
nand U3313 (N_3313,N_2697,N_2817);
nor U3314 (N_3314,N_3009,N_3007);
nand U3315 (N_3315,N_2862,N_3097);
or U3316 (N_3316,N_2941,N_2734);
and U3317 (N_3317,N_2945,N_3061);
nor U3318 (N_3318,N_2761,N_2671);
nor U3319 (N_3319,N_2551,N_2975);
and U3320 (N_3320,N_2932,N_3056);
nand U3321 (N_3321,N_2528,N_3109);
xnor U3322 (N_3322,N_2840,N_2584);
nand U3323 (N_3323,N_2989,N_2985);
and U3324 (N_3324,N_2823,N_3000);
nand U3325 (N_3325,N_2882,N_2651);
and U3326 (N_3326,N_3037,N_3028);
nor U3327 (N_3327,N_2971,N_2759);
xor U3328 (N_3328,N_2742,N_3030);
xnor U3329 (N_3329,N_2705,N_3057);
nand U3330 (N_3330,N_3094,N_2709);
xor U3331 (N_3331,N_3055,N_2764);
or U3332 (N_3332,N_2816,N_2916);
and U3333 (N_3333,N_2998,N_3011);
and U3334 (N_3334,N_2714,N_2898);
and U3335 (N_3335,N_3039,N_2765);
nor U3336 (N_3336,N_2979,N_2757);
or U3337 (N_3337,N_2907,N_3121);
xor U3338 (N_3338,N_3098,N_2928);
xor U3339 (N_3339,N_3018,N_3106);
and U3340 (N_3340,N_3015,N_2809);
nor U3341 (N_3341,N_2980,N_2931);
xnor U3342 (N_3342,N_2595,N_2586);
xnor U3343 (N_3343,N_2830,N_2696);
nand U3344 (N_3344,N_2852,N_3043);
nor U3345 (N_3345,N_3003,N_2827);
or U3346 (N_3346,N_2885,N_3072);
and U3347 (N_3347,N_2605,N_3076);
xor U3348 (N_3348,N_2768,N_3108);
and U3349 (N_3349,N_2633,N_2561);
and U3350 (N_3350,N_3114,N_2639);
and U3351 (N_3351,N_2803,N_2972);
nor U3352 (N_3352,N_2516,N_3064);
or U3353 (N_3353,N_2974,N_2685);
nor U3354 (N_3354,N_2617,N_2667);
nor U3355 (N_3355,N_2593,N_3049);
and U3356 (N_3356,N_2504,N_2969);
nand U3357 (N_3357,N_2648,N_2993);
and U3358 (N_3358,N_2655,N_2670);
xor U3359 (N_3359,N_3048,N_2623);
or U3360 (N_3360,N_2611,N_2968);
or U3361 (N_3361,N_2797,N_2779);
and U3362 (N_3362,N_2608,N_2688);
and U3363 (N_3363,N_3020,N_2961);
xor U3364 (N_3364,N_2854,N_2833);
nand U3365 (N_3365,N_3070,N_2541);
or U3366 (N_3366,N_3005,N_2599);
nor U3367 (N_3367,N_2851,N_2934);
nor U3368 (N_3368,N_2555,N_2579);
nand U3369 (N_3369,N_2557,N_2844);
and U3370 (N_3370,N_2715,N_2721);
and U3371 (N_3371,N_3124,N_2527);
nand U3372 (N_3372,N_2694,N_2656);
or U3373 (N_3373,N_2564,N_2877);
nand U3374 (N_3374,N_3054,N_2950);
or U3375 (N_3375,N_2951,N_2707);
or U3376 (N_3376,N_2841,N_2802);
nor U3377 (N_3377,N_2524,N_2960);
xnor U3378 (N_3378,N_3016,N_2729);
nor U3379 (N_3379,N_2727,N_2832);
xnor U3380 (N_3380,N_3036,N_2938);
or U3381 (N_3381,N_2647,N_3040);
xor U3382 (N_3382,N_2910,N_2749);
nand U3383 (N_3383,N_2732,N_2661);
and U3384 (N_3384,N_2724,N_2792);
nor U3385 (N_3385,N_2534,N_2520);
nand U3386 (N_3386,N_2638,N_2999);
or U3387 (N_3387,N_2834,N_2791);
or U3388 (N_3388,N_2680,N_2645);
xnor U3389 (N_3389,N_2601,N_2736);
nand U3390 (N_3390,N_2853,N_3110);
and U3391 (N_3391,N_2587,N_2831);
xor U3392 (N_3392,N_2929,N_2518);
nand U3393 (N_3393,N_2625,N_2569);
or U3394 (N_3394,N_2944,N_2917);
xor U3395 (N_3395,N_2869,N_2526);
nand U3396 (N_3396,N_3058,N_3051);
nand U3397 (N_3397,N_2702,N_2942);
xor U3398 (N_3398,N_2868,N_2771);
nand U3399 (N_3399,N_2507,N_2519);
xnor U3400 (N_3400,N_3052,N_3102);
xnor U3401 (N_3401,N_2556,N_3032);
xnor U3402 (N_3402,N_2635,N_2659);
or U3403 (N_3403,N_2856,N_2538);
and U3404 (N_3404,N_2698,N_3053);
xnor U3405 (N_3405,N_2808,N_2886);
or U3406 (N_3406,N_3078,N_3075);
xnor U3407 (N_3407,N_2773,N_3117);
nand U3408 (N_3408,N_2904,N_2731);
nor U3409 (N_3409,N_2863,N_2594);
nor U3410 (N_3410,N_2628,N_3101);
xnor U3411 (N_3411,N_2573,N_2892);
nand U3412 (N_3412,N_2745,N_2880);
nand U3413 (N_3413,N_3093,N_2943);
xor U3414 (N_3414,N_2946,N_2805);
nor U3415 (N_3415,N_2560,N_2585);
or U3416 (N_3416,N_2660,N_2784);
nor U3417 (N_3417,N_2621,N_2959);
nand U3418 (N_3418,N_2789,N_2788);
xnor U3419 (N_3419,N_2804,N_2554);
or U3420 (N_3420,N_2815,N_2889);
and U3421 (N_3421,N_2620,N_2567);
or U3422 (N_3422,N_3091,N_2977);
nor U3423 (N_3423,N_2806,N_3113);
nor U3424 (N_3424,N_2741,N_2988);
nand U3425 (N_3425,N_2743,N_3105);
nand U3426 (N_3426,N_2676,N_2807);
or U3427 (N_3427,N_3081,N_2626);
nand U3428 (N_3428,N_2995,N_3069);
nor U3429 (N_3429,N_3123,N_3004);
xor U3430 (N_3430,N_2566,N_2530);
xor U3431 (N_3431,N_2552,N_2850);
xor U3432 (N_3432,N_2503,N_2956);
or U3433 (N_3433,N_2935,N_2927);
xor U3434 (N_3434,N_2814,N_2926);
or U3435 (N_3435,N_2548,N_3041);
nand U3436 (N_3436,N_3112,N_2718);
nor U3437 (N_3437,N_2903,N_3121);
nor U3438 (N_3438,N_3101,N_2511);
nand U3439 (N_3439,N_2939,N_2693);
nand U3440 (N_3440,N_2810,N_2914);
nand U3441 (N_3441,N_3082,N_2717);
nand U3442 (N_3442,N_2964,N_2851);
nand U3443 (N_3443,N_2886,N_2814);
or U3444 (N_3444,N_2642,N_2552);
xnor U3445 (N_3445,N_2953,N_2745);
xor U3446 (N_3446,N_2915,N_2686);
xnor U3447 (N_3447,N_3124,N_2646);
or U3448 (N_3448,N_3090,N_2910);
nor U3449 (N_3449,N_2871,N_2985);
nor U3450 (N_3450,N_2756,N_2766);
and U3451 (N_3451,N_2742,N_2653);
nand U3452 (N_3452,N_2875,N_2835);
xnor U3453 (N_3453,N_2788,N_3076);
nand U3454 (N_3454,N_2722,N_2567);
and U3455 (N_3455,N_2841,N_2873);
xnor U3456 (N_3456,N_2517,N_2947);
nand U3457 (N_3457,N_3088,N_2902);
xnor U3458 (N_3458,N_3000,N_2955);
xnor U3459 (N_3459,N_2771,N_2967);
nor U3460 (N_3460,N_3114,N_2749);
nand U3461 (N_3461,N_2828,N_2688);
xnor U3462 (N_3462,N_2563,N_2716);
nand U3463 (N_3463,N_2568,N_2944);
xor U3464 (N_3464,N_3115,N_2778);
nand U3465 (N_3465,N_2958,N_2607);
and U3466 (N_3466,N_2729,N_2580);
or U3467 (N_3467,N_2621,N_3087);
and U3468 (N_3468,N_2925,N_2940);
or U3469 (N_3469,N_2815,N_2979);
nand U3470 (N_3470,N_2828,N_2563);
or U3471 (N_3471,N_3056,N_2567);
nor U3472 (N_3472,N_3044,N_2579);
nor U3473 (N_3473,N_2520,N_2704);
and U3474 (N_3474,N_2720,N_3022);
and U3475 (N_3475,N_2679,N_2814);
nor U3476 (N_3476,N_3060,N_2781);
xor U3477 (N_3477,N_2943,N_2961);
xnor U3478 (N_3478,N_2781,N_3009);
and U3479 (N_3479,N_2702,N_3082);
or U3480 (N_3480,N_2623,N_2645);
nor U3481 (N_3481,N_2520,N_2815);
nor U3482 (N_3482,N_2878,N_2920);
nand U3483 (N_3483,N_2515,N_3105);
nor U3484 (N_3484,N_2693,N_2653);
or U3485 (N_3485,N_2539,N_2699);
xnor U3486 (N_3486,N_2777,N_3011);
nand U3487 (N_3487,N_3007,N_2722);
xor U3488 (N_3488,N_2791,N_2732);
or U3489 (N_3489,N_2868,N_2653);
xnor U3490 (N_3490,N_2919,N_2806);
nor U3491 (N_3491,N_2527,N_2629);
nand U3492 (N_3492,N_2652,N_2700);
or U3493 (N_3493,N_3026,N_2729);
nor U3494 (N_3494,N_2735,N_2979);
xor U3495 (N_3495,N_2561,N_2803);
nor U3496 (N_3496,N_2632,N_3008);
or U3497 (N_3497,N_3073,N_2592);
or U3498 (N_3498,N_2786,N_2886);
nand U3499 (N_3499,N_2951,N_2831);
and U3500 (N_3500,N_3039,N_2547);
xor U3501 (N_3501,N_2510,N_2592);
nor U3502 (N_3502,N_2846,N_2985);
nor U3503 (N_3503,N_3043,N_2681);
nor U3504 (N_3504,N_3077,N_2984);
nand U3505 (N_3505,N_2673,N_2608);
nand U3506 (N_3506,N_2913,N_2533);
and U3507 (N_3507,N_2517,N_2869);
or U3508 (N_3508,N_3022,N_2958);
nor U3509 (N_3509,N_3074,N_2676);
or U3510 (N_3510,N_2732,N_2774);
nand U3511 (N_3511,N_3010,N_2846);
nand U3512 (N_3512,N_2848,N_2828);
or U3513 (N_3513,N_2708,N_2613);
nand U3514 (N_3514,N_2684,N_2833);
and U3515 (N_3515,N_2511,N_2562);
xnor U3516 (N_3516,N_3000,N_2918);
or U3517 (N_3517,N_2798,N_3061);
or U3518 (N_3518,N_2937,N_2682);
or U3519 (N_3519,N_3028,N_2687);
xor U3520 (N_3520,N_3052,N_2956);
and U3521 (N_3521,N_2768,N_2930);
or U3522 (N_3522,N_3041,N_3023);
xor U3523 (N_3523,N_2593,N_2622);
and U3524 (N_3524,N_2970,N_2529);
or U3525 (N_3525,N_3046,N_2557);
and U3526 (N_3526,N_2674,N_2963);
nand U3527 (N_3527,N_2912,N_2750);
or U3528 (N_3528,N_2864,N_3075);
or U3529 (N_3529,N_3093,N_2899);
nand U3530 (N_3530,N_2658,N_2515);
xnor U3531 (N_3531,N_2767,N_2532);
nand U3532 (N_3532,N_2624,N_3059);
nor U3533 (N_3533,N_2941,N_2628);
nor U3534 (N_3534,N_2995,N_2966);
nand U3535 (N_3535,N_2584,N_2651);
or U3536 (N_3536,N_2695,N_2749);
nor U3537 (N_3537,N_3024,N_2665);
or U3538 (N_3538,N_2562,N_3077);
nand U3539 (N_3539,N_2509,N_2784);
xnor U3540 (N_3540,N_2962,N_2646);
or U3541 (N_3541,N_2723,N_2815);
and U3542 (N_3542,N_2776,N_3038);
nand U3543 (N_3543,N_2812,N_2989);
xor U3544 (N_3544,N_2538,N_2821);
and U3545 (N_3545,N_2607,N_2952);
or U3546 (N_3546,N_2589,N_3098);
nor U3547 (N_3547,N_2791,N_2895);
nor U3548 (N_3548,N_2809,N_2776);
nor U3549 (N_3549,N_2531,N_3016);
or U3550 (N_3550,N_3074,N_2634);
and U3551 (N_3551,N_2920,N_2667);
and U3552 (N_3552,N_3025,N_3088);
xor U3553 (N_3553,N_2931,N_3085);
or U3554 (N_3554,N_2913,N_2801);
or U3555 (N_3555,N_3027,N_2515);
and U3556 (N_3556,N_3062,N_2566);
nand U3557 (N_3557,N_2782,N_3102);
nand U3558 (N_3558,N_3005,N_3060);
xnor U3559 (N_3559,N_2729,N_2650);
or U3560 (N_3560,N_3055,N_2687);
xnor U3561 (N_3561,N_3123,N_2626);
xor U3562 (N_3562,N_2645,N_2669);
nor U3563 (N_3563,N_2595,N_2804);
and U3564 (N_3564,N_2667,N_3095);
nor U3565 (N_3565,N_2875,N_2665);
nor U3566 (N_3566,N_2620,N_2529);
nand U3567 (N_3567,N_2955,N_3011);
and U3568 (N_3568,N_2997,N_2735);
xor U3569 (N_3569,N_2599,N_2987);
xnor U3570 (N_3570,N_2746,N_2814);
nor U3571 (N_3571,N_2864,N_2551);
nand U3572 (N_3572,N_2764,N_2707);
and U3573 (N_3573,N_2810,N_2530);
nor U3574 (N_3574,N_2505,N_2880);
xnor U3575 (N_3575,N_3012,N_2811);
nand U3576 (N_3576,N_2788,N_2828);
or U3577 (N_3577,N_2653,N_2752);
and U3578 (N_3578,N_2761,N_2623);
or U3579 (N_3579,N_2764,N_2978);
or U3580 (N_3580,N_2530,N_2506);
nand U3581 (N_3581,N_2913,N_2531);
nand U3582 (N_3582,N_2680,N_2543);
xor U3583 (N_3583,N_3039,N_3017);
xor U3584 (N_3584,N_2572,N_2772);
xnor U3585 (N_3585,N_3057,N_3103);
nor U3586 (N_3586,N_2744,N_3012);
xnor U3587 (N_3587,N_2960,N_2865);
xnor U3588 (N_3588,N_2542,N_3050);
or U3589 (N_3589,N_3022,N_3060);
xnor U3590 (N_3590,N_2650,N_2835);
nor U3591 (N_3591,N_2846,N_3077);
and U3592 (N_3592,N_2852,N_3096);
nor U3593 (N_3593,N_2787,N_3078);
nor U3594 (N_3594,N_2510,N_3003);
and U3595 (N_3595,N_2704,N_2713);
nor U3596 (N_3596,N_3006,N_2769);
or U3597 (N_3597,N_2960,N_2702);
nand U3598 (N_3598,N_2724,N_2785);
nor U3599 (N_3599,N_2951,N_2614);
and U3600 (N_3600,N_2640,N_2989);
xnor U3601 (N_3601,N_3049,N_2534);
nand U3602 (N_3602,N_3040,N_2922);
nor U3603 (N_3603,N_2641,N_2847);
and U3604 (N_3604,N_2604,N_2818);
nor U3605 (N_3605,N_3080,N_3118);
and U3606 (N_3606,N_2543,N_2710);
and U3607 (N_3607,N_2638,N_3039);
xor U3608 (N_3608,N_2866,N_2767);
xor U3609 (N_3609,N_3110,N_2713);
or U3610 (N_3610,N_2524,N_2523);
xnor U3611 (N_3611,N_2515,N_2861);
nand U3612 (N_3612,N_2729,N_2795);
and U3613 (N_3613,N_2765,N_2883);
and U3614 (N_3614,N_2640,N_2581);
xnor U3615 (N_3615,N_2689,N_2891);
or U3616 (N_3616,N_2636,N_3047);
and U3617 (N_3617,N_2870,N_2988);
or U3618 (N_3618,N_2963,N_2897);
nor U3619 (N_3619,N_3065,N_2762);
xor U3620 (N_3620,N_2645,N_2527);
or U3621 (N_3621,N_3068,N_3027);
or U3622 (N_3622,N_2539,N_2684);
nor U3623 (N_3623,N_3094,N_3068);
nor U3624 (N_3624,N_2723,N_2585);
or U3625 (N_3625,N_2723,N_2863);
and U3626 (N_3626,N_2929,N_3083);
or U3627 (N_3627,N_3076,N_2701);
or U3628 (N_3628,N_2807,N_2967);
or U3629 (N_3629,N_2911,N_3009);
or U3630 (N_3630,N_2953,N_3096);
nor U3631 (N_3631,N_2828,N_2886);
xnor U3632 (N_3632,N_2980,N_2903);
nand U3633 (N_3633,N_2606,N_2513);
and U3634 (N_3634,N_2792,N_2636);
and U3635 (N_3635,N_2680,N_2676);
nor U3636 (N_3636,N_3055,N_2932);
nor U3637 (N_3637,N_2748,N_2984);
nand U3638 (N_3638,N_2672,N_2870);
xnor U3639 (N_3639,N_2549,N_2738);
nand U3640 (N_3640,N_3009,N_2584);
or U3641 (N_3641,N_2901,N_3010);
or U3642 (N_3642,N_2653,N_2667);
nand U3643 (N_3643,N_2680,N_2714);
nand U3644 (N_3644,N_3000,N_2596);
nor U3645 (N_3645,N_2698,N_2736);
or U3646 (N_3646,N_2776,N_2945);
or U3647 (N_3647,N_2826,N_2810);
nor U3648 (N_3648,N_2842,N_2889);
nand U3649 (N_3649,N_2701,N_3120);
or U3650 (N_3650,N_2659,N_2535);
or U3651 (N_3651,N_2904,N_3104);
nor U3652 (N_3652,N_2911,N_2836);
and U3653 (N_3653,N_2599,N_3123);
and U3654 (N_3654,N_3009,N_2804);
and U3655 (N_3655,N_2638,N_2665);
or U3656 (N_3656,N_2565,N_3015);
nand U3657 (N_3657,N_3046,N_3074);
and U3658 (N_3658,N_2984,N_2969);
or U3659 (N_3659,N_2966,N_3061);
or U3660 (N_3660,N_2952,N_2977);
or U3661 (N_3661,N_2964,N_3121);
nor U3662 (N_3662,N_2947,N_2680);
and U3663 (N_3663,N_2777,N_2891);
xor U3664 (N_3664,N_2856,N_2630);
xnor U3665 (N_3665,N_2726,N_2655);
nor U3666 (N_3666,N_2877,N_2646);
nand U3667 (N_3667,N_2723,N_2891);
xor U3668 (N_3668,N_2966,N_3066);
xor U3669 (N_3669,N_2773,N_3064);
or U3670 (N_3670,N_2554,N_3105);
and U3671 (N_3671,N_2667,N_3056);
xor U3672 (N_3672,N_2624,N_2586);
nor U3673 (N_3673,N_2748,N_2857);
or U3674 (N_3674,N_2964,N_2523);
xnor U3675 (N_3675,N_3034,N_2985);
or U3676 (N_3676,N_2766,N_2759);
and U3677 (N_3677,N_2527,N_3057);
nor U3678 (N_3678,N_2915,N_2803);
nor U3679 (N_3679,N_2805,N_2581);
nand U3680 (N_3680,N_2915,N_3107);
or U3681 (N_3681,N_2613,N_2746);
nor U3682 (N_3682,N_2660,N_2876);
and U3683 (N_3683,N_2993,N_3042);
xor U3684 (N_3684,N_2838,N_2587);
or U3685 (N_3685,N_3061,N_2634);
nand U3686 (N_3686,N_2561,N_3105);
nor U3687 (N_3687,N_2556,N_2811);
and U3688 (N_3688,N_2965,N_2661);
xor U3689 (N_3689,N_2626,N_3031);
and U3690 (N_3690,N_2965,N_2794);
or U3691 (N_3691,N_2973,N_2963);
nand U3692 (N_3692,N_2568,N_2610);
nor U3693 (N_3693,N_2906,N_2812);
or U3694 (N_3694,N_3110,N_2981);
nand U3695 (N_3695,N_3104,N_2518);
or U3696 (N_3696,N_2567,N_2856);
nand U3697 (N_3697,N_2631,N_3093);
nand U3698 (N_3698,N_3058,N_2718);
and U3699 (N_3699,N_2546,N_2997);
xnor U3700 (N_3700,N_2736,N_3006);
xnor U3701 (N_3701,N_2947,N_3018);
and U3702 (N_3702,N_2757,N_3113);
nor U3703 (N_3703,N_2824,N_2743);
or U3704 (N_3704,N_2647,N_2573);
and U3705 (N_3705,N_3045,N_2507);
or U3706 (N_3706,N_3099,N_2979);
xor U3707 (N_3707,N_2617,N_2690);
xor U3708 (N_3708,N_3057,N_2844);
nor U3709 (N_3709,N_2578,N_2650);
nor U3710 (N_3710,N_2643,N_2988);
nand U3711 (N_3711,N_2546,N_2714);
or U3712 (N_3712,N_2833,N_2648);
and U3713 (N_3713,N_2981,N_2558);
nor U3714 (N_3714,N_2886,N_3007);
xor U3715 (N_3715,N_3035,N_2804);
xnor U3716 (N_3716,N_2809,N_2924);
and U3717 (N_3717,N_3100,N_3109);
nand U3718 (N_3718,N_3026,N_2643);
and U3719 (N_3719,N_2947,N_2808);
nor U3720 (N_3720,N_3107,N_2932);
nand U3721 (N_3721,N_2994,N_2595);
nor U3722 (N_3722,N_2517,N_2591);
or U3723 (N_3723,N_2521,N_2689);
and U3724 (N_3724,N_2859,N_2727);
nor U3725 (N_3725,N_2567,N_3087);
xnor U3726 (N_3726,N_2773,N_2747);
nand U3727 (N_3727,N_2650,N_3019);
or U3728 (N_3728,N_2602,N_2962);
xnor U3729 (N_3729,N_2596,N_3055);
xor U3730 (N_3730,N_3032,N_2683);
nor U3731 (N_3731,N_2585,N_2701);
nand U3732 (N_3732,N_2552,N_2525);
xnor U3733 (N_3733,N_2815,N_3061);
or U3734 (N_3734,N_2997,N_3074);
or U3735 (N_3735,N_2642,N_2678);
xor U3736 (N_3736,N_2662,N_2689);
nand U3737 (N_3737,N_2864,N_2720);
or U3738 (N_3738,N_2523,N_2864);
nand U3739 (N_3739,N_2586,N_3082);
or U3740 (N_3740,N_2947,N_2523);
and U3741 (N_3741,N_2537,N_2642);
nor U3742 (N_3742,N_2946,N_2830);
and U3743 (N_3743,N_2628,N_2543);
xnor U3744 (N_3744,N_2862,N_2506);
xnor U3745 (N_3745,N_2956,N_3082);
nand U3746 (N_3746,N_3101,N_3115);
nand U3747 (N_3747,N_2779,N_2954);
xor U3748 (N_3748,N_3017,N_3069);
nor U3749 (N_3749,N_2665,N_3055);
and U3750 (N_3750,N_3195,N_3355);
nand U3751 (N_3751,N_3424,N_3741);
xor U3752 (N_3752,N_3343,N_3464);
and U3753 (N_3753,N_3554,N_3188);
xor U3754 (N_3754,N_3176,N_3206);
and U3755 (N_3755,N_3604,N_3369);
nand U3756 (N_3756,N_3420,N_3517);
nor U3757 (N_3757,N_3238,N_3278);
nor U3758 (N_3758,N_3256,N_3286);
nand U3759 (N_3759,N_3461,N_3160);
and U3760 (N_3760,N_3483,N_3588);
xnor U3761 (N_3761,N_3512,N_3585);
nand U3762 (N_3762,N_3395,N_3387);
nand U3763 (N_3763,N_3510,N_3540);
or U3764 (N_3764,N_3684,N_3217);
and U3765 (N_3765,N_3391,N_3144);
xnor U3766 (N_3766,N_3600,N_3565);
nor U3767 (N_3767,N_3330,N_3676);
nor U3768 (N_3768,N_3629,N_3710);
or U3769 (N_3769,N_3735,N_3323);
or U3770 (N_3770,N_3563,N_3313);
nand U3771 (N_3771,N_3419,N_3739);
nor U3772 (N_3772,N_3263,N_3360);
and U3773 (N_3773,N_3380,N_3454);
nor U3774 (N_3774,N_3520,N_3605);
nor U3775 (N_3775,N_3322,N_3375);
nor U3776 (N_3776,N_3253,N_3610);
and U3777 (N_3777,N_3165,N_3426);
nor U3778 (N_3778,N_3132,N_3708);
nor U3779 (N_3779,N_3423,N_3244);
or U3780 (N_3780,N_3177,N_3243);
and U3781 (N_3781,N_3315,N_3574);
xor U3782 (N_3782,N_3357,N_3533);
nand U3783 (N_3783,N_3560,N_3449);
xnor U3784 (N_3784,N_3163,N_3185);
xnor U3785 (N_3785,N_3445,N_3466);
nand U3786 (N_3786,N_3523,N_3573);
xor U3787 (N_3787,N_3431,N_3478);
nand U3788 (N_3788,N_3641,N_3630);
xor U3789 (N_3789,N_3631,N_3361);
nor U3790 (N_3790,N_3499,N_3374);
nand U3791 (N_3791,N_3175,N_3743);
or U3792 (N_3792,N_3183,N_3309);
nand U3793 (N_3793,N_3715,N_3696);
xnor U3794 (N_3794,N_3521,N_3224);
nand U3795 (N_3795,N_3704,N_3548);
nand U3796 (N_3796,N_3151,N_3511);
nor U3797 (N_3797,N_3261,N_3486);
and U3798 (N_3798,N_3404,N_3685);
or U3799 (N_3799,N_3532,N_3683);
xor U3800 (N_3800,N_3658,N_3161);
or U3801 (N_3801,N_3410,N_3157);
or U3802 (N_3802,N_3535,N_3194);
or U3803 (N_3803,N_3666,N_3179);
xor U3804 (N_3804,N_3576,N_3158);
or U3805 (N_3805,N_3166,N_3267);
xnor U3806 (N_3806,N_3236,N_3377);
nor U3807 (N_3807,N_3342,N_3593);
xnor U3808 (N_3808,N_3366,N_3616);
and U3809 (N_3809,N_3341,N_3640);
and U3810 (N_3810,N_3694,N_3582);
nand U3811 (N_3811,N_3612,N_3692);
or U3812 (N_3812,N_3703,N_3442);
and U3813 (N_3813,N_3524,N_3452);
xor U3814 (N_3814,N_3264,N_3314);
nand U3815 (N_3815,N_3501,N_3526);
xnor U3816 (N_3816,N_3584,N_3212);
or U3817 (N_3817,N_3558,N_3348);
and U3818 (N_3818,N_3417,N_3411);
xnor U3819 (N_3819,N_3288,N_3407);
xor U3820 (N_3820,N_3648,N_3205);
nor U3821 (N_3821,N_3496,N_3713);
xnor U3822 (N_3822,N_3537,N_3399);
nor U3823 (N_3823,N_3642,N_3714);
nor U3824 (N_3824,N_3650,N_3497);
xnor U3825 (N_3825,N_3571,N_3699);
or U3826 (N_3826,N_3325,N_3637);
nor U3827 (N_3827,N_3663,N_3706);
or U3828 (N_3828,N_3262,N_3187);
xor U3829 (N_3829,N_3198,N_3277);
nor U3830 (N_3830,N_3339,N_3254);
or U3831 (N_3831,N_3638,N_3659);
or U3832 (N_3832,N_3636,N_3562);
or U3833 (N_3833,N_3207,N_3436);
nor U3834 (N_3834,N_3229,N_3724);
nor U3835 (N_3835,N_3733,N_3354);
or U3836 (N_3836,N_3586,N_3297);
and U3837 (N_3837,N_3285,N_3200);
nand U3838 (N_3838,N_3283,N_3709);
xnor U3839 (N_3839,N_3304,N_3271);
or U3840 (N_3840,N_3432,N_3580);
xor U3841 (N_3841,N_3422,N_3249);
xor U3842 (N_3842,N_3591,N_3418);
nor U3843 (N_3843,N_3317,N_3305);
and U3844 (N_3844,N_3279,N_3326);
and U3845 (N_3845,N_3492,N_3430);
xor U3846 (N_3846,N_3602,N_3572);
xnor U3847 (N_3847,N_3139,N_3196);
xor U3848 (N_3848,N_3172,N_3547);
and U3849 (N_3849,N_3351,N_3202);
xor U3850 (N_3850,N_3655,N_3570);
nand U3851 (N_3851,N_3583,N_3362);
or U3852 (N_3852,N_3346,N_3544);
nor U3853 (N_3853,N_3311,N_3579);
xor U3854 (N_3854,N_3656,N_3135);
nand U3855 (N_3855,N_3536,N_3748);
or U3856 (N_3856,N_3728,N_3258);
nand U3857 (N_3857,N_3514,N_3633);
xnor U3858 (N_3858,N_3551,N_3159);
nor U3859 (N_3859,N_3647,N_3552);
or U3860 (N_3860,N_3595,N_3654);
nor U3861 (N_3861,N_3401,N_3589);
nor U3862 (N_3862,N_3394,N_3414);
nand U3863 (N_3863,N_3193,N_3481);
or U3864 (N_3864,N_3259,N_3270);
xor U3865 (N_3865,N_3413,N_3503);
xor U3866 (N_3866,N_3664,N_3613);
nor U3867 (N_3867,N_3290,N_3458);
and U3868 (N_3868,N_3392,N_3722);
or U3869 (N_3869,N_3127,N_3251);
and U3870 (N_3870,N_3334,N_3332);
and U3871 (N_3871,N_3597,N_3191);
or U3872 (N_3872,N_3408,N_3303);
and U3873 (N_3873,N_3203,N_3624);
or U3874 (N_3874,N_3299,N_3336);
nor U3875 (N_3875,N_3367,N_3740);
and U3876 (N_3876,N_3467,N_3575);
and U3877 (N_3877,N_3566,N_3513);
or U3878 (N_3878,N_3321,N_3539);
nand U3879 (N_3879,N_3470,N_3555);
or U3880 (N_3880,N_3131,N_3718);
or U3881 (N_3881,N_3695,N_3670);
and U3882 (N_3882,N_3180,N_3538);
nand U3883 (N_3883,N_3310,N_3688);
or U3884 (N_3884,N_3620,N_3434);
xor U3885 (N_3885,N_3266,N_3462);
or U3886 (N_3886,N_3383,N_3247);
nor U3887 (N_3887,N_3686,N_3744);
nand U3888 (N_3888,N_3669,N_3644);
nand U3889 (N_3889,N_3156,N_3182);
and U3890 (N_3890,N_3292,N_3527);
nor U3891 (N_3891,N_3707,N_3437);
and U3892 (N_3892,N_3682,N_3427);
nor U3893 (N_3893,N_3371,N_3433);
nor U3894 (N_3894,N_3569,N_3701);
xor U3895 (N_3895,N_3468,N_3561);
xnor U3896 (N_3896,N_3646,N_3618);
nand U3897 (N_3897,N_3403,N_3316);
or U3898 (N_3898,N_3384,N_3596);
nand U3899 (N_3899,N_3729,N_3352);
xnor U3900 (N_3900,N_3528,N_3609);
nor U3901 (N_3901,N_3245,N_3518);
and U3902 (N_3902,N_3344,N_3214);
nor U3903 (N_3903,N_3439,N_3275);
nand U3904 (N_3904,N_3502,N_3170);
xor U3905 (N_3905,N_3747,N_3622);
and U3906 (N_3906,N_3730,N_3287);
or U3907 (N_3907,N_3665,N_3474);
and U3908 (N_3908,N_3498,N_3678);
nand U3909 (N_3909,N_3672,N_3661);
or U3910 (N_3910,N_3673,N_3737);
xnor U3911 (N_3911,N_3396,N_3276);
and U3912 (N_3912,N_3457,N_3577);
nand U3913 (N_3913,N_3643,N_3459);
nor U3914 (N_3914,N_3356,N_3363);
xnor U3915 (N_3915,N_3745,N_3429);
xnor U3916 (N_3916,N_3690,N_3142);
nand U3917 (N_3917,N_3705,N_3141);
xnor U3918 (N_3918,N_3746,N_3494);
nor U3919 (N_3919,N_3208,N_3308);
nor U3920 (N_3920,N_3649,N_3542);
and U3921 (N_3921,N_3397,N_3675);
xor U3922 (N_3922,N_3184,N_3485);
nand U3923 (N_3923,N_3329,N_3711);
nor U3924 (N_3924,N_3412,N_3252);
nor U3925 (N_3925,N_3226,N_3222);
nand U3926 (N_3926,N_3400,N_3280);
nand U3927 (N_3927,N_3509,N_3152);
nor U3928 (N_3928,N_3475,N_3409);
xnor U3929 (N_3929,N_3318,N_3164);
or U3930 (N_3930,N_3149,N_3534);
nand U3931 (N_3931,N_3712,N_3134);
nor U3932 (N_3932,N_3625,N_3438);
xor U3933 (N_3933,N_3189,N_3385);
nor U3934 (N_3934,N_3697,N_3140);
nand U3935 (N_3935,N_3353,N_3289);
nand U3936 (N_3936,N_3136,N_3578);
xnor U3937 (N_3937,N_3328,N_3463);
nand U3938 (N_3938,N_3220,N_3153);
and U3939 (N_3939,N_3441,N_3607);
xnor U3940 (N_3940,N_3133,N_3626);
and U3941 (N_3941,N_3530,N_3443);
and U3942 (N_3942,N_3240,N_3347);
or U3943 (N_3943,N_3716,N_3300);
or U3944 (N_3944,N_3233,N_3549);
nor U3945 (N_3945,N_3508,N_3568);
xor U3946 (N_3946,N_3691,N_3564);
nor U3947 (N_3947,N_3386,N_3448);
and U3948 (N_3948,N_3720,N_3615);
or U3949 (N_3949,N_3681,N_3199);
nand U3950 (N_3950,N_3250,N_3307);
nor U3951 (N_3951,N_3210,N_3365);
nand U3952 (N_3952,N_3320,N_3456);
xor U3953 (N_3953,N_3465,N_3405);
nor U3954 (N_3954,N_3679,N_3627);
or U3955 (N_3955,N_3450,N_3333);
nor U3956 (N_3956,N_3487,N_3306);
xnor U3957 (N_3957,N_3192,N_3702);
or U3958 (N_3958,N_3186,N_3639);
and U3959 (N_3959,N_3378,N_3484);
nand U3960 (N_3960,N_3628,N_3234);
xor U3961 (N_3961,N_3274,N_3345);
nand U3962 (N_3962,N_3213,N_3265);
and U3963 (N_3963,N_3125,N_3145);
nor U3964 (N_3964,N_3653,N_3143);
xor U3965 (N_3965,N_3727,N_3293);
nor U3966 (N_3966,N_3446,N_3359);
nor U3967 (N_3967,N_3382,N_3340);
xnor U3968 (N_3968,N_3489,N_3657);
and U3969 (N_3969,N_3298,N_3368);
xor U3970 (N_3970,N_3215,N_3389);
nand U3971 (N_3971,N_3693,N_3594);
nand U3972 (N_3972,N_3301,N_3324);
nand U3973 (N_3973,N_3331,N_3668);
and U3974 (N_3974,N_3327,N_3651);
nor U3975 (N_3975,N_3621,N_3617);
and U3976 (N_3976,N_3557,N_3381);
nand U3977 (N_3977,N_3272,N_3398);
xnor U3978 (N_3978,N_3689,N_3662);
xnor U3979 (N_3979,N_3230,N_3455);
or U3980 (N_3980,N_3227,N_3137);
nand U3981 (N_3981,N_3599,N_3505);
and U3982 (N_3982,N_3169,N_3519);
nor U3983 (N_3983,N_3338,N_3723);
and U3984 (N_3984,N_3126,N_3491);
or U3985 (N_3985,N_3241,N_3260);
xnor U3986 (N_3986,N_3268,N_3614);
nand U3987 (N_3987,N_3736,N_3129);
nor U3988 (N_3988,N_3171,N_3543);
nand U3989 (N_3989,N_3529,N_3674);
nand U3990 (N_3990,N_3516,N_3531);
nand U3991 (N_3991,N_3294,N_3592);
and U3992 (N_3992,N_3619,N_3319);
or U3993 (N_3993,N_3225,N_3372);
nor U3994 (N_3994,N_3601,N_3598);
nand U3995 (N_3995,N_3731,N_3553);
xnor U3996 (N_3996,N_3635,N_3216);
nand U3997 (N_3997,N_3482,N_3393);
nor U3998 (N_3998,N_3416,N_3373);
nor U3999 (N_3999,N_3608,N_3201);
and U4000 (N_4000,N_3209,N_3239);
nand U4001 (N_4001,N_3173,N_3721);
xnor U4002 (N_4002,N_3645,N_3559);
or U4003 (N_4003,N_3364,N_3506);
or U4004 (N_4004,N_3273,N_3504);
xnor U4005 (N_4005,N_3477,N_3734);
or U4006 (N_4006,N_3232,N_3507);
or U4007 (N_4007,N_3379,N_3219);
and U4008 (N_4008,N_3660,N_3223);
xnor U4009 (N_4009,N_3302,N_3550);
and U4010 (N_4010,N_3130,N_3178);
xor U4011 (N_4011,N_3444,N_3128);
or U4012 (N_4012,N_3556,N_3235);
or U4013 (N_4013,N_3228,N_3738);
xnor U4014 (N_4014,N_3337,N_3488);
xnor U4015 (N_4015,N_3146,N_3221);
and U4016 (N_4016,N_3447,N_3358);
nand U4017 (N_4017,N_3680,N_3719);
nor U4018 (N_4018,N_3632,N_3567);
nand U4019 (N_4019,N_3671,N_3269);
and U4020 (N_4020,N_3204,N_3197);
nand U4021 (N_4021,N_3147,N_3652);
nor U4022 (N_4022,N_3495,N_3296);
nor U4023 (N_4023,N_3623,N_3291);
nor U4024 (N_4024,N_3546,N_3473);
nand U4025 (N_4025,N_3242,N_3402);
or U4026 (N_4026,N_3376,N_3606);
or U4027 (N_4027,N_3148,N_3425);
or U4028 (N_4028,N_3515,N_3218);
nand U4029 (N_4029,N_3282,N_3611);
and U4030 (N_4030,N_3155,N_3168);
nand U4031 (N_4031,N_3541,N_3154);
nand U4032 (N_4032,N_3435,N_3237);
nand U4033 (N_4033,N_3174,N_3388);
or U4034 (N_4034,N_3248,N_3479);
xnor U4035 (N_4035,N_3732,N_3469);
nor U4036 (N_4036,N_3749,N_3350);
or U4037 (N_4037,N_3698,N_3742);
nand U4038 (N_4038,N_3390,N_3167);
xor U4039 (N_4039,N_3717,N_3525);
nand U4040 (N_4040,N_3370,N_3590);
nor U4041 (N_4041,N_3150,N_3677);
xor U4042 (N_4042,N_3255,N_3472);
or U4043 (N_4043,N_3725,N_3460);
or U4044 (N_4044,N_3522,N_3490);
nor U4045 (N_4045,N_3421,N_3284);
or U4046 (N_4046,N_3246,N_3428);
nand U4047 (N_4047,N_3211,N_3295);
xor U4048 (N_4048,N_3726,N_3581);
nor U4049 (N_4049,N_3471,N_3493);
nor U4050 (N_4050,N_3500,N_3700);
and U4051 (N_4051,N_3312,N_3634);
nor U4052 (N_4052,N_3476,N_3281);
nor U4053 (N_4053,N_3667,N_3545);
nand U4054 (N_4054,N_3480,N_3406);
nor U4055 (N_4055,N_3687,N_3451);
and U4056 (N_4056,N_3603,N_3440);
and U4057 (N_4057,N_3138,N_3181);
xor U4058 (N_4058,N_3231,N_3415);
xnor U4059 (N_4059,N_3335,N_3190);
and U4060 (N_4060,N_3453,N_3162);
nand U4061 (N_4061,N_3587,N_3257);
xor U4062 (N_4062,N_3349,N_3659);
xor U4063 (N_4063,N_3506,N_3421);
xor U4064 (N_4064,N_3428,N_3131);
and U4065 (N_4065,N_3447,N_3266);
nor U4066 (N_4066,N_3678,N_3407);
or U4067 (N_4067,N_3695,N_3312);
and U4068 (N_4068,N_3356,N_3720);
and U4069 (N_4069,N_3474,N_3335);
nand U4070 (N_4070,N_3289,N_3343);
nand U4071 (N_4071,N_3470,N_3305);
and U4072 (N_4072,N_3494,N_3406);
nand U4073 (N_4073,N_3290,N_3289);
nor U4074 (N_4074,N_3353,N_3204);
xor U4075 (N_4075,N_3681,N_3687);
and U4076 (N_4076,N_3316,N_3571);
nor U4077 (N_4077,N_3382,N_3621);
nor U4078 (N_4078,N_3738,N_3572);
or U4079 (N_4079,N_3564,N_3271);
nor U4080 (N_4080,N_3522,N_3373);
nand U4081 (N_4081,N_3588,N_3525);
nand U4082 (N_4082,N_3521,N_3655);
or U4083 (N_4083,N_3397,N_3226);
and U4084 (N_4084,N_3414,N_3557);
nor U4085 (N_4085,N_3569,N_3174);
nor U4086 (N_4086,N_3368,N_3182);
or U4087 (N_4087,N_3455,N_3722);
nor U4088 (N_4088,N_3741,N_3654);
nand U4089 (N_4089,N_3607,N_3478);
and U4090 (N_4090,N_3223,N_3550);
nand U4091 (N_4091,N_3167,N_3447);
xnor U4092 (N_4092,N_3371,N_3627);
nand U4093 (N_4093,N_3464,N_3136);
nor U4094 (N_4094,N_3153,N_3308);
xnor U4095 (N_4095,N_3549,N_3740);
or U4096 (N_4096,N_3497,N_3323);
or U4097 (N_4097,N_3599,N_3345);
nor U4098 (N_4098,N_3659,N_3367);
nor U4099 (N_4099,N_3528,N_3204);
xor U4100 (N_4100,N_3742,N_3192);
or U4101 (N_4101,N_3745,N_3358);
or U4102 (N_4102,N_3680,N_3287);
nor U4103 (N_4103,N_3385,N_3390);
nor U4104 (N_4104,N_3388,N_3709);
or U4105 (N_4105,N_3172,N_3701);
xnor U4106 (N_4106,N_3744,N_3236);
xor U4107 (N_4107,N_3630,N_3410);
xor U4108 (N_4108,N_3608,N_3268);
nand U4109 (N_4109,N_3423,N_3692);
and U4110 (N_4110,N_3293,N_3248);
xnor U4111 (N_4111,N_3362,N_3593);
and U4112 (N_4112,N_3531,N_3518);
or U4113 (N_4113,N_3720,N_3204);
or U4114 (N_4114,N_3245,N_3651);
nor U4115 (N_4115,N_3628,N_3618);
nor U4116 (N_4116,N_3331,N_3143);
or U4117 (N_4117,N_3460,N_3540);
nor U4118 (N_4118,N_3693,N_3366);
nand U4119 (N_4119,N_3259,N_3233);
and U4120 (N_4120,N_3175,N_3629);
nand U4121 (N_4121,N_3462,N_3485);
xnor U4122 (N_4122,N_3531,N_3513);
nor U4123 (N_4123,N_3398,N_3744);
nor U4124 (N_4124,N_3619,N_3735);
xor U4125 (N_4125,N_3634,N_3501);
nor U4126 (N_4126,N_3497,N_3460);
or U4127 (N_4127,N_3728,N_3171);
xor U4128 (N_4128,N_3474,N_3731);
nand U4129 (N_4129,N_3701,N_3679);
nor U4130 (N_4130,N_3732,N_3417);
nor U4131 (N_4131,N_3674,N_3212);
xor U4132 (N_4132,N_3603,N_3655);
nand U4133 (N_4133,N_3414,N_3438);
xnor U4134 (N_4134,N_3312,N_3291);
xnor U4135 (N_4135,N_3154,N_3471);
nor U4136 (N_4136,N_3262,N_3224);
and U4137 (N_4137,N_3365,N_3639);
nor U4138 (N_4138,N_3380,N_3186);
xor U4139 (N_4139,N_3289,N_3385);
xor U4140 (N_4140,N_3151,N_3373);
xnor U4141 (N_4141,N_3341,N_3370);
or U4142 (N_4142,N_3377,N_3659);
xor U4143 (N_4143,N_3448,N_3591);
or U4144 (N_4144,N_3190,N_3488);
nor U4145 (N_4145,N_3707,N_3555);
nand U4146 (N_4146,N_3703,N_3559);
xor U4147 (N_4147,N_3670,N_3744);
nor U4148 (N_4148,N_3246,N_3417);
nor U4149 (N_4149,N_3267,N_3455);
or U4150 (N_4150,N_3749,N_3588);
xnor U4151 (N_4151,N_3204,N_3573);
nand U4152 (N_4152,N_3641,N_3346);
nor U4153 (N_4153,N_3244,N_3516);
or U4154 (N_4154,N_3574,N_3344);
nor U4155 (N_4155,N_3545,N_3207);
nand U4156 (N_4156,N_3711,N_3646);
nand U4157 (N_4157,N_3394,N_3676);
nor U4158 (N_4158,N_3633,N_3461);
nor U4159 (N_4159,N_3639,N_3364);
or U4160 (N_4160,N_3212,N_3164);
xor U4161 (N_4161,N_3623,N_3577);
or U4162 (N_4162,N_3668,N_3442);
nand U4163 (N_4163,N_3294,N_3601);
xor U4164 (N_4164,N_3480,N_3600);
xnor U4165 (N_4165,N_3149,N_3203);
or U4166 (N_4166,N_3382,N_3728);
xnor U4167 (N_4167,N_3498,N_3721);
xor U4168 (N_4168,N_3628,N_3310);
or U4169 (N_4169,N_3543,N_3594);
and U4170 (N_4170,N_3232,N_3744);
or U4171 (N_4171,N_3672,N_3408);
nand U4172 (N_4172,N_3475,N_3294);
nor U4173 (N_4173,N_3278,N_3174);
or U4174 (N_4174,N_3345,N_3546);
or U4175 (N_4175,N_3590,N_3672);
and U4176 (N_4176,N_3601,N_3523);
or U4177 (N_4177,N_3667,N_3512);
xor U4178 (N_4178,N_3717,N_3278);
xnor U4179 (N_4179,N_3565,N_3550);
xnor U4180 (N_4180,N_3131,N_3531);
or U4181 (N_4181,N_3212,N_3597);
xnor U4182 (N_4182,N_3182,N_3511);
xnor U4183 (N_4183,N_3657,N_3272);
or U4184 (N_4184,N_3340,N_3642);
nor U4185 (N_4185,N_3151,N_3612);
nor U4186 (N_4186,N_3514,N_3612);
and U4187 (N_4187,N_3333,N_3380);
nand U4188 (N_4188,N_3377,N_3349);
or U4189 (N_4189,N_3341,N_3149);
nand U4190 (N_4190,N_3265,N_3151);
xnor U4191 (N_4191,N_3457,N_3305);
nand U4192 (N_4192,N_3213,N_3669);
nor U4193 (N_4193,N_3255,N_3491);
and U4194 (N_4194,N_3334,N_3134);
nor U4195 (N_4195,N_3208,N_3214);
or U4196 (N_4196,N_3452,N_3237);
and U4197 (N_4197,N_3381,N_3440);
and U4198 (N_4198,N_3606,N_3702);
or U4199 (N_4199,N_3312,N_3475);
and U4200 (N_4200,N_3636,N_3606);
xor U4201 (N_4201,N_3141,N_3185);
xnor U4202 (N_4202,N_3220,N_3511);
nor U4203 (N_4203,N_3670,N_3211);
xnor U4204 (N_4204,N_3181,N_3637);
xor U4205 (N_4205,N_3256,N_3234);
nand U4206 (N_4206,N_3220,N_3237);
or U4207 (N_4207,N_3322,N_3667);
xor U4208 (N_4208,N_3290,N_3277);
nand U4209 (N_4209,N_3374,N_3244);
and U4210 (N_4210,N_3472,N_3191);
nor U4211 (N_4211,N_3661,N_3437);
xnor U4212 (N_4212,N_3660,N_3432);
or U4213 (N_4213,N_3456,N_3253);
and U4214 (N_4214,N_3244,N_3291);
nor U4215 (N_4215,N_3606,N_3545);
xnor U4216 (N_4216,N_3599,N_3199);
xnor U4217 (N_4217,N_3354,N_3684);
nand U4218 (N_4218,N_3369,N_3464);
xnor U4219 (N_4219,N_3292,N_3330);
or U4220 (N_4220,N_3322,N_3733);
xnor U4221 (N_4221,N_3505,N_3275);
nor U4222 (N_4222,N_3171,N_3247);
or U4223 (N_4223,N_3222,N_3338);
or U4224 (N_4224,N_3462,N_3172);
and U4225 (N_4225,N_3250,N_3318);
or U4226 (N_4226,N_3429,N_3274);
nand U4227 (N_4227,N_3242,N_3683);
and U4228 (N_4228,N_3679,N_3371);
or U4229 (N_4229,N_3469,N_3427);
and U4230 (N_4230,N_3269,N_3172);
and U4231 (N_4231,N_3424,N_3744);
nor U4232 (N_4232,N_3440,N_3443);
nor U4233 (N_4233,N_3145,N_3685);
nand U4234 (N_4234,N_3554,N_3662);
and U4235 (N_4235,N_3260,N_3469);
nand U4236 (N_4236,N_3737,N_3557);
xnor U4237 (N_4237,N_3661,N_3393);
nand U4238 (N_4238,N_3533,N_3634);
and U4239 (N_4239,N_3416,N_3453);
nor U4240 (N_4240,N_3701,N_3652);
xnor U4241 (N_4241,N_3672,N_3603);
xnor U4242 (N_4242,N_3465,N_3179);
nor U4243 (N_4243,N_3717,N_3651);
or U4244 (N_4244,N_3507,N_3497);
xnor U4245 (N_4245,N_3298,N_3322);
xnor U4246 (N_4246,N_3450,N_3575);
xnor U4247 (N_4247,N_3526,N_3658);
xor U4248 (N_4248,N_3236,N_3166);
and U4249 (N_4249,N_3264,N_3503);
nand U4250 (N_4250,N_3211,N_3429);
xor U4251 (N_4251,N_3584,N_3577);
and U4252 (N_4252,N_3451,N_3336);
or U4253 (N_4253,N_3622,N_3685);
nor U4254 (N_4254,N_3260,N_3367);
xor U4255 (N_4255,N_3344,N_3135);
nor U4256 (N_4256,N_3565,N_3551);
or U4257 (N_4257,N_3463,N_3233);
or U4258 (N_4258,N_3560,N_3634);
and U4259 (N_4259,N_3650,N_3207);
xor U4260 (N_4260,N_3240,N_3158);
and U4261 (N_4261,N_3139,N_3739);
and U4262 (N_4262,N_3709,N_3253);
or U4263 (N_4263,N_3324,N_3304);
nand U4264 (N_4264,N_3563,N_3279);
or U4265 (N_4265,N_3626,N_3383);
nor U4266 (N_4266,N_3638,N_3416);
and U4267 (N_4267,N_3236,N_3237);
xnor U4268 (N_4268,N_3667,N_3323);
nand U4269 (N_4269,N_3730,N_3212);
or U4270 (N_4270,N_3294,N_3398);
xnor U4271 (N_4271,N_3424,N_3675);
or U4272 (N_4272,N_3571,N_3221);
nor U4273 (N_4273,N_3527,N_3558);
xnor U4274 (N_4274,N_3547,N_3284);
and U4275 (N_4275,N_3406,N_3529);
xor U4276 (N_4276,N_3633,N_3641);
nor U4277 (N_4277,N_3264,N_3298);
and U4278 (N_4278,N_3624,N_3190);
or U4279 (N_4279,N_3333,N_3568);
nand U4280 (N_4280,N_3276,N_3471);
nor U4281 (N_4281,N_3567,N_3631);
nand U4282 (N_4282,N_3709,N_3583);
nor U4283 (N_4283,N_3560,N_3233);
or U4284 (N_4284,N_3358,N_3193);
and U4285 (N_4285,N_3575,N_3413);
and U4286 (N_4286,N_3438,N_3733);
nand U4287 (N_4287,N_3363,N_3721);
nor U4288 (N_4288,N_3191,N_3397);
nand U4289 (N_4289,N_3698,N_3681);
xor U4290 (N_4290,N_3406,N_3309);
xnor U4291 (N_4291,N_3565,N_3678);
or U4292 (N_4292,N_3732,N_3547);
xor U4293 (N_4293,N_3462,N_3675);
nand U4294 (N_4294,N_3564,N_3651);
xnor U4295 (N_4295,N_3190,N_3528);
xor U4296 (N_4296,N_3289,N_3136);
nand U4297 (N_4297,N_3242,N_3622);
xnor U4298 (N_4298,N_3407,N_3232);
nor U4299 (N_4299,N_3592,N_3320);
xor U4300 (N_4300,N_3687,N_3524);
or U4301 (N_4301,N_3598,N_3399);
xnor U4302 (N_4302,N_3181,N_3202);
or U4303 (N_4303,N_3681,N_3626);
xnor U4304 (N_4304,N_3324,N_3541);
nor U4305 (N_4305,N_3561,N_3446);
nor U4306 (N_4306,N_3397,N_3524);
xor U4307 (N_4307,N_3656,N_3234);
nand U4308 (N_4308,N_3190,N_3436);
nor U4309 (N_4309,N_3604,N_3359);
xnor U4310 (N_4310,N_3464,N_3689);
or U4311 (N_4311,N_3303,N_3537);
xnor U4312 (N_4312,N_3615,N_3211);
or U4313 (N_4313,N_3474,N_3386);
and U4314 (N_4314,N_3701,N_3292);
or U4315 (N_4315,N_3242,N_3510);
nand U4316 (N_4316,N_3452,N_3360);
xnor U4317 (N_4317,N_3656,N_3686);
nor U4318 (N_4318,N_3230,N_3442);
nor U4319 (N_4319,N_3252,N_3410);
or U4320 (N_4320,N_3193,N_3205);
or U4321 (N_4321,N_3258,N_3514);
nor U4322 (N_4322,N_3633,N_3304);
nand U4323 (N_4323,N_3706,N_3707);
and U4324 (N_4324,N_3567,N_3354);
xnor U4325 (N_4325,N_3266,N_3551);
nand U4326 (N_4326,N_3367,N_3517);
and U4327 (N_4327,N_3369,N_3324);
nand U4328 (N_4328,N_3512,N_3341);
nor U4329 (N_4329,N_3258,N_3178);
nand U4330 (N_4330,N_3230,N_3440);
nand U4331 (N_4331,N_3428,N_3721);
nor U4332 (N_4332,N_3459,N_3351);
xnor U4333 (N_4333,N_3624,N_3508);
and U4334 (N_4334,N_3249,N_3450);
or U4335 (N_4335,N_3687,N_3680);
xor U4336 (N_4336,N_3412,N_3163);
and U4337 (N_4337,N_3161,N_3704);
nor U4338 (N_4338,N_3197,N_3354);
and U4339 (N_4339,N_3528,N_3155);
and U4340 (N_4340,N_3451,N_3130);
nor U4341 (N_4341,N_3537,N_3244);
xnor U4342 (N_4342,N_3693,N_3582);
nand U4343 (N_4343,N_3443,N_3303);
or U4344 (N_4344,N_3537,N_3593);
nor U4345 (N_4345,N_3677,N_3304);
nand U4346 (N_4346,N_3383,N_3720);
nor U4347 (N_4347,N_3437,N_3666);
or U4348 (N_4348,N_3496,N_3351);
nor U4349 (N_4349,N_3171,N_3339);
and U4350 (N_4350,N_3346,N_3575);
or U4351 (N_4351,N_3719,N_3665);
or U4352 (N_4352,N_3745,N_3528);
nand U4353 (N_4353,N_3295,N_3431);
nand U4354 (N_4354,N_3505,N_3694);
xnor U4355 (N_4355,N_3268,N_3665);
or U4356 (N_4356,N_3488,N_3305);
and U4357 (N_4357,N_3382,N_3377);
nor U4358 (N_4358,N_3622,N_3624);
nand U4359 (N_4359,N_3476,N_3529);
nor U4360 (N_4360,N_3152,N_3580);
nor U4361 (N_4361,N_3698,N_3240);
or U4362 (N_4362,N_3682,N_3171);
or U4363 (N_4363,N_3267,N_3308);
nor U4364 (N_4364,N_3566,N_3272);
and U4365 (N_4365,N_3707,N_3655);
nand U4366 (N_4366,N_3404,N_3306);
xor U4367 (N_4367,N_3716,N_3684);
or U4368 (N_4368,N_3525,N_3501);
xor U4369 (N_4369,N_3162,N_3313);
and U4370 (N_4370,N_3610,N_3724);
nand U4371 (N_4371,N_3520,N_3515);
xnor U4372 (N_4372,N_3554,N_3244);
nor U4373 (N_4373,N_3452,N_3488);
and U4374 (N_4374,N_3545,N_3375);
xnor U4375 (N_4375,N_3988,N_3887);
nor U4376 (N_4376,N_3774,N_4225);
and U4377 (N_4377,N_4035,N_4199);
or U4378 (N_4378,N_4257,N_4325);
and U4379 (N_4379,N_4269,N_4373);
xor U4380 (N_4380,N_3868,N_3943);
or U4381 (N_4381,N_3779,N_4064);
and U4382 (N_4382,N_3948,N_3944);
nor U4383 (N_4383,N_4371,N_4060);
xnor U4384 (N_4384,N_4326,N_4022);
nand U4385 (N_4385,N_3980,N_3938);
xnor U4386 (N_4386,N_4366,N_4043);
or U4387 (N_4387,N_4249,N_4331);
and U4388 (N_4388,N_4195,N_3947);
xor U4389 (N_4389,N_4251,N_3959);
or U4390 (N_4390,N_3768,N_4115);
nand U4391 (N_4391,N_3782,N_4224);
and U4392 (N_4392,N_4023,N_4092);
or U4393 (N_4393,N_4038,N_3850);
and U4394 (N_4394,N_3998,N_3916);
and U4395 (N_4395,N_4059,N_3780);
and U4396 (N_4396,N_4200,N_3917);
and U4397 (N_4397,N_4279,N_3922);
xnor U4398 (N_4398,N_4363,N_4046);
nor U4399 (N_4399,N_4079,N_4024);
xnor U4400 (N_4400,N_3974,N_3890);
nand U4401 (N_4401,N_4278,N_3940);
and U4402 (N_4402,N_4283,N_4179);
or U4403 (N_4403,N_4147,N_4328);
or U4404 (N_4404,N_4051,N_3787);
xor U4405 (N_4405,N_4004,N_4314);
nand U4406 (N_4406,N_4333,N_4086);
or U4407 (N_4407,N_4361,N_3790);
or U4408 (N_4408,N_3800,N_4159);
nand U4409 (N_4409,N_3818,N_4360);
nand U4410 (N_4410,N_4210,N_4223);
nand U4411 (N_4411,N_4134,N_3759);
or U4412 (N_4412,N_3777,N_3860);
nand U4413 (N_4413,N_4213,N_4356);
or U4414 (N_4414,N_3976,N_3880);
or U4415 (N_4415,N_4012,N_3961);
or U4416 (N_4416,N_4364,N_3793);
xnor U4417 (N_4417,N_3865,N_4015);
nor U4418 (N_4418,N_4300,N_4165);
and U4419 (N_4419,N_4085,N_3760);
and U4420 (N_4420,N_4353,N_4172);
nor U4421 (N_4421,N_3762,N_4139);
xnor U4422 (N_4422,N_4002,N_3897);
nand U4423 (N_4423,N_3789,N_4344);
nand U4424 (N_4424,N_4112,N_4266);
xor U4425 (N_4425,N_4233,N_4161);
nand U4426 (N_4426,N_3799,N_3968);
nor U4427 (N_4427,N_4070,N_3978);
and U4428 (N_4428,N_3870,N_4011);
and U4429 (N_4429,N_4080,N_3776);
or U4430 (N_4430,N_4227,N_3775);
and U4431 (N_4431,N_3771,N_4183);
nand U4432 (N_4432,N_3927,N_3894);
nand U4433 (N_4433,N_4054,N_4262);
nor U4434 (N_4434,N_4310,N_4191);
nand U4435 (N_4435,N_4355,N_3813);
xor U4436 (N_4436,N_3994,N_4194);
or U4437 (N_4437,N_3820,N_4126);
nor U4438 (N_4438,N_3846,N_3791);
or U4439 (N_4439,N_4350,N_4319);
nor U4440 (N_4440,N_4274,N_3911);
nand U4441 (N_4441,N_4248,N_4349);
nor U4442 (N_4442,N_4055,N_4313);
and U4443 (N_4443,N_3814,N_3839);
nand U4444 (N_4444,N_3951,N_3769);
or U4445 (N_4445,N_3928,N_4317);
and U4446 (N_4446,N_4261,N_4323);
nand U4447 (N_4447,N_4304,N_3979);
or U4448 (N_4448,N_4288,N_4107);
nor U4449 (N_4449,N_3995,N_3907);
or U4450 (N_4450,N_4268,N_4184);
and U4451 (N_4451,N_4169,N_3908);
nand U4452 (N_4452,N_4127,N_4050);
and U4453 (N_4453,N_3822,N_3902);
or U4454 (N_4454,N_4132,N_4216);
and U4455 (N_4455,N_4287,N_4186);
xor U4456 (N_4456,N_3990,N_3874);
xnor U4457 (N_4457,N_4252,N_4007);
or U4458 (N_4458,N_3946,N_4357);
xnor U4459 (N_4459,N_3861,N_4263);
nand U4460 (N_4460,N_3784,N_3914);
xor U4461 (N_4461,N_4187,N_3854);
and U4462 (N_4462,N_4280,N_3832);
nor U4463 (N_4463,N_3877,N_4155);
or U4464 (N_4464,N_4009,N_4005);
xor U4465 (N_4465,N_4207,N_3882);
or U4466 (N_4466,N_4352,N_3953);
nand U4467 (N_4467,N_4163,N_4048);
xor U4468 (N_4468,N_4108,N_4359);
and U4469 (N_4469,N_3954,N_4220);
xor U4470 (N_4470,N_3815,N_3848);
and U4471 (N_4471,N_3862,N_3801);
and U4472 (N_4472,N_3767,N_4081);
nor U4473 (N_4473,N_4197,N_4094);
nor U4474 (N_4474,N_4222,N_4236);
or U4475 (N_4475,N_3852,N_3925);
nand U4476 (N_4476,N_4158,N_4201);
or U4477 (N_4477,N_4311,N_4069);
and U4478 (N_4478,N_3888,N_3824);
or U4479 (N_4479,N_3991,N_4109);
and U4480 (N_4480,N_3772,N_4296);
or U4481 (N_4481,N_4097,N_4075);
or U4482 (N_4482,N_3872,N_3964);
and U4483 (N_4483,N_4273,N_4321);
or U4484 (N_4484,N_4206,N_3881);
or U4485 (N_4485,N_4088,N_4343);
and U4486 (N_4486,N_4071,N_4167);
nand U4487 (N_4487,N_4175,N_4276);
nor U4488 (N_4488,N_4334,N_4026);
nand U4489 (N_4489,N_3817,N_4341);
and U4490 (N_4490,N_4302,N_4033);
xnor U4491 (N_4491,N_4250,N_3984);
nor U4492 (N_4492,N_3807,N_4111);
or U4493 (N_4493,N_4282,N_3905);
nand U4494 (N_4494,N_4131,N_4087);
and U4495 (N_4495,N_4299,N_3755);
and U4496 (N_4496,N_3786,N_3886);
or U4497 (N_4497,N_4133,N_3924);
and U4498 (N_4498,N_3836,N_4077);
nand U4499 (N_4499,N_4370,N_4255);
xor U4500 (N_4500,N_3898,N_4148);
nor U4501 (N_4501,N_4156,N_4078);
and U4502 (N_4502,N_4093,N_3828);
nand U4503 (N_4503,N_4157,N_4217);
nand U4504 (N_4504,N_3867,N_3950);
nand U4505 (N_4505,N_4259,N_3983);
or U4506 (N_4506,N_3831,N_3751);
nand U4507 (N_4507,N_4219,N_4149);
or U4508 (N_4508,N_3834,N_4198);
and U4509 (N_4509,N_4138,N_3972);
nand U4510 (N_4510,N_3986,N_4053);
xor U4511 (N_4511,N_4245,N_4083);
nand U4512 (N_4512,N_3830,N_4190);
nand U4513 (N_4513,N_4332,N_3941);
and U4514 (N_4514,N_3891,N_4162);
nor U4515 (N_4515,N_3802,N_4065);
or U4516 (N_4516,N_3765,N_4253);
or U4517 (N_4517,N_3921,N_3808);
or U4518 (N_4518,N_4020,N_4120);
or U4519 (N_4519,N_3781,N_3931);
xor U4520 (N_4520,N_3838,N_4034);
and U4521 (N_4521,N_3909,N_3884);
nor U4522 (N_4522,N_3812,N_4119);
nor U4523 (N_4523,N_3809,N_3858);
xor U4524 (N_4524,N_4042,N_3923);
or U4525 (N_4525,N_4368,N_4286);
and U4526 (N_4526,N_4056,N_3840);
nand U4527 (N_4527,N_4105,N_3956);
and U4528 (N_4528,N_3811,N_3845);
xor U4529 (N_4529,N_4298,N_4218);
or U4530 (N_4530,N_4256,N_4058);
and U4531 (N_4531,N_4303,N_3883);
and U4532 (N_4532,N_3826,N_4312);
xnor U4533 (N_4533,N_3949,N_3837);
and U4534 (N_4534,N_4141,N_3999);
and U4535 (N_4535,N_3764,N_4103);
nor U4536 (N_4536,N_4072,N_4211);
nand U4537 (N_4537,N_4137,N_4171);
nand U4538 (N_4538,N_3859,N_3933);
and U4539 (N_4539,N_3942,N_4045);
xor U4540 (N_4540,N_4128,N_4084);
and U4541 (N_4541,N_3847,N_4316);
and U4542 (N_4542,N_4315,N_3778);
nand U4543 (N_4543,N_4052,N_3993);
nand U4544 (N_4544,N_3900,N_4068);
nor U4545 (N_4545,N_3920,N_3821);
or U4546 (N_4546,N_4322,N_4293);
nand U4547 (N_4547,N_4180,N_3798);
or U4548 (N_4548,N_4102,N_4168);
nor U4549 (N_4549,N_4150,N_3997);
nand U4550 (N_4550,N_3875,N_4308);
nand U4551 (N_4551,N_4151,N_3992);
xor U4552 (N_4552,N_3969,N_4208);
or U4553 (N_4553,N_4044,N_4099);
or U4554 (N_4554,N_3981,N_4057);
nand U4555 (N_4555,N_4289,N_3878);
xnor U4556 (N_4556,N_3932,N_3970);
and U4557 (N_4557,N_4265,N_4135);
nor U4558 (N_4558,N_3975,N_3803);
or U4559 (N_4559,N_4113,N_4309);
nor U4560 (N_4560,N_4152,N_3756);
xor U4561 (N_4561,N_3792,N_4267);
xor U4562 (N_4562,N_4330,N_3804);
and U4563 (N_4563,N_3855,N_4041);
nand U4564 (N_4564,N_3987,N_3757);
nand U4565 (N_4565,N_4241,N_4346);
and U4566 (N_4566,N_4324,N_3904);
xnor U4567 (N_4567,N_4095,N_4008);
and U4568 (N_4568,N_4067,N_4305);
and U4569 (N_4569,N_3788,N_4226);
xnor U4570 (N_4570,N_4030,N_4329);
nand U4571 (N_4571,N_3844,N_3752);
or U4572 (N_4572,N_3849,N_4284);
nand U4573 (N_4573,N_3758,N_3753);
nand U4574 (N_4574,N_3971,N_3977);
xor U4575 (N_4575,N_3885,N_3982);
or U4576 (N_4576,N_4039,N_4181);
nor U4577 (N_4577,N_4114,N_4285);
xnor U4578 (N_4578,N_3952,N_4367);
nor U4579 (N_4579,N_4027,N_4215);
nor U4580 (N_4580,N_4320,N_4117);
nand U4581 (N_4581,N_3829,N_3973);
nor U4582 (N_4582,N_3816,N_3823);
nand U4583 (N_4583,N_3843,N_4238);
nor U4584 (N_4584,N_3879,N_4010);
or U4585 (N_4585,N_4337,N_3825);
nand U4586 (N_4586,N_3985,N_4205);
xor U4587 (N_4587,N_4176,N_3841);
nand U4588 (N_4588,N_4028,N_4096);
nor U4589 (N_4589,N_3945,N_4232);
nand U4590 (N_4590,N_4202,N_4244);
nor U4591 (N_4591,N_4275,N_3856);
nand U4592 (N_4592,N_4212,N_3842);
nand U4593 (N_4593,N_4348,N_4374);
nor U4594 (N_4594,N_4091,N_4237);
xnor U4595 (N_4595,N_3853,N_3957);
or U4596 (N_4596,N_3866,N_4170);
nor U4597 (N_4597,N_4240,N_3750);
nor U4598 (N_4598,N_3889,N_4017);
nand U4599 (N_4599,N_3773,N_3919);
or U4600 (N_4600,N_4228,N_4369);
xnor U4601 (N_4601,N_3851,N_3763);
xnor U4602 (N_4602,N_3958,N_4264);
xor U4603 (N_4603,N_3901,N_4076);
nor U4604 (N_4604,N_4189,N_4047);
xnor U4605 (N_4605,N_4182,N_4136);
xor U4606 (N_4606,N_3937,N_4318);
xor U4607 (N_4607,N_4339,N_4101);
and U4608 (N_4608,N_4082,N_4291);
and U4609 (N_4609,N_4365,N_4106);
and U4610 (N_4610,N_3963,N_4014);
nor U4611 (N_4611,N_4307,N_4025);
or U4612 (N_4612,N_4243,N_4290);
nand U4613 (N_4613,N_3939,N_3873);
nand U4614 (N_4614,N_3918,N_4142);
or U4615 (N_4615,N_4254,N_3934);
nand U4616 (N_4616,N_4063,N_3864);
nor U4617 (N_4617,N_4089,N_4049);
nor U4618 (N_4618,N_3915,N_4016);
nand U4619 (N_4619,N_3871,N_4340);
and U4620 (N_4620,N_4153,N_3766);
and U4621 (N_4621,N_3827,N_4140);
and U4622 (N_4622,N_4110,N_4090);
xor U4623 (N_4623,N_4196,N_4021);
and U4624 (N_4624,N_4164,N_4229);
nand U4625 (N_4625,N_4029,N_4272);
or U4626 (N_4626,N_3926,N_4301);
and U4627 (N_4627,N_3796,N_4347);
and U4628 (N_4628,N_3930,N_4338);
xnor U4629 (N_4629,N_4239,N_3895);
nand U4630 (N_4630,N_4116,N_4281);
nand U4631 (N_4631,N_4297,N_4271);
xor U4632 (N_4632,N_4258,N_3869);
nor U4633 (N_4633,N_4098,N_4154);
and U4634 (N_4634,N_4124,N_3896);
and U4635 (N_4635,N_3770,N_3794);
or U4636 (N_4636,N_4032,N_4061);
nand U4637 (N_4637,N_4335,N_3783);
xnor U4638 (N_4638,N_4174,N_4351);
nand U4639 (N_4639,N_3965,N_3960);
or U4640 (N_4640,N_4003,N_3899);
and U4641 (N_4641,N_3966,N_3893);
nor U4642 (N_4642,N_3955,N_3929);
or U4643 (N_4643,N_4294,N_4292);
nand U4644 (N_4644,N_4129,N_4062);
xnor U4645 (N_4645,N_3906,N_4372);
nand U4646 (N_4646,N_4230,N_4100);
nor U4647 (N_4647,N_4345,N_4234);
nor U4648 (N_4648,N_4122,N_4177);
nor U4649 (N_4649,N_4277,N_4066);
and U4650 (N_4650,N_4362,N_4235);
or U4651 (N_4651,N_4203,N_4146);
nor U4652 (N_4652,N_4242,N_4246);
and U4653 (N_4653,N_3806,N_4221);
or U4654 (N_4654,N_4000,N_3967);
and U4655 (N_4655,N_3935,N_4358);
or U4656 (N_4656,N_4342,N_4354);
or U4657 (N_4657,N_3785,N_4144);
nor U4658 (N_4658,N_4036,N_3910);
or U4659 (N_4659,N_4193,N_3833);
or U4660 (N_4660,N_3962,N_4121);
nor U4661 (N_4661,N_4192,N_4037);
nand U4662 (N_4662,N_4214,N_4130);
nand U4663 (N_4663,N_4160,N_3805);
and U4664 (N_4664,N_4125,N_3936);
or U4665 (N_4665,N_4073,N_4031);
xnor U4666 (N_4666,N_4019,N_3754);
xor U4667 (N_4667,N_4006,N_4118);
or U4668 (N_4668,N_4173,N_4270);
xor U4669 (N_4669,N_4247,N_3903);
nor U4670 (N_4670,N_4327,N_3863);
or U4671 (N_4671,N_4306,N_4209);
nand U4672 (N_4672,N_4013,N_4143);
nor U4673 (N_4673,N_3819,N_3810);
nor U4674 (N_4674,N_3989,N_3795);
nand U4675 (N_4675,N_4231,N_3876);
nor U4676 (N_4676,N_4104,N_4295);
xor U4677 (N_4677,N_4040,N_3913);
or U4678 (N_4678,N_4145,N_3761);
xnor U4679 (N_4679,N_4260,N_4074);
nor U4680 (N_4680,N_3835,N_3857);
xnor U4681 (N_4681,N_4018,N_4166);
nand U4682 (N_4682,N_4204,N_4188);
and U4683 (N_4683,N_3996,N_3892);
or U4684 (N_4684,N_3912,N_4123);
nor U4685 (N_4685,N_3797,N_4185);
and U4686 (N_4686,N_4336,N_4178);
nor U4687 (N_4687,N_4001,N_4163);
nor U4688 (N_4688,N_4005,N_3933);
and U4689 (N_4689,N_3849,N_3855);
nand U4690 (N_4690,N_4140,N_3950);
or U4691 (N_4691,N_4223,N_4164);
or U4692 (N_4692,N_3982,N_4364);
nor U4693 (N_4693,N_3913,N_3821);
nor U4694 (N_4694,N_3793,N_4369);
nand U4695 (N_4695,N_3904,N_4188);
xor U4696 (N_4696,N_4160,N_3913);
xnor U4697 (N_4697,N_4184,N_4225);
nor U4698 (N_4698,N_3982,N_3863);
nand U4699 (N_4699,N_3894,N_3875);
xor U4700 (N_4700,N_4014,N_3753);
or U4701 (N_4701,N_3956,N_3856);
nand U4702 (N_4702,N_3809,N_4003);
xor U4703 (N_4703,N_3798,N_4270);
nand U4704 (N_4704,N_4265,N_3847);
xnor U4705 (N_4705,N_3955,N_4342);
nand U4706 (N_4706,N_4257,N_4104);
nand U4707 (N_4707,N_3824,N_4239);
nor U4708 (N_4708,N_4265,N_4297);
xnor U4709 (N_4709,N_4222,N_4235);
nor U4710 (N_4710,N_4374,N_4265);
or U4711 (N_4711,N_4215,N_4022);
and U4712 (N_4712,N_4227,N_4166);
and U4713 (N_4713,N_4323,N_3791);
nor U4714 (N_4714,N_4260,N_3905);
xor U4715 (N_4715,N_4037,N_3905);
xor U4716 (N_4716,N_4048,N_3942);
nand U4717 (N_4717,N_4307,N_4014);
nor U4718 (N_4718,N_4142,N_4317);
nor U4719 (N_4719,N_3869,N_3909);
and U4720 (N_4720,N_4348,N_3978);
nor U4721 (N_4721,N_4278,N_4067);
xnor U4722 (N_4722,N_3778,N_3790);
xor U4723 (N_4723,N_4223,N_3805);
xor U4724 (N_4724,N_4172,N_3777);
nand U4725 (N_4725,N_3930,N_4166);
nor U4726 (N_4726,N_3843,N_4085);
or U4727 (N_4727,N_4191,N_3764);
xor U4728 (N_4728,N_4095,N_3779);
xnor U4729 (N_4729,N_3856,N_4246);
nor U4730 (N_4730,N_4154,N_4036);
or U4731 (N_4731,N_3772,N_4204);
nand U4732 (N_4732,N_3957,N_4153);
and U4733 (N_4733,N_4014,N_4147);
nand U4734 (N_4734,N_3819,N_3955);
and U4735 (N_4735,N_3905,N_3858);
or U4736 (N_4736,N_3969,N_4119);
nor U4737 (N_4737,N_4350,N_3817);
and U4738 (N_4738,N_4284,N_4154);
xor U4739 (N_4739,N_4008,N_3946);
xnor U4740 (N_4740,N_4307,N_4213);
nand U4741 (N_4741,N_4263,N_3930);
or U4742 (N_4742,N_4174,N_3907);
and U4743 (N_4743,N_3790,N_4003);
xnor U4744 (N_4744,N_3874,N_4204);
and U4745 (N_4745,N_3940,N_4196);
or U4746 (N_4746,N_4206,N_4275);
or U4747 (N_4747,N_4341,N_4178);
nor U4748 (N_4748,N_4007,N_4020);
xor U4749 (N_4749,N_4066,N_3839);
or U4750 (N_4750,N_4312,N_3935);
nand U4751 (N_4751,N_3754,N_4267);
or U4752 (N_4752,N_3894,N_4072);
or U4753 (N_4753,N_3759,N_4288);
xor U4754 (N_4754,N_4038,N_4182);
and U4755 (N_4755,N_3806,N_3780);
and U4756 (N_4756,N_3955,N_3751);
nor U4757 (N_4757,N_3954,N_4259);
xnor U4758 (N_4758,N_4096,N_4327);
nor U4759 (N_4759,N_4012,N_3787);
nand U4760 (N_4760,N_4227,N_4356);
nor U4761 (N_4761,N_4013,N_4260);
xor U4762 (N_4762,N_4364,N_3880);
nor U4763 (N_4763,N_3834,N_4331);
or U4764 (N_4764,N_4112,N_4040);
or U4765 (N_4765,N_3856,N_3977);
or U4766 (N_4766,N_3821,N_3864);
nor U4767 (N_4767,N_4192,N_4302);
or U4768 (N_4768,N_4226,N_4140);
nand U4769 (N_4769,N_4266,N_3915);
nand U4770 (N_4770,N_4096,N_3840);
and U4771 (N_4771,N_3933,N_4315);
and U4772 (N_4772,N_4331,N_4158);
nor U4773 (N_4773,N_3771,N_3795);
nor U4774 (N_4774,N_4064,N_4073);
xnor U4775 (N_4775,N_3790,N_4166);
and U4776 (N_4776,N_4180,N_3816);
nor U4777 (N_4777,N_4358,N_4141);
or U4778 (N_4778,N_3787,N_3878);
and U4779 (N_4779,N_4177,N_3918);
xnor U4780 (N_4780,N_3849,N_4134);
and U4781 (N_4781,N_4117,N_4146);
or U4782 (N_4782,N_4214,N_3940);
nor U4783 (N_4783,N_4333,N_4043);
nand U4784 (N_4784,N_4262,N_3804);
and U4785 (N_4785,N_3832,N_4161);
and U4786 (N_4786,N_4063,N_4126);
and U4787 (N_4787,N_4154,N_4113);
nor U4788 (N_4788,N_3939,N_3867);
and U4789 (N_4789,N_4347,N_3926);
and U4790 (N_4790,N_4299,N_4268);
and U4791 (N_4791,N_3907,N_4013);
or U4792 (N_4792,N_4007,N_3879);
or U4793 (N_4793,N_3796,N_4289);
nand U4794 (N_4794,N_4160,N_4336);
or U4795 (N_4795,N_4010,N_3999);
nor U4796 (N_4796,N_4031,N_3811);
xnor U4797 (N_4797,N_3779,N_4206);
nand U4798 (N_4798,N_4161,N_4240);
nor U4799 (N_4799,N_3800,N_4151);
nor U4800 (N_4800,N_3840,N_3921);
nor U4801 (N_4801,N_4320,N_4091);
and U4802 (N_4802,N_4046,N_4281);
and U4803 (N_4803,N_4240,N_4323);
and U4804 (N_4804,N_3807,N_4282);
xnor U4805 (N_4805,N_3820,N_4131);
nand U4806 (N_4806,N_4099,N_3941);
nor U4807 (N_4807,N_3854,N_4369);
and U4808 (N_4808,N_4053,N_4253);
xnor U4809 (N_4809,N_4207,N_4221);
xnor U4810 (N_4810,N_4246,N_3972);
xnor U4811 (N_4811,N_4029,N_3938);
and U4812 (N_4812,N_4334,N_3810);
xor U4813 (N_4813,N_4171,N_3956);
xnor U4814 (N_4814,N_4089,N_4311);
nand U4815 (N_4815,N_4372,N_4119);
nand U4816 (N_4816,N_3953,N_4031);
xnor U4817 (N_4817,N_4255,N_4203);
nor U4818 (N_4818,N_4121,N_3913);
and U4819 (N_4819,N_4313,N_4351);
xnor U4820 (N_4820,N_4373,N_3826);
nand U4821 (N_4821,N_4153,N_4198);
xor U4822 (N_4822,N_3894,N_4259);
or U4823 (N_4823,N_4159,N_4153);
and U4824 (N_4824,N_3810,N_4049);
nor U4825 (N_4825,N_3938,N_4239);
or U4826 (N_4826,N_4319,N_4217);
or U4827 (N_4827,N_3781,N_4304);
and U4828 (N_4828,N_4154,N_3872);
xor U4829 (N_4829,N_3999,N_3843);
nand U4830 (N_4830,N_3887,N_4078);
nand U4831 (N_4831,N_4361,N_4060);
and U4832 (N_4832,N_4184,N_3826);
nand U4833 (N_4833,N_4209,N_4174);
nor U4834 (N_4834,N_3836,N_4136);
nor U4835 (N_4835,N_3912,N_3985);
and U4836 (N_4836,N_4350,N_4344);
xnor U4837 (N_4837,N_4064,N_4332);
nand U4838 (N_4838,N_3752,N_3952);
and U4839 (N_4839,N_4277,N_4157);
or U4840 (N_4840,N_4003,N_3880);
or U4841 (N_4841,N_4231,N_3773);
xnor U4842 (N_4842,N_3760,N_4181);
and U4843 (N_4843,N_4056,N_3796);
xnor U4844 (N_4844,N_3810,N_3751);
xnor U4845 (N_4845,N_4182,N_4347);
xor U4846 (N_4846,N_4150,N_4090);
and U4847 (N_4847,N_4032,N_3758);
and U4848 (N_4848,N_3796,N_4263);
xnor U4849 (N_4849,N_4012,N_4069);
nor U4850 (N_4850,N_4119,N_3848);
nand U4851 (N_4851,N_3881,N_3863);
nor U4852 (N_4852,N_4214,N_3791);
nor U4853 (N_4853,N_4188,N_4241);
nor U4854 (N_4854,N_4206,N_4104);
nand U4855 (N_4855,N_3934,N_4150);
nand U4856 (N_4856,N_4170,N_4105);
or U4857 (N_4857,N_4057,N_4296);
xor U4858 (N_4858,N_4164,N_3922);
nand U4859 (N_4859,N_3782,N_3981);
xnor U4860 (N_4860,N_4089,N_4257);
xor U4861 (N_4861,N_4224,N_3830);
and U4862 (N_4862,N_4035,N_4081);
or U4863 (N_4863,N_4306,N_3957);
and U4864 (N_4864,N_4329,N_4155);
or U4865 (N_4865,N_4073,N_4251);
nand U4866 (N_4866,N_3960,N_4004);
nand U4867 (N_4867,N_4051,N_4117);
and U4868 (N_4868,N_3904,N_3979);
xnor U4869 (N_4869,N_3879,N_3906);
nor U4870 (N_4870,N_3944,N_4201);
or U4871 (N_4871,N_3904,N_4004);
nor U4872 (N_4872,N_4185,N_4370);
nor U4873 (N_4873,N_4312,N_3851);
nor U4874 (N_4874,N_3864,N_4210);
nand U4875 (N_4875,N_3840,N_4065);
xnor U4876 (N_4876,N_3852,N_3889);
xor U4877 (N_4877,N_3937,N_3871);
xor U4878 (N_4878,N_3966,N_4286);
nand U4879 (N_4879,N_4291,N_3889);
or U4880 (N_4880,N_4266,N_3787);
nand U4881 (N_4881,N_4233,N_3921);
or U4882 (N_4882,N_4078,N_4221);
xnor U4883 (N_4883,N_3864,N_4045);
nor U4884 (N_4884,N_4094,N_3879);
nor U4885 (N_4885,N_3918,N_4141);
or U4886 (N_4886,N_3885,N_3945);
nand U4887 (N_4887,N_3839,N_4295);
and U4888 (N_4888,N_3885,N_4290);
and U4889 (N_4889,N_3997,N_4113);
nand U4890 (N_4890,N_4258,N_3831);
nand U4891 (N_4891,N_4275,N_4054);
and U4892 (N_4892,N_4255,N_3905);
or U4893 (N_4893,N_4132,N_4133);
and U4894 (N_4894,N_4253,N_4236);
xnor U4895 (N_4895,N_4171,N_3823);
and U4896 (N_4896,N_3894,N_3791);
and U4897 (N_4897,N_4084,N_4032);
or U4898 (N_4898,N_4013,N_4012);
or U4899 (N_4899,N_4202,N_4229);
and U4900 (N_4900,N_3906,N_3776);
xnor U4901 (N_4901,N_4222,N_3833);
and U4902 (N_4902,N_4023,N_3846);
and U4903 (N_4903,N_4024,N_4229);
nand U4904 (N_4904,N_3762,N_4054);
nor U4905 (N_4905,N_4200,N_3989);
nor U4906 (N_4906,N_4117,N_3856);
nor U4907 (N_4907,N_3967,N_3845);
xor U4908 (N_4908,N_3890,N_3969);
nor U4909 (N_4909,N_3939,N_4216);
and U4910 (N_4910,N_3939,N_4223);
nand U4911 (N_4911,N_3972,N_3768);
or U4912 (N_4912,N_3755,N_4259);
or U4913 (N_4913,N_3880,N_3965);
or U4914 (N_4914,N_4208,N_4305);
xor U4915 (N_4915,N_3987,N_3841);
and U4916 (N_4916,N_3948,N_3994);
nand U4917 (N_4917,N_3856,N_4180);
and U4918 (N_4918,N_4315,N_4324);
xor U4919 (N_4919,N_4318,N_4072);
or U4920 (N_4920,N_4243,N_3819);
nor U4921 (N_4921,N_3762,N_4021);
or U4922 (N_4922,N_4121,N_4352);
nand U4923 (N_4923,N_3826,N_4151);
and U4924 (N_4924,N_4238,N_4051);
xnor U4925 (N_4925,N_4079,N_3919);
and U4926 (N_4926,N_4271,N_4326);
nand U4927 (N_4927,N_4300,N_4156);
nor U4928 (N_4928,N_4327,N_3825);
xnor U4929 (N_4929,N_3931,N_4193);
or U4930 (N_4930,N_4247,N_3834);
nand U4931 (N_4931,N_4328,N_3877);
or U4932 (N_4932,N_3769,N_3842);
and U4933 (N_4933,N_3911,N_4195);
xor U4934 (N_4934,N_3889,N_3821);
and U4935 (N_4935,N_4012,N_4121);
nand U4936 (N_4936,N_3797,N_4134);
and U4937 (N_4937,N_4019,N_4083);
and U4938 (N_4938,N_4215,N_3880);
nand U4939 (N_4939,N_4003,N_4247);
or U4940 (N_4940,N_4010,N_3769);
nand U4941 (N_4941,N_4263,N_4289);
or U4942 (N_4942,N_4352,N_4239);
nand U4943 (N_4943,N_4000,N_4019);
and U4944 (N_4944,N_4133,N_4059);
nor U4945 (N_4945,N_4147,N_4250);
nor U4946 (N_4946,N_4099,N_4308);
nor U4947 (N_4947,N_3794,N_4334);
nor U4948 (N_4948,N_3865,N_4280);
nor U4949 (N_4949,N_4315,N_4302);
nor U4950 (N_4950,N_3937,N_4209);
nor U4951 (N_4951,N_3844,N_3951);
and U4952 (N_4952,N_4218,N_3956);
xnor U4953 (N_4953,N_3832,N_3822);
nand U4954 (N_4954,N_3857,N_4334);
nand U4955 (N_4955,N_4258,N_4072);
and U4956 (N_4956,N_3839,N_4084);
nand U4957 (N_4957,N_3919,N_4145);
or U4958 (N_4958,N_3926,N_3982);
nor U4959 (N_4959,N_4105,N_4144);
and U4960 (N_4960,N_3786,N_3781);
or U4961 (N_4961,N_4122,N_3991);
nor U4962 (N_4962,N_4261,N_4346);
and U4963 (N_4963,N_3784,N_4254);
nor U4964 (N_4964,N_3927,N_3903);
or U4965 (N_4965,N_4223,N_3767);
nand U4966 (N_4966,N_4085,N_3856);
and U4967 (N_4967,N_3918,N_3903);
or U4968 (N_4968,N_3765,N_4289);
and U4969 (N_4969,N_4184,N_3918);
xnor U4970 (N_4970,N_4194,N_4122);
xnor U4971 (N_4971,N_4229,N_3773);
nor U4972 (N_4972,N_4064,N_4290);
or U4973 (N_4973,N_3922,N_3988);
or U4974 (N_4974,N_4128,N_3827);
and U4975 (N_4975,N_3803,N_3888);
nand U4976 (N_4976,N_4032,N_3985);
nor U4977 (N_4977,N_3776,N_4094);
and U4978 (N_4978,N_4105,N_3984);
nand U4979 (N_4979,N_3998,N_3896);
or U4980 (N_4980,N_4090,N_4064);
or U4981 (N_4981,N_4137,N_4108);
or U4982 (N_4982,N_4337,N_3813);
nor U4983 (N_4983,N_4224,N_3878);
and U4984 (N_4984,N_3986,N_4185);
nor U4985 (N_4985,N_4067,N_4113);
xor U4986 (N_4986,N_3939,N_4355);
or U4987 (N_4987,N_4240,N_4340);
nand U4988 (N_4988,N_3890,N_4223);
xnor U4989 (N_4989,N_4252,N_4003);
and U4990 (N_4990,N_4342,N_3819);
and U4991 (N_4991,N_4359,N_4068);
nor U4992 (N_4992,N_3781,N_4332);
nor U4993 (N_4993,N_3966,N_4303);
nand U4994 (N_4994,N_3949,N_4145);
and U4995 (N_4995,N_3979,N_4049);
or U4996 (N_4996,N_4092,N_3902);
or U4997 (N_4997,N_3997,N_4299);
and U4998 (N_4998,N_4261,N_4071);
nor U4999 (N_4999,N_4293,N_3888);
nor U5000 (N_5000,N_4817,N_4636);
nor U5001 (N_5001,N_4395,N_4989);
xnor U5002 (N_5002,N_4597,N_4965);
xnor U5003 (N_5003,N_4766,N_4957);
or U5004 (N_5004,N_4670,N_4833);
or U5005 (N_5005,N_4708,N_4583);
nand U5006 (N_5006,N_4585,N_4401);
and U5007 (N_5007,N_4468,N_4623);
nor U5008 (N_5008,N_4855,N_4629);
nor U5009 (N_5009,N_4725,N_4621);
and U5010 (N_5010,N_4896,N_4776);
or U5011 (N_5011,N_4720,N_4757);
xor U5012 (N_5012,N_4609,N_4922);
nand U5013 (N_5013,N_4536,N_4642);
and U5014 (N_5014,N_4506,N_4400);
and U5015 (N_5015,N_4494,N_4984);
xor U5016 (N_5016,N_4594,N_4836);
and U5017 (N_5017,N_4414,N_4684);
xnor U5018 (N_5018,N_4691,N_4527);
or U5019 (N_5019,N_4813,N_4412);
nand U5020 (N_5020,N_4473,N_4688);
or U5021 (N_5021,N_4744,N_4978);
nor U5022 (N_5022,N_4849,N_4971);
xor U5023 (N_5023,N_4674,N_4445);
nand U5024 (N_5024,N_4552,N_4747);
xnor U5025 (N_5025,N_4694,N_4808);
xnor U5026 (N_5026,N_4386,N_4469);
or U5027 (N_5027,N_4596,N_4668);
nand U5028 (N_5028,N_4772,N_4475);
nor U5029 (N_5029,N_4943,N_4441);
or U5030 (N_5030,N_4826,N_4915);
or U5031 (N_5031,N_4431,N_4570);
xnor U5032 (N_5032,N_4900,N_4483);
nor U5033 (N_5033,N_4793,N_4550);
xnor U5034 (N_5034,N_4759,N_4852);
nor U5035 (N_5035,N_4589,N_4437);
xor U5036 (N_5036,N_4860,N_4798);
and U5037 (N_5037,N_4937,N_4549);
xor U5038 (N_5038,N_4819,N_4880);
xor U5039 (N_5039,N_4627,N_4731);
and U5040 (N_5040,N_4985,N_4661);
or U5041 (N_5041,N_4887,N_4663);
or U5042 (N_5042,N_4422,N_4418);
nand U5043 (N_5043,N_4804,N_4940);
nor U5044 (N_5044,N_4909,N_4561);
xor U5045 (N_5045,N_4548,N_4509);
and U5046 (N_5046,N_4812,N_4498);
and U5047 (N_5047,N_4396,N_4917);
and U5048 (N_5048,N_4768,N_4814);
or U5049 (N_5049,N_4767,N_4873);
nor U5050 (N_5050,N_4877,N_4902);
xor U5051 (N_5051,N_4955,N_4925);
and U5052 (N_5052,N_4695,N_4683);
or U5053 (N_5053,N_4923,N_4921);
and U5054 (N_5054,N_4635,N_4480);
xor U5055 (N_5055,N_4500,N_4894);
nand U5056 (N_5056,N_4547,N_4779);
xor U5057 (N_5057,N_4998,N_4610);
and U5058 (N_5058,N_4775,N_4493);
nand U5059 (N_5059,N_4528,N_4736);
nor U5060 (N_5060,N_4618,N_4903);
and U5061 (N_5061,N_4600,N_4620);
nand U5062 (N_5062,N_4639,N_4750);
and U5063 (N_5063,N_4944,N_4789);
nor U5064 (N_5064,N_4898,N_4869);
nor U5065 (N_5065,N_4387,N_4686);
or U5066 (N_5066,N_4790,N_4444);
nand U5067 (N_5067,N_4490,N_4477);
xnor U5068 (N_5068,N_4861,N_4999);
nand U5069 (N_5069,N_4590,N_4533);
or U5070 (N_5070,N_4541,N_4572);
nor U5071 (N_5071,N_4384,N_4435);
or U5072 (N_5072,N_4728,N_4713);
nand U5073 (N_5073,N_4593,N_4739);
nor U5074 (N_5074,N_4843,N_4946);
nor U5075 (N_5075,N_4993,N_4913);
nand U5076 (N_5076,N_4613,N_4931);
nor U5077 (N_5077,N_4619,N_4914);
nand U5078 (N_5078,N_4941,N_4862);
or U5079 (N_5079,N_4390,N_4553);
nand U5080 (N_5080,N_4377,N_4942);
and U5081 (N_5081,N_4632,N_4979);
nand U5082 (N_5082,N_4425,N_4457);
or U5083 (N_5083,N_4587,N_4936);
nor U5084 (N_5084,N_4835,N_4781);
and U5085 (N_5085,N_4696,N_4465);
and U5086 (N_5086,N_4823,N_4928);
nor U5087 (N_5087,N_4563,N_4889);
xnor U5088 (N_5088,N_4950,N_4973);
or U5089 (N_5089,N_4540,N_4727);
and U5090 (N_5090,N_4774,N_4615);
or U5091 (N_5091,N_4487,N_4641);
xnor U5092 (N_5092,N_4910,N_4565);
xnor U5093 (N_5093,N_4482,N_4901);
nand U5094 (N_5094,N_4949,N_4994);
nand U5095 (N_5095,N_4771,N_4741);
and U5096 (N_5096,N_4648,N_4452);
nor U5097 (N_5097,N_4612,N_4983);
nand U5098 (N_5098,N_4375,N_4522);
and U5099 (N_5099,N_4420,N_4970);
nor U5100 (N_5100,N_4885,N_4962);
nor U5101 (N_5101,N_4729,N_4893);
or U5102 (N_5102,N_4640,N_4968);
or U5103 (N_5103,N_4464,N_4599);
xor U5104 (N_5104,N_4568,N_4912);
or U5105 (N_5105,N_4508,N_4748);
xnor U5106 (N_5106,N_4433,N_4577);
nand U5107 (N_5107,N_4758,N_4625);
and U5108 (N_5108,N_4530,N_4899);
xnor U5109 (N_5109,N_4669,N_4637);
nand U5110 (N_5110,N_4542,N_4388);
nand U5111 (N_5111,N_4537,N_4831);
or U5112 (N_5112,N_4996,N_4918);
nor U5113 (N_5113,N_4939,N_4408);
nand U5114 (N_5114,N_4990,N_4700);
nand U5115 (N_5115,N_4959,N_4545);
and U5116 (N_5116,N_4461,N_4822);
xor U5117 (N_5117,N_4491,N_4709);
nand U5118 (N_5118,N_4643,N_4379);
nand U5119 (N_5119,N_4551,N_4672);
or U5120 (N_5120,N_4692,N_4543);
nand U5121 (N_5121,N_4714,N_4966);
or U5122 (N_5122,N_4829,N_4956);
nand U5123 (N_5123,N_4484,N_4850);
nand U5124 (N_5124,N_4571,N_4438);
nor U5125 (N_5125,N_4876,N_4719);
or U5126 (N_5126,N_4389,N_4488);
nor U5127 (N_5127,N_4821,N_4449);
xnor U5128 (N_5128,N_4846,N_4559);
nor U5129 (N_5129,N_4872,N_4825);
or U5130 (N_5130,N_4578,N_4690);
xnor U5131 (N_5131,N_4385,N_4888);
nand U5132 (N_5132,N_4398,N_4754);
or U5133 (N_5133,N_4782,N_4424);
and U5134 (N_5134,N_4534,N_4702);
or U5135 (N_5135,N_4497,N_4697);
nor U5136 (N_5136,N_4864,N_4575);
or U5137 (N_5137,N_4574,N_4626);
nor U5138 (N_5138,N_4582,N_4809);
nand U5139 (N_5139,N_4410,N_4638);
nand U5140 (N_5140,N_4718,N_4448);
xnor U5141 (N_5141,N_4785,N_4816);
nor U5142 (N_5142,N_4988,N_4603);
nand U5143 (N_5143,N_4791,N_4611);
and U5144 (N_5144,N_4751,N_4908);
nand U5145 (N_5145,N_4711,N_4838);
nand U5146 (N_5146,N_4505,N_4411);
or U5147 (N_5147,N_4832,N_4980);
or U5148 (N_5148,N_4617,N_4556);
or U5149 (N_5149,N_4870,N_4932);
or U5150 (N_5150,N_4586,N_4907);
nand U5151 (N_5151,N_4397,N_4967);
or U5152 (N_5152,N_4800,N_4780);
or U5153 (N_5153,N_4515,N_4476);
nor U5154 (N_5154,N_4777,N_4699);
and U5155 (N_5155,N_4704,N_4830);
and U5156 (N_5156,N_4453,N_4976);
nand U5157 (N_5157,N_4404,N_4419);
nand U5158 (N_5158,N_4882,N_4981);
nor U5159 (N_5159,N_4646,N_4383);
or U5160 (N_5160,N_4847,N_4681);
nor U5161 (N_5161,N_4992,N_4742);
nor U5162 (N_5162,N_4687,N_4558);
nor U5163 (N_5163,N_4701,N_4502);
xnor U5164 (N_5164,N_4824,N_4656);
or U5165 (N_5165,N_4698,N_4724);
xnor U5166 (N_5166,N_4975,N_4666);
xor U5167 (N_5167,N_4866,N_4733);
or U5168 (N_5168,N_4455,N_4394);
and U5169 (N_5169,N_4529,N_4693);
or U5170 (N_5170,N_4730,N_4952);
and U5171 (N_5171,N_4763,N_4427);
xor U5172 (N_5172,N_4446,N_4470);
nand U5173 (N_5173,N_4871,N_4749);
nor U5174 (N_5174,N_4562,N_4512);
nor U5175 (N_5175,N_4517,N_4428);
or U5176 (N_5176,N_4972,N_4659);
nor U5177 (N_5177,N_4647,N_4867);
xnor U5178 (N_5178,N_4839,N_4507);
or U5179 (N_5179,N_4991,N_4679);
nor U5180 (N_5180,N_4525,N_4521);
nand U5181 (N_5181,N_4716,N_4503);
or U5182 (N_5182,N_4710,N_4868);
xor U5183 (N_5183,N_4454,N_4496);
nand U5184 (N_5184,N_4891,N_4608);
and U5185 (N_5185,N_4840,N_4706);
nor U5186 (N_5186,N_4649,N_4426);
or U5187 (N_5187,N_4675,N_4924);
nor U5188 (N_5188,N_4634,N_4853);
nor U5189 (N_5189,N_4795,N_4818);
and U5190 (N_5190,N_4930,N_4462);
nor U5191 (N_5191,N_4986,N_4409);
nand U5192 (N_5192,N_4858,N_4654);
or U5193 (N_5193,N_4606,N_4743);
nor U5194 (N_5194,N_4598,N_4566);
and U5195 (N_5195,N_4671,N_4665);
and U5196 (N_5196,N_4960,N_4844);
or U5197 (N_5197,N_4653,N_4879);
and U5198 (N_5198,N_4805,N_4680);
nand U5199 (N_5199,N_4514,N_4682);
nor U5200 (N_5200,N_4841,N_4874);
xor U5201 (N_5201,N_4532,N_4450);
nand U5202 (N_5202,N_4953,N_4756);
and U5203 (N_5203,N_4746,N_4581);
xnor U5204 (N_5204,N_4792,N_4467);
and U5205 (N_5205,N_4905,N_4784);
nor U5206 (N_5206,N_4616,N_4633);
or U5207 (N_5207,N_4655,N_4740);
nand U5208 (N_5208,N_4607,N_4745);
or U5209 (N_5209,N_4604,N_4723);
nor U5210 (N_5210,N_4519,N_4510);
xnor U5211 (N_5211,N_4715,N_4660);
or U5212 (N_5212,N_4883,N_4753);
and U5213 (N_5213,N_4624,N_4391);
xor U5214 (N_5214,N_4834,N_4760);
nor U5215 (N_5215,N_4657,N_4458);
nor U5216 (N_5216,N_4752,N_4995);
nor U5217 (N_5217,N_4828,N_4544);
and U5218 (N_5218,N_4920,N_4897);
nor U5219 (N_5219,N_4380,N_4938);
and U5220 (N_5220,N_4429,N_4906);
xnor U5221 (N_5221,N_4851,N_4630);
and U5222 (N_5222,N_4765,N_4837);
nand U5223 (N_5223,N_4778,N_4678);
xor U5224 (N_5224,N_4403,N_4459);
xnor U5225 (N_5225,N_4531,N_4685);
xnor U5226 (N_5226,N_4854,N_4886);
or U5227 (N_5227,N_4423,N_4602);
nor U5228 (N_5228,N_4413,N_4927);
nand U5229 (N_5229,N_4788,N_4492);
and U5230 (N_5230,N_4722,N_4416);
nand U5231 (N_5231,N_4584,N_4667);
xnor U5232 (N_5232,N_4764,N_4463);
nor U5233 (N_5233,N_4875,N_4474);
or U5234 (N_5234,N_4399,N_4878);
nor U5235 (N_5235,N_4721,N_4555);
nand U5236 (N_5236,N_4755,N_4436);
nor U5237 (N_5237,N_4762,N_4689);
nand U5238 (N_5238,N_4892,N_4554);
or U5239 (N_5239,N_4523,N_4734);
nor U5240 (N_5240,N_4485,N_4948);
nor U5241 (N_5241,N_4895,N_4859);
nor U5242 (N_5242,N_4439,N_4863);
xor U5243 (N_5243,N_4479,N_4430);
nand U5244 (N_5244,N_4732,N_4472);
nand U5245 (N_5245,N_4890,N_4440);
or U5246 (N_5246,N_4415,N_4803);
nor U5247 (N_5247,N_4707,N_4495);
nor U5248 (N_5248,N_4443,N_4567);
nand U5249 (N_5249,N_4802,N_4478);
and U5250 (N_5250,N_4934,N_4376);
and U5251 (N_5251,N_4576,N_4539);
xor U5252 (N_5252,N_4442,N_4964);
xor U5253 (N_5253,N_4499,N_4884);
and U5254 (N_5254,N_4526,N_4622);
or U5255 (N_5255,N_4588,N_4865);
and U5256 (N_5256,N_4974,N_4712);
nand U5257 (N_5257,N_4489,N_4511);
or U5258 (N_5258,N_4662,N_4518);
nand U5259 (N_5259,N_4857,N_4773);
nor U5260 (N_5260,N_4579,N_4806);
nor U5261 (N_5261,N_4726,N_4848);
nor U5262 (N_5262,N_4947,N_4796);
xnor U5263 (N_5263,N_4801,N_4392);
and U5264 (N_5264,N_4538,N_4516);
and U5265 (N_5265,N_4969,N_4378);
or U5266 (N_5266,N_4820,N_4770);
xor U5267 (N_5267,N_4651,N_4845);
and U5268 (N_5268,N_4735,N_4504);
or U5269 (N_5269,N_4569,N_4524);
and U5270 (N_5270,N_4811,N_4520);
and U5271 (N_5271,N_4807,N_4580);
nor U5272 (N_5272,N_4881,N_4460);
and U5273 (N_5273,N_4573,N_4402);
nor U5274 (N_5274,N_4393,N_4977);
xnor U5275 (N_5275,N_4560,N_4815);
nand U5276 (N_5276,N_4787,N_4447);
nand U5277 (N_5277,N_4929,N_4381);
nor U5278 (N_5278,N_4595,N_4513);
xnor U5279 (N_5279,N_4631,N_4963);
nand U5280 (N_5280,N_4456,N_4958);
nand U5281 (N_5281,N_4933,N_4501);
nand U5282 (N_5282,N_4961,N_4451);
xor U5283 (N_5283,N_4856,N_4591);
nor U5284 (N_5284,N_4557,N_4601);
and U5285 (N_5285,N_4405,N_4904);
or U5286 (N_5286,N_4650,N_4919);
nand U5287 (N_5287,N_4481,N_4794);
or U5288 (N_5288,N_4717,N_4644);
or U5289 (N_5289,N_4676,N_4738);
nand U5290 (N_5290,N_4471,N_4592);
nor U5291 (N_5291,N_4466,N_4926);
nor U5292 (N_5292,N_4769,N_4421);
nor U5293 (N_5293,N_4673,N_4614);
nor U5294 (N_5294,N_4783,N_4786);
nand U5295 (N_5295,N_4382,N_4703);
nor U5296 (N_5296,N_4705,N_4417);
nor U5297 (N_5297,N_4799,N_4546);
and U5298 (N_5298,N_4564,N_4842);
xor U5299 (N_5299,N_4997,N_4737);
and U5300 (N_5300,N_4664,N_4652);
xnor U5301 (N_5301,N_4987,N_4982);
xor U5302 (N_5302,N_4677,N_4797);
or U5303 (N_5303,N_4911,N_4407);
or U5304 (N_5304,N_4628,N_4954);
and U5305 (N_5305,N_4935,N_4951);
or U5306 (N_5306,N_4761,N_4605);
or U5307 (N_5307,N_4916,N_4432);
xor U5308 (N_5308,N_4406,N_4535);
nand U5309 (N_5309,N_4945,N_4434);
nand U5310 (N_5310,N_4827,N_4645);
nor U5311 (N_5311,N_4486,N_4658);
or U5312 (N_5312,N_4810,N_4407);
nor U5313 (N_5313,N_4770,N_4666);
and U5314 (N_5314,N_4412,N_4674);
and U5315 (N_5315,N_4573,N_4842);
or U5316 (N_5316,N_4455,N_4811);
or U5317 (N_5317,N_4681,N_4843);
nand U5318 (N_5318,N_4451,N_4996);
or U5319 (N_5319,N_4616,N_4718);
or U5320 (N_5320,N_4437,N_4950);
or U5321 (N_5321,N_4974,N_4836);
and U5322 (N_5322,N_4396,N_4646);
or U5323 (N_5323,N_4842,N_4506);
nor U5324 (N_5324,N_4555,N_4930);
and U5325 (N_5325,N_4510,N_4593);
nor U5326 (N_5326,N_4494,N_4543);
and U5327 (N_5327,N_4958,N_4498);
nand U5328 (N_5328,N_4523,N_4949);
or U5329 (N_5329,N_4460,N_4759);
xnor U5330 (N_5330,N_4677,N_4739);
nor U5331 (N_5331,N_4794,N_4665);
nor U5332 (N_5332,N_4870,N_4786);
xnor U5333 (N_5333,N_4466,N_4984);
nor U5334 (N_5334,N_4828,N_4712);
nand U5335 (N_5335,N_4428,N_4750);
xor U5336 (N_5336,N_4667,N_4717);
xor U5337 (N_5337,N_4511,N_4833);
or U5338 (N_5338,N_4631,N_4889);
nor U5339 (N_5339,N_4733,N_4605);
nor U5340 (N_5340,N_4966,N_4565);
nand U5341 (N_5341,N_4527,N_4465);
nor U5342 (N_5342,N_4872,N_4561);
xor U5343 (N_5343,N_4714,N_4893);
and U5344 (N_5344,N_4545,N_4806);
nor U5345 (N_5345,N_4564,N_4925);
nand U5346 (N_5346,N_4465,N_4415);
or U5347 (N_5347,N_4562,N_4685);
xor U5348 (N_5348,N_4760,N_4780);
nand U5349 (N_5349,N_4826,N_4426);
xor U5350 (N_5350,N_4524,N_4970);
nand U5351 (N_5351,N_4731,N_4658);
xnor U5352 (N_5352,N_4502,N_4908);
nand U5353 (N_5353,N_4600,N_4881);
xnor U5354 (N_5354,N_4676,N_4503);
nor U5355 (N_5355,N_4628,N_4973);
or U5356 (N_5356,N_4927,N_4645);
or U5357 (N_5357,N_4385,N_4584);
and U5358 (N_5358,N_4561,N_4955);
and U5359 (N_5359,N_4610,N_4409);
nor U5360 (N_5360,N_4678,N_4562);
and U5361 (N_5361,N_4886,N_4792);
xor U5362 (N_5362,N_4829,N_4820);
xor U5363 (N_5363,N_4790,N_4746);
xnor U5364 (N_5364,N_4743,N_4479);
and U5365 (N_5365,N_4789,N_4475);
and U5366 (N_5366,N_4952,N_4551);
or U5367 (N_5367,N_4983,N_4771);
nor U5368 (N_5368,N_4499,N_4921);
nor U5369 (N_5369,N_4432,N_4555);
nand U5370 (N_5370,N_4745,N_4866);
nand U5371 (N_5371,N_4585,N_4745);
xor U5372 (N_5372,N_4541,N_4524);
and U5373 (N_5373,N_4458,N_4876);
and U5374 (N_5374,N_4678,N_4843);
or U5375 (N_5375,N_4837,N_4656);
or U5376 (N_5376,N_4513,N_4729);
or U5377 (N_5377,N_4886,N_4734);
and U5378 (N_5378,N_4458,N_4440);
nor U5379 (N_5379,N_4844,N_4490);
xnor U5380 (N_5380,N_4960,N_4984);
xor U5381 (N_5381,N_4487,N_4407);
nor U5382 (N_5382,N_4456,N_4655);
and U5383 (N_5383,N_4459,N_4775);
xnor U5384 (N_5384,N_4520,N_4720);
nor U5385 (N_5385,N_4694,N_4834);
nor U5386 (N_5386,N_4574,N_4489);
or U5387 (N_5387,N_4724,N_4818);
nand U5388 (N_5388,N_4637,N_4537);
xor U5389 (N_5389,N_4502,N_4919);
nand U5390 (N_5390,N_4405,N_4532);
and U5391 (N_5391,N_4957,N_4735);
or U5392 (N_5392,N_4939,N_4511);
nor U5393 (N_5393,N_4624,N_4817);
and U5394 (N_5394,N_4680,N_4440);
and U5395 (N_5395,N_4598,N_4915);
or U5396 (N_5396,N_4526,N_4743);
or U5397 (N_5397,N_4984,N_4470);
nand U5398 (N_5398,N_4677,N_4524);
and U5399 (N_5399,N_4766,N_4543);
nand U5400 (N_5400,N_4464,N_4527);
nand U5401 (N_5401,N_4646,N_4612);
nand U5402 (N_5402,N_4805,N_4511);
nor U5403 (N_5403,N_4902,N_4760);
xor U5404 (N_5404,N_4473,N_4784);
and U5405 (N_5405,N_4737,N_4780);
or U5406 (N_5406,N_4725,N_4867);
nand U5407 (N_5407,N_4768,N_4540);
nand U5408 (N_5408,N_4808,N_4397);
or U5409 (N_5409,N_4717,N_4804);
and U5410 (N_5410,N_4573,N_4820);
xor U5411 (N_5411,N_4821,N_4561);
or U5412 (N_5412,N_4501,N_4924);
nor U5413 (N_5413,N_4500,N_4595);
xnor U5414 (N_5414,N_4671,N_4438);
nand U5415 (N_5415,N_4878,N_4720);
and U5416 (N_5416,N_4858,N_4394);
nor U5417 (N_5417,N_4521,N_4457);
nand U5418 (N_5418,N_4461,N_4672);
nand U5419 (N_5419,N_4961,N_4968);
nand U5420 (N_5420,N_4951,N_4633);
or U5421 (N_5421,N_4811,N_4944);
xor U5422 (N_5422,N_4921,N_4612);
and U5423 (N_5423,N_4987,N_4888);
nand U5424 (N_5424,N_4964,N_4921);
nor U5425 (N_5425,N_4378,N_4815);
nor U5426 (N_5426,N_4755,N_4771);
or U5427 (N_5427,N_4795,N_4946);
nand U5428 (N_5428,N_4456,N_4781);
nor U5429 (N_5429,N_4766,N_4616);
or U5430 (N_5430,N_4457,N_4706);
and U5431 (N_5431,N_4814,N_4482);
nand U5432 (N_5432,N_4867,N_4780);
nand U5433 (N_5433,N_4552,N_4825);
nor U5434 (N_5434,N_4731,N_4602);
or U5435 (N_5435,N_4787,N_4398);
nand U5436 (N_5436,N_4891,N_4887);
nor U5437 (N_5437,N_4557,N_4597);
or U5438 (N_5438,N_4628,N_4885);
or U5439 (N_5439,N_4630,N_4762);
nor U5440 (N_5440,N_4839,N_4973);
nand U5441 (N_5441,N_4415,N_4933);
xor U5442 (N_5442,N_4556,N_4809);
xor U5443 (N_5443,N_4412,N_4835);
nor U5444 (N_5444,N_4824,N_4862);
and U5445 (N_5445,N_4910,N_4748);
xnor U5446 (N_5446,N_4989,N_4579);
xor U5447 (N_5447,N_4837,N_4914);
and U5448 (N_5448,N_4877,N_4862);
and U5449 (N_5449,N_4513,N_4705);
or U5450 (N_5450,N_4637,N_4643);
or U5451 (N_5451,N_4894,N_4724);
or U5452 (N_5452,N_4622,N_4418);
xnor U5453 (N_5453,N_4560,N_4770);
nand U5454 (N_5454,N_4721,N_4611);
xnor U5455 (N_5455,N_4957,N_4732);
xnor U5456 (N_5456,N_4970,N_4402);
nor U5457 (N_5457,N_4530,N_4464);
xnor U5458 (N_5458,N_4656,N_4937);
and U5459 (N_5459,N_4476,N_4545);
nor U5460 (N_5460,N_4829,N_4594);
nand U5461 (N_5461,N_4406,N_4548);
or U5462 (N_5462,N_4948,N_4911);
or U5463 (N_5463,N_4414,N_4524);
or U5464 (N_5464,N_4950,N_4668);
or U5465 (N_5465,N_4501,N_4643);
nor U5466 (N_5466,N_4962,N_4896);
nor U5467 (N_5467,N_4488,N_4948);
or U5468 (N_5468,N_4901,N_4725);
nand U5469 (N_5469,N_4950,N_4454);
or U5470 (N_5470,N_4540,N_4861);
and U5471 (N_5471,N_4891,N_4927);
nand U5472 (N_5472,N_4507,N_4673);
or U5473 (N_5473,N_4674,N_4679);
nor U5474 (N_5474,N_4479,N_4863);
nor U5475 (N_5475,N_4955,N_4418);
nand U5476 (N_5476,N_4691,N_4950);
nor U5477 (N_5477,N_4436,N_4932);
nand U5478 (N_5478,N_4899,N_4770);
xnor U5479 (N_5479,N_4454,N_4860);
xor U5480 (N_5480,N_4655,N_4499);
xnor U5481 (N_5481,N_4954,N_4493);
nand U5482 (N_5482,N_4822,N_4538);
or U5483 (N_5483,N_4387,N_4734);
and U5484 (N_5484,N_4815,N_4671);
nor U5485 (N_5485,N_4931,N_4974);
nor U5486 (N_5486,N_4516,N_4735);
and U5487 (N_5487,N_4375,N_4533);
xor U5488 (N_5488,N_4730,N_4910);
and U5489 (N_5489,N_4987,N_4411);
xnor U5490 (N_5490,N_4419,N_4521);
nand U5491 (N_5491,N_4740,N_4648);
or U5492 (N_5492,N_4460,N_4604);
nand U5493 (N_5493,N_4961,N_4802);
nand U5494 (N_5494,N_4480,N_4986);
xnor U5495 (N_5495,N_4930,N_4785);
or U5496 (N_5496,N_4438,N_4940);
and U5497 (N_5497,N_4589,N_4381);
xnor U5498 (N_5498,N_4821,N_4555);
nand U5499 (N_5499,N_4430,N_4580);
xor U5500 (N_5500,N_4783,N_4713);
nor U5501 (N_5501,N_4956,N_4849);
or U5502 (N_5502,N_4979,N_4722);
or U5503 (N_5503,N_4467,N_4869);
nand U5504 (N_5504,N_4764,N_4667);
nor U5505 (N_5505,N_4490,N_4744);
xor U5506 (N_5506,N_4810,N_4880);
and U5507 (N_5507,N_4683,N_4523);
nand U5508 (N_5508,N_4825,N_4990);
and U5509 (N_5509,N_4688,N_4474);
xor U5510 (N_5510,N_4458,N_4576);
nand U5511 (N_5511,N_4492,N_4560);
nor U5512 (N_5512,N_4522,N_4944);
nor U5513 (N_5513,N_4411,N_4891);
or U5514 (N_5514,N_4611,N_4399);
xnor U5515 (N_5515,N_4498,N_4983);
nor U5516 (N_5516,N_4671,N_4854);
nor U5517 (N_5517,N_4758,N_4832);
or U5518 (N_5518,N_4681,N_4863);
nor U5519 (N_5519,N_4794,N_4844);
or U5520 (N_5520,N_4653,N_4945);
nor U5521 (N_5521,N_4478,N_4897);
nor U5522 (N_5522,N_4602,N_4966);
and U5523 (N_5523,N_4730,N_4630);
or U5524 (N_5524,N_4677,N_4586);
nand U5525 (N_5525,N_4806,N_4695);
nand U5526 (N_5526,N_4873,N_4695);
and U5527 (N_5527,N_4497,N_4946);
xnor U5528 (N_5528,N_4460,N_4867);
xnor U5529 (N_5529,N_4745,N_4698);
and U5530 (N_5530,N_4605,N_4497);
xnor U5531 (N_5531,N_4805,N_4825);
and U5532 (N_5532,N_4689,N_4754);
nor U5533 (N_5533,N_4471,N_4541);
or U5534 (N_5534,N_4408,N_4451);
or U5535 (N_5535,N_4631,N_4608);
nor U5536 (N_5536,N_4894,N_4631);
and U5537 (N_5537,N_4821,N_4629);
nand U5538 (N_5538,N_4857,N_4466);
or U5539 (N_5539,N_4874,N_4537);
and U5540 (N_5540,N_4382,N_4815);
nor U5541 (N_5541,N_4941,N_4810);
nand U5542 (N_5542,N_4992,N_4870);
nor U5543 (N_5543,N_4498,N_4707);
xnor U5544 (N_5544,N_4447,N_4605);
and U5545 (N_5545,N_4882,N_4523);
or U5546 (N_5546,N_4661,N_4569);
and U5547 (N_5547,N_4906,N_4673);
nand U5548 (N_5548,N_4830,N_4739);
or U5549 (N_5549,N_4691,N_4941);
xor U5550 (N_5550,N_4974,N_4532);
xor U5551 (N_5551,N_4396,N_4753);
nor U5552 (N_5552,N_4823,N_4875);
nor U5553 (N_5553,N_4512,N_4419);
and U5554 (N_5554,N_4754,N_4777);
xor U5555 (N_5555,N_4894,N_4924);
nor U5556 (N_5556,N_4678,N_4810);
xor U5557 (N_5557,N_4765,N_4614);
nand U5558 (N_5558,N_4649,N_4942);
nor U5559 (N_5559,N_4710,N_4574);
nor U5560 (N_5560,N_4550,N_4667);
nor U5561 (N_5561,N_4861,N_4772);
xnor U5562 (N_5562,N_4859,N_4887);
and U5563 (N_5563,N_4860,N_4886);
xnor U5564 (N_5564,N_4459,N_4409);
or U5565 (N_5565,N_4421,N_4649);
nand U5566 (N_5566,N_4646,N_4402);
and U5567 (N_5567,N_4771,N_4394);
nor U5568 (N_5568,N_4664,N_4942);
nor U5569 (N_5569,N_4907,N_4855);
nand U5570 (N_5570,N_4519,N_4412);
or U5571 (N_5571,N_4555,N_4403);
or U5572 (N_5572,N_4828,N_4982);
and U5573 (N_5573,N_4464,N_4655);
nor U5574 (N_5574,N_4581,N_4534);
and U5575 (N_5575,N_4777,N_4955);
xor U5576 (N_5576,N_4701,N_4715);
nand U5577 (N_5577,N_4891,N_4458);
nor U5578 (N_5578,N_4558,N_4581);
and U5579 (N_5579,N_4430,N_4699);
nand U5580 (N_5580,N_4575,N_4515);
or U5581 (N_5581,N_4584,N_4767);
and U5582 (N_5582,N_4879,N_4779);
nand U5583 (N_5583,N_4724,N_4759);
or U5584 (N_5584,N_4747,N_4516);
or U5585 (N_5585,N_4453,N_4985);
xnor U5586 (N_5586,N_4405,N_4670);
xor U5587 (N_5587,N_4929,N_4411);
or U5588 (N_5588,N_4975,N_4430);
xnor U5589 (N_5589,N_4967,N_4676);
nand U5590 (N_5590,N_4495,N_4570);
nor U5591 (N_5591,N_4649,N_4776);
or U5592 (N_5592,N_4854,N_4856);
or U5593 (N_5593,N_4812,N_4486);
or U5594 (N_5594,N_4782,N_4571);
and U5595 (N_5595,N_4931,N_4493);
nor U5596 (N_5596,N_4880,N_4545);
or U5597 (N_5597,N_4675,N_4912);
or U5598 (N_5598,N_4564,N_4424);
xnor U5599 (N_5599,N_4644,N_4721);
nor U5600 (N_5600,N_4894,N_4527);
xnor U5601 (N_5601,N_4446,N_4849);
or U5602 (N_5602,N_4657,N_4453);
nor U5603 (N_5603,N_4509,N_4698);
nand U5604 (N_5604,N_4737,N_4718);
nand U5605 (N_5605,N_4458,N_4725);
or U5606 (N_5606,N_4803,N_4858);
nand U5607 (N_5607,N_4714,N_4540);
or U5608 (N_5608,N_4769,N_4818);
nor U5609 (N_5609,N_4902,N_4436);
nand U5610 (N_5610,N_4869,N_4466);
or U5611 (N_5611,N_4996,N_4861);
nand U5612 (N_5612,N_4948,N_4960);
nor U5613 (N_5613,N_4776,N_4766);
xnor U5614 (N_5614,N_4417,N_4750);
nand U5615 (N_5615,N_4545,N_4713);
or U5616 (N_5616,N_4778,N_4542);
nor U5617 (N_5617,N_4907,N_4641);
and U5618 (N_5618,N_4833,N_4939);
and U5619 (N_5619,N_4467,N_4460);
or U5620 (N_5620,N_4981,N_4690);
nor U5621 (N_5621,N_4426,N_4914);
nand U5622 (N_5622,N_4746,N_4813);
and U5623 (N_5623,N_4891,N_4823);
or U5624 (N_5624,N_4934,N_4573);
or U5625 (N_5625,N_5317,N_5063);
or U5626 (N_5626,N_5068,N_5495);
xor U5627 (N_5627,N_5203,N_5428);
or U5628 (N_5628,N_5041,N_5486);
or U5629 (N_5629,N_5544,N_5419);
and U5630 (N_5630,N_5248,N_5366);
nand U5631 (N_5631,N_5214,N_5226);
xor U5632 (N_5632,N_5255,N_5208);
and U5633 (N_5633,N_5001,N_5605);
and U5634 (N_5634,N_5302,N_5073);
and U5635 (N_5635,N_5092,N_5039);
and U5636 (N_5636,N_5450,N_5612);
nor U5637 (N_5637,N_5078,N_5115);
nand U5638 (N_5638,N_5426,N_5123);
and U5639 (N_5639,N_5021,N_5119);
nand U5640 (N_5640,N_5615,N_5326);
xnor U5641 (N_5641,N_5154,N_5582);
nand U5642 (N_5642,N_5029,N_5146);
and U5643 (N_5643,N_5310,N_5571);
nor U5644 (N_5644,N_5246,N_5179);
and U5645 (N_5645,N_5237,N_5077);
and U5646 (N_5646,N_5249,N_5431);
nand U5647 (N_5647,N_5169,N_5409);
nand U5648 (N_5648,N_5532,N_5329);
and U5649 (N_5649,N_5555,N_5177);
or U5650 (N_5650,N_5332,N_5057);
xnor U5651 (N_5651,N_5480,N_5309);
nand U5652 (N_5652,N_5586,N_5066);
nor U5653 (N_5653,N_5053,N_5090);
nand U5654 (N_5654,N_5410,N_5412);
and U5655 (N_5655,N_5254,N_5566);
or U5656 (N_5656,N_5405,N_5079);
or U5657 (N_5657,N_5181,N_5100);
or U5658 (N_5658,N_5272,N_5402);
xnor U5659 (N_5659,N_5304,N_5084);
nand U5660 (N_5660,N_5472,N_5393);
nand U5661 (N_5661,N_5505,N_5368);
xnor U5662 (N_5662,N_5104,N_5502);
nand U5663 (N_5663,N_5099,N_5551);
nor U5664 (N_5664,N_5245,N_5250);
nor U5665 (N_5665,N_5175,N_5506);
xor U5666 (N_5666,N_5618,N_5478);
or U5667 (N_5667,N_5383,N_5578);
nor U5668 (N_5668,N_5596,N_5442);
and U5669 (N_5669,N_5599,N_5269);
nand U5670 (N_5670,N_5305,N_5318);
nor U5671 (N_5671,N_5377,N_5388);
and U5672 (N_5672,N_5430,N_5363);
nor U5673 (N_5673,N_5474,N_5518);
xnor U5674 (N_5674,N_5024,N_5496);
xnor U5675 (N_5675,N_5244,N_5213);
or U5676 (N_5676,N_5341,N_5315);
nand U5677 (N_5677,N_5313,N_5488);
and U5678 (N_5678,N_5439,N_5286);
nor U5679 (N_5679,N_5219,N_5270);
nor U5680 (N_5680,N_5008,N_5593);
or U5681 (N_5681,N_5441,N_5065);
nand U5682 (N_5682,N_5414,N_5209);
and U5683 (N_5683,N_5183,N_5359);
nand U5684 (N_5684,N_5344,N_5278);
or U5685 (N_5685,N_5295,N_5462);
nor U5686 (N_5686,N_5493,N_5477);
xnor U5687 (N_5687,N_5266,N_5314);
and U5688 (N_5688,N_5561,N_5260);
nor U5689 (N_5689,N_5171,N_5095);
and U5690 (N_5690,N_5563,N_5576);
and U5691 (N_5691,N_5547,N_5355);
xor U5692 (N_5692,N_5490,N_5413);
nor U5693 (N_5693,N_5469,N_5613);
nor U5694 (N_5694,N_5558,N_5030);
xor U5695 (N_5695,N_5500,N_5225);
nor U5696 (N_5696,N_5550,N_5097);
nor U5697 (N_5697,N_5150,N_5281);
and U5698 (N_5698,N_5386,N_5407);
nor U5699 (N_5699,N_5299,N_5149);
nor U5700 (N_5700,N_5070,N_5617);
and U5701 (N_5701,N_5607,N_5156);
and U5702 (N_5702,N_5044,N_5301);
xnor U5703 (N_5703,N_5257,N_5610);
xnor U5704 (N_5704,N_5180,N_5433);
nor U5705 (N_5705,N_5212,N_5290);
and U5706 (N_5706,N_5148,N_5522);
nand U5707 (N_5707,N_5193,N_5583);
or U5708 (N_5708,N_5381,N_5394);
nand U5709 (N_5709,N_5015,N_5273);
or U5710 (N_5710,N_5492,N_5619);
and U5711 (N_5711,N_5062,N_5198);
nand U5712 (N_5712,N_5006,N_5334);
xnor U5713 (N_5713,N_5235,N_5320);
or U5714 (N_5714,N_5539,N_5350);
nor U5715 (N_5715,N_5423,N_5293);
xor U5716 (N_5716,N_5113,N_5398);
and U5717 (N_5717,N_5598,N_5467);
nor U5718 (N_5718,N_5157,N_5542);
nor U5719 (N_5719,N_5517,N_5601);
or U5720 (N_5720,N_5087,N_5076);
nor U5721 (N_5721,N_5312,N_5515);
or U5722 (N_5722,N_5373,N_5534);
nor U5723 (N_5723,N_5138,N_5168);
nand U5724 (N_5724,N_5139,N_5155);
nand U5725 (N_5725,N_5436,N_5448);
or U5726 (N_5726,N_5222,N_5173);
nor U5727 (N_5727,N_5161,N_5404);
and U5728 (N_5728,N_5470,N_5557);
nand U5729 (N_5729,N_5365,N_5590);
or U5730 (N_5730,N_5485,N_5098);
nor U5731 (N_5731,N_5567,N_5553);
nor U5732 (N_5732,N_5252,N_5352);
nor U5733 (N_5733,N_5579,N_5584);
xor U5734 (N_5734,N_5476,N_5487);
and U5735 (N_5735,N_5536,N_5292);
or U5736 (N_5736,N_5336,N_5415);
or U5737 (N_5737,N_5004,N_5562);
xnor U5738 (N_5738,N_5162,N_5459);
or U5739 (N_5739,N_5112,N_5242);
or U5740 (N_5740,N_5570,N_5125);
nor U5741 (N_5741,N_5201,N_5159);
xor U5742 (N_5742,N_5220,N_5240);
xor U5743 (N_5743,N_5014,N_5211);
or U5744 (N_5744,N_5444,N_5075);
nand U5745 (N_5745,N_5432,N_5274);
and U5746 (N_5746,N_5338,N_5446);
nand U5747 (N_5747,N_5483,N_5569);
nand U5748 (N_5748,N_5568,N_5460);
or U5749 (N_5749,N_5587,N_5330);
nor U5750 (N_5750,N_5121,N_5559);
and U5751 (N_5751,N_5323,N_5424);
and U5752 (N_5752,N_5058,N_5306);
and U5753 (N_5753,N_5140,N_5549);
nand U5754 (N_5754,N_5507,N_5069);
nand U5755 (N_5755,N_5316,N_5376);
and U5756 (N_5756,N_5083,N_5117);
and U5757 (N_5757,N_5283,N_5061);
nand U5758 (N_5758,N_5481,N_5333);
nand U5759 (N_5759,N_5452,N_5353);
nand U5760 (N_5760,N_5543,N_5210);
or U5761 (N_5761,N_5133,N_5253);
nor U5762 (N_5762,N_5199,N_5124);
xor U5763 (N_5763,N_5294,N_5527);
nor U5764 (N_5764,N_5554,N_5538);
and U5765 (N_5765,N_5378,N_5205);
or U5766 (N_5766,N_5552,N_5565);
nor U5767 (N_5767,N_5375,N_5367);
nand U5768 (N_5768,N_5064,N_5319);
and U5769 (N_5769,N_5331,N_5230);
nand U5770 (N_5770,N_5546,N_5611);
or U5771 (N_5771,N_5231,N_5429);
or U5772 (N_5772,N_5497,N_5608);
nor U5773 (N_5773,N_5042,N_5003);
xnor U5774 (N_5774,N_5200,N_5166);
xnor U5775 (N_5775,N_5389,N_5624);
nor U5776 (N_5776,N_5132,N_5144);
xnor U5777 (N_5777,N_5287,N_5580);
nand U5778 (N_5778,N_5277,N_5342);
nor U5779 (N_5779,N_5581,N_5236);
nand U5780 (N_5780,N_5228,N_5167);
or U5781 (N_5781,N_5108,N_5120);
and U5782 (N_5782,N_5056,N_5118);
xnor U5783 (N_5783,N_5498,N_5002);
nor U5784 (N_5784,N_5371,N_5384);
or U5785 (N_5785,N_5597,N_5267);
nand U5786 (N_5786,N_5060,N_5466);
xor U5787 (N_5787,N_5036,N_5229);
nand U5788 (N_5788,N_5202,N_5455);
nand U5789 (N_5789,N_5296,N_5545);
xnor U5790 (N_5790,N_5501,N_5526);
nand U5791 (N_5791,N_5391,N_5513);
or U5792 (N_5792,N_5013,N_5028);
or U5793 (N_5793,N_5390,N_5592);
nor U5794 (N_5794,N_5195,N_5408);
and U5795 (N_5795,N_5454,N_5122);
nand U5796 (N_5796,N_5279,N_5461);
nand U5797 (N_5797,N_5000,N_5052);
nor U5798 (N_5798,N_5018,N_5143);
and U5799 (N_5799,N_5129,N_5349);
nand U5800 (N_5800,N_5434,N_5145);
nor U5801 (N_5801,N_5465,N_5085);
or U5802 (N_5802,N_5172,N_5094);
xnor U5803 (N_5803,N_5622,N_5241);
or U5804 (N_5804,N_5114,N_5616);
xor U5805 (N_5805,N_5548,N_5457);
or U5806 (N_5806,N_5512,N_5354);
nand U5807 (N_5807,N_5223,N_5300);
or U5808 (N_5808,N_5417,N_5298);
xnor U5809 (N_5809,N_5324,N_5445);
and U5810 (N_5810,N_5268,N_5131);
and U5811 (N_5811,N_5110,N_5401);
or U5812 (N_5812,N_5089,N_5535);
nor U5813 (N_5813,N_5288,N_5449);
and U5814 (N_5814,N_5016,N_5251);
nand U5815 (N_5815,N_5456,N_5479);
and U5816 (N_5816,N_5186,N_5604);
nand U5817 (N_5817,N_5380,N_5468);
or U5818 (N_5818,N_5010,N_5007);
xnor U5819 (N_5819,N_5361,N_5032);
nor U5820 (N_5820,N_5348,N_5484);
or U5821 (N_5821,N_5372,N_5050);
or U5822 (N_5822,N_5392,N_5239);
xor U5823 (N_5823,N_5182,N_5174);
nand U5824 (N_5824,N_5343,N_5285);
and U5825 (N_5825,N_5422,N_5093);
nor U5826 (N_5826,N_5303,N_5152);
xnor U5827 (N_5827,N_5047,N_5033);
or U5828 (N_5828,N_5369,N_5311);
nor U5829 (N_5829,N_5102,N_5051);
nor U5830 (N_5830,N_5564,N_5351);
and U5831 (N_5831,N_5510,N_5126);
or U5832 (N_5832,N_5594,N_5588);
and U5833 (N_5833,N_5280,N_5227);
nor U5834 (N_5834,N_5074,N_5530);
nor U5835 (N_5835,N_5308,N_5247);
or U5836 (N_5836,N_5447,N_5482);
nand U5837 (N_5837,N_5435,N_5101);
or U5838 (N_5838,N_5040,N_5185);
nand U5839 (N_5839,N_5284,N_5215);
and U5840 (N_5840,N_5071,N_5556);
xor U5841 (N_5841,N_5504,N_5086);
or U5842 (N_5842,N_5012,N_5491);
nor U5843 (N_5843,N_5081,N_5560);
and U5844 (N_5844,N_5216,N_5259);
nand U5845 (N_5845,N_5163,N_5537);
nand U5846 (N_5846,N_5623,N_5463);
nor U5847 (N_5847,N_5147,N_5233);
and U5848 (N_5848,N_5489,N_5356);
or U5849 (N_5849,N_5027,N_5525);
xor U5850 (N_5850,N_5475,N_5243);
nor U5851 (N_5851,N_5382,N_5346);
xor U5852 (N_5852,N_5443,N_5011);
or U5853 (N_5853,N_5282,N_5595);
nor U5854 (N_5854,N_5509,N_5049);
nor U5855 (N_5855,N_5606,N_5358);
or U5856 (N_5856,N_5023,N_5031);
or U5857 (N_5857,N_5364,N_5048);
nor U5858 (N_5858,N_5141,N_5204);
nand U5859 (N_5859,N_5196,N_5418);
and U5860 (N_5860,N_5406,N_5153);
or U5861 (N_5861,N_5059,N_5528);
and U5862 (N_5862,N_5025,N_5337);
nor U5863 (N_5863,N_5524,N_5322);
nor U5864 (N_5864,N_5494,N_5135);
or U5865 (N_5865,N_5009,N_5178);
or U5866 (N_5866,N_5207,N_5043);
and U5867 (N_5867,N_5054,N_5503);
nor U5868 (N_5868,N_5573,N_5116);
nand U5869 (N_5869,N_5109,N_5022);
nor U5870 (N_5870,N_5519,N_5221);
nor U5871 (N_5871,N_5575,N_5345);
nor U5872 (N_5872,N_5357,N_5464);
or U5873 (N_5873,N_5327,N_5194);
or U5874 (N_5874,N_5411,N_5265);
xor U5875 (N_5875,N_5034,N_5238);
or U5876 (N_5876,N_5335,N_5451);
xnor U5877 (N_5877,N_5275,N_5020);
nand U5878 (N_5878,N_5165,N_5160);
and U5879 (N_5879,N_5111,N_5609);
or U5880 (N_5880,N_5105,N_5264);
or U5881 (N_5881,N_5420,N_5514);
nor U5882 (N_5882,N_5440,N_5262);
and U5883 (N_5883,N_5256,N_5387);
nand U5884 (N_5884,N_5602,N_5072);
or U5885 (N_5885,N_5499,N_5055);
xnor U5886 (N_5886,N_5427,N_5137);
or U5887 (N_5887,N_5385,N_5589);
or U5888 (N_5888,N_5523,N_5176);
or U5889 (N_5889,N_5471,N_5276);
nand U5890 (N_5890,N_5019,N_5026);
nand U5891 (N_5891,N_5614,N_5164);
nor U5892 (N_5892,N_5421,N_5045);
nand U5893 (N_5893,N_5192,N_5263);
xor U5894 (N_5894,N_5189,N_5458);
or U5895 (N_5895,N_5080,N_5271);
nand U5896 (N_5896,N_5520,N_5107);
nor U5897 (N_5897,N_5621,N_5397);
or U5898 (N_5898,N_5142,N_5425);
xor U5899 (N_5899,N_5516,N_5151);
xnor U5900 (N_5900,N_5374,N_5037);
or U5901 (N_5901,N_5188,N_5218);
nand U5902 (N_5902,N_5191,N_5603);
nand U5903 (N_5903,N_5325,N_5158);
and U5904 (N_5904,N_5379,N_5184);
nor U5905 (N_5905,N_5591,N_5396);
or U5906 (N_5906,N_5321,N_5170);
nor U5907 (N_5907,N_5291,N_5134);
nand U5908 (N_5908,N_5339,N_5533);
xor U5909 (N_5909,N_5400,N_5258);
nor U5910 (N_5910,N_5541,N_5046);
nor U5911 (N_5911,N_5197,N_5473);
xnor U5912 (N_5912,N_5261,N_5370);
nor U5913 (N_5913,N_5360,N_5540);
nor U5914 (N_5914,N_5600,N_5307);
nor U5915 (N_5915,N_5127,N_5082);
nor U5916 (N_5916,N_5574,N_5620);
nor U5917 (N_5917,N_5005,N_5395);
nor U5918 (N_5918,N_5416,N_5224);
or U5919 (N_5919,N_5130,N_5088);
xnor U5920 (N_5920,N_5437,N_5232);
nor U5921 (N_5921,N_5399,N_5187);
nand U5922 (N_5922,N_5585,N_5521);
xnor U5923 (N_5923,N_5096,N_5340);
nand U5924 (N_5924,N_5511,N_5328);
and U5925 (N_5925,N_5289,N_5217);
xnor U5926 (N_5926,N_5136,N_5453);
nor U5927 (N_5927,N_5508,N_5106);
xor U5928 (N_5928,N_5531,N_5038);
nand U5929 (N_5929,N_5067,N_5128);
and U5930 (N_5930,N_5438,N_5017);
xnor U5931 (N_5931,N_5206,N_5577);
nand U5932 (N_5932,N_5403,N_5572);
nor U5933 (N_5933,N_5362,N_5529);
nor U5934 (N_5934,N_5190,N_5347);
or U5935 (N_5935,N_5297,N_5035);
xnor U5936 (N_5936,N_5091,N_5234);
nand U5937 (N_5937,N_5103,N_5485);
xor U5938 (N_5938,N_5130,N_5393);
or U5939 (N_5939,N_5474,N_5096);
or U5940 (N_5940,N_5398,N_5446);
nand U5941 (N_5941,N_5073,N_5524);
nand U5942 (N_5942,N_5150,N_5499);
nand U5943 (N_5943,N_5037,N_5372);
nor U5944 (N_5944,N_5241,N_5285);
xor U5945 (N_5945,N_5498,N_5404);
or U5946 (N_5946,N_5035,N_5064);
and U5947 (N_5947,N_5237,N_5384);
and U5948 (N_5948,N_5411,N_5231);
and U5949 (N_5949,N_5093,N_5591);
or U5950 (N_5950,N_5551,N_5318);
or U5951 (N_5951,N_5457,N_5509);
and U5952 (N_5952,N_5531,N_5277);
or U5953 (N_5953,N_5388,N_5102);
or U5954 (N_5954,N_5389,N_5099);
or U5955 (N_5955,N_5401,N_5620);
and U5956 (N_5956,N_5304,N_5381);
nand U5957 (N_5957,N_5320,N_5095);
or U5958 (N_5958,N_5350,N_5542);
and U5959 (N_5959,N_5427,N_5170);
xnor U5960 (N_5960,N_5570,N_5236);
xnor U5961 (N_5961,N_5267,N_5394);
nand U5962 (N_5962,N_5592,N_5467);
or U5963 (N_5963,N_5253,N_5103);
xnor U5964 (N_5964,N_5296,N_5613);
or U5965 (N_5965,N_5535,N_5621);
nand U5966 (N_5966,N_5562,N_5512);
xor U5967 (N_5967,N_5298,N_5173);
nor U5968 (N_5968,N_5105,N_5259);
nand U5969 (N_5969,N_5146,N_5174);
nand U5970 (N_5970,N_5596,N_5283);
and U5971 (N_5971,N_5155,N_5527);
nor U5972 (N_5972,N_5224,N_5086);
or U5973 (N_5973,N_5160,N_5609);
xor U5974 (N_5974,N_5581,N_5296);
nand U5975 (N_5975,N_5376,N_5234);
and U5976 (N_5976,N_5269,N_5133);
and U5977 (N_5977,N_5044,N_5199);
nand U5978 (N_5978,N_5073,N_5534);
nor U5979 (N_5979,N_5600,N_5065);
and U5980 (N_5980,N_5110,N_5268);
nand U5981 (N_5981,N_5480,N_5325);
nor U5982 (N_5982,N_5078,N_5087);
or U5983 (N_5983,N_5263,N_5136);
xor U5984 (N_5984,N_5293,N_5161);
xor U5985 (N_5985,N_5114,N_5298);
nor U5986 (N_5986,N_5390,N_5219);
or U5987 (N_5987,N_5501,N_5255);
nand U5988 (N_5988,N_5621,N_5327);
and U5989 (N_5989,N_5420,N_5528);
nor U5990 (N_5990,N_5051,N_5260);
xor U5991 (N_5991,N_5109,N_5108);
xnor U5992 (N_5992,N_5224,N_5450);
and U5993 (N_5993,N_5229,N_5282);
or U5994 (N_5994,N_5158,N_5622);
and U5995 (N_5995,N_5599,N_5610);
nand U5996 (N_5996,N_5530,N_5043);
nor U5997 (N_5997,N_5025,N_5043);
or U5998 (N_5998,N_5238,N_5550);
and U5999 (N_5999,N_5196,N_5534);
and U6000 (N_6000,N_5217,N_5325);
and U6001 (N_6001,N_5034,N_5416);
nor U6002 (N_6002,N_5204,N_5269);
nor U6003 (N_6003,N_5106,N_5017);
and U6004 (N_6004,N_5024,N_5224);
nand U6005 (N_6005,N_5247,N_5496);
or U6006 (N_6006,N_5223,N_5183);
or U6007 (N_6007,N_5395,N_5144);
nand U6008 (N_6008,N_5586,N_5142);
nand U6009 (N_6009,N_5478,N_5594);
and U6010 (N_6010,N_5354,N_5085);
nand U6011 (N_6011,N_5374,N_5096);
nor U6012 (N_6012,N_5554,N_5331);
nand U6013 (N_6013,N_5326,N_5433);
xor U6014 (N_6014,N_5319,N_5297);
nand U6015 (N_6015,N_5599,N_5142);
xor U6016 (N_6016,N_5394,N_5197);
and U6017 (N_6017,N_5016,N_5201);
nor U6018 (N_6018,N_5487,N_5207);
xnor U6019 (N_6019,N_5143,N_5463);
or U6020 (N_6020,N_5594,N_5297);
xnor U6021 (N_6021,N_5336,N_5466);
xnor U6022 (N_6022,N_5167,N_5209);
and U6023 (N_6023,N_5481,N_5503);
nand U6024 (N_6024,N_5446,N_5367);
xor U6025 (N_6025,N_5322,N_5299);
nand U6026 (N_6026,N_5290,N_5035);
or U6027 (N_6027,N_5404,N_5084);
nand U6028 (N_6028,N_5175,N_5086);
and U6029 (N_6029,N_5267,N_5234);
xor U6030 (N_6030,N_5286,N_5567);
or U6031 (N_6031,N_5337,N_5262);
xor U6032 (N_6032,N_5425,N_5578);
nor U6033 (N_6033,N_5502,N_5248);
nand U6034 (N_6034,N_5575,N_5092);
xor U6035 (N_6035,N_5094,N_5567);
and U6036 (N_6036,N_5400,N_5393);
xor U6037 (N_6037,N_5135,N_5439);
or U6038 (N_6038,N_5580,N_5307);
or U6039 (N_6039,N_5542,N_5411);
nand U6040 (N_6040,N_5384,N_5421);
xnor U6041 (N_6041,N_5601,N_5118);
nand U6042 (N_6042,N_5405,N_5271);
nand U6043 (N_6043,N_5198,N_5355);
nor U6044 (N_6044,N_5602,N_5518);
xnor U6045 (N_6045,N_5048,N_5597);
or U6046 (N_6046,N_5406,N_5211);
nor U6047 (N_6047,N_5047,N_5621);
and U6048 (N_6048,N_5303,N_5101);
xnor U6049 (N_6049,N_5550,N_5546);
and U6050 (N_6050,N_5073,N_5431);
nand U6051 (N_6051,N_5335,N_5156);
nor U6052 (N_6052,N_5161,N_5186);
or U6053 (N_6053,N_5609,N_5615);
nor U6054 (N_6054,N_5410,N_5101);
nand U6055 (N_6055,N_5002,N_5189);
xnor U6056 (N_6056,N_5101,N_5183);
nor U6057 (N_6057,N_5536,N_5048);
or U6058 (N_6058,N_5449,N_5489);
xnor U6059 (N_6059,N_5566,N_5518);
nor U6060 (N_6060,N_5021,N_5057);
nand U6061 (N_6061,N_5196,N_5297);
xnor U6062 (N_6062,N_5440,N_5335);
nand U6063 (N_6063,N_5485,N_5124);
and U6064 (N_6064,N_5578,N_5376);
or U6065 (N_6065,N_5049,N_5271);
and U6066 (N_6066,N_5314,N_5623);
and U6067 (N_6067,N_5048,N_5238);
and U6068 (N_6068,N_5163,N_5114);
or U6069 (N_6069,N_5247,N_5094);
nand U6070 (N_6070,N_5231,N_5126);
and U6071 (N_6071,N_5047,N_5237);
or U6072 (N_6072,N_5159,N_5503);
and U6073 (N_6073,N_5376,N_5153);
and U6074 (N_6074,N_5491,N_5457);
xor U6075 (N_6075,N_5477,N_5335);
nor U6076 (N_6076,N_5438,N_5300);
xor U6077 (N_6077,N_5468,N_5303);
nor U6078 (N_6078,N_5199,N_5014);
nand U6079 (N_6079,N_5562,N_5246);
and U6080 (N_6080,N_5365,N_5152);
and U6081 (N_6081,N_5307,N_5079);
and U6082 (N_6082,N_5154,N_5486);
and U6083 (N_6083,N_5128,N_5081);
and U6084 (N_6084,N_5099,N_5108);
and U6085 (N_6085,N_5544,N_5179);
or U6086 (N_6086,N_5272,N_5528);
xor U6087 (N_6087,N_5072,N_5554);
nor U6088 (N_6088,N_5009,N_5064);
nand U6089 (N_6089,N_5154,N_5193);
and U6090 (N_6090,N_5222,N_5614);
or U6091 (N_6091,N_5507,N_5068);
and U6092 (N_6092,N_5407,N_5482);
xnor U6093 (N_6093,N_5126,N_5117);
nand U6094 (N_6094,N_5268,N_5181);
nand U6095 (N_6095,N_5015,N_5617);
nand U6096 (N_6096,N_5492,N_5482);
nor U6097 (N_6097,N_5596,N_5211);
nor U6098 (N_6098,N_5574,N_5007);
or U6099 (N_6099,N_5542,N_5330);
xnor U6100 (N_6100,N_5219,N_5332);
and U6101 (N_6101,N_5395,N_5269);
nand U6102 (N_6102,N_5362,N_5264);
xnor U6103 (N_6103,N_5137,N_5055);
nor U6104 (N_6104,N_5388,N_5225);
or U6105 (N_6105,N_5501,N_5514);
and U6106 (N_6106,N_5296,N_5378);
nand U6107 (N_6107,N_5208,N_5607);
xor U6108 (N_6108,N_5175,N_5525);
and U6109 (N_6109,N_5191,N_5003);
or U6110 (N_6110,N_5427,N_5450);
and U6111 (N_6111,N_5559,N_5295);
nor U6112 (N_6112,N_5288,N_5209);
nand U6113 (N_6113,N_5492,N_5373);
nand U6114 (N_6114,N_5391,N_5606);
xnor U6115 (N_6115,N_5362,N_5262);
or U6116 (N_6116,N_5612,N_5335);
or U6117 (N_6117,N_5505,N_5610);
nor U6118 (N_6118,N_5096,N_5284);
nand U6119 (N_6119,N_5260,N_5497);
and U6120 (N_6120,N_5203,N_5138);
or U6121 (N_6121,N_5219,N_5461);
nor U6122 (N_6122,N_5389,N_5128);
or U6123 (N_6123,N_5226,N_5014);
xnor U6124 (N_6124,N_5285,N_5191);
and U6125 (N_6125,N_5218,N_5420);
and U6126 (N_6126,N_5287,N_5348);
xor U6127 (N_6127,N_5098,N_5304);
nor U6128 (N_6128,N_5085,N_5041);
nand U6129 (N_6129,N_5085,N_5383);
nand U6130 (N_6130,N_5198,N_5527);
or U6131 (N_6131,N_5313,N_5553);
or U6132 (N_6132,N_5275,N_5556);
and U6133 (N_6133,N_5061,N_5075);
nor U6134 (N_6134,N_5543,N_5038);
nand U6135 (N_6135,N_5028,N_5046);
or U6136 (N_6136,N_5199,N_5285);
nand U6137 (N_6137,N_5090,N_5505);
nand U6138 (N_6138,N_5598,N_5601);
xor U6139 (N_6139,N_5064,N_5362);
and U6140 (N_6140,N_5298,N_5513);
and U6141 (N_6141,N_5499,N_5202);
and U6142 (N_6142,N_5557,N_5520);
or U6143 (N_6143,N_5014,N_5324);
or U6144 (N_6144,N_5028,N_5280);
nand U6145 (N_6145,N_5048,N_5417);
nor U6146 (N_6146,N_5295,N_5303);
xnor U6147 (N_6147,N_5229,N_5479);
and U6148 (N_6148,N_5075,N_5372);
nand U6149 (N_6149,N_5306,N_5121);
or U6150 (N_6150,N_5465,N_5099);
nor U6151 (N_6151,N_5550,N_5157);
xor U6152 (N_6152,N_5218,N_5203);
nor U6153 (N_6153,N_5107,N_5236);
and U6154 (N_6154,N_5095,N_5012);
and U6155 (N_6155,N_5563,N_5121);
nor U6156 (N_6156,N_5391,N_5589);
xnor U6157 (N_6157,N_5260,N_5574);
and U6158 (N_6158,N_5343,N_5005);
nand U6159 (N_6159,N_5153,N_5270);
xor U6160 (N_6160,N_5353,N_5498);
or U6161 (N_6161,N_5114,N_5290);
and U6162 (N_6162,N_5399,N_5259);
nor U6163 (N_6163,N_5123,N_5237);
nor U6164 (N_6164,N_5401,N_5080);
nor U6165 (N_6165,N_5364,N_5508);
nor U6166 (N_6166,N_5364,N_5422);
or U6167 (N_6167,N_5175,N_5458);
or U6168 (N_6168,N_5568,N_5076);
nor U6169 (N_6169,N_5156,N_5308);
or U6170 (N_6170,N_5488,N_5103);
xnor U6171 (N_6171,N_5595,N_5217);
or U6172 (N_6172,N_5533,N_5383);
nor U6173 (N_6173,N_5404,N_5245);
nor U6174 (N_6174,N_5188,N_5051);
or U6175 (N_6175,N_5169,N_5015);
or U6176 (N_6176,N_5433,N_5011);
and U6177 (N_6177,N_5178,N_5562);
nor U6178 (N_6178,N_5019,N_5587);
nand U6179 (N_6179,N_5104,N_5342);
nand U6180 (N_6180,N_5463,N_5564);
nor U6181 (N_6181,N_5112,N_5265);
nand U6182 (N_6182,N_5051,N_5515);
or U6183 (N_6183,N_5320,N_5406);
and U6184 (N_6184,N_5107,N_5454);
xnor U6185 (N_6185,N_5392,N_5262);
and U6186 (N_6186,N_5283,N_5004);
or U6187 (N_6187,N_5389,N_5120);
or U6188 (N_6188,N_5243,N_5007);
xnor U6189 (N_6189,N_5149,N_5612);
nor U6190 (N_6190,N_5471,N_5432);
xnor U6191 (N_6191,N_5182,N_5038);
nor U6192 (N_6192,N_5560,N_5622);
nor U6193 (N_6193,N_5521,N_5424);
xnor U6194 (N_6194,N_5279,N_5434);
nand U6195 (N_6195,N_5061,N_5587);
nor U6196 (N_6196,N_5067,N_5432);
or U6197 (N_6197,N_5321,N_5322);
nor U6198 (N_6198,N_5166,N_5514);
and U6199 (N_6199,N_5134,N_5323);
xnor U6200 (N_6200,N_5230,N_5007);
or U6201 (N_6201,N_5045,N_5083);
or U6202 (N_6202,N_5194,N_5167);
or U6203 (N_6203,N_5355,N_5585);
nor U6204 (N_6204,N_5004,N_5274);
or U6205 (N_6205,N_5124,N_5271);
nor U6206 (N_6206,N_5008,N_5267);
and U6207 (N_6207,N_5365,N_5382);
xnor U6208 (N_6208,N_5397,N_5583);
nand U6209 (N_6209,N_5409,N_5490);
xor U6210 (N_6210,N_5362,N_5110);
and U6211 (N_6211,N_5081,N_5506);
or U6212 (N_6212,N_5323,N_5545);
or U6213 (N_6213,N_5448,N_5012);
or U6214 (N_6214,N_5387,N_5519);
and U6215 (N_6215,N_5138,N_5512);
and U6216 (N_6216,N_5352,N_5306);
nor U6217 (N_6217,N_5122,N_5005);
xnor U6218 (N_6218,N_5507,N_5033);
nand U6219 (N_6219,N_5293,N_5144);
and U6220 (N_6220,N_5093,N_5509);
and U6221 (N_6221,N_5322,N_5158);
xnor U6222 (N_6222,N_5457,N_5012);
or U6223 (N_6223,N_5431,N_5055);
and U6224 (N_6224,N_5297,N_5614);
nor U6225 (N_6225,N_5075,N_5348);
nand U6226 (N_6226,N_5456,N_5357);
or U6227 (N_6227,N_5404,N_5024);
nand U6228 (N_6228,N_5084,N_5080);
nand U6229 (N_6229,N_5187,N_5035);
xor U6230 (N_6230,N_5611,N_5088);
or U6231 (N_6231,N_5326,N_5493);
nor U6232 (N_6232,N_5023,N_5294);
and U6233 (N_6233,N_5343,N_5304);
and U6234 (N_6234,N_5583,N_5537);
or U6235 (N_6235,N_5015,N_5008);
or U6236 (N_6236,N_5606,N_5544);
nor U6237 (N_6237,N_5397,N_5439);
nor U6238 (N_6238,N_5116,N_5618);
nand U6239 (N_6239,N_5481,N_5312);
or U6240 (N_6240,N_5460,N_5398);
nand U6241 (N_6241,N_5461,N_5058);
xnor U6242 (N_6242,N_5136,N_5138);
nand U6243 (N_6243,N_5061,N_5241);
xor U6244 (N_6244,N_5018,N_5008);
xor U6245 (N_6245,N_5260,N_5355);
or U6246 (N_6246,N_5328,N_5004);
nand U6247 (N_6247,N_5296,N_5130);
or U6248 (N_6248,N_5241,N_5349);
nor U6249 (N_6249,N_5566,N_5301);
xnor U6250 (N_6250,N_6180,N_6138);
or U6251 (N_6251,N_5680,N_5979);
and U6252 (N_6252,N_5674,N_5995);
nand U6253 (N_6253,N_6012,N_5791);
nand U6254 (N_6254,N_6190,N_5795);
nor U6255 (N_6255,N_5780,N_6169);
nand U6256 (N_6256,N_6183,N_6021);
and U6257 (N_6257,N_5818,N_6049);
nand U6258 (N_6258,N_6130,N_5944);
and U6259 (N_6259,N_5851,N_6038);
nor U6260 (N_6260,N_6092,N_5881);
xnor U6261 (N_6261,N_6058,N_5732);
or U6262 (N_6262,N_5776,N_5855);
or U6263 (N_6263,N_6240,N_6152);
nor U6264 (N_6264,N_5648,N_5894);
xnor U6265 (N_6265,N_5629,N_6026);
nor U6266 (N_6266,N_5999,N_5840);
nor U6267 (N_6267,N_5889,N_5811);
and U6268 (N_6268,N_5789,N_5736);
xor U6269 (N_6269,N_6193,N_5774);
nand U6270 (N_6270,N_5842,N_5691);
and U6271 (N_6271,N_5934,N_6024);
xor U6272 (N_6272,N_5800,N_5793);
nor U6273 (N_6273,N_6128,N_6001);
nor U6274 (N_6274,N_5782,N_5830);
and U6275 (N_6275,N_5985,N_6159);
nand U6276 (N_6276,N_5667,N_5743);
or U6277 (N_6277,N_6062,N_5824);
nor U6278 (N_6278,N_5775,N_5849);
nand U6279 (N_6279,N_5844,N_5873);
xnor U6280 (N_6280,N_6247,N_5837);
and U6281 (N_6281,N_5910,N_5801);
and U6282 (N_6282,N_6084,N_6151);
nand U6283 (N_6283,N_5929,N_5927);
or U6284 (N_6284,N_6003,N_5703);
and U6285 (N_6285,N_5988,N_5947);
nor U6286 (N_6286,N_5865,N_5933);
nand U6287 (N_6287,N_5996,N_6132);
or U6288 (N_6288,N_5870,N_5816);
nor U6289 (N_6289,N_6039,N_6223);
and U6290 (N_6290,N_5841,N_6107);
and U6291 (N_6291,N_5746,N_5852);
xnor U6292 (N_6292,N_5652,N_6077);
or U6293 (N_6293,N_5978,N_6019);
xnor U6294 (N_6294,N_5712,N_5874);
nor U6295 (N_6295,N_5903,N_6002);
nor U6296 (N_6296,N_6164,N_6185);
nand U6297 (N_6297,N_5670,N_6233);
nor U6298 (N_6298,N_5863,N_5964);
nand U6299 (N_6299,N_5750,N_5945);
and U6300 (N_6300,N_5812,N_5633);
nand U6301 (N_6301,N_5992,N_5970);
or U6302 (N_6302,N_6086,N_5885);
xor U6303 (N_6303,N_5734,N_6141);
and U6304 (N_6304,N_6199,N_5936);
or U6305 (N_6305,N_5883,N_5913);
or U6306 (N_6306,N_5857,N_5848);
and U6307 (N_6307,N_6133,N_5876);
nand U6308 (N_6308,N_5636,N_5815);
nand U6309 (N_6309,N_5639,N_5668);
and U6310 (N_6310,N_5861,N_6103);
xnor U6311 (N_6311,N_6112,N_5696);
or U6312 (N_6312,N_5896,N_5882);
or U6313 (N_6313,N_5958,N_6027);
or U6314 (N_6314,N_5659,N_6249);
nor U6315 (N_6315,N_6129,N_6165);
xor U6316 (N_6316,N_6192,N_5845);
xnor U6317 (N_6317,N_5950,N_6120);
and U6318 (N_6318,N_6235,N_6025);
nand U6319 (N_6319,N_6007,N_5969);
xor U6320 (N_6320,N_6031,N_6110);
nand U6321 (N_6321,N_5737,N_5955);
and U6322 (N_6322,N_6217,N_6010);
or U6323 (N_6323,N_5854,N_6045);
nor U6324 (N_6324,N_6176,N_6149);
nor U6325 (N_6325,N_5713,N_6237);
xnor U6326 (N_6326,N_5898,N_5693);
or U6327 (N_6327,N_6234,N_5821);
nor U6328 (N_6328,N_5905,N_6067);
nand U6329 (N_6329,N_5654,N_5688);
nor U6330 (N_6330,N_6232,N_6136);
nor U6331 (N_6331,N_6211,N_5627);
nor U6332 (N_6332,N_6071,N_6078);
xnor U6333 (N_6333,N_6108,N_6059);
or U6334 (N_6334,N_5904,N_6150);
xor U6335 (N_6335,N_6040,N_6171);
or U6336 (N_6336,N_5959,N_5822);
nor U6337 (N_6337,N_6097,N_6061);
xor U6338 (N_6338,N_5798,N_5866);
or U6339 (N_6339,N_5957,N_6032);
and U6340 (N_6340,N_6218,N_5990);
xor U6341 (N_6341,N_5707,N_5642);
and U6342 (N_6342,N_6029,N_5856);
xor U6343 (N_6343,N_6013,N_5725);
nand U6344 (N_6344,N_5804,N_5867);
and U6345 (N_6345,N_5901,N_5980);
and U6346 (N_6346,N_5912,N_6083);
and U6347 (N_6347,N_6053,N_5790);
nor U6348 (N_6348,N_6056,N_5831);
xor U6349 (N_6349,N_5635,N_6225);
or U6350 (N_6350,N_5781,N_6178);
xnor U6351 (N_6351,N_6048,N_6207);
and U6352 (N_6352,N_5838,N_6115);
or U6353 (N_6353,N_5679,N_6091);
and U6354 (N_6354,N_6198,N_6119);
xor U6355 (N_6355,N_5653,N_6157);
nand U6356 (N_6356,N_6009,N_6008);
xor U6357 (N_6357,N_6182,N_5993);
and U6358 (N_6358,N_5983,N_5968);
nand U6359 (N_6359,N_6022,N_5987);
and U6360 (N_6360,N_5665,N_6096);
or U6361 (N_6361,N_5641,N_5808);
or U6362 (N_6362,N_5926,N_5777);
nor U6363 (N_6363,N_6065,N_5711);
or U6364 (N_6364,N_6172,N_5917);
nor U6365 (N_6365,N_5788,N_5739);
or U6366 (N_6366,N_5714,N_5891);
nor U6367 (N_6367,N_6095,N_5833);
xnor U6368 (N_6368,N_5689,N_5986);
nand U6369 (N_6369,N_6005,N_5690);
and U6370 (N_6370,N_6014,N_5643);
and U6371 (N_6371,N_6208,N_5864);
xnor U6372 (N_6372,N_5723,N_5890);
xor U6373 (N_6373,N_5759,N_5631);
xor U6374 (N_6374,N_5902,N_5735);
nor U6375 (N_6375,N_6194,N_5971);
nor U6376 (N_6376,N_6105,N_5839);
nand U6377 (N_6377,N_5930,N_5975);
nand U6378 (N_6378,N_5915,N_5880);
xor U6379 (N_6379,N_5662,N_5697);
or U6380 (N_6380,N_5892,N_5819);
or U6381 (N_6381,N_5906,N_6134);
xor U6382 (N_6382,N_5731,N_5921);
or U6383 (N_6383,N_5708,N_5922);
nor U6384 (N_6384,N_5692,N_6188);
nor U6385 (N_6385,N_5757,N_6226);
nand U6386 (N_6386,N_5802,N_6050);
or U6387 (N_6387,N_6229,N_6156);
nand U6388 (N_6388,N_5813,N_6135);
nand U6389 (N_6389,N_5722,N_6241);
and U6390 (N_6390,N_6201,N_5686);
and U6391 (N_6391,N_5721,N_5710);
or U6392 (N_6392,N_5756,N_6139);
xnor U6393 (N_6393,N_6230,N_6142);
xnor U6394 (N_6394,N_6051,N_5687);
nand U6395 (N_6395,N_5733,N_5773);
nand U6396 (N_6396,N_6227,N_5650);
and U6397 (N_6397,N_5871,N_5893);
and U6398 (N_6398,N_5860,N_5884);
xor U6399 (N_6399,N_6028,N_5656);
xor U6400 (N_6400,N_5799,N_5977);
and U6401 (N_6401,N_6044,N_6042);
and U6402 (N_6402,N_5754,N_6148);
and U6403 (N_6403,N_5942,N_5684);
nor U6404 (N_6404,N_5651,N_5677);
and U6405 (N_6405,N_6126,N_5869);
or U6406 (N_6406,N_5786,N_6212);
nand U6407 (N_6407,N_6203,N_5760);
xnor U6408 (N_6408,N_6189,N_5628);
nand U6409 (N_6409,N_5796,N_5729);
and U6410 (N_6410,N_5909,N_5836);
nor U6411 (N_6411,N_6098,N_5744);
nor U6412 (N_6412,N_5761,N_5937);
nand U6413 (N_6413,N_6043,N_5853);
nand U6414 (N_6414,N_5973,N_6113);
xor U6415 (N_6415,N_5718,N_5850);
nand U6416 (N_6416,N_6236,N_5742);
or U6417 (N_6417,N_5803,N_5899);
or U6418 (N_6418,N_5875,N_5982);
xnor U6419 (N_6419,N_5728,N_5724);
nand U6420 (N_6420,N_6166,N_6036);
nand U6421 (N_6421,N_6089,N_5877);
or U6422 (N_6422,N_6041,N_5814);
or U6423 (N_6423,N_6163,N_5868);
xnor U6424 (N_6424,N_5961,N_5946);
nand U6425 (N_6425,N_6175,N_5784);
nand U6426 (N_6426,N_5655,N_6161);
and U6427 (N_6427,N_6106,N_5626);
nand U6428 (N_6428,N_5768,N_5705);
xnor U6429 (N_6429,N_5741,N_6206);
xnor U6430 (N_6430,N_6220,N_6079);
nor U6431 (N_6431,N_6131,N_5956);
xnor U6432 (N_6432,N_6076,N_5829);
xnor U6433 (N_6433,N_6145,N_5663);
nand U6434 (N_6434,N_5704,N_5785);
nor U6435 (N_6435,N_6093,N_5716);
xor U6436 (N_6436,N_6243,N_5991);
nand U6437 (N_6437,N_5952,N_5630);
xnor U6438 (N_6438,N_6085,N_5758);
nor U6439 (N_6439,N_5751,N_5787);
and U6440 (N_6440,N_5770,N_6124);
nor U6441 (N_6441,N_5632,N_6052);
and U6442 (N_6442,N_6057,N_5657);
xor U6443 (N_6443,N_5954,N_6087);
xor U6444 (N_6444,N_5694,N_5888);
nand U6445 (N_6445,N_6070,N_5911);
or U6446 (N_6446,N_6162,N_6155);
nor U6447 (N_6447,N_6147,N_6094);
nor U6448 (N_6448,N_5805,N_5698);
and U6449 (N_6449,N_6143,N_5939);
nor U6450 (N_6450,N_5681,N_5682);
or U6451 (N_6451,N_6099,N_5963);
nand U6452 (N_6452,N_6210,N_5706);
nand U6453 (N_6453,N_6101,N_5972);
nand U6454 (N_6454,N_5685,N_5951);
or U6455 (N_6455,N_5932,N_5726);
and U6456 (N_6456,N_5807,N_5820);
and U6457 (N_6457,N_5678,N_6231);
and U6458 (N_6458,N_5660,N_6018);
or U6459 (N_6459,N_5778,N_6090);
xnor U6460 (N_6460,N_6011,N_5923);
nor U6461 (N_6461,N_5900,N_5645);
nor U6462 (N_6462,N_6023,N_6200);
and U6463 (N_6463,N_5753,N_6248);
and U6464 (N_6464,N_6184,N_5749);
nor U6465 (N_6465,N_5826,N_6088);
xor U6466 (N_6466,N_5717,N_6004);
or U6467 (N_6467,N_5797,N_5938);
or U6468 (N_6468,N_6000,N_6037);
nand U6469 (N_6469,N_5727,N_5994);
or U6470 (N_6470,N_5772,N_6158);
or U6471 (N_6471,N_5981,N_5638);
xor U6472 (N_6472,N_5740,N_6006);
nand U6473 (N_6473,N_5962,N_6046);
nor U6474 (N_6474,N_6196,N_6244);
xor U6475 (N_6475,N_6239,N_5715);
or U6476 (N_6476,N_5872,N_6238);
and U6477 (N_6477,N_5918,N_6213);
nand U6478 (N_6478,N_5832,N_6117);
nand U6479 (N_6479,N_5916,N_6063);
nor U6480 (N_6480,N_5919,N_6020);
nand U6481 (N_6481,N_6137,N_5771);
or U6482 (N_6482,N_5658,N_5779);
nor U6483 (N_6483,N_6104,N_5908);
and U6484 (N_6484,N_6109,N_5755);
nand U6485 (N_6485,N_5646,N_5664);
nor U6486 (N_6486,N_6122,N_6174);
xnor U6487 (N_6487,N_6246,N_6173);
xnor U6488 (N_6488,N_6082,N_5669);
and U6489 (N_6489,N_6202,N_5752);
nand U6490 (N_6490,N_6222,N_5738);
and U6491 (N_6491,N_6214,N_5859);
and U6492 (N_6492,N_6160,N_5763);
or U6493 (N_6493,N_5720,N_6035);
and U6494 (N_6494,N_5823,N_6060);
xor U6495 (N_6495,N_6015,N_6216);
and U6496 (N_6496,N_6205,N_6195);
xor U6497 (N_6497,N_6219,N_5666);
or U6498 (N_6498,N_6034,N_5640);
xnor U6499 (N_6499,N_6017,N_6170);
nand U6500 (N_6500,N_5960,N_5809);
xor U6501 (N_6501,N_6181,N_6073);
xor U6502 (N_6502,N_5943,N_5997);
xnor U6503 (N_6503,N_5675,N_6197);
nor U6504 (N_6504,N_6047,N_5817);
nand U6505 (N_6505,N_5941,N_6221);
xor U6506 (N_6506,N_6114,N_5827);
nand U6507 (N_6507,N_5794,N_5701);
nand U6508 (N_6508,N_5767,N_6016);
or U6509 (N_6509,N_6154,N_6167);
or U6510 (N_6510,N_6074,N_5966);
xor U6511 (N_6511,N_5907,N_6186);
xnor U6512 (N_6512,N_6153,N_6204);
nor U6513 (N_6513,N_5948,N_5649);
and U6514 (N_6514,N_5719,N_6191);
and U6515 (N_6515,N_5953,N_5924);
nor U6516 (N_6516,N_6066,N_6127);
and U6517 (N_6517,N_5935,N_5676);
or U6518 (N_6518,N_6179,N_6054);
or U6519 (N_6519,N_5846,N_5745);
or U6520 (N_6520,N_5644,N_5984);
nor U6521 (N_6521,N_5862,N_5765);
nor U6522 (N_6522,N_6102,N_5895);
or U6523 (N_6523,N_5747,N_6069);
and U6524 (N_6524,N_5858,N_5835);
nand U6525 (N_6525,N_6030,N_5783);
and U6526 (N_6526,N_5928,N_5730);
nor U6527 (N_6527,N_5967,N_5843);
xor U6528 (N_6528,N_5931,N_6080);
xor U6529 (N_6529,N_5637,N_6100);
nor U6530 (N_6530,N_5764,N_6144);
xnor U6531 (N_6531,N_6121,N_5810);
nor U6532 (N_6532,N_5847,N_5709);
nand U6533 (N_6533,N_6081,N_5702);
xnor U6534 (N_6534,N_6146,N_6125);
and U6535 (N_6535,N_5683,N_6118);
and U6536 (N_6536,N_5949,N_5828);
nor U6537 (N_6537,N_6242,N_5625);
and U6538 (N_6538,N_5748,N_5887);
and U6539 (N_6539,N_5965,N_5886);
nand U6540 (N_6540,N_5914,N_5806);
xnor U6541 (N_6541,N_5879,N_5998);
or U6542 (N_6542,N_6228,N_6072);
nand U6543 (N_6543,N_6168,N_5920);
nor U6544 (N_6544,N_5762,N_6123);
and U6545 (N_6545,N_5834,N_5792);
and U6546 (N_6546,N_6245,N_5671);
nand U6547 (N_6547,N_6140,N_6068);
nand U6548 (N_6548,N_5672,N_5878);
and U6549 (N_6549,N_6055,N_6033);
xor U6550 (N_6550,N_5974,N_5647);
and U6551 (N_6551,N_6111,N_6224);
nand U6552 (N_6552,N_5925,N_5700);
xor U6553 (N_6553,N_5695,N_6187);
or U6554 (N_6554,N_6215,N_5766);
nor U6555 (N_6555,N_5661,N_6116);
and U6556 (N_6556,N_6177,N_5940);
nand U6557 (N_6557,N_5825,N_5673);
or U6558 (N_6558,N_6064,N_6209);
nor U6559 (N_6559,N_5634,N_6075);
nand U6560 (N_6560,N_5976,N_5989);
and U6561 (N_6561,N_5699,N_5897);
and U6562 (N_6562,N_5769,N_6030);
nor U6563 (N_6563,N_5759,N_5996);
nor U6564 (N_6564,N_6064,N_6196);
nor U6565 (N_6565,N_6096,N_5966);
and U6566 (N_6566,N_5635,N_5881);
or U6567 (N_6567,N_5997,N_5932);
nand U6568 (N_6568,N_6208,N_5956);
xnor U6569 (N_6569,N_6051,N_5679);
or U6570 (N_6570,N_5987,N_6218);
and U6571 (N_6571,N_5670,N_5950);
or U6572 (N_6572,N_6124,N_5705);
xnor U6573 (N_6573,N_5831,N_5914);
nor U6574 (N_6574,N_5628,N_5839);
nor U6575 (N_6575,N_5877,N_5683);
nor U6576 (N_6576,N_6203,N_6077);
or U6577 (N_6577,N_6216,N_6205);
or U6578 (N_6578,N_5704,N_6004);
or U6579 (N_6579,N_5921,N_5695);
or U6580 (N_6580,N_6058,N_5930);
or U6581 (N_6581,N_5730,N_6016);
xor U6582 (N_6582,N_5656,N_6200);
nor U6583 (N_6583,N_5915,N_6085);
nor U6584 (N_6584,N_5885,N_5998);
or U6585 (N_6585,N_5814,N_5819);
or U6586 (N_6586,N_6231,N_5669);
and U6587 (N_6587,N_6028,N_6241);
xnor U6588 (N_6588,N_6042,N_6086);
or U6589 (N_6589,N_6142,N_5692);
and U6590 (N_6590,N_6140,N_5679);
nor U6591 (N_6591,N_6125,N_6070);
nor U6592 (N_6592,N_6143,N_5917);
nand U6593 (N_6593,N_5910,N_5947);
or U6594 (N_6594,N_5692,N_6214);
and U6595 (N_6595,N_6202,N_5861);
nand U6596 (N_6596,N_5981,N_5945);
and U6597 (N_6597,N_5631,N_6125);
or U6598 (N_6598,N_5890,N_5647);
and U6599 (N_6599,N_6208,N_6102);
nand U6600 (N_6600,N_6213,N_6161);
nor U6601 (N_6601,N_5795,N_5829);
nor U6602 (N_6602,N_6223,N_6182);
nor U6603 (N_6603,N_5664,N_5950);
and U6604 (N_6604,N_5845,N_6202);
nand U6605 (N_6605,N_5638,N_6199);
or U6606 (N_6606,N_6205,N_5636);
or U6607 (N_6607,N_6028,N_5653);
xnor U6608 (N_6608,N_6137,N_5909);
nand U6609 (N_6609,N_5881,N_5705);
or U6610 (N_6610,N_5739,N_5758);
nand U6611 (N_6611,N_6008,N_5888);
and U6612 (N_6612,N_5719,N_5696);
nor U6613 (N_6613,N_5957,N_6054);
nand U6614 (N_6614,N_5932,N_6010);
nor U6615 (N_6615,N_5704,N_5692);
nand U6616 (N_6616,N_6101,N_5941);
nor U6617 (N_6617,N_5712,N_5727);
xor U6618 (N_6618,N_5662,N_5729);
and U6619 (N_6619,N_5731,N_5837);
and U6620 (N_6620,N_6092,N_6002);
and U6621 (N_6621,N_6148,N_6100);
nand U6622 (N_6622,N_5895,N_6039);
and U6623 (N_6623,N_5900,N_6150);
nor U6624 (N_6624,N_5919,N_6189);
xor U6625 (N_6625,N_5710,N_6054);
xnor U6626 (N_6626,N_5810,N_6241);
nand U6627 (N_6627,N_5835,N_5975);
xor U6628 (N_6628,N_6229,N_6157);
nand U6629 (N_6629,N_5952,N_6055);
xor U6630 (N_6630,N_5698,N_5941);
or U6631 (N_6631,N_6243,N_6189);
nor U6632 (N_6632,N_5895,N_5993);
and U6633 (N_6633,N_6153,N_5747);
xor U6634 (N_6634,N_6028,N_5989);
nor U6635 (N_6635,N_5971,N_5671);
xor U6636 (N_6636,N_5769,N_5880);
nor U6637 (N_6637,N_6211,N_6179);
or U6638 (N_6638,N_5713,N_5778);
nor U6639 (N_6639,N_5825,N_5728);
nor U6640 (N_6640,N_6117,N_5684);
xnor U6641 (N_6641,N_6069,N_5761);
or U6642 (N_6642,N_5762,N_6113);
xor U6643 (N_6643,N_5926,N_5975);
and U6644 (N_6644,N_5749,N_5689);
and U6645 (N_6645,N_5633,N_5754);
xnor U6646 (N_6646,N_6105,N_5908);
nor U6647 (N_6647,N_5832,N_5646);
and U6648 (N_6648,N_5698,N_5858);
nor U6649 (N_6649,N_5863,N_6112);
and U6650 (N_6650,N_5817,N_6040);
nor U6651 (N_6651,N_6133,N_5648);
and U6652 (N_6652,N_5949,N_5697);
or U6653 (N_6653,N_6061,N_5966);
or U6654 (N_6654,N_6001,N_5880);
and U6655 (N_6655,N_6244,N_6248);
and U6656 (N_6656,N_5718,N_6000);
xnor U6657 (N_6657,N_6184,N_6134);
and U6658 (N_6658,N_6020,N_6178);
or U6659 (N_6659,N_6208,N_6040);
and U6660 (N_6660,N_5633,N_5871);
or U6661 (N_6661,N_6156,N_6163);
xor U6662 (N_6662,N_6085,N_5714);
and U6663 (N_6663,N_5948,N_5863);
nand U6664 (N_6664,N_5963,N_5823);
and U6665 (N_6665,N_5875,N_6124);
or U6666 (N_6666,N_5713,N_5658);
or U6667 (N_6667,N_6111,N_6235);
nor U6668 (N_6668,N_6013,N_5934);
xor U6669 (N_6669,N_5694,N_5970);
and U6670 (N_6670,N_5689,N_5863);
and U6671 (N_6671,N_5904,N_6033);
xnor U6672 (N_6672,N_6079,N_6157);
nor U6673 (N_6673,N_6246,N_5688);
xnor U6674 (N_6674,N_5653,N_6180);
nor U6675 (N_6675,N_5736,N_5995);
or U6676 (N_6676,N_5691,N_5753);
and U6677 (N_6677,N_5844,N_5697);
nand U6678 (N_6678,N_5985,N_6051);
or U6679 (N_6679,N_5699,N_5652);
or U6680 (N_6680,N_6217,N_5866);
nor U6681 (N_6681,N_5695,N_6142);
xnor U6682 (N_6682,N_5672,N_6107);
or U6683 (N_6683,N_6140,N_5902);
xnor U6684 (N_6684,N_5926,N_5994);
xor U6685 (N_6685,N_5646,N_5984);
xor U6686 (N_6686,N_5778,N_5918);
and U6687 (N_6687,N_5651,N_6234);
xor U6688 (N_6688,N_5996,N_5818);
and U6689 (N_6689,N_5839,N_5927);
nor U6690 (N_6690,N_5959,N_5839);
nor U6691 (N_6691,N_5964,N_5668);
and U6692 (N_6692,N_6192,N_6242);
or U6693 (N_6693,N_6096,N_6160);
or U6694 (N_6694,N_5640,N_5944);
or U6695 (N_6695,N_5728,N_5749);
nor U6696 (N_6696,N_5933,N_6163);
and U6697 (N_6697,N_6103,N_6061);
or U6698 (N_6698,N_5974,N_5758);
or U6699 (N_6699,N_6075,N_6244);
nand U6700 (N_6700,N_6086,N_5773);
xor U6701 (N_6701,N_5968,N_5863);
xor U6702 (N_6702,N_6210,N_6109);
nor U6703 (N_6703,N_5987,N_5663);
and U6704 (N_6704,N_6124,N_5983);
and U6705 (N_6705,N_6245,N_6047);
nand U6706 (N_6706,N_5830,N_6118);
or U6707 (N_6707,N_5984,N_6078);
and U6708 (N_6708,N_5770,N_5789);
nor U6709 (N_6709,N_5914,N_6010);
xor U6710 (N_6710,N_5769,N_5756);
and U6711 (N_6711,N_6006,N_5934);
nor U6712 (N_6712,N_5890,N_6160);
nor U6713 (N_6713,N_6113,N_6109);
nor U6714 (N_6714,N_6209,N_5730);
xnor U6715 (N_6715,N_5647,N_5939);
and U6716 (N_6716,N_5886,N_5778);
nand U6717 (N_6717,N_6191,N_5878);
or U6718 (N_6718,N_5773,N_5862);
nor U6719 (N_6719,N_5985,N_5799);
nor U6720 (N_6720,N_6122,N_5850);
nor U6721 (N_6721,N_5657,N_5961);
nand U6722 (N_6722,N_5993,N_5916);
nor U6723 (N_6723,N_5679,N_5974);
xor U6724 (N_6724,N_6151,N_6171);
xor U6725 (N_6725,N_5647,N_5803);
or U6726 (N_6726,N_6079,N_5631);
nor U6727 (N_6727,N_5699,N_6053);
and U6728 (N_6728,N_6244,N_5795);
and U6729 (N_6729,N_5981,N_6195);
xnor U6730 (N_6730,N_6199,N_5953);
or U6731 (N_6731,N_5862,N_5780);
or U6732 (N_6732,N_5813,N_5831);
or U6733 (N_6733,N_6232,N_6243);
or U6734 (N_6734,N_5736,N_5967);
nand U6735 (N_6735,N_5999,N_5869);
xnor U6736 (N_6736,N_5847,N_6023);
xor U6737 (N_6737,N_6067,N_5928);
and U6738 (N_6738,N_6076,N_6162);
or U6739 (N_6739,N_6234,N_5836);
or U6740 (N_6740,N_5637,N_6186);
nand U6741 (N_6741,N_5853,N_6139);
xor U6742 (N_6742,N_6190,N_5884);
and U6743 (N_6743,N_5984,N_5935);
or U6744 (N_6744,N_5947,N_6164);
or U6745 (N_6745,N_6144,N_5687);
or U6746 (N_6746,N_5950,N_5791);
or U6747 (N_6747,N_5781,N_5728);
or U6748 (N_6748,N_6006,N_5676);
nand U6749 (N_6749,N_6146,N_6201);
and U6750 (N_6750,N_6146,N_6156);
nor U6751 (N_6751,N_5778,N_5934);
and U6752 (N_6752,N_6048,N_6164);
xor U6753 (N_6753,N_5753,N_5799);
nand U6754 (N_6754,N_5662,N_5907);
nor U6755 (N_6755,N_6015,N_5767);
nand U6756 (N_6756,N_6156,N_6154);
or U6757 (N_6757,N_5819,N_6046);
nor U6758 (N_6758,N_6020,N_5705);
nor U6759 (N_6759,N_5767,N_5638);
or U6760 (N_6760,N_6150,N_5786);
xor U6761 (N_6761,N_5841,N_6014);
nand U6762 (N_6762,N_6078,N_5964);
xnor U6763 (N_6763,N_5900,N_5861);
or U6764 (N_6764,N_6015,N_5741);
nand U6765 (N_6765,N_6240,N_5993);
nand U6766 (N_6766,N_6133,N_5920);
nand U6767 (N_6767,N_5918,N_5705);
nand U6768 (N_6768,N_6119,N_6245);
and U6769 (N_6769,N_5830,N_6075);
and U6770 (N_6770,N_5808,N_5742);
nor U6771 (N_6771,N_6121,N_5935);
or U6772 (N_6772,N_6152,N_5803);
xnor U6773 (N_6773,N_6121,N_5665);
and U6774 (N_6774,N_6052,N_6153);
nor U6775 (N_6775,N_5681,N_5960);
xor U6776 (N_6776,N_5736,N_6207);
xnor U6777 (N_6777,N_6136,N_5952);
nor U6778 (N_6778,N_6119,N_5884);
nand U6779 (N_6779,N_6126,N_5853);
or U6780 (N_6780,N_5849,N_5797);
and U6781 (N_6781,N_5947,N_6081);
or U6782 (N_6782,N_6236,N_5987);
or U6783 (N_6783,N_5673,N_5888);
nand U6784 (N_6784,N_6177,N_6037);
and U6785 (N_6785,N_6127,N_5822);
or U6786 (N_6786,N_5982,N_6214);
or U6787 (N_6787,N_5989,N_6155);
nor U6788 (N_6788,N_6227,N_5670);
and U6789 (N_6789,N_5856,N_5972);
and U6790 (N_6790,N_6119,N_6122);
nor U6791 (N_6791,N_5972,N_5784);
nand U6792 (N_6792,N_5968,N_5912);
or U6793 (N_6793,N_6003,N_6231);
xor U6794 (N_6794,N_5934,N_5638);
nand U6795 (N_6795,N_5800,N_6184);
nand U6796 (N_6796,N_5705,N_6119);
and U6797 (N_6797,N_5670,N_6214);
and U6798 (N_6798,N_5771,N_5869);
or U6799 (N_6799,N_6132,N_5648);
xor U6800 (N_6800,N_5780,N_5734);
and U6801 (N_6801,N_5697,N_5666);
and U6802 (N_6802,N_5917,N_6150);
nor U6803 (N_6803,N_5747,N_5878);
or U6804 (N_6804,N_5800,N_5666);
xor U6805 (N_6805,N_5813,N_5734);
nand U6806 (N_6806,N_5694,N_6120);
or U6807 (N_6807,N_5857,N_5986);
xnor U6808 (N_6808,N_6139,N_5789);
nor U6809 (N_6809,N_6205,N_5831);
nor U6810 (N_6810,N_6223,N_5875);
and U6811 (N_6811,N_6051,N_5907);
and U6812 (N_6812,N_6093,N_6166);
xnor U6813 (N_6813,N_6239,N_6008);
or U6814 (N_6814,N_6019,N_5659);
nor U6815 (N_6815,N_5861,N_6106);
and U6816 (N_6816,N_5790,N_5833);
nor U6817 (N_6817,N_6012,N_5686);
nor U6818 (N_6818,N_6161,N_6217);
nand U6819 (N_6819,N_5966,N_5974);
nor U6820 (N_6820,N_6155,N_5936);
or U6821 (N_6821,N_5701,N_5784);
xnor U6822 (N_6822,N_6014,N_5698);
xnor U6823 (N_6823,N_6239,N_6193);
xnor U6824 (N_6824,N_5977,N_5776);
xnor U6825 (N_6825,N_6135,N_6158);
or U6826 (N_6826,N_6227,N_6135);
nor U6827 (N_6827,N_5756,N_6109);
xnor U6828 (N_6828,N_5907,N_5667);
xnor U6829 (N_6829,N_5881,N_6024);
nor U6830 (N_6830,N_5694,N_5698);
xor U6831 (N_6831,N_5715,N_5890);
nand U6832 (N_6832,N_5708,N_6026);
or U6833 (N_6833,N_5853,N_5714);
and U6834 (N_6834,N_5736,N_6021);
or U6835 (N_6835,N_6164,N_5840);
and U6836 (N_6836,N_6172,N_5645);
xor U6837 (N_6837,N_5896,N_6036);
xor U6838 (N_6838,N_5743,N_5909);
nor U6839 (N_6839,N_6138,N_6243);
or U6840 (N_6840,N_5944,N_5822);
or U6841 (N_6841,N_5718,N_5651);
nand U6842 (N_6842,N_6243,N_5898);
and U6843 (N_6843,N_6112,N_5862);
xor U6844 (N_6844,N_5654,N_6243);
nor U6845 (N_6845,N_5670,N_6016);
nand U6846 (N_6846,N_5755,N_5725);
or U6847 (N_6847,N_5856,N_5703);
nor U6848 (N_6848,N_5686,N_5849);
xnor U6849 (N_6849,N_5961,N_5827);
or U6850 (N_6850,N_5670,N_5889);
nand U6851 (N_6851,N_5866,N_5763);
and U6852 (N_6852,N_5651,N_6119);
xor U6853 (N_6853,N_5865,N_5688);
or U6854 (N_6854,N_5738,N_5940);
nor U6855 (N_6855,N_5741,N_5860);
xor U6856 (N_6856,N_6034,N_6155);
and U6857 (N_6857,N_5860,N_5629);
xnor U6858 (N_6858,N_6146,N_6111);
xnor U6859 (N_6859,N_6103,N_6011);
xnor U6860 (N_6860,N_5787,N_6154);
xor U6861 (N_6861,N_5915,N_6001);
nand U6862 (N_6862,N_6194,N_6220);
nor U6863 (N_6863,N_5749,N_6082);
nor U6864 (N_6864,N_5783,N_5843);
nor U6865 (N_6865,N_5928,N_6052);
nand U6866 (N_6866,N_5952,N_5870);
or U6867 (N_6867,N_5718,N_5768);
xnor U6868 (N_6868,N_5649,N_5774);
xnor U6869 (N_6869,N_6082,N_6216);
and U6870 (N_6870,N_5676,N_6228);
xnor U6871 (N_6871,N_6002,N_6198);
and U6872 (N_6872,N_6204,N_5712);
and U6873 (N_6873,N_5839,N_6182);
and U6874 (N_6874,N_6144,N_5815);
and U6875 (N_6875,N_6474,N_6823);
xnor U6876 (N_6876,N_6802,N_6760);
xnor U6877 (N_6877,N_6560,N_6275);
or U6878 (N_6878,N_6464,N_6412);
xnor U6879 (N_6879,N_6840,N_6589);
xor U6880 (N_6880,N_6576,N_6253);
and U6881 (N_6881,N_6652,N_6252);
nor U6882 (N_6882,N_6684,N_6870);
nand U6883 (N_6883,N_6538,N_6422);
or U6884 (N_6884,N_6764,N_6563);
nand U6885 (N_6885,N_6740,N_6264);
nand U6886 (N_6886,N_6721,N_6568);
or U6887 (N_6887,N_6796,N_6536);
nor U6888 (N_6888,N_6733,N_6850);
nand U6889 (N_6889,N_6393,N_6537);
nand U6890 (N_6890,N_6809,N_6778);
or U6891 (N_6891,N_6658,N_6487);
nand U6892 (N_6892,N_6411,N_6403);
nand U6893 (N_6893,N_6857,N_6708);
nand U6894 (N_6894,N_6803,N_6626);
and U6895 (N_6895,N_6799,N_6292);
nand U6896 (N_6896,N_6552,N_6797);
xnor U6897 (N_6897,N_6468,N_6871);
nand U6898 (N_6898,N_6754,N_6620);
xnor U6899 (N_6899,N_6414,N_6299);
xor U6900 (N_6900,N_6842,N_6555);
and U6901 (N_6901,N_6387,N_6565);
nand U6902 (N_6902,N_6305,N_6321);
or U6903 (N_6903,N_6274,N_6451);
or U6904 (N_6904,N_6250,N_6661);
nor U6905 (N_6905,N_6499,N_6470);
nand U6906 (N_6906,N_6746,N_6554);
or U6907 (N_6907,N_6456,N_6849);
xor U6908 (N_6908,N_6744,N_6524);
or U6909 (N_6909,N_6587,N_6636);
nor U6910 (N_6910,N_6279,N_6435);
xor U6911 (N_6911,N_6845,N_6611);
nor U6912 (N_6912,N_6651,N_6289);
xor U6913 (N_6913,N_6779,N_6866);
or U6914 (N_6914,N_6262,N_6263);
nor U6915 (N_6915,N_6790,N_6513);
nand U6916 (N_6916,N_6401,N_6362);
or U6917 (N_6917,N_6710,N_6374);
or U6918 (N_6918,N_6697,N_6415);
and U6919 (N_6919,N_6325,N_6514);
and U6920 (N_6920,N_6859,N_6648);
nor U6921 (N_6921,N_6404,N_6357);
xnor U6922 (N_6922,N_6476,N_6699);
nand U6923 (N_6923,N_6670,N_6315);
nor U6924 (N_6924,N_6682,N_6355);
or U6925 (N_6925,N_6787,N_6356);
and U6926 (N_6926,N_6344,N_6496);
nand U6927 (N_6927,N_6542,N_6314);
xnor U6928 (N_6928,N_6388,N_6707);
and U6929 (N_6929,N_6385,N_6724);
or U6930 (N_6930,N_6869,N_6683);
and U6931 (N_6931,N_6711,N_6632);
nand U6932 (N_6932,N_6265,N_6665);
or U6933 (N_6933,N_6532,N_6286);
xnor U6934 (N_6934,N_6704,N_6295);
nor U6935 (N_6935,N_6527,N_6692);
nand U6936 (N_6936,N_6772,N_6360);
xor U6937 (N_6937,N_6719,N_6328);
nand U6938 (N_6938,N_6425,N_6673);
xnor U6939 (N_6939,N_6591,N_6465);
or U6940 (N_6940,N_6864,N_6348);
and U6941 (N_6941,N_6698,N_6580);
nor U6942 (N_6942,N_6291,N_6742);
and U6943 (N_6943,N_6782,N_6773);
nor U6944 (N_6944,N_6266,N_6624);
and U6945 (N_6945,N_6302,N_6256);
nand U6946 (N_6946,N_6353,N_6569);
or U6947 (N_6947,N_6361,N_6607);
nor U6948 (N_6948,N_6585,N_6383);
or U6949 (N_6949,N_6453,N_6440);
and U6950 (N_6950,N_6556,N_6365);
nand U6951 (N_6951,N_6756,N_6812);
xnor U6952 (N_6952,N_6418,N_6493);
and U6953 (N_6953,N_6592,N_6805);
nor U6954 (N_6954,N_6663,N_6660);
and U6955 (N_6955,N_6480,N_6460);
and U6956 (N_6956,N_6371,N_6529);
and U6957 (N_6957,N_6329,N_6509);
or U6958 (N_6958,N_6798,N_6466);
or U6959 (N_6959,N_6351,N_6479);
xnor U6960 (N_6960,N_6874,N_6449);
nor U6961 (N_6961,N_6590,N_6347);
nand U6962 (N_6962,N_6671,N_6814);
nor U6963 (N_6963,N_6800,N_6410);
nand U6964 (N_6964,N_6689,N_6614);
nor U6965 (N_6965,N_6825,N_6553);
xor U6966 (N_6966,N_6285,N_6852);
or U6967 (N_6967,N_6830,N_6276);
nor U6968 (N_6968,N_6306,N_6310);
or U6969 (N_6969,N_6363,N_6455);
nor U6970 (N_6970,N_6766,N_6714);
or U6971 (N_6971,N_6584,N_6337);
or U6972 (N_6972,N_6722,N_6634);
or U6973 (N_6973,N_6327,N_6577);
and U6974 (N_6974,N_6533,N_6441);
or U6975 (N_6975,N_6511,N_6677);
nor U6976 (N_6976,N_6503,N_6531);
xnor U6977 (N_6977,N_6312,N_6428);
nor U6978 (N_6978,N_6816,N_6848);
nor U6979 (N_6979,N_6405,N_6561);
nor U6980 (N_6980,N_6334,N_6281);
or U6981 (N_6981,N_6437,N_6745);
and U6982 (N_6982,N_6856,N_6617);
xnor U6983 (N_6983,N_6844,N_6622);
nor U6984 (N_6984,N_6776,N_6510);
nor U6985 (N_6985,N_6432,N_6725);
and U6986 (N_6986,N_6434,N_6680);
or U6987 (N_6987,N_6873,N_6627);
nor U6988 (N_6988,N_6333,N_6841);
and U6989 (N_6989,N_6446,N_6332);
xor U6990 (N_6990,N_6581,N_6664);
and U6991 (N_6991,N_6442,N_6559);
nand U6992 (N_6992,N_6280,N_6331);
nand U6993 (N_6993,N_6349,N_6278);
xnor U6994 (N_6994,N_6458,N_6420);
or U6995 (N_6995,N_6540,N_6771);
or U6996 (N_6996,N_6753,N_6260);
nand U6997 (N_6997,N_6792,N_6755);
xnor U6998 (N_6998,N_6322,N_6400);
nor U6999 (N_6999,N_6272,N_6588);
nor U7000 (N_7000,N_6716,N_6583);
nor U7001 (N_7001,N_6346,N_6824);
nand U7002 (N_7002,N_6427,N_6702);
and U7003 (N_7003,N_6390,N_6368);
nand U7004 (N_7004,N_6734,N_6489);
nand U7005 (N_7005,N_6439,N_6619);
nand U7006 (N_7006,N_6855,N_6737);
nand U7007 (N_7007,N_6654,N_6429);
xor U7008 (N_7008,N_6597,N_6567);
or U7009 (N_7009,N_6793,N_6598);
xor U7010 (N_7010,N_6681,N_6727);
or U7011 (N_7011,N_6672,N_6547);
xnor U7012 (N_7012,N_6463,N_6609);
nand U7013 (N_7013,N_6720,N_6638);
or U7014 (N_7014,N_6775,N_6821);
and U7015 (N_7015,N_6695,N_6324);
xnor U7016 (N_7016,N_6837,N_6717);
and U7017 (N_7017,N_6731,N_6625);
nand U7018 (N_7018,N_6288,N_6656);
xor U7019 (N_7019,N_6868,N_6606);
and U7020 (N_7020,N_6522,N_6495);
nand U7021 (N_7021,N_6646,N_6732);
xor U7022 (N_7022,N_6574,N_6340);
or U7023 (N_7023,N_6718,N_6501);
nor U7024 (N_7024,N_6573,N_6795);
nand U7025 (N_7025,N_6558,N_6688);
xor U7026 (N_7026,N_6623,N_6268);
xor U7027 (N_7027,N_6743,N_6467);
nor U7028 (N_7028,N_6438,N_6788);
or U7029 (N_7029,N_6398,N_6525);
nor U7030 (N_7030,N_6271,N_6251);
or U7031 (N_7031,N_6596,N_6369);
nand U7032 (N_7032,N_6431,N_6486);
nand U7033 (N_7033,N_6535,N_6748);
nand U7034 (N_7034,N_6762,N_6785);
or U7035 (N_7035,N_6655,N_6381);
nand U7036 (N_7036,N_6639,N_6594);
xor U7037 (N_7037,N_6863,N_6784);
nand U7038 (N_7038,N_6459,N_6818);
nor U7039 (N_7039,N_6872,N_6804);
or U7040 (N_7040,N_6336,N_6450);
nand U7041 (N_7041,N_6701,N_6502);
or U7042 (N_7042,N_6444,N_6736);
or U7043 (N_7043,N_6436,N_6354);
and U7044 (N_7044,N_6515,N_6382);
nor U7045 (N_7045,N_6578,N_6657);
nand U7046 (N_7046,N_6376,N_6696);
nand U7047 (N_7047,N_6575,N_6300);
xor U7048 (N_7048,N_6618,N_6367);
or U7049 (N_7049,N_6723,N_6423);
nand U7050 (N_7050,N_6297,N_6603);
xor U7051 (N_7051,N_6323,N_6482);
or U7052 (N_7052,N_6298,N_6497);
nand U7053 (N_7053,N_6526,N_6506);
xnor U7054 (N_7054,N_6765,N_6786);
or U7055 (N_7055,N_6508,N_6811);
and U7056 (N_7056,N_6339,N_6666);
nand U7057 (N_7057,N_6481,N_6758);
xor U7058 (N_7058,N_6254,N_6473);
and U7059 (N_7059,N_6582,N_6330);
and U7060 (N_7060,N_6518,N_6301);
nor U7061 (N_7061,N_6320,N_6649);
xor U7062 (N_7062,N_6676,N_6342);
xnor U7063 (N_7063,N_6426,N_6570);
nor U7064 (N_7064,N_6548,N_6728);
nor U7065 (N_7065,N_6392,N_6386);
or U7066 (N_7066,N_6685,N_6512);
nor U7067 (N_7067,N_6507,N_6359);
and U7068 (N_7068,N_6729,N_6551);
nand U7069 (N_7069,N_6546,N_6862);
xor U7070 (N_7070,N_6396,N_6579);
xnor U7071 (N_7071,N_6693,N_6806);
or U7072 (N_7072,N_6421,N_6475);
nand U7073 (N_7073,N_6854,N_6599);
or U7074 (N_7074,N_6366,N_6621);
nor U7075 (N_7075,N_6452,N_6308);
and U7076 (N_7076,N_6377,N_6601);
xor U7077 (N_7077,N_6703,N_6768);
nand U7078 (N_7078,N_6832,N_6303);
nand U7079 (N_7079,N_6774,N_6761);
nand U7080 (N_7080,N_6541,N_6343);
nor U7081 (N_7081,N_6759,N_6307);
nor U7082 (N_7082,N_6605,N_6491);
xor U7083 (N_7083,N_6447,N_6813);
xor U7084 (N_7084,N_6678,N_6726);
xnor U7085 (N_7085,N_6822,N_6853);
nor U7086 (N_7086,N_6416,N_6640);
xor U7087 (N_7087,N_6741,N_6494);
and U7088 (N_7088,N_6647,N_6397);
and U7089 (N_7089,N_6867,N_6687);
xor U7090 (N_7090,N_6642,N_6767);
nand U7091 (N_7091,N_6738,N_6523);
or U7092 (N_7092,N_6549,N_6282);
or U7093 (N_7093,N_6408,N_6375);
nand U7094 (N_7094,N_6338,N_6694);
or U7095 (N_7095,N_6739,N_6690);
xnor U7096 (N_7096,N_6769,N_6828);
xor U7097 (N_7097,N_6613,N_6443);
nor U7098 (N_7098,N_6835,N_6600);
nor U7099 (N_7099,N_6630,N_6808);
and U7100 (N_7100,N_6820,N_6372);
and U7101 (N_7101,N_6571,N_6335);
xor U7102 (N_7102,N_6843,N_6662);
nor U7103 (N_7103,N_6653,N_6311);
xor U7104 (N_7104,N_6261,N_6545);
nor U7105 (N_7105,N_6277,N_6430);
xor U7106 (N_7106,N_6750,N_6604);
nor U7107 (N_7107,N_6516,N_6419);
and U7108 (N_7108,N_6586,N_6394);
xnor U7109 (N_7109,N_6273,N_6564);
nor U7110 (N_7110,N_6602,N_6500);
nand U7111 (N_7111,N_6341,N_6712);
or U7112 (N_7112,N_6608,N_6316);
nand U7113 (N_7113,N_6395,N_6829);
nand U7114 (N_7114,N_6705,N_6478);
xnor U7115 (N_7115,N_6294,N_6259);
nand U7116 (N_7116,N_6833,N_6402);
and U7117 (N_7117,N_6817,N_6424);
nand U7118 (N_7118,N_6836,N_6783);
or U7119 (N_7119,N_6706,N_6700);
or U7120 (N_7120,N_6629,N_6448);
xnor U7121 (N_7121,N_6650,N_6675);
nor U7122 (N_7122,N_6409,N_6757);
nand U7123 (N_7123,N_6645,N_6407);
xor U7124 (N_7124,N_6637,N_6490);
xnor U7125 (N_7125,N_6378,N_6595);
xor U7126 (N_7126,N_6815,N_6257);
nand U7127 (N_7127,N_6807,N_6296);
xor U7128 (N_7128,N_6631,N_6370);
or U7129 (N_7129,N_6484,N_6319);
and U7130 (N_7130,N_6287,N_6454);
or U7131 (N_7131,N_6827,N_6667);
and U7132 (N_7132,N_6747,N_6794);
nand U7133 (N_7133,N_6643,N_6462);
nand U7134 (N_7134,N_6483,N_6635);
nor U7135 (N_7135,N_6399,N_6530);
nor U7136 (N_7136,N_6358,N_6612);
nand U7137 (N_7137,N_6528,N_6544);
or U7138 (N_7138,N_6477,N_6749);
xor U7139 (N_7139,N_6520,N_6610);
xnor U7140 (N_7140,N_6615,N_6679);
nand U7141 (N_7141,N_6593,N_6364);
xnor U7142 (N_7142,N_6770,N_6838);
nand U7143 (N_7143,N_6566,N_6686);
xnor U7144 (N_7144,N_6290,N_6391);
and U7145 (N_7145,N_6457,N_6534);
nor U7146 (N_7146,N_6819,N_6669);
nand U7147 (N_7147,N_6562,N_6269);
and U7148 (N_7148,N_6735,N_6791);
nor U7149 (N_7149,N_6293,N_6270);
xor U7150 (N_7150,N_6846,N_6267);
xnor U7151 (N_7151,N_6550,N_6860);
and U7152 (N_7152,N_6763,N_6709);
xnor U7153 (N_7153,N_6413,N_6461);
xnor U7154 (N_7154,N_6557,N_6539);
nor U7155 (N_7155,N_6752,N_6644);
xnor U7156 (N_7156,N_6839,N_6313);
nor U7157 (N_7157,N_6668,N_6380);
nand U7158 (N_7158,N_6831,N_6826);
xnor U7159 (N_7159,N_6345,N_6781);
or U7160 (N_7160,N_6352,N_6674);
and U7161 (N_7161,N_6284,N_6713);
and U7162 (N_7162,N_6801,N_6505);
nor U7163 (N_7163,N_6572,N_6730);
nor U7164 (N_7164,N_6751,N_6258);
xnor U7165 (N_7165,N_6858,N_6659);
xor U7166 (N_7166,N_6304,N_6789);
or U7167 (N_7167,N_6847,N_6488);
or U7168 (N_7168,N_6384,N_6255);
or U7169 (N_7169,N_6445,N_6715);
and U7170 (N_7170,N_6691,N_6326);
xnor U7171 (N_7171,N_6317,N_6472);
nor U7172 (N_7172,N_6641,N_6318);
nand U7173 (N_7173,N_6373,N_6471);
or U7174 (N_7174,N_6633,N_6543);
and U7175 (N_7175,N_6389,N_6616);
or U7176 (N_7176,N_6834,N_6417);
or U7177 (N_7177,N_6350,N_6517);
and U7178 (N_7178,N_6469,N_6406);
xor U7179 (N_7179,N_6810,N_6433);
and U7180 (N_7180,N_6521,N_6519);
xor U7181 (N_7181,N_6498,N_6851);
or U7182 (N_7182,N_6861,N_6628);
xor U7183 (N_7183,N_6485,N_6777);
and U7184 (N_7184,N_6865,N_6780);
or U7185 (N_7185,N_6492,N_6283);
and U7186 (N_7186,N_6379,N_6309);
nand U7187 (N_7187,N_6504,N_6310);
xor U7188 (N_7188,N_6655,N_6657);
and U7189 (N_7189,N_6837,N_6297);
or U7190 (N_7190,N_6496,N_6690);
xor U7191 (N_7191,N_6336,N_6657);
nor U7192 (N_7192,N_6488,N_6427);
xnor U7193 (N_7193,N_6445,N_6689);
nor U7194 (N_7194,N_6451,N_6533);
and U7195 (N_7195,N_6806,N_6553);
nand U7196 (N_7196,N_6674,N_6718);
or U7197 (N_7197,N_6574,N_6667);
and U7198 (N_7198,N_6463,N_6802);
xnor U7199 (N_7199,N_6546,N_6674);
nor U7200 (N_7200,N_6826,N_6382);
or U7201 (N_7201,N_6441,N_6520);
or U7202 (N_7202,N_6587,N_6738);
xor U7203 (N_7203,N_6782,N_6860);
and U7204 (N_7204,N_6786,N_6250);
nand U7205 (N_7205,N_6311,N_6316);
nor U7206 (N_7206,N_6412,N_6324);
nor U7207 (N_7207,N_6781,N_6459);
and U7208 (N_7208,N_6319,N_6273);
and U7209 (N_7209,N_6802,N_6805);
and U7210 (N_7210,N_6254,N_6853);
nor U7211 (N_7211,N_6614,N_6432);
and U7212 (N_7212,N_6745,N_6606);
or U7213 (N_7213,N_6354,N_6630);
nor U7214 (N_7214,N_6337,N_6680);
nand U7215 (N_7215,N_6711,N_6433);
nand U7216 (N_7216,N_6259,N_6600);
or U7217 (N_7217,N_6454,N_6473);
and U7218 (N_7218,N_6256,N_6463);
or U7219 (N_7219,N_6782,N_6367);
nand U7220 (N_7220,N_6403,N_6454);
and U7221 (N_7221,N_6258,N_6686);
nand U7222 (N_7222,N_6324,N_6573);
nor U7223 (N_7223,N_6421,N_6873);
nand U7224 (N_7224,N_6646,N_6596);
xor U7225 (N_7225,N_6864,N_6297);
and U7226 (N_7226,N_6292,N_6725);
or U7227 (N_7227,N_6293,N_6654);
nor U7228 (N_7228,N_6412,N_6549);
nand U7229 (N_7229,N_6760,N_6831);
and U7230 (N_7230,N_6582,N_6300);
nand U7231 (N_7231,N_6795,N_6683);
nand U7232 (N_7232,N_6615,N_6744);
or U7233 (N_7233,N_6763,N_6470);
or U7234 (N_7234,N_6534,N_6460);
nor U7235 (N_7235,N_6723,N_6874);
xor U7236 (N_7236,N_6853,N_6860);
or U7237 (N_7237,N_6550,N_6521);
nor U7238 (N_7238,N_6523,N_6531);
nand U7239 (N_7239,N_6829,N_6765);
nand U7240 (N_7240,N_6714,N_6399);
nand U7241 (N_7241,N_6426,N_6319);
xor U7242 (N_7242,N_6643,N_6390);
and U7243 (N_7243,N_6706,N_6688);
or U7244 (N_7244,N_6297,N_6289);
or U7245 (N_7245,N_6714,N_6293);
or U7246 (N_7246,N_6613,N_6457);
and U7247 (N_7247,N_6603,N_6729);
and U7248 (N_7248,N_6257,N_6704);
and U7249 (N_7249,N_6838,N_6702);
nand U7250 (N_7250,N_6580,N_6791);
or U7251 (N_7251,N_6614,N_6767);
or U7252 (N_7252,N_6258,N_6687);
nand U7253 (N_7253,N_6836,N_6323);
nand U7254 (N_7254,N_6755,N_6693);
or U7255 (N_7255,N_6260,N_6695);
and U7256 (N_7256,N_6329,N_6577);
xnor U7257 (N_7257,N_6293,N_6702);
or U7258 (N_7258,N_6851,N_6355);
nand U7259 (N_7259,N_6534,N_6707);
xnor U7260 (N_7260,N_6428,N_6744);
or U7261 (N_7261,N_6594,N_6526);
nor U7262 (N_7262,N_6856,N_6272);
and U7263 (N_7263,N_6451,N_6302);
nand U7264 (N_7264,N_6787,N_6529);
nand U7265 (N_7265,N_6772,N_6749);
xor U7266 (N_7266,N_6601,N_6367);
xor U7267 (N_7267,N_6821,N_6582);
xor U7268 (N_7268,N_6400,N_6682);
xor U7269 (N_7269,N_6529,N_6279);
nor U7270 (N_7270,N_6475,N_6337);
or U7271 (N_7271,N_6476,N_6744);
nand U7272 (N_7272,N_6862,N_6748);
and U7273 (N_7273,N_6376,N_6728);
nor U7274 (N_7274,N_6824,N_6745);
nor U7275 (N_7275,N_6864,N_6482);
or U7276 (N_7276,N_6739,N_6405);
nor U7277 (N_7277,N_6778,N_6796);
and U7278 (N_7278,N_6665,N_6439);
xnor U7279 (N_7279,N_6491,N_6562);
and U7280 (N_7280,N_6372,N_6426);
xor U7281 (N_7281,N_6605,N_6503);
nand U7282 (N_7282,N_6449,N_6765);
nand U7283 (N_7283,N_6591,N_6857);
xnor U7284 (N_7284,N_6613,N_6285);
or U7285 (N_7285,N_6291,N_6833);
and U7286 (N_7286,N_6490,N_6555);
nor U7287 (N_7287,N_6722,N_6304);
nor U7288 (N_7288,N_6432,N_6645);
nor U7289 (N_7289,N_6481,N_6662);
and U7290 (N_7290,N_6676,N_6752);
nand U7291 (N_7291,N_6677,N_6691);
nor U7292 (N_7292,N_6410,N_6545);
xnor U7293 (N_7293,N_6287,N_6752);
xor U7294 (N_7294,N_6704,N_6860);
nor U7295 (N_7295,N_6604,N_6379);
or U7296 (N_7296,N_6314,N_6312);
xnor U7297 (N_7297,N_6265,N_6530);
and U7298 (N_7298,N_6252,N_6583);
nand U7299 (N_7299,N_6716,N_6669);
nor U7300 (N_7300,N_6792,N_6396);
nor U7301 (N_7301,N_6756,N_6751);
nand U7302 (N_7302,N_6801,N_6484);
nor U7303 (N_7303,N_6756,N_6517);
nor U7304 (N_7304,N_6477,N_6482);
nand U7305 (N_7305,N_6682,N_6508);
and U7306 (N_7306,N_6541,N_6252);
nor U7307 (N_7307,N_6579,N_6635);
nand U7308 (N_7308,N_6829,N_6259);
nor U7309 (N_7309,N_6328,N_6653);
nor U7310 (N_7310,N_6512,N_6450);
and U7311 (N_7311,N_6847,N_6558);
nand U7312 (N_7312,N_6442,N_6738);
and U7313 (N_7313,N_6426,N_6754);
or U7314 (N_7314,N_6783,N_6811);
and U7315 (N_7315,N_6861,N_6577);
and U7316 (N_7316,N_6750,N_6786);
nand U7317 (N_7317,N_6810,N_6425);
nor U7318 (N_7318,N_6755,N_6860);
and U7319 (N_7319,N_6490,N_6642);
nand U7320 (N_7320,N_6854,N_6519);
nor U7321 (N_7321,N_6263,N_6487);
nand U7322 (N_7322,N_6455,N_6292);
or U7323 (N_7323,N_6678,N_6389);
nor U7324 (N_7324,N_6850,N_6599);
xnor U7325 (N_7325,N_6845,N_6412);
or U7326 (N_7326,N_6309,N_6700);
and U7327 (N_7327,N_6803,N_6710);
nand U7328 (N_7328,N_6553,N_6529);
or U7329 (N_7329,N_6440,N_6562);
or U7330 (N_7330,N_6394,N_6458);
nand U7331 (N_7331,N_6369,N_6419);
or U7332 (N_7332,N_6319,N_6404);
nor U7333 (N_7333,N_6279,N_6338);
nor U7334 (N_7334,N_6478,N_6330);
or U7335 (N_7335,N_6660,N_6833);
and U7336 (N_7336,N_6400,N_6804);
or U7337 (N_7337,N_6372,N_6343);
nand U7338 (N_7338,N_6630,N_6552);
xor U7339 (N_7339,N_6758,N_6651);
or U7340 (N_7340,N_6394,N_6390);
and U7341 (N_7341,N_6294,N_6836);
and U7342 (N_7342,N_6440,N_6334);
nor U7343 (N_7343,N_6400,N_6526);
xnor U7344 (N_7344,N_6407,N_6847);
and U7345 (N_7345,N_6364,N_6324);
xnor U7346 (N_7346,N_6754,N_6319);
nor U7347 (N_7347,N_6529,N_6483);
and U7348 (N_7348,N_6516,N_6253);
xor U7349 (N_7349,N_6525,N_6661);
or U7350 (N_7350,N_6871,N_6745);
and U7351 (N_7351,N_6486,N_6282);
nor U7352 (N_7352,N_6775,N_6719);
xnor U7353 (N_7353,N_6403,N_6286);
xor U7354 (N_7354,N_6254,N_6586);
and U7355 (N_7355,N_6751,N_6327);
or U7356 (N_7356,N_6457,N_6873);
or U7357 (N_7357,N_6364,N_6392);
and U7358 (N_7358,N_6542,N_6769);
nand U7359 (N_7359,N_6297,N_6649);
nor U7360 (N_7360,N_6390,N_6433);
xor U7361 (N_7361,N_6466,N_6838);
nor U7362 (N_7362,N_6385,N_6689);
nor U7363 (N_7363,N_6681,N_6687);
or U7364 (N_7364,N_6451,N_6398);
xnor U7365 (N_7365,N_6648,N_6420);
nor U7366 (N_7366,N_6664,N_6365);
nor U7367 (N_7367,N_6355,N_6416);
nor U7368 (N_7368,N_6408,N_6539);
and U7369 (N_7369,N_6849,N_6498);
nand U7370 (N_7370,N_6647,N_6652);
nor U7371 (N_7371,N_6571,N_6728);
xnor U7372 (N_7372,N_6702,N_6707);
or U7373 (N_7373,N_6323,N_6569);
nor U7374 (N_7374,N_6669,N_6414);
xor U7375 (N_7375,N_6591,N_6370);
or U7376 (N_7376,N_6387,N_6293);
nor U7377 (N_7377,N_6569,N_6543);
and U7378 (N_7378,N_6869,N_6544);
nand U7379 (N_7379,N_6817,N_6680);
and U7380 (N_7380,N_6668,N_6549);
nor U7381 (N_7381,N_6348,N_6369);
and U7382 (N_7382,N_6416,N_6338);
nand U7383 (N_7383,N_6712,N_6540);
xnor U7384 (N_7384,N_6318,N_6560);
xor U7385 (N_7385,N_6491,N_6683);
nand U7386 (N_7386,N_6463,N_6286);
or U7387 (N_7387,N_6446,N_6360);
nor U7388 (N_7388,N_6592,N_6715);
nor U7389 (N_7389,N_6652,N_6745);
xor U7390 (N_7390,N_6270,N_6532);
or U7391 (N_7391,N_6694,N_6807);
and U7392 (N_7392,N_6405,N_6449);
nand U7393 (N_7393,N_6645,N_6745);
nor U7394 (N_7394,N_6711,N_6552);
or U7395 (N_7395,N_6579,N_6870);
or U7396 (N_7396,N_6584,N_6757);
xnor U7397 (N_7397,N_6747,N_6659);
nand U7398 (N_7398,N_6457,N_6274);
nor U7399 (N_7399,N_6369,N_6796);
nor U7400 (N_7400,N_6312,N_6265);
nor U7401 (N_7401,N_6670,N_6399);
nor U7402 (N_7402,N_6665,N_6299);
nand U7403 (N_7403,N_6259,N_6718);
nor U7404 (N_7404,N_6816,N_6461);
nand U7405 (N_7405,N_6449,N_6850);
nor U7406 (N_7406,N_6306,N_6263);
xnor U7407 (N_7407,N_6298,N_6674);
or U7408 (N_7408,N_6821,N_6839);
nand U7409 (N_7409,N_6839,N_6792);
xnor U7410 (N_7410,N_6432,N_6436);
xnor U7411 (N_7411,N_6757,N_6504);
or U7412 (N_7412,N_6793,N_6794);
or U7413 (N_7413,N_6762,N_6419);
nor U7414 (N_7414,N_6864,N_6645);
or U7415 (N_7415,N_6384,N_6563);
nand U7416 (N_7416,N_6785,N_6544);
xor U7417 (N_7417,N_6719,N_6817);
or U7418 (N_7418,N_6347,N_6831);
or U7419 (N_7419,N_6362,N_6696);
and U7420 (N_7420,N_6275,N_6385);
xor U7421 (N_7421,N_6855,N_6685);
xnor U7422 (N_7422,N_6735,N_6658);
or U7423 (N_7423,N_6786,N_6793);
nor U7424 (N_7424,N_6335,N_6811);
nand U7425 (N_7425,N_6474,N_6696);
and U7426 (N_7426,N_6525,N_6772);
nand U7427 (N_7427,N_6578,N_6821);
nand U7428 (N_7428,N_6262,N_6723);
xnor U7429 (N_7429,N_6750,N_6399);
or U7430 (N_7430,N_6723,N_6259);
nor U7431 (N_7431,N_6764,N_6631);
and U7432 (N_7432,N_6394,N_6342);
nand U7433 (N_7433,N_6468,N_6252);
xor U7434 (N_7434,N_6824,N_6292);
nand U7435 (N_7435,N_6280,N_6419);
xnor U7436 (N_7436,N_6272,N_6645);
xnor U7437 (N_7437,N_6320,N_6849);
nand U7438 (N_7438,N_6792,N_6535);
or U7439 (N_7439,N_6824,N_6641);
xor U7440 (N_7440,N_6747,N_6538);
and U7441 (N_7441,N_6637,N_6778);
xnor U7442 (N_7442,N_6578,N_6543);
nor U7443 (N_7443,N_6282,N_6661);
nor U7444 (N_7444,N_6318,N_6738);
or U7445 (N_7445,N_6517,N_6853);
nand U7446 (N_7446,N_6329,N_6756);
or U7447 (N_7447,N_6472,N_6364);
nand U7448 (N_7448,N_6766,N_6404);
or U7449 (N_7449,N_6444,N_6730);
nand U7450 (N_7450,N_6727,N_6660);
and U7451 (N_7451,N_6322,N_6682);
or U7452 (N_7452,N_6842,N_6854);
nand U7453 (N_7453,N_6662,N_6635);
or U7454 (N_7454,N_6610,N_6835);
or U7455 (N_7455,N_6867,N_6806);
and U7456 (N_7456,N_6802,N_6776);
nand U7457 (N_7457,N_6465,N_6311);
xnor U7458 (N_7458,N_6415,N_6625);
xor U7459 (N_7459,N_6836,N_6478);
nor U7460 (N_7460,N_6677,N_6628);
or U7461 (N_7461,N_6541,N_6402);
xnor U7462 (N_7462,N_6433,N_6435);
xor U7463 (N_7463,N_6495,N_6464);
or U7464 (N_7464,N_6313,N_6743);
or U7465 (N_7465,N_6372,N_6752);
and U7466 (N_7466,N_6785,N_6645);
xnor U7467 (N_7467,N_6443,N_6580);
nand U7468 (N_7468,N_6714,N_6408);
xnor U7469 (N_7469,N_6464,N_6473);
nor U7470 (N_7470,N_6694,N_6490);
nand U7471 (N_7471,N_6617,N_6458);
and U7472 (N_7472,N_6496,N_6270);
nor U7473 (N_7473,N_6534,N_6577);
and U7474 (N_7474,N_6858,N_6800);
or U7475 (N_7475,N_6335,N_6341);
nor U7476 (N_7476,N_6709,N_6856);
and U7477 (N_7477,N_6348,N_6796);
or U7478 (N_7478,N_6686,N_6487);
or U7479 (N_7479,N_6323,N_6530);
and U7480 (N_7480,N_6321,N_6374);
nor U7481 (N_7481,N_6460,N_6763);
or U7482 (N_7482,N_6651,N_6418);
and U7483 (N_7483,N_6279,N_6772);
nand U7484 (N_7484,N_6729,N_6776);
or U7485 (N_7485,N_6336,N_6603);
and U7486 (N_7486,N_6712,N_6475);
nor U7487 (N_7487,N_6702,N_6691);
or U7488 (N_7488,N_6604,N_6484);
xor U7489 (N_7489,N_6293,N_6839);
xnor U7490 (N_7490,N_6477,N_6467);
nand U7491 (N_7491,N_6426,N_6490);
xnor U7492 (N_7492,N_6677,N_6736);
and U7493 (N_7493,N_6687,N_6713);
and U7494 (N_7494,N_6704,N_6857);
and U7495 (N_7495,N_6713,N_6654);
xnor U7496 (N_7496,N_6657,N_6741);
or U7497 (N_7497,N_6514,N_6464);
nor U7498 (N_7498,N_6777,N_6725);
or U7499 (N_7499,N_6350,N_6781);
or U7500 (N_7500,N_7001,N_7223);
nor U7501 (N_7501,N_7179,N_7258);
and U7502 (N_7502,N_7371,N_7076);
or U7503 (N_7503,N_7364,N_6928);
nor U7504 (N_7504,N_7286,N_7447);
nand U7505 (N_7505,N_6984,N_7302);
nor U7506 (N_7506,N_7180,N_7226);
xnor U7507 (N_7507,N_7466,N_7003);
or U7508 (N_7508,N_7240,N_6967);
nor U7509 (N_7509,N_7341,N_7314);
nor U7510 (N_7510,N_7396,N_7196);
nor U7511 (N_7511,N_7279,N_7126);
or U7512 (N_7512,N_6931,N_7122);
nand U7513 (N_7513,N_7351,N_7113);
or U7514 (N_7514,N_7084,N_6917);
nand U7515 (N_7515,N_7205,N_7343);
nand U7516 (N_7516,N_7170,N_7451);
nand U7517 (N_7517,N_6882,N_7441);
xor U7518 (N_7518,N_7337,N_7212);
nor U7519 (N_7519,N_7339,N_7317);
nand U7520 (N_7520,N_6976,N_7164);
and U7521 (N_7521,N_7020,N_7190);
or U7522 (N_7522,N_7008,N_7292);
nand U7523 (N_7523,N_7407,N_7257);
nand U7524 (N_7524,N_7499,N_7335);
nand U7525 (N_7525,N_7347,N_7215);
or U7526 (N_7526,N_7024,N_7022);
nand U7527 (N_7527,N_7385,N_7108);
and U7528 (N_7528,N_7038,N_7181);
or U7529 (N_7529,N_7394,N_7437);
and U7530 (N_7530,N_7442,N_7333);
xor U7531 (N_7531,N_7231,N_7019);
nor U7532 (N_7532,N_7141,N_7493);
nand U7533 (N_7533,N_7117,N_7089);
or U7534 (N_7534,N_7267,N_7209);
nand U7535 (N_7535,N_7206,N_7485);
and U7536 (N_7536,N_6956,N_7046);
nand U7537 (N_7537,N_6914,N_7112);
nor U7538 (N_7538,N_7497,N_7092);
nor U7539 (N_7539,N_7438,N_7390);
and U7540 (N_7540,N_7366,N_7289);
nand U7541 (N_7541,N_7102,N_6909);
or U7542 (N_7542,N_7430,N_7344);
xnor U7543 (N_7543,N_6966,N_7176);
xnor U7544 (N_7544,N_7077,N_7406);
xnor U7545 (N_7545,N_7210,N_7177);
nor U7546 (N_7546,N_6968,N_7266);
xor U7547 (N_7547,N_7027,N_7376);
xnor U7548 (N_7548,N_7080,N_7250);
or U7549 (N_7549,N_6959,N_6972);
and U7550 (N_7550,N_7489,N_7459);
and U7551 (N_7551,N_6985,N_6905);
and U7552 (N_7552,N_6901,N_7326);
or U7553 (N_7553,N_7203,N_7247);
or U7554 (N_7554,N_6925,N_7048);
and U7555 (N_7555,N_7373,N_6918);
xor U7556 (N_7556,N_7241,N_7290);
nor U7557 (N_7557,N_7086,N_6915);
and U7558 (N_7558,N_6963,N_7152);
xor U7559 (N_7559,N_7197,N_6937);
and U7560 (N_7560,N_6907,N_7041);
nor U7561 (N_7561,N_7032,N_7487);
and U7562 (N_7562,N_7349,N_7051);
and U7563 (N_7563,N_7370,N_7475);
and U7564 (N_7564,N_6981,N_7011);
or U7565 (N_7565,N_7356,N_7143);
and U7566 (N_7566,N_6897,N_6975);
nor U7567 (N_7567,N_7061,N_7418);
or U7568 (N_7568,N_7060,N_7204);
nor U7569 (N_7569,N_7228,N_6886);
and U7570 (N_7570,N_7275,N_6900);
xor U7571 (N_7571,N_6879,N_6932);
nand U7572 (N_7572,N_7098,N_7220);
and U7573 (N_7573,N_7105,N_7276);
or U7574 (N_7574,N_7156,N_7169);
nand U7575 (N_7575,N_6883,N_7272);
and U7576 (N_7576,N_6916,N_7194);
and U7577 (N_7577,N_7382,N_7303);
xor U7578 (N_7578,N_6934,N_7054);
or U7579 (N_7579,N_7449,N_6933);
or U7580 (N_7580,N_7414,N_7182);
nand U7581 (N_7581,N_7053,N_7118);
xor U7582 (N_7582,N_7318,N_7386);
nor U7583 (N_7583,N_7033,N_7191);
nor U7584 (N_7584,N_7184,N_7433);
nand U7585 (N_7585,N_7104,N_6876);
nand U7586 (N_7586,N_7288,N_7448);
nor U7587 (N_7587,N_7144,N_7171);
xor U7588 (N_7588,N_7109,N_7021);
xnor U7589 (N_7589,N_6941,N_7026);
xnor U7590 (N_7590,N_7238,N_7149);
and U7591 (N_7591,N_7012,N_7165);
nor U7592 (N_7592,N_7239,N_7101);
nor U7593 (N_7593,N_7100,N_7132);
nor U7594 (N_7594,N_7476,N_7484);
nor U7595 (N_7595,N_7235,N_7013);
and U7596 (N_7596,N_7059,N_7273);
or U7597 (N_7597,N_7178,N_7488);
and U7598 (N_7598,N_6908,N_7455);
and U7599 (N_7599,N_7221,N_6880);
nand U7600 (N_7600,N_7227,N_7408);
nor U7601 (N_7601,N_7157,N_6919);
nand U7602 (N_7602,N_7047,N_7062);
or U7603 (N_7603,N_7262,N_7270);
xor U7604 (N_7604,N_7265,N_7103);
xnor U7605 (N_7605,N_7316,N_7444);
xnor U7606 (N_7606,N_7142,N_6904);
xnor U7607 (N_7607,N_7417,N_7123);
nor U7608 (N_7608,N_7049,N_7342);
and U7609 (N_7609,N_7137,N_7387);
and U7610 (N_7610,N_7055,N_7261);
nor U7611 (N_7611,N_6877,N_6993);
nor U7612 (N_7612,N_7116,N_7357);
or U7613 (N_7613,N_7217,N_7065);
xnor U7614 (N_7614,N_7378,N_7461);
nor U7615 (N_7615,N_7242,N_7007);
nor U7616 (N_7616,N_6962,N_7307);
xor U7617 (N_7617,N_7148,N_6930);
and U7618 (N_7618,N_7355,N_7099);
nand U7619 (N_7619,N_6983,N_7078);
or U7620 (N_7620,N_6978,N_7293);
and U7621 (N_7621,N_7374,N_7167);
or U7622 (N_7622,N_7482,N_7473);
nor U7623 (N_7623,N_6952,N_7070);
nor U7624 (N_7624,N_7249,N_6960);
nand U7625 (N_7625,N_7398,N_7492);
and U7626 (N_7626,N_6923,N_7480);
or U7627 (N_7627,N_7000,N_7134);
xor U7628 (N_7628,N_6958,N_7395);
and U7629 (N_7629,N_7229,N_7338);
nor U7630 (N_7630,N_7224,N_7006);
xnor U7631 (N_7631,N_7172,N_7423);
xnor U7632 (N_7632,N_7422,N_7346);
nand U7633 (N_7633,N_7068,N_7236);
xor U7634 (N_7634,N_6935,N_7472);
or U7635 (N_7635,N_7151,N_7133);
xor U7636 (N_7636,N_7067,N_7173);
xor U7637 (N_7637,N_7413,N_6986);
nand U7638 (N_7638,N_7427,N_7491);
xnor U7639 (N_7639,N_7363,N_6954);
and U7640 (N_7640,N_6940,N_7096);
and U7641 (N_7641,N_7309,N_7158);
xor U7642 (N_7642,N_7434,N_7034);
xor U7643 (N_7643,N_7478,N_7463);
nand U7644 (N_7644,N_7028,N_7120);
nor U7645 (N_7645,N_7277,N_6944);
xnor U7646 (N_7646,N_7097,N_7345);
xnor U7647 (N_7647,N_7075,N_6903);
xor U7648 (N_7648,N_7446,N_6911);
nor U7649 (N_7649,N_7439,N_6949);
nor U7650 (N_7650,N_7160,N_6996);
and U7651 (N_7651,N_6979,N_7017);
nand U7652 (N_7652,N_7256,N_6957);
nor U7653 (N_7653,N_7403,N_7308);
nand U7654 (N_7654,N_7232,N_7321);
nor U7655 (N_7655,N_7009,N_7483);
nor U7656 (N_7656,N_7271,N_7029);
and U7657 (N_7657,N_6999,N_7411);
xor U7658 (N_7658,N_7083,N_6946);
or U7659 (N_7659,N_7297,N_6898);
or U7660 (N_7660,N_7090,N_7462);
and U7661 (N_7661,N_7018,N_7107);
nor U7662 (N_7662,N_7243,N_7136);
xnor U7663 (N_7663,N_6938,N_7052);
xnor U7664 (N_7664,N_7435,N_7336);
nor U7665 (N_7665,N_6955,N_7031);
nand U7666 (N_7666,N_6973,N_7058);
xnor U7667 (N_7667,N_7352,N_7319);
xor U7668 (N_7668,N_7081,N_7381);
and U7669 (N_7669,N_6910,N_7340);
xnor U7670 (N_7670,N_7495,N_7313);
nand U7671 (N_7671,N_7150,N_6939);
and U7672 (N_7672,N_7311,N_7274);
nor U7673 (N_7673,N_7044,N_6922);
xor U7674 (N_7674,N_7372,N_7332);
xnor U7675 (N_7675,N_7004,N_7071);
or U7676 (N_7676,N_7014,N_7079);
or U7677 (N_7677,N_7384,N_7399);
and U7678 (N_7678,N_7361,N_7379);
xor U7679 (N_7679,N_7131,N_7481);
nor U7680 (N_7680,N_7025,N_7207);
or U7681 (N_7681,N_7329,N_6961);
nor U7682 (N_7682,N_7404,N_7425);
or U7683 (N_7683,N_7436,N_7320);
nand U7684 (N_7684,N_6991,N_7431);
or U7685 (N_7685,N_7416,N_7278);
and U7686 (N_7686,N_7315,N_6893);
xnor U7687 (N_7687,N_7216,N_7168);
nor U7688 (N_7688,N_7082,N_6950);
xor U7689 (N_7689,N_7244,N_7036);
nand U7690 (N_7690,N_6990,N_7260);
and U7691 (N_7691,N_7063,N_7147);
nand U7692 (N_7692,N_7002,N_7045);
and U7693 (N_7693,N_7299,N_6936);
and U7694 (N_7694,N_6974,N_7193);
nand U7695 (N_7695,N_6943,N_7445);
or U7696 (N_7696,N_7305,N_7187);
or U7697 (N_7697,N_6989,N_7095);
or U7698 (N_7698,N_7405,N_7400);
and U7699 (N_7699,N_7354,N_7331);
nand U7700 (N_7700,N_7312,N_7469);
and U7701 (N_7701,N_7161,N_7353);
or U7702 (N_7702,N_7456,N_7162);
nor U7703 (N_7703,N_7454,N_7284);
or U7704 (N_7704,N_7073,N_7375);
nor U7705 (N_7705,N_7085,N_7415);
or U7706 (N_7706,N_7300,N_7135);
nand U7707 (N_7707,N_6927,N_6929);
xnor U7708 (N_7708,N_7237,N_7129);
nor U7709 (N_7709,N_7155,N_7016);
and U7710 (N_7710,N_7233,N_7072);
xnor U7711 (N_7711,N_7367,N_7200);
or U7712 (N_7712,N_7380,N_7470);
nor U7713 (N_7713,N_7474,N_7296);
or U7714 (N_7714,N_7124,N_6894);
nand U7715 (N_7715,N_7183,N_6947);
nand U7716 (N_7716,N_7139,N_7424);
nor U7717 (N_7717,N_6902,N_7348);
or U7718 (N_7718,N_6913,N_7056);
and U7719 (N_7719,N_7304,N_7057);
nand U7720 (N_7720,N_7254,N_7285);
nor U7721 (N_7721,N_7291,N_7467);
and U7722 (N_7722,N_7443,N_7263);
nand U7723 (N_7723,N_7298,N_7490);
xor U7724 (N_7724,N_7130,N_6920);
xor U7725 (N_7725,N_7030,N_7219);
xnor U7726 (N_7726,N_7213,N_7410);
or U7727 (N_7727,N_7163,N_7377);
xor U7728 (N_7728,N_6884,N_7259);
nand U7729 (N_7729,N_6887,N_6896);
nand U7730 (N_7730,N_7330,N_7214);
xnor U7731 (N_7731,N_7429,N_7005);
or U7732 (N_7732,N_7397,N_7322);
xor U7733 (N_7733,N_7360,N_7106);
and U7734 (N_7734,N_7440,N_7428);
and U7735 (N_7735,N_7039,N_7010);
xnor U7736 (N_7736,N_7269,N_7283);
nand U7737 (N_7737,N_6926,N_7460);
and U7738 (N_7738,N_7409,N_7218);
and U7739 (N_7739,N_7211,N_7121);
nor U7740 (N_7740,N_7458,N_7225);
xor U7741 (N_7741,N_7393,N_7392);
nand U7742 (N_7742,N_6965,N_7419);
and U7743 (N_7743,N_7175,N_7230);
and U7744 (N_7744,N_6982,N_7362);
xnor U7745 (N_7745,N_7234,N_7325);
xnor U7746 (N_7746,N_7365,N_7185);
nand U7747 (N_7747,N_7281,N_7401);
and U7748 (N_7748,N_7119,N_6912);
nand U7749 (N_7749,N_7094,N_6994);
and U7750 (N_7750,N_6942,N_7264);
and U7751 (N_7751,N_6892,N_7093);
xor U7752 (N_7752,N_7208,N_7383);
nand U7753 (N_7753,N_7452,N_7159);
nand U7754 (N_7754,N_7468,N_7245);
nor U7755 (N_7755,N_7388,N_7268);
nand U7756 (N_7756,N_6881,N_7138);
nand U7757 (N_7757,N_7328,N_7023);
xnor U7758 (N_7758,N_7153,N_7323);
nor U7759 (N_7759,N_6977,N_7091);
nand U7760 (N_7760,N_7301,N_6899);
xor U7761 (N_7761,N_6924,N_6891);
nand U7762 (N_7762,N_7402,N_7146);
or U7763 (N_7763,N_7035,N_7192);
nor U7764 (N_7764,N_7471,N_7222);
xor U7765 (N_7765,N_7464,N_7140);
xnor U7766 (N_7766,N_6921,N_7453);
xnor U7767 (N_7767,N_7465,N_7253);
xnor U7768 (N_7768,N_6980,N_6889);
xor U7769 (N_7769,N_7199,N_7115);
and U7770 (N_7770,N_6885,N_7043);
or U7771 (N_7771,N_6997,N_6888);
nor U7772 (N_7772,N_7064,N_7069);
or U7773 (N_7773,N_7479,N_7477);
or U7774 (N_7774,N_7358,N_7040);
nor U7775 (N_7775,N_7334,N_6988);
and U7776 (N_7776,N_7486,N_6970);
nand U7777 (N_7777,N_7450,N_7127);
or U7778 (N_7778,N_7350,N_6969);
nor U7779 (N_7779,N_6890,N_7294);
xnor U7780 (N_7780,N_6992,N_7498);
nor U7781 (N_7781,N_7457,N_6906);
nor U7782 (N_7782,N_7110,N_7306);
nand U7783 (N_7783,N_7015,N_7186);
nand U7784 (N_7784,N_7421,N_7426);
and U7785 (N_7785,N_6953,N_7202);
nor U7786 (N_7786,N_7412,N_7327);
nor U7787 (N_7787,N_7246,N_6998);
or U7788 (N_7788,N_7188,N_7496);
xnor U7789 (N_7789,N_7391,N_7114);
nor U7790 (N_7790,N_7252,N_7111);
and U7791 (N_7791,N_6945,N_7066);
nor U7792 (N_7792,N_7174,N_7074);
and U7793 (N_7793,N_7166,N_7195);
or U7794 (N_7794,N_7287,N_6964);
nor U7795 (N_7795,N_6948,N_7145);
xnor U7796 (N_7796,N_7125,N_7050);
or U7797 (N_7797,N_7432,N_7282);
xnor U7798 (N_7798,N_7189,N_7369);
nor U7799 (N_7799,N_7201,N_7128);
or U7800 (N_7800,N_6971,N_7295);
xor U7801 (N_7801,N_7280,N_7310);
nand U7802 (N_7802,N_6878,N_6995);
nand U7803 (N_7803,N_7248,N_7494);
and U7804 (N_7804,N_7037,N_7251);
or U7805 (N_7805,N_7255,N_6987);
or U7806 (N_7806,N_7042,N_7198);
nor U7807 (N_7807,N_7359,N_7389);
or U7808 (N_7808,N_7368,N_7087);
xor U7809 (N_7809,N_7154,N_6951);
or U7810 (N_7810,N_7088,N_6875);
nor U7811 (N_7811,N_6895,N_7324);
nand U7812 (N_7812,N_7420,N_7362);
and U7813 (N_7813,N_7254,N_7347);
xor U7814 (N_7814,N_7228,N_7280);
and U7815 (N_7815,N_7379,N_6955);
or U7816 (N_7816,N_7198,N_7391);
and U7817 (N_7817,N_7192,N_6968);
nor U7818 (N_7818,N_7279,N_7066);
nor U7819 (N_7819,N_7270,N_7385);
or U7820 (N_7820,N_7395,N_6971);
xnor U7821 (N_7821,N_7342,N_7290);
nor U7822 (N_7822,N_7031,N_7150);
xor U7823 (N_7823,N_7461,N_6887);
or U7824 (N_7824,N_6966,N_7010);
or U7825 (N_7825,N_6942,N_7383);
or U7826 (N_7826,N_7237,N_7007);
xnor U7827 (N_7827,N_7094,N_6922);
and U7828 (N_7828,N_7021,N_7449);
xor U7829 (N_7829,N_7188,N_7443);
xor U7830 (N_7830,N_6981,N_7184);
xnor U7831 (N_7831,N_7010,N_6931);
nor U7832 (N_7832,N_7156,N_7415);
and U7833 (N_7833,N_6943,N_7209);
nand U7834 (N_7834,N_6945,N_7152);
or U7835 (N_7835,N_7394,N_7460);
nor U7836 (N_7836,N_7036,N_7364);
and U7837 (N_7837,N_7060,N_7266);
or U7838 (N_7838,N_7044,N_7375);
and U7839 (N_7839,N_6888,N_7242);
xor U7840 (N_7840,N_7071,N_7030);
nor U7841 (N_7841,N_7145,N_7030);
nor U7842 (N_7842,N_7239,N_6963);
and U7843 (N_7843,N_7417,N_7421);
and U7844 (N_7844,N_7478,N_7229);
nor U7845 (N_7845,N_7265,N_7099);
or U7846 (N_7846,N_7472,N_7009);
and U7847 (N_7847,N_7300,N_7067);
and U7848 (N_7848,N_7326,N_7398);
or U7849 (N_7849,N_7397,N_7369);
or U7850 (N_7850,N_7367,N_7231);
nand U7851 (N_7851,N_7247,N_6946);
or U7852 (N_7852,N_7053,N_7239);
nand U7853 (N_7853,N_7149,N_6941);
nor U7854 (N_7854,N_7185,N_7007);
nor U7855 (N_7855,N_7107,N_7493);
xnor U7856 (N_7856,N_7476,N_7368);
nor U7857 (N_7857,N_6918,N_6915);
xnor U7858 (N_7858,N_7238,N_7152);
nand U7859 (N_7859,N_7404,N_7062);
and U7860 (N_7860,N_7386,N_6892);
nor U7861 (N_7861,N_7162,N_7231);
nor U7862 (N_7862,N_7283,N_7142);
or U7863 (N_7863,N_7197,N_7460);
xor U7864 (N_7864,N_7156,N_7194);
xor U7865 (N_7865,N_6885,N_7064);
xor U7866 (N_7866,N_7315,N_7105);
nand U7867 (N_7867,N_7214,N_7144);
or U7868 (N_7868,N_7216,N_7369);
or U7869 (N_7869,N_7072,N_7168);
and U7870 (N_7870,N_7307,N_7167);
nor U7871 (N_7871,N_7260,N_6972);
nand U7872 (N_7872,N_7248,N_7138);
xnor U7873 (N_7873,N_7103,N_7423);
nor U7874 (N_7874,N_7341,N_7292);
nor U7875 (N_7875,N_6943,N_7468);
and U7876 (N_7876,N_6893,N_7361);
or U7877 (N_7877,N_6926,N_7238);
nor U7878 (N_7878,N_6886,N_7219);
and U7879 (N_7879,N_7491,N_7113);
nand U7880 (N_7880,N_7073,N_7422);
or U7881 (N_7881,N_6923,N_7320);
xnor U7882 (N_7882,N_7017,N_7021);
xor U7883 (N_7883,N_7430,N_6957);
nand U7884 (N_7884,N_7217,N_7240);
or U7885 (N_7885,N_7366,N_7183);
and U7886 (N_7886,N_7019,N_7053);
nor U7887 (N_7887,N_6877,N_6936);
or U7888 (N_7888,N_6960,N_7304);
nand U7889 (N_7889,N_7190,N_7282);
and U7890 (N_7890,N_7472,N_7125);
and U7891 (N_7891,N_7284,N_7380);
nand U7892 (N_7892,N_7188,N_7430);
and U7893 (N_7893,N_6971,N_6887);
nand U7894 (N_7894,N_7146,N_7128);
nand U7895 (N_7895,N_7343,N_7201);
or U7896 (N_7896,N_7229,N_7040);
and U7897 (N_7897,N_7176,N_7071);
nand U7898 (N_7898,N_6956,N_7083);
and U7899 (N_7899,N_7139,N_7171);
xor U7900 (N_7900,N_7314,N_7115);
and U7901 (N_7901,N_7256,N_7329);
and U7902 (N_7902,N_7121,N_6910);
xor U7903 (N_7903,N_7097,N_7103);
nand U7904 (N_7904,N_7440,N_6964);
and U7905 (N_7905,N_6947,N_7257);
or U7906 (N_7906,N_6956,N_7360);
and U7907 (N_7907,N_7270,N_7124);
or U7908 (N_7908,N_7382,N_7022);
nand U7909 (N_7909,N_6954,N_7088);
nand U7910 (N_7910,N_7242,N_7096);
and U7911 (N_7911,N_7478,N_7489);
nor U7912 (N_7912,N_7440,N_6882);
nand U7913 (N_7913,N_7061,N_6955);
nand U7914 (N_7914,N_7045,N_6896);
and U7915 (N_7915,N_6990,N_7438);
and U7916 (N_7916,N_7132,N_6938);
nand U7917 (N_7917,N_7394,N_7221);
or U7918 (N_7918,N_7113,N_6991);
xor U7919 (N_7919,N_6974,N_7377);
or U7920 (N_7920,N_7259,N_6987);
and U7921 (N_7921,N_6935,N_7251);
or U7922 (N_7922,N_7340,N_7177);
or U7923 (N_7923,N_7497,N_7428);
nor U7924 (N_7924,N_7097,N_7334);
nand U7925 (N_7925,N_7465,N_7221);
nor U7926 (N_7926,N_7244,N_7489);
and U7927 (N_7927,N_7363,N_6962);
and U7928 (N_7928,N_7260,N_6920);
and U7929 (N_7929,N_7134,N_7454);
or U7930 (N_7930,N_7036,N_6966);
and U7931 (N_7931,N_7347,N_7362);
or U7932 (N_7932,N_7409,N_7254);
or U7933 (N_7933,N_7332,N_7213);
and U7934 (N_7934,N_7210,N_7028);
nand U7935 (N_7935,N_7491,N_7259);
and U7936 (N_7936,N_6975,N_7022);
nand U7937 (N_7937,N_7156,N_7374);
nor U7938 (N_7938,N_7295,N_6993);
nand U7939 (N_7939,N_7006,N_6993);
nand U7940 (N_7940,N_7172,N_6925);
or U7941 (N_7941,N_7345,N_6934);
and U7942 (N_7942,N_7294,N_7193);
nand U7943 (N_7943,N_7428,N_7424);
nand U7944 (N_7944,N_7374,N_7010);
xnor U7945 (N_7945,N_7192,N_6985);
xor U7946 (N_7946,N_6978,N_7223);
xor U7947 (N_7947,N_7092,N_7030);
and U7948 (N_7948,N_7409,N_7217);
and U7949 (N_7949,N_7303,N_7445);
nor U7950 (N_7950,N_6952,N_7422);
xnor U7951 (N_7951,N_7088,N_7087);
or U7952 (N_7952,N_7053,N_7237);
nand U7953 (N_7953,N_7140,N_7484);
nor U7954 (N_7954,N_7435,N_6953);
or U7955 (N_7955,N_7170,N_7227);
or U7956 (N_7956,N_6917,N_6906);
and U7957 (N_7957,N_7208,N_7162);
nor U7958 (N_7958,N_7442,N_6983);
nand U7959 (N_7959,N_7174,N_6909);
nand U7960 (N_7960,N_7292,N_7251);
nand U7961 (N_7961,N_7400,N_7174);
nor U7962 (N_7962,N_7351,N_7380);
nor U7963 (N_7963,N_7123,N_7375);
nor U7964 (N_7964,N_7100,N_7417);
xnor U7965 (N_7965,N_6938,N_6900);
nor U7966 (N_7966,N_6946,N_7453);
xor U7967 (N_7967,N_6924,N_7462);
or U7968 (N_7968,N_7049,N_7005);
xnor U7969 (N_7969,N_6922,N_7101);
xor U7970 (N_7970,N_6901,N_7026);
xor U7971 (N_7971,N_7387,N_7142);
nand U7972 (N_7972,N_7116,N_7468);
nor U7973 (N_7973,N_7456,N_7284);
nand U7974 (N_7974,N_6945,N_7292);
nand U7975 (N_7975,N_6996,N_7453);
nand U7976 (N_7976,N_7375,N_7253);
or U7977 (N_7977,N_7266,N_7330);
nand U7978 (N_7978,N_7176,N_7432);
or U7979 (N_7979,N_7323,N_6878);
or U7980 (N_7980,N_7121,N_7188);
nor U7981 (N_7981,N_7187,N_7316);
or U7982 (N_7982,N_7078,N_7476);
nor U7983 (N_7983,N_7160,N_7495);
xnor U7984 (N_7984,N_7237,N_6937);
or U7985 (N_7985,N_7062,N_7387);
or U7986 (N_7986,N_6922,N_7250);
nor U7987 (N_7987,N_7264,N_7389);
nor U7988 (N_7988,N_7132,N_7237);
nand U7989 (N_7989,N_7307,N_7443);
nand U7990 (N_7990,N_7264,N_7372);
nor U7991 (N_7991,N_6938,N_7006);
nor U7992 (N_7992,N_7151,N_6915);
nand U7993 (N_7993,N_7146,N_6903);
nand U7994 (N_7994,N_6985,N_7188);
nor U7995 (N_7995,N_7364,N_7381);
or U7996 (N_7996,N_7035,N_7417);
xnor U7997 (N_7997,N_7395,N_7098);
or U7998 (N_7998,N_7429,N_7312);
or U7999 (N_7999,N_7076,N_7151);
or U8000 (N_8000,N_7258,N_7211);
and U8001 (N_8001,N_7094,N_7288);
nor U8002 (N_8002,N_7151,N_7343);
and U8003 (N_8003,N_7466,N_7297);
and U8004 (N_8004,N_7476,N_7426);
and U8005 (N_8005,N_7390,N_7477);
nor U8006 (N_8006,N_6911,N_7358);
or U8007 (N_8007,N_7467,N_7430);
or U8008 (N_8008,N_7118,N_7056);
or U8009 (N_8009,N_6965,N_7264);
xnor U8010 (N_8010,N_7384,N_7491);
nand U8011 (N_8011,N_7033,N_7077);
nand U8012 (N_8012,N_6965,N_6946);
xnor U8013 (N_8013,N_7033,N_7410);
nand U8014 (N_8014,N_6929,N_7185);
nor U8015 (N_8015,N_7256,N_7033);
and U8016 (N_8016,N_7002,N_7088);
nand U8017 (N_8017,N_7365,N_7204);
xnor U8018 (N_8018,N_7167,N_7151);
nor U8019 (N_8019,N_6996,N_7081);
nor U8020 (N_8020,N_6902,N_6907);
and U8021 (N_8021,N_7121,N_7106);
xor U8022 (N_8022,N_7343,N_7093);
xor U8023 (N_8023,N_6886,N_6922);
or U8024 (N_8024,N_7190,N_7441);
and U8025 (N_8025,N_7074,N_6945);
and U8026 (N_8026,N_7068,N_7173);
and U8027 (N_8027,N_6918,N_7403);
xnor U8028 (N_8028,N_6935,N_7266);
and U8029 (N_8029,N_7043,N_7448);
and U8030 (N_8030,N_6955,N_7186);
and U8031 (N_8031,N_7317,N_7154);
and U8032 (N_8032,N_7081,N_7271);
xnor U8033 (N_8033,N_7466,N_7034);
and U8034 (N_8034,N_7025,N_7438);
nand U8035 (N_8035,N_7050,N_7070);
xnor U8036 (N_8036,N_7113,N_6902);
and U8037 (N_8037,N_7471,N_6902);
nand U8038 (N_8038,N_7394,N_7087);
or U8039 (N_8039,N_7477,N_7392);
or U8040 (N_8040,N_7440,N_7199);
and U8041 (N_8041,N_7004,N_7054);
nor U8042 (N_8042,N_7378,N_7410);
nand U8043 (N_8043,N_7348,N_7237);
nand U8044 (N_8044,N_7187,N_7313);
nand U8045 (N_8045,N_7309,N_7440);
xor U8046 (N_8046,N_7398,N_7177);
xnor U8047 (N_8047,N_7049,N_7278);
nand U8048 (N_8048,N_7409,N_7450);
xnor U8049 (N_8049,N_7375,N_7216);
xnor U8050 (N_8050,N_7346,N_7275);
nor U8051 (N_8051,N_6908,N_7016);
nand U8052 (N_8052,N_7228,N_6963);
xnor U8053 (N_8053,N_7046,N_7335);
xnor U8054 (N_8054,N_7122,N_7139);
nor U8055 (N_8055,N_7271,N_7091);
nand U8056 (N_8056,N_7433,N_7393);
and U8057 (N_8057,N_7448,N_7166);
nand U8058 (N_8058,N_7286,N_7432);
nor U8059 (N_8059,N_6889,N_7214);
xor U8060 (N_8060,N_7137,N_7256);
or U8061 (N_8061,N_6898,N_7095);
and U8062 (N_8062,N_7048,N_7390);
xnor U8063 (N_8063,N_7314,N_7480);
and U8064 (N_8064,N_7457,N_7190);
and U8065 (N_8065,N_7067,N_7372);
nand U8066 (N_8066,N_6935,N_7056);
or U8067 (N_8067,N_7154,N_6914);
or U8068 (N_8068,N_7178,N_7353);
nand U8069 (N_8069,N_6971,N_7042);
nor U8070 (N_8070,N_7456,N_7059);
nor U8071 (N_8071,N_7280,N_7383);
and U8072 (N_8072,N_7113,N_7028);
and U8073 (N_8073,N_7458,N_7399);
nor U8074 (N_8074,N_7129,N_7071);
and U8075 (N_8075,N_7100,N_6982);
nor U8076 (N_8076,N_7105,N_7332);
and U8077 (N_8077,N_7391,N_7423);
nand U8078 (N_8078,N_7471,N_7156);
or U8079 (N_8079,N_7333,N_7413);
xnor U8080 (N_8080,N_7213,N_7170);
or U8081 (N_8081,N_7233,N_7410);
or U8082 (N_8082,N_7492,N_7308);
xnor U8083 (N_8083,N_6938,N_6888);
xnor U8084 (N_8084,N_7408,N_7198);
or U8085 (N_8085,N_7384,N_6959);
xor U8086 (N_8086,N_7324,N_7079);
and U8087 (N_8087,N_7285,N_6979);
nand U8088 (N_8088,N_6906,N_7019);
xor U8089 (N_8089,N_7398,N_7025);
nand U8090 (N_8090,N_6950,N_7016);
nand U8091 (N_8091,N_7282,N_7398);
or U8092 (N_8092,N_7291,N_7390);
nor U8093 (N_8093,N_7315,N_7132);
or U8094 (N_8094,N_7168,N_6923);
and U8095 (N_8095,N_7138,N_7140);
nand U8096 (N_8096,N_7491,N_6878);
nor U8097 (N_8097,N_6962,N_7316);
xor U8098 (N_8098,N_7183,N_6975);
and U8099 (N_8099,N_7178,N_6890);
nand U8100 (N_8100,N_7162,N_6979);
or U8101 (N_8101,N_7150,N_7350);
nor U8102 (N_8102,N_7365,N_7226);
nand U8103 (N_8103,N_7277,N_7241);
or U8104 (N_8104,N_6995,N_7387);
or U8105 (N_8105,N_6962,N_7110);
nor U8106 (N_8106,N_7363,N_7179);
or U8107 (N_8107,N_7236,N_7382);
nand U8108 (N_8108,N_7106,N_7051);
nand U8109 (N_8109,N_7420,N_7368);
or U8110 (N_8110,N_7470,N_7404);
nand U8111 (N_8111,N_7160,N_7020);
nor U8112 (N_8112,N_6889,N_6923);
xnor U8113 (N_8113,N_7410,N_6898);
nand U8114 (N_8114,N_6977,N_6971);
nand U8115 (N_8115,N_7282,N_7407);
nor U8116 (N_8116,N_6915,N_7336);
xnor U8117 (N_8117,N_6944,N_7255);
nor U8118 (N_8118,N_6890,N_7135);
and U8119 (N_8119,N_6984,N_7416);
or U8120 (N_8120,N_7135,N_7125);
nand U8121 (N_8121,N_6929,N_6931);
nor U8122 (N_8122,N_7303,N_6893);
or U8123 (N_8123,N_6909,N_7355);
nor U8124 (N_8124,N_6961,N_7310);
xnor U8125 (N_8125,N_7995,N_7690);
or U8126 (N_8126,N_8072,N_7919);
xnor U8127 (N_8127,N_7842,N_7816);
nand U8128 (N_8128,N_8109,N_7519);
nand U8129 (N_8129,N_7797,N_7939);
nor U8130 (N_8130,N_7825,N_8055);
and U8131 (N_8131,N_8098,N_7695);
or U8132 (N_8132,N_8089,N_7853);
xnor U8133 (N_8133,N_8012,N_7955);
and U8134 (N_8134,N_7879,N_7624);
nor U8135 (N_8135,N_8119,N_8000);
xor U8136 (N_8136,N_8014,N_8095);
and U8137 (N_8137,N_7608,N_7888);
or U8138 (N_8138,N_7947,N_7691);
xnor U8139 (N_8139,N_8084,N_8011);
nand U8140 (N_8140,N_7874,N_7904);
and U8141 (N_8141,N_7882,N_7654);
nand U8142 (N_8142,N_7872,N_7633);
nor U8143 (N_8143,N_8066,N_7595);
xnor U8144 (N_8144,N_8035,N_7546);
nor U8145 (N_8145,N_8013,N_7584);
xnor U8146 (N_8146,N_7764,N_7547);
xor U8147 (N_8147,N_7524,N_8123);
or U8148 (N_8148,N_7986,N_7731);
xnor U8149 (N_8149,N_7861,N_7589);
nor U8150 (N_8150,N_8042,N_7532);
xor U8151 (N_8151,N_7761,N_7693);
and U8152 (N_8152,N_7940,N_7614);
and U8153 (N_8153,N_7854,N_7709);
nand U8154 (N_8154,N_7970,N_8043);
and U8155 (N_8155,N_8063,N_7605);
nand U8156 (N_8156,N_7634,N_8031);
and U8157 (N_8157,N_7735,N_7609);
or U8158 (N_8158,N_7907,N_8053);
xnor U8159 (N_8159,N_7616,N_7680);
xor U8160 (N_8160,N_8106,N_7728);
xnor U8161 (N_8161,N_7617,N_7933);
xnor U8162 (N_8162,N_7581,N_7583);
nand U8163 (N_8163,N_7769,N_8114);
and U8164 (N_8164,N_7507,N_7977);
xor U8165 (N_8165,N_8080,N_7619);
or U8166 (N_8166,N_7674,N_8033);
or U8167 (N_8167,N_7618,N_8096);
nor U8168 (N_8168,N_7500,N_7530);
nor U8169 (N_8169,N_7664,N_7596);
nor U8170 (N_8170,N_7850,N_8024);
xor U8171 (N_8171,N_7648,N_7705);
xor U8172 (N_8172,N_8026,N_7629);
xor U8173 (N_8173,N_7949,N_7673);
nand U8174 (N_8174,N_7972,N_7672);
xnor U8175 (N_8175,N_7578,N_8107);
nand U8176 (N_8176,N_7716,N_8056);
nor U8177 (N_8177,N_7717,N_8082);
and U8178 (N_8178,N_7649,N_7537);
and U8179 (N_8179,N_7739,N_7545);
xnor U8180 (N_8180,N_7815,N_7784);
nand U8181 (N_8181,N_7892,N_7699);
or U8182 (N_8182,N_7833,N_7975);
xor U8183 (N_8183,N_7756,N_7909);
xor U8184 (N_8184,N_7794,N_7754);
xnor U8185 (N_8185,N_7561,N_7568);
xnor U8186 (N_8186,N_7708,N_7718);
or U8187 (N_8187,N_8087,N_7788);
and U8188 (N_8188,N_7598,N_7987);
and U8189 (N_8189,N_7566,N_7508);
and U8190 (N_8190,N_7540,N_8081);
nor U8191 (N_8191,N_7623,N_7526);
nor U8192 (N_8192,N_7963,N_7979);
and U8193 (N_8193,N_8067,N_7518);
or U8194 (N_8194,N_8021,N_7948);
xor U8195 (N_8195,N_8105,N_7553);
xnor U8196 (N_8196,N_7538,N_7936);
xnor U8197 (N_8197,N_8102,N_7625);
nand U8198 (N_8198,N_7604,N_7533);
nand U8199 (N_8199,N_7509,N_8112);
nand U8200 (N_8200,N_8009,N_7849);
or U8201 (N_8201,N_7851,N_7787);
nand U8202 (N_8202,N_7505,N_7594);
nor U8203 (N_8203,N_7704,N_7783);
or U8204 (N_8204,N_7801,N_7841);
nand U8205 (N_8205,N_7657,N_7750);
nand U8206 (N_8206,N_8097,N_7539);
and U8207 (N_8207,N_8025,N_8037);
nor U8208 (N_8208,N_7820,N_7791);
and U8209 (N_8209,N_7582,N_7786);
nand U8210 (N_8210,N_7865,N_7744);
nor U8211 (N_8211,N_7817,N_7610);
nor U8212 (N_8212,N_7682,N_7562);
nand U8213 (N_8213,N_7757,N_7698);
nand U8214 (N_8214,N_8069,N_7550);
xor U8215 (N_8215,N_7800,N_7721);
nor U8216 (N_8216,N_7703,N_7994);
and U8217 (N_8217,N_8070,N_7593);
xnor U8218 (N_8218,N_8005,N_7501);
and U8219 (N_8219,N_7517,N_7910);
or U8220 (N_8220,N_7762,N_7962);
nor U8221 (N_8221,N_7809,N_7782);
or U8222 (N_8222,N_8007,N_7966);
or U8223 (N_8223,N_7871,N_7636);
and U8224 (N_8224,N_7603,N_7645);
nor U8225 (N_8225,N_7938,N_7821);
nor U8226 (N_8226,N_7920,N_7732);
and U8227 (N_8227,N_7643,N_8077);
nand U8228 (N_8228,N_7612,N_7544);
nand U8229 (N_8229,N_7510,N_7707);
xor U8230 (N_8230,N_8004,N_7844);
or U8231 (N_8231,N_7881,N_7776);
xor U8232 (N_8232,N_7671,N_8113);
xor U8233 (N_8233,N_7552,N_7777);
xnor U8234 (N_8234,N_7795,N_8027);
nor U8235 (N_8235,N_7734,N_7831);
nand U8236 (N_8236,N_7845,N_7869);
or U8237 (N_8237,N_7893,N_7846);
nand U8238 (N_8238,N_7516,N_7745);
nor U8239 (N_8239,N_7567,N_7676);
and U8240 (N_8240,N_7529,N_7912);
and U8241 (N_8241,N_8029,N_7923);
or U8242 (N_8242,N_7549,N_7944);
or U8243 (N_8243,N_8022,N_7958);
nor U8244 (N_8244,N_7890,N_7760);
or U8245 (N_8245,N_7806,N_8120);
nor U8246 (N_8246,N_8046,N_7733);
and U8247 (N_8247,N_7860,N_7915);
and U8248 (N_8248,N_7719,N_7635);
nor U8249 (N_8249,N_7896,N_7875);
or U8250 (N_8250,N_7902,N_7922);
or U8251 (N_8251,N_7889,N_7985);
xor U8252 (N_8252,N_7993,N_8051);
and U8253 (N_8253,N_7931,N_8038);
or U8254 (N_8254,N_8085,N_7877);
nand U8255 (N_8255,N_7813,N_7651);
nor U8256 (N_8256,N_7864,N_8121);
and U8257 (N_8257,N_7688,N_7961);
and U8258 (N_8258,N_7627,N_8094);
and U8259 (N_8259,N_8086,N_7670);
nor U8260 (N_8260,N_7686,N_7639);
and U8261 (N_8261,N_7789,N_7836);
and U8262 (N_8262,N_7863,N_8091);
nor U8263 (N_8263,N_7675,N_7577);
or U8264 (N_8264,N_7973,N_8036);
xnor U8265 (N_8265,N_7918,N_7590);
and U8266 (N_8266,N_8048,N_7752);
xor U8267 (N_8267,N_7997,N_7711);
and U8268 (N_8268,N_7662,N_7576);
or U8269 (N_8269,N_7701,N_8061);
xnor U8270 (N_8270,N_7870,N_7681);
nand U8271 (N_8271,N_7978,N_8079);
or U8272 (N_8272,N_7823,N_7942);
or U8273 (N_8273,N_8003,N_7878);
nor U8274 (N_8274,N_7677,N_7747);
xnor U8275 (N_8275,N_7883,N_7937);
and U8276 (N_8276,N_7905,N_8078);
and U8277 (N_8277,N_7725,N_8088);
nand U8278 (N_8278,N_7655,N_8068);
xor U8279 (N_8279,N_7683,N_7876);
or U8280 (N_8280,N_7988,N_7900);
nand U8281 (N_8281,N_7687,N_7780);
nand U8282 (N_8282,N_7571,N_7775);
nand U8283 (N_8283,N_7724,N_7886);
xor U8284 (N_8284,N_7898,N_8058);
xnor U8285 (N_8285,N_7897,N_7781);
nor U8286 (N_8286,N_7990,N_7976);
xnor U8287 (N_8287,N_7785,N_8059);
and U8288 (N_8288,N_7950,N_7765);
xor U8289 (N_8289,N_7513,N_8032);
nand U8290 (N_8290,N_7965,N_7759);
or U8291 (N_8291,N_7723,N_7790);
xnor U8292 (N_8292,N_7726,N_8075);
and U8293 (N_8293,N_7826,N_7514);
xnor U8294 (N_8294,N_7715,N_7894);
nor U8295 (N_8295,N_7586,N_8001);
xor U8296 (N_8296,N_7588,N_7722);
xnor U8297 (N_8297,N_8040,N_7521);
and U8298 (N_8298,N_8062,N_7697);
and U8299 (N_8299,N_7702,N_7758);
nand U8300 (N_8300,N_7984,N_7660);
or U8301 (N_8301,N_7793,N_7502);
xnor U8302 (N_8302,N_7968,N_7742);
and U8303 (N_8303,N_7525,N_7749);
or U8304 (N_8304,N_8010,N_8045);
xnor U8305 (N_8305,N_7601,N_7555);
and U8306 (N_8306,N_7741,N_7773);
or U8307 (N_8307,N_7903,N_7527);
xnor U8308 (N_8308,N_7585,N_7934);
or U8309 (N_8309,N_7796,N_7641);
nand U8310 (N_8310,N_7906,N_8101);
xor U8311 (N_8311,N_8060,N_7637);
or U8312 (N_8312,N_7969,N_7504);
nor U8313 (N_8313,N_8049,N_7859);
or U8314 (N_8314,N_7650,N_7798);
xor U8315 (N_8315,N_7692,N_7587);
nand U8316 (N_8316,N_8071,N_7925);
xnor U8317 (N_8317,N_7679,N_7974);
and U8318 (N_8318,N_7843,N_8116);
xnor U8319 (N_8319,N_7822,N_7522);
nor U8320 (N_8320,N_7819,N_7803);
xor U8321 (N_8321,N_7964,N_7929);
and U8322 (N_8322,N_7631,N_7827);
or U8323 (N_8323,N_7712,N_7740);
nor U8324 (N_8324,N_7930,N_7792);
nand U8325 (N_8325,N_7511,N_7512);
nand U8326 (N_8326,N_7710,N_7808);
or U8327 (N_8327,N_7943,N_7957);
nand U8328 (N_8328,N_7835,N_7613);
xor U8329 (N_8329,N_8050,N_7572);
xnor U8330 (N_8330,N_7506,N_8076);
nor U8331 (N_8331,N_7981,N_7829);
or U8332 (N_8332,N_8044,N_7980);
or U8333 (N_8333,N_8028,N_7768);
or U8334 (N_8334,N_7996,N_7927);
or U8335 (N_8335,N_8052,N_8111);
and U8336 (N_8336,N_7563,N_7665);
or U8337 (N_8337,N_7659,N_7812);
and U8338 (N_8338,N_8090,N_7954);
xnor U8339 (N_8339,N_7736,N_7873);
or U8340 (N_8340,N_7630,N_8118);
or U8341 (N_8341,N_7998,N_7989);
nor U8342 (N_8342,N_7602,N_8015);
or U8343 (N_8343,N_7621,N_7622);
nand U8344 (N_8344,N_7620,N_7811);
xor U8345 (N_8345,N_7945,N_7983);
nand U8346 (N_8346,N_7535,N_8117);
and U8347 (N_8347,N_7579,N_7556);
xor U8348 (N_8348,N_8100,N_7606);
or U8349 (N_8349,N_7548,N_7678);
or U8350 (N_8350,N_7884,N_7696);
or U8351 (N_8351,N_7600,N_7607);
nand U8352 (N_8352,N_7971,N_7916);
or U8353 (N_8353,N_8034,N_7531);
or U8354 (N_8354,N_7838,N_8016);
nor U8355 (N_8355,N_7810,N_7684);
nand U8356 (N_8356,N_7862,N_7661);
xor U8357 (N_8357,N_7644,N_7828);
nor U8358 (N_8358,N_7951,N_7564);
or U8359 (N_8359,N_7685,N_7592);
nor U8360 (N_8360,N_7834,N_7580);
nor U8361 (N_8361,N_7774,N_7557);
and U8362 (N_8362,N_7528,N_7541);
nand U8363 (N_8363,N_7959,N_7523);
nor U8364 (N_8364,N_7652,N_7559);
xnor U8365 (N_8365,N_8093,N_7867);
xor U8366 (N_8366,N_7840,N_7642);
xor U8367 (N_8367,N_8073,N_7799);
or U8368 (N_8368,N_7667,N_8064);
nor U8369 (N_8369,N_8115,N_7766);
nand U8370 (N_8370,N_7727,N_7771);
nand U8371 (N_8371,N_7668,N_7669);
or U8372 (N_8372,N_7899,N_7772);
or U8373 (N_8373,N_8002,N_7573);
nor U8374 (N_8374,N_7536,N_7615);
xor U8375 (N_8375,N_7730,N_8065);
or U8376 (N_8376,N_7830,N_7991);
xor U8377 (N_8377,N_7720,N_7554);
xor U8378 (N_8378,N_7926,N_7856);
nand U8379 (N_8379,N_7713,N_7611);
nor U8380 (N_8380,N_8054,N_7914);
and U8381 (N_8381,N_8017,N_8083);
and U8382 (N_8382,N_8041,N_7880);
xnor U8383 (N_8383,N_7852,N_7542);
nand U8384 (N_8384,N_7558,N_7839);
or U8385 (N_8385,N_7628,N_7767);
nand U8386 (N_8386,N_8110,N_7913);
nand U8387 (N_8387,N_7700,N_7520);
xor U8388 (N_8388,N_7814,N_7551);
nor U8389 (N_8389,N_7515,N_8103);
and U8390 (N_8390,N_7917,N_8039);
nand U8391 (N_8391,N_7921,N_7737);
xor U8392 (N_8392,N_7807,N_8057);
or U8393 (N_8393,N_8108,N_7967);
nor U8394 (N_8394,N_7658,N_7887);
nand U8395 (N_8395,N_7847,N_7848);
xnor U8396 (N_8396,N_7908,N_7818);
nor U8397 (N_8397,N_8019,N_7560);
nor U8398 (N_8398,N_8023,N_7569);
nor U8399 (N_8399,N_7743,N_7632);
and U8400 (N_8400,N_7802,N_7666);
nor U8401 (N_8401,N_7953,N_7729);
nand U8402 (N_8402,N_7770,N_7960);
and U8403 (N_8403,N_7924,N_7946);
nor U8404 (N_8404,N_7982,N_7779);
or U8405 (N_8405,N_7857,N_7575);
or U8406 (N_8406,N_7778,N_7868);
and U8407 (N_8407,N_7640,N_7748);
or U8408 (N_8408,N_7753,N_8006);
nor U8409 (N_8409,N_8008,N_7565);
or U8410 (N_8410,N_8124,N_7574);
nand U8411 (N_8411,N_7503,N_7999);
nand U8412 (N_8412,N_7738,N_7932);
and U8413 (N_8413,N_8020,N_7638);
xnor U8414 (N_8414,N_8122,N_7824);
nor U8415 (N_8415,N_7689,N_8104);
xnor U8416 (N_8416,N_7706,N_7837);
xor U8417 (N_8417,N_7885,N_8092);
and U8418 (N_8418,N_7694,N_7992);
nor U8419 (N_8419,N_7866,N_7891);
and U8420 (N_8420,N_7597,N_7832);
or U8421 (N_8421,N_7763,N_7928);
or U8422 (N_8422,N_7591,N_7911);
nand U8423 (N_8423,N_8047,N_7855);
nor U8424 (N_8424,N_8018,N_7646);
or U8425 (N_8425,N_8099,N_7626);
or U8426 (N_8426,N_8030,N_7956);
xor U8427 (N_8427,N_7746,N_7653);
nor U8428 (N_8428,N_7543,N_7570);
and U8429 (N_8429,N_7804,N_7941);
nand U8430 (N_8430,N_7895,N_7858);
and U8431 (N_8431,N_7751,N_7952);
nor U8432 (N_8432,N_7935,N_7714);
nand U8433 (N_8433,N_7755,N_8074);
xor U8434 (N_8434,N_7663,N_7534);
and U8435 (N_8435,N_7901,N_7647);
and U8436 (N_8436,N_7656,N_7599);
nand U8437 (N_8437,N_7805,N_8110);
and U8438 (N_8438,N_7947,N_7833);
or U8439 (N_8439,N_8112,N_7817);
or U8440 (N_8440,N_8010,N_7956);
nor U8441 (N_8441,N_7619,N_7796);
xnor U8442 (N_8442,N_7825,N_7547);
xor U8443 (N_8443,N_7672,N_7966);
or U8444 (N_8444,N_7770,N_7705);
nand U8445 (N_8445,N_8106,N_7547);
and U8446 (N_8446,N_7760,N_7814);
xor U8447 (N_8447,N_7895,N_7683);
and U8448 (N_8448,N_7927,N_7748);
nor U8449 (N_8449,N_7524,N_7710);
and U8450 (N_8450,N_7778,N_7553);
or U8451 (N_8451,N_8105,N_7837);
or U8452 (N_8452,N_7709,N_7827);
nor U8453 (N_8453,N_7994,N_7996);
and U8454 (N_8454,N_7867,N_7709);
and U8455 (N_8455,N_7569,N_7656);
and U8456 (N_8456,N_8025,N_8101);
xor U8457 (N_8457,N_7559,N_7644);
xor U8458 (N_8458,N_7753,N_7650);
xor U8459 (N_8459,N_7938,N_7597);
xor U8460 (N_8460,N_8027,N_7564);
nand U8461 (N_8461,N_7923,N_8054);
or U8462 (N_8462,N_8032,N_7890);
xnor U8463 (N_8463,N_7655,N_8088);
and U8464 (N_8464,N_7762,N_7628);
nand U8465 (N_8465,N_7633,N_7986);
nand U8466 (N_8466,N_7578,N_7612);
or U8467 (N_8467,N_7972,N_7891);
nand U8468 (N_8468,N_7934,N_7885);
and U8469 (N_8469,N_8075,N_7514);
xnor U8470 (N_8470,N_8014,N_7801);
or U8471 (N_8471,N_7557,N_7773);
nor U8472 (N_8472,N_7566,N_7711);
nor U8473 (N_8473,N_7658,N_7763);
xnor U8474 (N_8474,N_7742,N_7589);
nand U8475 (N_8475,N_7834,N_7941);
nor U8476 (N_8476,N_7692,N_7854);
xnor U8477 (N_8477,N_7741,N_7552);
or U8478 (N_8478,N_7731,N_7613);
or U8479 (N_8479,N_7718,N_7763);
or U8480 (N_8480,N_7737,N_7520);
and U8481 (N_8481,N_7756,N_7920);
nor U8482 (N_8482,N_7591,N_7717);
nand U8483 (N_8483,N_8023,N_7915);
nor U8484 (N_8484,N_7957,N_7887);
nand U8485 (N_8485,N_7676,N_7969);
xnor U8486 (N_8486,N_8089,N_8043);
nand U8487 (N_8487,N_7629,N_8008);
xor U8488 (N_8488,N_8115,N_8063);
nand U8489 (N_8489,N_8008,N_8122);
or U8490 (N_8490,N_7853,N_8083);
and U8491 (N_8491,N_7510,N_7978);
and U8492 (N_8492,N_7684,N_7873);
xnor U8493 (N_8493,N_7520,N_8053);
xnor U8494 (N_8494,N_8090,N_7553);
and U8495 (N_8495,N_8119,N_7908);
nand U8496 (N_8496,N_8032,N_7844);
nor U8497 (N_8497,N_7911,N_7843);
or U8498 (N_8498,N_7515,N_8102);
xor U8499 (N_8499,N_7566,N_8092);
xor U8500 (N_8500,N_7602,N_7801);
and U8501 (N_8501,N_8059,N_7503);
xnor U8502 (N_8502,N_7954,N_8081);
nand U8503 (N_8503,N_7941,N_7895);
or U8504 (N_8504,N_7644,N_7941);
or U8505 (N_8505,N_7869,N_7666);
nor U8506 (N_8506,N_8012,N_8020);
nand U8507 (N_8507,N_7774,N_7758);
and U8508 (N_8508,N_7588,N_8029);
xnor U8509 (N_8509,N_7912,N_7558);
nand U8510 (N_8510,N_7943,N_7597);
or U8511 (N_8511,N_7895,N_7954);
and U8512 (N_8512,N_7891,N_7722);
and U8513 (N_8513,N_7954,N_7969);
or U8514 (N_8514,N_7925,N_7783);
nand U8515 (N_8515,N_8067,N_7522);
xor U8516 (N_8516,N_8099,N_7589);
nor U8517 (N_8517,N_7729,N_7956);
nor U8518 (N_8518,N_7749,N_8054);
xor U8519 (N_8519,N_7887,N_7541);
nor U8520 (N_8520,N_7749,N_8041);
or U8521 (N_8521,N_7964,N_7799);
xor U8522 (N_8522,N_7667,N_8082);
or U8523 (N_8523,N_8025,N_7613);
nor U8524 (N_8524,N_7913,N_7936);
xnor U8525 (N_8525,N_7765,N_8050);
nand U8526 (N_8526,N_7619,N_8117);
and U8527 (N_8527,N_7718,N_8097);
nor U8528 (N_8528,N_7777,N_8095);
nand U8529 (N_8529,N_7701,N_7545);
and U8530 (N_8530,N_7604,N_7843);
xnor U8531 (N_8531,N_7516,N_7703);
nor U8532 (N_8532,N_8037,N_7982);
nand U8533 (N_8533,N_7590,N_7683);
xnor U8534 (N_8534,N_7991,N_7790);
or U8535 (N_8535,N_7764,N_7849);
xor U8536 (N_8536,N_7852,N_7732);
and U8537 (N_8537,N_8021,N_7533);
and U8538 (N_8538,N_7820,N_8081);
nor U8539 (N_8539,N_7938,N_8102);
nor U8540 (N_8540,N_8039,N_8003);
or U8541 (N_8541,N_8000,N_7531);
or U8542 (N_8542,N_7946,N_7560);
nand U8543 (N_8543,N_8074,N_7632);
or U8544 (N_8544,N_8001,N_7607);
nand U8545 (N_8545,N_7653,N_7683);
nand U8546 (N_8546,N_7514,N_7692);
xnor U8547 (N_8547,N_7731,N_7957);
nor U8548 (N_8548,N_7688,N_7573);
or U8549 (N_8549,N_8000,N_7912);
or U8550 (N_8550,N_7991,N_7587);
nor U8551 (N_8551,N_7956,N_8112);
nor U8552 (N_8552,N_7538,N_7921);
xor U8553 (N_8553,N_7511,N_7861);
or U8554 (N_8554,N_7898,N_7864);
nand U8555 (N_8555,N_7955,N_8065);
or U8556 (N_8556,N_8050,N_7734);
and U8557 (N_8557,N_7625,N_7584);
nand U8558 (N_8558,N_7936,N_7753);
and U8559 (N_8559,N_7709,N_7965);
nor U8560 (N_8560,N_7616,N_7777);
or U8561 (N_8561,N_8009,N_7733);
nand U8562 (N_8562,N_8003,N_7635);
nor U8563 (N_8563,N_7841,N_7614);
xor U8564 (N_8564,N_7614,N_7933);
nor U8565 (N_8565,N_8069,N_7600);
or U8566 (N_8566,N_7743,N_7951);
and U8567 (N_8567,N_7712,N_7663);
and U8568 (N_8568,N_7730,N_8119);
nor U8569 (N_8569,N_7914,N_7981);
or U8570 (N_8570,N_8087,N_7953);
or U8571 (N_8571,N_7503,N_8115);
nand U8572 (N_8572,N_7960,N_7837);
nand U8573 (N_8573,N_7993,N_7949);
and U8574 (N_8574,N_7817,N_7679);
nand U8575 (N_8575,N_7590,N_7796);
or U8576 (N_8576,N_7698,N_7862);
and U8577 (N_8577,N_8017,N_7926);
and U8578 (N_8578,N_8040,N_7671);
or U8579 (N_8579,N_8052,N_7516);
xnor U8580 (N_8580,N_7978,N_7718);
xor U8581 (N_8581,N_8060,N_7567);
and U8582 (N_8582,N_7620,N_7831);
or U8583 (N_8583,N_7795,N_8098);
nand U8584 (N_8584,N_7964,N_7717);
and U8585 (N_8585,N_8000,N_8097);
or U8586 (N_8586,N_7642,N_7908);
nor U8587 (N_8587,N_7540,N_7522);
or U8588 (N_8588,N_8019,N_7563);
nand U8589 (N_8589,N_7907,N_7936);
xor U8590 (N_8590,N_7930,N_7655);
and U8591 (N_8591,N_8024,N_7683);
or U8592 (N_8592,N_7801,N_7607);
nor U8593 (N_8593,N_7694,N_7940);
nand U8594 (N_8594,N_7988,N_7879);
nor U8595 (N_8595,N_7512,N_7877);
or U8596 (N_8596,N_8099,N_7871);
and U8597 (N_8597,N_8097,N_7746);
xnor U8598 (N_8598,N_7515,N_7711);
or U8599 (N_8599,N_8035,N_7689);
nand U8600 (N_8600,N_7624,N_7930);
nand U8601 (N_8601,N_7706,N_8001);
xnor U8602 (N_8602,N_7519,N_7618);
xnor U8603 (N_8603,N_8071,N_7661);
nand U8604 (N_8604,N_7855,N_7929);
xor U8605 (N_8605,N_7579,N_7535);
nor U8606 (N_8606,N_8123,N_7733);
nand U8607 (N_8607,N_7593,N_7703);
xor U8608 (N_8608,N_7795,N_7819);
or U8609 (N_8609,N_7972,N_7645);
nor U8610 (N_8610,N_7518,N_7914);
xor U8611 (N_8611,N_7825,N_7530);
and U8612 (N_8612,N_8011,N_7711);
nor U8613 (N_8613,N_8123,N_7665);
or U8614 (N_8614,N_7852,N_7668);
nand U8615 (N_8615,N_7648,N_7843);
xor U8616 (N_8616,N_7777,N_7702);
and U8617 (N_8617,N_7847,N_8118);
and U8618 (N_8618,N_7618,N_7872);
xnor U8619 (N_8619,N_7935,N_8031);
and U8620 (N_8620,N_8102,N_7760);
xnor U8621 (N_8621,N_7553,N_7502);
and U8622 (N_8622,N_7976,N_7928);
nor U8623 (N_8623,N_8045,N_7947);
or U8624 (N_8624,N_7507,N_7707);
nand U8625 (N_8625,N_8085,N_7686);
nand U8626 (N_8626,N_7748,N_7827);
xor U8627 (N_8627,N_7731,N_7745);
nor U8628 (N_8628,N_8032,N_7833);
and U8629 (N_8629,N_7667,N_7581);
or U8630 (N_8630,N_7887,N_7539);
nor U8631 (N_8631,N_7903,N_7696);
xor U8632 (N_8632,N_7852,N_7610);
nand U8633 (N_8633,N_7539,N_8063);
nor U8634 (N_8634,N_7759,N_7812);
xnor U8635 (N_8635,N_7973,N_7934);
nand U8636 (N_8636,N_7799,N_7666);
nand U8637 (N_8637,N_7711,N_7612);
and U8638 (N_8638,N_7756,N_7609);
nor U8639 (N_8639,N_7598,N_7922);
nand U8640 (N_8640,N_7624,N_8017);
nor U8641 (N_8641,N_7533,N_7858);
xnor U8642 (N_8642,N_7872,N_7512);
or U8643 (N_8643,N_7892,N_7805);
or U8644 (N_8644,N_7535,N_8044);
or U8645 (N_8645,N_7782,N_7912);
or U8646 (N_8646,N_7803,N_7962);
nor U8647 (N_8647,N_7839,N_7967);
or U8648 (N_8648,N_7784,N_7611);
nor U8649 (N_8649,N_7565,N_7523);
xor U8650 (N_8650,N_7591,N_7539);
nand U8651 (N_8651,N_7783,N_8095);
nand U8652 (N_8652,N_7976,N_7912);
or U8653 (N_8653,N_8074,N_7945);
nand U8654 (N_8654,N_7803,N_7850);
xor U8655 (N_8655,N_7557,N_7602);
xor U8656 (N_8656,N_8107,N_7810);
nor U8657 (N_8657,N_7798,N_7575);
nor U8658 (N_8658,N_7557,N_7668);
or U8659 (N_8659,N_7663,N_7605);
nor U8660 (N_8660,N_7581,N_7968);
and U8661 (N_8661,N_7610,N_7972);
xnor U8662 (N_8662,N_7881,N_7962);
or U8663 (N_8663,N_8022,N_7923);
nand U8664 (N_8664,N_7866,N_7733);
xnor U8665 (N_8665,N_7759,N_8119);
nor U8666 (N_8666,N_7666,N_7572);
or U8667 (N_8667,N_7887,N_7515);
or U8668 (N_8668,N_7790,N_7797);
nand U8669 (N_8669,N_7857,N_7961);
and U8670 (N_8670,N_7514,N_7747);
nand U8671 (N_8671,N_7827,N_7938);
and U8672 (N_8672,N_8084,N_8007);
nand U8673 (N_8673,N_8011,N_7586);
xnor U8674 (N_8674,N_7842,N_7811);
nor U8675 (N_8675,N_7902,N_8116);
xor U8676 (N_8676,N_8114,N_8124);
nor U8677 (N_8677,N_7961,N_7683);
xnor U8678 (N_8678,N_7573,N_7831);
nor U8679 (N_8679,N_7720,N_7865);
and U8680 (N_8680,N_7949,N_8038);
xnor U8681 (N_8681,N_8081,N_7799);
or U8682 (N_8682,N_7529,N_7968);
nor U8683 (N_8683,N_7773,N_7837);
or U8684 (N_8684,N_7832,N_7825);
or U8685 (N_8685,N_7845,N_7799);
nand U8686 (N_8686,N_7573,N_8070);
nor U8687 (N_8687,N_7734,N_7965);
or U8688 (N_8688,N_7635,N_7528);
nand U8689 (N_8689,N_8065,N_7883);
nand U8690 (N_8690,N_7732,N_7558);
nand U8691 (N_8691,N_7556,N_7797);
nor U8692 (N_8692,N_8049,N_7685);
nand U8693 (N_8693,N_7971,N_7893);
and U8694 (N_8694,N_7966,N_7833);
nor U8695 (N_8695,N_7521,N_8074);
and U8696 (N_8696,N_8121,N_7886);
or U8697 (N_8697,N_7863,N_7795);
or U8698 (N_8698,N_7841,N_7548);
nand U8699 (N_8699,N_7597,N_7853);
nand U8700 (N_8700,N_7532,N_7624);
or U8701 (N_8701,N_7706,N_7627);
nand U8702 (N_8702,N_7689,N_7846);
or U8703 (N_8703,N_7503,N_8027);
or U8704 (N_8704,N_7656,N_7826);
or U8705 (N_8705,N_7642,N_8061);
nand U8706 (N_8706,N_7743,N_8048);
and U8707 (N_8707,N_7720,N_8081);
nor U8708 (N_8708,N_7887,N_7741);
nor U8709 (N_8709,N_7661,N_8079);
nand U8710 (N_8710,N_7692,N_7825);
or U8711 (N_8711,N_7796,N_7668);
and U8712 (N_8712,N_7929,N_7885);
xnor U8713 (N_8713,N_7585,N_7973);
xnor U8714 (N_8714,N_8010,N_7976);
or U8715 (N_8715,N_7594,N_7616);
nand U8716 (N_8716,N_7735,N_8079);
and U8717 (N_8717,N_8026,N_7534);
and U8718 (N_8718,N_7686,N_7812);
xor U8719 (N_8719,N_7889,N_8011);
xor U8720 (N_8720,N_7878,N_7789);
nor U8721 (N_8721,N_8106,N_7730);
nand U8722 (N_8722,N_7575,N_8056);
and U8723 (N_8723,N_7932,N_7662);
or U8724 (N_8724,N_8094,N_8052);
and U8725 (N_8725,N_7665,N_7896);
and U8726 (N_8726,N_7864,N_7508);
nand U8727 (N_8727,N_7511,N_7883);
and U8728 (N_8728,N_7770,N_7804);
nor U8729 (N_8729,N_7586,N_7972);
xor U8730 (N_8730,N_7625,N_7867);
xor U8731 (N_8731,N_7598,N_7730);
or U8732 (N_8732,N_8026,N_7529);
xnor U8733 (N_8733,N_7598,N_7812);
nor U8734 (N_8734,N_7690,N_7565);
or U8735 (N_8735,N_8090,N_8117);
nor U8736 (N_8736,N_7677,N_7606);
and U8737 (N_8737,N_7618,N_7513);
nor U8738 (N_8738,N_7862,N_7642);
xor U8739 (N_8739,N_7601,N_7678);
or U8740 (N_8740,N_7945,N_7542);
xnor U8741 (N_8741,N_7742,N_8078);
and U8742 (N_8742,N_7982,N_7605);
nor U8743 (N_8743,N_8020,N_7940);
and U8744 (N_8744,N_7953,N_7697);
or U8745 (N_8745,N_7900,N_7688);
xor U8746 (N_8746,N_7570,N_7746);
and U8747 (N_8747,N_7880,N_7971);
xor U8748 (N_8748,N_7625,N_7838);
xnor U8749 (N_8749,N_7623,N_8124);
or U8750 (N_8750,N_8638,N_8640);
nor U8751 (N_8751,N_8460,N_8248);
nand U8752 (N_8752,N_8571,N_8481);
xnor U8753 (N_8753,N_8564,N_8729);
or U8754 (N_8754,N_8332,N_8441);
nand U8755 (N_8755,N_8280,N_8498);
and U8756 (N_8756,N_8695,N_8524);
or U8757 (N_8757,N_8644,N_8488);
nor U8758 (N_8758,N_8643,N_8664);
nor U8759 (N_8759,N_8514,N_8509);
xnor U8760 (N_8760,N_8297,N_8518);
xnor U8761 (N_8761,N_8631,N_8499);
and U8762 (N_8762,N_8741,N_8195);
or U8763 (N_8763,N_8550,N_8412);
nand U8764 (N_8764,N_8503,N_8272);
and U8765 (N_8765,N_8600,N_8344);
xnor U8766 (N_8766,N_8579,N_8671);
xor U8767 (N_8767,N_8372,N_8164);
nor U8768 (N_8768,N_8743,N_8725);
and U8769 (N_8769,N_8511,N_8526);
nor U8770 (N_8770,N_8167,N_8217);
or U8771 (N_8771,N_8396,N_8668);
nand U8772 (N_8772,N_8383,N_8458);
xnor U8773 (N_8773,N_8491,N_8284);
nor U8774 (N_8774,N_8206,N_8733);
nor U8775 (N_8775,N_8457,N_8483);
xor U8776 (N_8776,N_8288,N_8180);
or U8777 (N_8777,N_8392,N_8692);
and U8778 (N_8778,N_8727,N_8429);
or U8779 (N_8779,N_8447,N_8724);
and U8780 (N_8780,N_8565,N_8740);
or U8781 (N_8781,N_8494,N_8232);
nand U8782 (N_8782,N_8475,N_8282);
and U8783 (N_8783,N_8278,N_8188);
nor U8784 (N_8784,N_8165,N_8463);
nand U8785 (N_8785,N_8318,N_8127);
nor U8786 (N_8786,N_8723,N_8647);
nor U8787 (N_8787,N_8251,N_8194);
and U8788 (N_8788,N_8615,N_8354);
xnor U8789 (N_8789,N_8225,N_8694);
xor U8790 (N_8790,N_8701,N_8140);
or U8791 (N_8791,N_8350,N_8489);
nor U8792 (N_8792,N_8566,N_8128);
nand U8793 (N_8793,N_8618,N_8697);
or U8794 (N_8794,N_8577,N_8541);
and U8795 (N_8795,N_8530,N_8185);
nor U8796 (N_8796,N_8472,N_8339);
nor U8797 (N_8797,N_8490,N_8135);
or U8798 (N_8798,N_8540,N_8146);
and U8799 (N_8799,N_8721,N_8163);
nor U8800 (N_8800,N_8734,N_8404);
and U8801 (N_8801,N_8269,N_8560);
and U8802 (N_8802,N_8663,N_8744);
nand U8803 (N_8803,N_8656,N_8190);
nor U8804 (N_8804,N_8289,N_8270);
nand U8805 (N_8805,N_8608,N_8374);
nand U8806 (N_8806,N_8448,N_8262);
xnor U8807 (N_8807,N_8479,N_8314);
nor U8808 (N_8808,N_8258,N_8287);
xor U8809 (N_8809,N_8731,N_8405);
or U8810 (N_8810,N_8214,N_8415);
or U8811 (N_8811,N_8634,N_8425);
or U8812 (N_8812,N_8604,N_8516);
and U8813 (N_8813,N_8547,N_8500);
nor U8814 (N_8814,N_8179,N_8141);
xnor U8815 (N_8815,N_8279,N_8598);
and U8816 (N_8816,N_8584,N_8655);
nand U8817 (N_8817,N_8613,N_8702);
and U8818 (N_8818,N_8726,N_8574);
nand U8819 (N_8819,N_8482,N_8402);
nand U8820 (N_8820,N_8535,N_8310);
nand U8821 (N_8821,N_8485,N_8267);
nor U8822 (N_8822,N_8271,N_8421);
nand U8823 (N_8823,N_8543,N_8477);
nand U8824 (N_8824,N_8224,N_8522);
nand U8825 (N_8825,N_8196,N_8384);
or U8826 (N_8826,N_8456,N_8276);
xnor U8827 (N_8827,N_8192,N_8698);
nor U8828 (N_8828,N_8567,N_8432);
nor U8829 (N_8829,N_8238,N_8520);
or U8830 (N_8830,N_8747,N_8667);
or U8831 (N_8831,N_8294,N_8342);
nand U8832 (N_8832,N_8242,N_8126);
or U8833 (N_8833,N_8394,N_8635);
nor U8834 (N_8834,N_8557,N_8470);
nor U8835 (N_8835,N_8673,N_8260);
nand U8836 (N_8836,N_8245,N_8411);
and U8837 (N_8837,N_8437,N_8320);
xnor U8838 (N_8838,N_8606,N_8221);
nand U8839 (N_8839,N_8544,N_8610);
or U8840 (N_8840,N_8220,N_8501);
or U8841 (N_8841,N_8469,N_8597);
nor U8842 (N_8842,N_8665,N_8235);
and U8843 (N_8843,N_8476,N_8704);
nand U8844 (N_8844,N_8317,N_8409);
nand U8845 (N_8845,N_8125,N_8473);
or U8846 (N_8846,N_8393,N_8707);
or U8847 (N_8847,N_8202,N_8308);
nand U8848 (N_8848,N_8453,N_8601);
nand U8849 (N_8849,N_8418,N_8433);
nor U8850 (N_8850,N_8528,N_8609);
or U8851 (N_8851,N_8705,N_8537);
and U8852 (N_8852,N_8681,N_8546);
nor U8853 (N_8853,N_8373,N_8395);
nor U8854 (N_8854,N_8134,N_8171);
xor U8855 (N_8855,N_8335,N_8653);
nand U8856 (N_8856,N_8486,N_8385);
nand U8857 (N_8857,N_8145,N_8716);
xor U8858 (N_8858,N_8328,N_8617);
or U8859 (N_8859,N_8382,N_8711);
or U8860 (N_8860,N_8302,N_8348);
nand U8861 (N_8861,N_8728,N_8438);
xnor U8862 (N_8862,N_8474,N_8714);
or U8863 (N_8863,N_8508,N_8155);
nor U8864 (N_8864,N_8417,N_8230);
nand U8865 (N_8865,N_8419,N_8131);
or U8866 (N_8866,N_8675,N_8264);
nor U8867 (N_8867,N_8151,N_8642);
or U8868 (N_8868,N_8246,N_8403);
or U8869 (N_8869,N_8170,N_8215);
nand U8870 (N_8870,N_8158,N_8523);
or U8871 (N_8871,N_8575,N_8172);
xnor U8872 (N_8872,N_8515,N_8189);
nor U8873 (N_8873,N_8391,N_8661);
nor U8874 (N_8874,N_8678,N_8381);
xor U8875 (N_8875,N_8371,N_8588);
nand U8876 (N_8876,N_8710,N_8651);
or U8877 (N_8877,N_8130,N_8532);
nor U8878 (N_8878,N_8378,N_8748);
and U8879 (N_8879,N_8362,N_8298);
or U8880 (N_8880,N_8676,N_8311);
xor U8881 (N_8881,N_8177,N_8495);
nand U8882 (N_8882,N_8589,N_8338);
nand U8883 (N_8883,N_8507,N_8413);
nor U8884 (N_8884,N_8454,N_8693);
and U8885 (N_8885,N_8504,N_8237);
or U8886 (N_8886,N_8244,N_8273);
and U8887 (N_8887,N_8205,N_8330);
xor U8888 (N_8888,N_8129,N_8305);
xnor U8889 (N_8889,N_8347,N_8444);
nand U8890 (N_8890,N_8443,N_8626);
xor U8891 (N_8891,N_8706,N_8623);
and U8892 (N_8892,N_8569,N_8228);
nand U8893 (N_8893,N_8505,N_8236);
nand U8894 (N_8894,N_8720,N_8239);
xor U8895 (N_8895,N_8277,N_8183);
and U8896 (N_8896,N_8401,N_8343);
nor U8897 (N_8897,N_8534,N_8380);
xor U8898 (N_8898,N_8138,N_8416);
nand U8899 (N_8899,N_8556,N_8240);
and U8900 (N_8900,N_8687,N_8708);
xor U8901 (N_8901,N_8684,N_8349);
or U8902 (N_8902,N_8386,N_8573);
xor U8903 (N_8903,N_8191,N_8536);
nand U8904 (N_8904,N_8266,N_8558);
and U8905 (N_8905,N_8683,N_8434);
or U8906 (N_8906,N_8545,N_8559);
and U8907 (N_8907,N_8178,N_8680);
nor U8908 (N_8908,N_8468,N_8324);
and U8909 (N_8909,N_8529,N_8493);
or U8910 (N_8910,N_8148,N_8738);
nor U8911 (N_8911,N_8492,N_8149);
or U8912 (N_8912,N_8351,N_8739);
nand U8913 (N_8913,N_8737,N_8531);
and U8914 (N_8914,N_8690,N_8363);
nor U8915 (N_8915,N_8719,N_8285);
or U8916 (N_8916,N_8592,N_8465);
nand U8917 (N_8917,N_8227,N_8368);
or U8918 (N_8918,N_8315,N_8630);
or U8919 (N_8919,N_8322,N_8143);
nand U8920 (N_8920,N_8358,N_8268);
nor U8921 (N_8921,N_8625,N_8576);
xor U8922 (N_8922,N_8677,N_8387);
and U8923 (N_8923,N_8436,N_8639);
nand U8924 (N_8924,N_8636,N_8650);
and U8925 (N_8925,N_8612,N_8410);
and U8926 (N_8926,N_8223,N_8641);
xor U8927 (N_8927,N_8341,N_8517);
nand U8928 (N_8928,N_8337,N_8548);
xor U8929 (N_8929,N_8309,N_8319);
and U8930 (N_8930,N_8388,N_8554);
nor U8931 (N_8931,N_8658,N_8250);
nor U8932 (N_8932,N_8602,N_8208);
or U8933 (N_8933,N_8255,N_8611);
or U8934 (N_8934,N_8484,N_8355);
xnor U8935 (N_8935,N_8399,N_8583);
nor U8936 (N_8936,N_8231,N_8136);
nand U8937 (N_8937,N_8539,N_8274);
nand U8938 (N_8938,N_8718,N_8291);
or U8939 (N_8939,N_8137,N_8591);
or U8940 (N_8940,N_8201,N_8464);
or U8941 (N_8941,N_8323,N_8506);
nor U8942 (N_8942,N_8519,N_8749);
and U8943 (N_8943,N_8281,N_8229);
or U8944 (N_8944,N_8379,N_8159);
or U8945 (N_8945,N_8203,N_8513);
and U8946 (N_8946,N_8166,N_8459);
and U8947 (N_8947,N_8478,N_8397);
and U8948 (N_8948,N_8450,N_8357);
or U8949 (N_8949,N_8301,N_8629);
nand U8950 (N_8950,N_8367,N_8426);
nand U8951 (N_8951,N_8722,N_8686);
xnor U8952 (N_8952,N_8712,N_8161);
and U8953 (N_8953,N_8263,N_8376);
xor U8954 (N_8954,N_8660,N_8637);
and U8955 (N_8955,N_8209,N_8585);
nor U8956 (N_8956,N_8624,N_8699);
or U8957 (N_8957,N_8168,N_8745);
nor U8958 (N_8958,N_8197,N_8207);
nand U8959 (N_8959,N_8688,N_8746);
xnor U8960 (N_8960,N_8552,N_8295);
nor U8961 (N_8961,N_8709,N_8646);
or U8962 (N_8962,N_8497,N_8461);
or U8963 (N_8963,N_8480,N_8157);
or U8964 (N_8964,N_8654,N_8241);
xor U8965 (N_8965,N_8369,N_8353);
or U8966 (N_8966,N_8657,N_8153);
nand U8967 (N_8967,N_8445,N_8252);
nand U8968 (N_8968,N_8213,N_8533);
nand U8969 (N_8969,N_8304,N_8147);
nor U8970 (N_8970,N_8312,N_8572);
or U8971 (N_8971,N_8621,N_8423);
nand U8972 (N_8972,N_8696,N_8570);
and U8973 (N_8973,N_8561,N_8555);
or U8974 (N_8974,N_8682,N_8595);
and U8975 (N_8975,N_8648,N_8669);
and U8976 (N_8976,N_8184,N_8150);
or U8977 (N_8977,N_8259,N_8133);
nor U8978 (N_8978,N_8303,N_8605);
nand U8979 (N_8979,N_8587,N_8487);
nand U8980 (N_8980,N_8175,N_8300);
nand U8981 (N_8981,N_8512,N_8193);
xor U8982 (N_8982,N_8685,N_8689);
nand U8983 (N_8983,N_8226,N_8527);
or U8984 (N_8984,N_8132,N_8510);
xor U8985 (N_8985,N_8521,N_8538);
nand U8986 (N_8986,N_8292,N_8365);
nor U8987 (N_8987,N_8306,N_8551);
and U8988 (N_8988,N_8139,N_8359);
xor U8989 (N_8989,N_8286,N_8340);
xor U8990 (N_8990,N_8216,N_8662);
nor U8991 (N_8991,N_8649,N_8496);
nor U8992 (N_8992,N_8700,N_8222);
nand U8993 (N_8993,N_8607,N_8442);
xnor U8994 (N_8994,N_8451,N_8666);
and U8995 (N_8995,N_8582,N_8406);
nor U8996 (N_8996,N_8389,N_8691);
and U8997 (N_8997,N_8254,N_8326);
xnor U8998 (N_8998,N_8243,N_8400);
and U8999 (N_8999,N_8174,N_8449);
nor U9000 (N_9000,N_8169,N_8659);
xor U9001 (N_9001,N_8614,N_8603);
and U9002 (N_9002,N_8346,N_8742);
nor U9003 (N_9003,N_8253,N_8173);
nor U9004 (N_9004,N_8211,N_8703);
xor U9005 (N_9005,N_8334,N_8176);
and U9006 (N_9006,N_8435,N_8290);
nand U9007 (N_9007,N_8452,N_8462);
nand U9008 (N_9008,N_8265,N_8553);
xnor U9009 (N_9009,N_8333,N_8313);
or U9010 (N_9010,N_8502,N_8307);
nand U9011 (N_9011,N_8275,N_8200);
nand U9012 (N_9012,N_8212,N_8420);
or U9013 (N_9013,N_8210,N_8632);
nor U9014 (N_9014,N_8622,N_8366);
and U9015 (N_9015,N_8455,N_8471);
nor U9016 (N_9016,N_8336,N_8542);
nor U9017 (N_9017,N_8467,N_8331);
nand U9018 (N_9018,N_8233,N_8428);
or U9019 (N_9019,N_8590,N_8652);
nor U9020 (N_9020,N_8620,N_8407);
nand U9021 (N_9021,N_8616,N_8356);
nor U9022 (N_9022,N_8594,N_8431);
or U9023 (N_9023,N_8439,N_8321);
xnor U9024 (N_9024,N_8142,N_8736);
nand U9025 (N_9025,N_8525,N_8144);
or U9026 (N_9026,N_8593,N_8364);
nor U9027 (N_9027,N_8581,N_8586);
xor U9028 (N_9028,N_8627,N_8345);
xnor U9029 (N_9029,N_8293,N_8257);
nor U9030 (N_9030,N_8735,N_8563);
or U9031 (N_9031,N_8329,N_8633);
nor U9032 (N_9032,N_8199,N_8218);
or U9033 (N_9033,N_8361,N_8562);
nand U9034 (N_9034,N_8296,N_8152);
xor U9035 (N_9035,N_8619,N_8549);
nor U9036 (N_9036,N_8580,N_8568);
nand U9037 (N_9037,N_8717,N_8670);
xor U9038 (N_9038,N_8408,N_8249);
nand U9039 (N_9039,N_8261,N_8596);
nor U9040 (N_9040,N_8219,N_8360);
and U9041 (N_9041,N_8299,N_8713);
or U9042 (N_9042,N_8352,N_8446);
xor U9043 (N_9043,N_8377,N_8679);
nor U9044 (N_9044,N_8427,N_8645);
xor U9045 (N_9045,N_8316,N_8283);
xor U9046 (N_9046,N_8370,N_8187);
xor U9047 (N_9047,N_8162,N_8398);
xnor U9048 (N_9048,N_8422,N_8715);
nand U9049 (N_9049,N_8414,N_8674);
or U9050 (N_9050,N_8154,N_8256);
nor U9051 (N_9051,N_8181,N_8204);
and U9052 (N_9052,N_8198,N_8730);
nand U9053 (N_9053,N_8160,N_8390);
xor U9054 (N_9054,N_8234,N_8186);
and U9055 (N_9055,N_8578,N_8325);
nand U9056 (N_9056,N_8430,N_8628);
xnor U9057 (N_9057,N_8247,N_8424);
nor U9058 (N_9058,N_8375,N_8599);
nand U9059 (N_9059,N_8672,N_8182);
or U9060 (N_9060,N_8732,N_8327);
or U9061 (N_9061,N_8156,N_8440);
or U9062 (N_9062,N_8466,N_8702);
xnor U9063 (N_9063,N_8695,N_8339);
xor U9064 (N_9064,N_8695,N_8320);
nand U9065 (N_9065,N_8302,N_8749);
and U9066 (N_9066,N_8580,N_8493);
nand U9067 (N_9067,N_8334,N_8342);
or U9068 (N_9068,N_8512,N_8131);
nand U9069 (N_9069,N_8525,N_8705);
nand U9070 (N_9070,N_8187,N_8476);
and U9071 (N_9071,N_8277,N_8528);
xnor U9072 (N_9072,N_8445,N_8261);
or U9073 (N_9073,N_8557,N_8646);
nor U9074 (N_9074,N_8317,N_8455);
nand U9075 (N_9075,N_8327,N_8383);
xor U9076 (N_9076,N_8401,N_8544);
nor U9077 (N_9077,N_8725,N_8616);
or U9078 (N_9078,N_8510,N_8306);
and U9079 (N_9079,N_8315,N_8150);
nor U9080 (N_9080,N_8215,N_8725);
and U9081 (N_9081,N_8230,N_8160);
xor U9082 (N_9082,N_8435,N_8324);
nand U9083 (N_9083,N_8633,N_8342);
nor U9084 (N_9084,N_8547,N_8415);
or U9085 (N_9085,N_8427,N_8349);
or U9086 (N_9086,N_8131,N_8466);
nand U9087 (N_9087,N_8146,N_8660);
xor U9088 (N_9088,N_8309,N_8462);
or U9089 (N_9089,N_8237,N_8266);
and U9090 (N_9090,N_8566,N_8383);
nand U9091 (N_9091,N_8390,N_8182);
or U9092 (N_9092,N_8689,N_8691);
and U9093 (N_9093,N_8718,N_8359);
or U9094 (N_9094,N_8646,N_8213);
and U9095 (N_9095,N_8317,N_8454);
and U9096 (N_9096,N_8615,N_8282);
nor U9097 (N_9097,N_8212,N_8342);
xor U9098 (N_9098,N_8657,N_8442);
xor U9099 (N_9099,N_8340,N_8349);
and U9100 (N_9100,N_8368,N_8471);
nor U9101 (N_9101,N_8738,N_8624);
or U9102 (N_9102,N_8575,N_8175);
nand U9103 (N_9103,N_8665,N_8731);
xor U9104 (N_9104,N_8612,N_8260);
xnor U9105 (N_9105,N_8126,N_8226);
nor U9106 (N_9106,N_8724,N_8548);
or U9107 (N_9107,N_8648,N_8473);
xnor U9108 (N_9108,N_8126,N_8170);
and U9109 (N_9109,N_8175,N_8387);
xnor U9110 (N_9110,N_8472,N_8740);
nor U9111 (N_9111,N_8141,N_8486);
xor U9112 (N_9112,N_8621,N_8545);
or U9113 (N_9113,N_8331,N_8303);
nand U9114 (N_9114,N_8707,N_8195);
or U9115 (N_9115,N_8671,N_8503);
or U9116 (N_9116,N_8268,N_8183);
or U9117 (N_9117,N_8191,N_8145);
nor U9118 (N_9118,N_8666,N_8689);
nand U9119 (N_9119,N_8401,N_8499);
xnor U9120 (N_9120,N_8422,N_8449);
nor U9121 (N_9121,N_8615,N_8335);
xnor U9122 (N_9122,N_8222,N_8497);
or U9123 (N_9123,N_8374,N_8520);
or U9124 (N_9124,N_8494,N_8527);
xnor U9125 (N_9125,N_8238,N_8190);
nor U9126 (N_9126,N_8352,N_8170);
nand U9127 (N_9127,N_8528,N_8536);
or U9128 (N_9128,N_8280,N_8196);
and U9129 (N_9129,N_8294,N_8488);
xnor U9130 (N_9130,N_8435,N_8478);
or U9131 (N_9131,N_8229,N_8608);
nor U9132 (N_9132,N_8277,N_8469);
nor U9133 (N_9133,N_8625,N_8275);
and U9134 (N_9134,N_8699,N_8414);
or U9135 (N_9135,N_8325,N_8449);
nand U9136 (N_9136,N_8650,N_8490);
nand U9137 (N_9137,N_8331,N_8573);
and U9138 (N_9138,N_8522,N_8242);
and U9139 (N_9139,N_8255,N_8389);
xor U9140 (N_9140,N_8157,N_8216);
or U9141 (N_9141,N_8450,N_8326);
or U9142 (N_9142,N_8686,N_8325);
nand U9143 (N_9143,N_8650,N_8711);
xor U9144 (N_9144,N_8664,N_8131);
nor U9145 (N_9145,N_8497,N_8500);
and U9146 (N_9146,N_8718,N_8217);
nor U9147 (N_9147,N_8328,N_8431);
and U9148 (N_9148,N_8680,N_8186);
nor U9149 (N_9149,N_8423,N_8163);
or U9150 (N_9150,N_8224,N_8145);
nor U9151 (N_9151,N_8175,N_8345);
xnor U9152 (N_9152,N_8721,N_8459);
or U9153 (N_9153,N_8354,N_8427);
or U9154 (N_9154,N_8528,N_8342);
or U9155 (N_9155,N_8388,N_8745);
or U9156 (N_9156,N_8272,N_8184);
and U9157 (N_9157,N_8175,N_8343);
nand U9158 (N_9158,N_8629,N_8532);
and U9159 (N_9159,N_8546,N_8247);
or U9160 (N_9160,N_8344,N_8650);
nor U9161 (N_9161,N_8494,N_8368);
xor U9162 (N_9162,N_8306,N_8303);
and U9163 (N_9163,N_8382,N_8743);
xnor U9164 (N_9164,N_8516,N_8433);
and U9165 (N_9165,N_8396,N_8469);
xnor U9166 (N_9166,N_8398,N_8247);
or U9167 (N_9167,N_8346,N_8183);
xor U9168 (N_9168,N_8608,N_8289);
nand U9169 (N_9169,N_8739,N_8591);
nand U9170 (N_9170,N_8201,N_8150);
nand U9171 (N_9171,N_8588,N_8725);
nor U9172 (N_9172,N_8235,N_8213);
or U9173 (N_9173,N_8471,N_8321);
nor U9174 (N_9174,N_8726,N_8546);
nor U9175 (N_9175,N_8126,N_8379);
and U9176 (N_9176,N_8607,N_8419);
xor U9177 (N_9177,N_8272,N_8425);
xnor U9178 (N_9178,N_8428,N_8389);
or U9179 (N_9179,N_8178,N_8467);
nor U9180 (N_9180,N_8713,N_8168);
nor U9181 (N_9181,N_8605,N_8744);
xnor U9182 (N_9182,N_8716,N_8628);
or U9183 (N_9183,N_8158,N_8482);
and U9184 (N_9184,N_8747,N_8566);
nor U9185 (N_9185,N_8295,N_8598);
and U9186 (N_9186,N_8206,N_8745);
nor U9187 (N_9187,N_8554,N_8164);
or U9188 (N_9188,N_8649,N_8192);
nor U9189 (N_9189,N_8633,N_8627);
and U9190 (N_9190,N_8550,N_8658);
or U9191 (N_9191,N_8379,N_8275);
or U9192 (N_9192,N_8321,N_8552);
xor U9193 (N_9193,N_8490,N_8347);
nor U9194 (N_9194,N_8747,N_8520);
nand U9195 (N_9195,N_8182,N_8632);
nor U9196 (N_9196,N_8256,N_8183);
or U9197 (N_9197,N_8498,N_8622);
nor U9198 (N_9198,N_8316,N_8415);
or U9199 (N_9199,N_8627,N_8311);
nand U9200 (N_9200,N_8644,N_8410);
and U9201 (N_9201,N_8410,N_8664);
nor U9202 (N_9202,N_8172,N_8290);
xnor U9203 (N_9203,N_8486,N_8455);
xor U9204 (N_9204,N_8158,N_8716);
xnor U9205 (N_9205,N_8210,N_8478);
nand U9206 (N_9206,N_8666,N_8329);
xnor U9207 (N_9207,N_8662,N_8233);
and U9208 (N_9208,N_8466,N_8399);
xor U9209 (N_9209,N_8706,N_8410);
and U9210 (N_9210,N_8303,N_8364);
nor U9211 (N_9211,N_8624,N_8742);
and U9212 (N_9212,N_8423,N_8591);
and U9213 (N_9213,N_8125,N_8573);
and U9214 (N_9214,N_8166,N_8521);
or U9215 (N_9215,N_8331,N_8516);
and U9216 (N_9216,N_8130,N_8174);
xnor U9217 (N_9217,N_8165,N_8136);
or U9218 (N_9218,N_8638,N_8565);
xor U9219 (N_9219,N_8659,N_8232);
and U9220 (N_9220,N_8342,N_8496);
nor U9221 (N_9221,N_8580,N_8273);
nand U9222 (N_9222,N_8278,N_8393);
or U9223 (N_9223,N_8650,N_8683);
xnor U9224 (N_9224,N_8735,N_8686);
nor U9225 (N_9225,N_8145,N_8333);
and U9226 (N_9226,N_8467,N_8358);
nand U9227 (N_9227,N_8382,N_8343);
nand U9228 (N_9228,N_8440,N_8554);
nand U9229 (N_9229,N_8672,N_8273);
and U9230 (N_9230,N_8126,N_8141);
nor U9231 (N_9231,N_8418,N_8226);
and U9232 (N_9232,N_8680,N_8375);
nor U9233 (N_9233,N_8462,N_8329);
nand U9234 (N_9234,N_8584,N_8606);
nor U9235 (N_9235,N_8319,N_8688);
nor U9236 (N_9236,N_8676,N_8378);
nand U9237 (N_9237,N_8564,N_8230);
nand U9238 (N_9238,N_8524,N_8446);
and U9239 (N_9239,N_8162,N_8522);
xor U9240 (N_9240,N_8256,N_8363);
nor U9241 (N_9241,N_8278,N_8681);
xor U9242 (N_9242,N_8339,N_8406);
or U9243 (N_9243,N_8129,N_8374);
or U9244 (N_9244,N_8198,N_8391);
nand U9245 (N_9245,N_8196,N_8535);
or U9246 (N_9246,N_8191,N_8589);
nand U9247 (N_9247,N_8540,N_8597);
and U9248 (N_9248,N_8193,N_8603);
or U9249 (N_9249,N_8602,N_8262);
or U9250 (N_9250,N_8139,N_8660);
nand U9251 (N_9251,N_8177,N_8367);
nand U9252 (N_9252,N_8379,N_8361);
or U9253 (N_9253,N_8545,N_8486);
and U9254 (N_9254,N_8513,N_8439);
nor U9255 (N_9255,N_8152,N_8714);
and U9256 (N_9256,N_8385,N_8358);
xor U9257 (N_9257,N_8605,N_8264);
and U9258 (N_9258,N_8495,N_8683);
nor U9259 (N_9259,N_8743,N_8152);
xor U9260 (N_9260,N_8588,N_8420);
and U9261 (N_9261,N_8579,N_8736);
xor U9262 (N_9262,N_8492,N_8724);
nor U9263 (N_9263,N_8493,N_8415);
xnor U9264 (N_9264,N_8587,N_8638);
nand U9265 (N_9265,N_8347,N_8473);
xor U9266 (N_9266,N_8150,N_8464);
and U9267 (N_9267,N_8582,N_8623);
nor U9268 (N_9268,N_8261,N_8302);
and U9269 (N_9269,N_8571,N_8680);
nand U9270 (N_9270,N_8670,N_8315);
nor U9271 (N_9271,N_8183,N_8514);
or U9272 (N_9272,N_8229,N_8474);
nand U9273 (N_9273,N_8134,N_8624);
nand U9274 (N_9274,N_8177,N_8414);
nand U9275 (N_9275,N_8360,N_8131);
xor U9276 (N_9276,N_8448,N_8449);
nor U9277 (N_9277,N_8155,N_8355);
nor U9278 (N_9278,N_8302,N_8412);
nor U9279 (N_9279,N_8149,N_8388);
or U9280 (N_9280,N_8307,N_8567);
or U9281 (N_9281,N_8194,N_8655);
and U9282 (N_9282,N_8271,N_8568);
nand U9283 (N_9283,N_8490,N_8396);
or U9284 (N_9284,N_8211,N_8335);
nand U9285 (N_9285,N_8236,N_8511);
and U9286 (N_9286,N_8489,N_8214);
and U9287 (N_9287,N_8309,N_8745);
nor U9288 (N_9288,N_8350,N_8695);
or U9289 (N_9289,N_8186,N_8275);
and U9290 (N_9290,N_8364,N_8143);
nand U9291 (N_9291,N_8595,N_8148);
xor U9292 (N_9292,N_8341,N_8307);
xor U9293 (N_9293,N_8210,N_8670);
nor U9294 (N_9294,N_8288,N_8690);
xnor U9295 (N_9295,N_8287,N_8474);
and U9296 (N_9296,N_8728,N_8213);
or U9297 (N_9297,N_8250,N_8286);
nor U9298 (N_9298,N_8727,N_8558);
and U9299 (N_9299,N_8508,N_8647);
and U9300 (N_9300,N_8263,N_8352);
nor U9301 (N_9301,N_8694,N_8555);
nor U9302 (N_9302,N_8686,N_8201);
nor U9303 (N_9303,N_8685,N_8472);
xnor U9304 (N_9304,N_8488,N_8742);
xor U9305 (N_9305,N_8282,N_8416);
nand U9306 (N_9306,N_8749,N_8552);
nor U9307 (N_9307,N_8709,N_8483);
nor U9308 (N_9308,N_8333,N_8365);
nand U9309 (N_9309,N_8289,N_8162);
and U9310 (N_9310,N_8639,N_8127);
or U9311 (N_9311,N_8310,N_8400);
nand U9312 (N_9312,N_8481,N_8518);
nor U9313 (N_9313,N_8133,N_8733);
and U9314 (N_9314,N_8563,N_8293);
and U9315 (N_9315,N_8281,N_8214);
and U9316 (N_9316,N_8298,N_8567);
nand U9317 (N_9317,N_8367,N_8640);
nand U9318 (N_9318,N_8155,N_8247);
nand U9319 (N_9319,N_8553,N_8368);
nor U9320 (N_9320,N_8355,N_8247);
xnor U9321 (N_9321,N_8406,N_8639);
and U9322 (N_9322,N_8329,N_8727);
or U9323 (N_9323,N_8348,N_8670);
xnor U9324 (N_9324,N_8248,N_8737);
xnor U9325 (N_9325,N_8273,N_8518);
nor U9326 (N_9326,N_8262,N_8520);
or U9327 (N_9327,N_8131,N_8297);
and U9328 (N_9328,N_8492,N_8467);
or U9329 (N_9329,N_8279,N_8344);
xnor U9330 (N_9330,N_8421,N_8347);
nand U9331 (N_9331,N_8463,N_8627);
nor U9332 (N_9332,N_8149,N_8736);
or U9333 (N_9333,N_8677,N_8193);
nand U9334 (N_9334,N_8706,N_8604);
or U9335 (N_9335,N_8247,N_8544);
nor U9336 (N_9336,N_8669,N_8171);
xnor U9337 (N_9337,N_8580,N_8514);
or U9338 (N_9338,N_8423,N_8729);
xor U9339 (N_9339,N_8268,N_8675);
or U9340 (N_9340,N_8354,N_8696);
nor U9341 (N_9341,N_8264,N_8428);
or U9342 (N_9342,N_8711,N_8376);
nor U9343 (N_9343,N_8402,N_8347);
or U9344 (N_9344,N_8554,N_8193);
or U9345 (N_9345,N_8642,N_8227);
nor U9346 (N_9346,N_8434,N_8581);
and U9347 (N_9347,N_8490,N_8264);
nand U9348 (N_9348,N_8584,N_8439);
or U9349 (N_9349,N_8380,N_8659);
nor U9350 (N_9350,N_8200,N_8660);
nand U9351 (N_9351,N_8257,N_8215);
and U9352 (N_9352,N_8705,N_8483);
xnor U9353 (N_9353,N_8677,N_8513);
nor U9354 (N_9354,N_8565,N_8129);
nor U9355 (N_9355,N_8427,N_8614);
nor U9356 (N_9356,N_8327,N_8687);
or U9357 (N_9357,N_8433,N_8484);
xnor U9358 (N_9358,N_8638,N_8644);
or U9359 (N_9359,N_8286,N_8246);
and U9360 (N_9360,N_8704,N_8508);
xor U9361 (N_9361,N_8422,N_8200);
nor U9362 (N_9362,N_8173,N_8275);
xor U9363 (N_9363,N_8356,N_8145);
or U9364 (N_9364,N_8216,N_8171);
or U9365 (N_9365,N_8740,N_8362);
nand U9366 (N_9366,N_8466,N_8667);
nor U9367 (N_9367,N_8274,N_8191);
and U9368 (N_9368,N_8173,N_8661);
nor U9369 (N_9369,N_8348,N_8154);
or U9370 (N_9370,N_8312,N_8316);
nand U9371 (N_9371,N_8211,N_8492);
xor U9372 (N_9372,N_8435,N_8660);
and U9373 (N_9373,N_8502,N_8146);
and U9374 (N_9374,N_8193,N_8370);
or U9375 (N_9375,N_8973,N_9190);
or U9376 (N_9376,N_8787,N_9252);
nand U9377 (N_9377,N_9038,N_9076);
nand U9378 (N_9378,N_9058,N_9176);
or U9379 (N_9379,N_8944,N_9001);
or U9380 (N_9380,N_8956,N_8836);
nand U9381 (N_9381,N_9238,N_9141);
and U9382 (N_9382,N_8792,N_9102);
and U9383 (N_9383,N_9042,N_9000);
xnor U9384 (N_9384,N_9148,N_9059);
or U9385 (N_9385,N_9025,N_8757);
xor U9386 (N_9386,N_9245,N_8919);
nand U9387 (N_9387,N_9033,N_8863);
and U9388 (N_9388,N_9039,N_9302);
nand U9389 (N_9389,N_9047,N_9103);
nor U9390 (N_9390,N_9088,N_9065);
and U9391 (N_9391,N_9143,N_9149);
nor U9392 (N_9392,N_9250,N_9355);
nor U9393 (N_9393,N_9136,N_9134);
or U9394 (N_9394,N_9184,N_9101);
or U9395 (N_9395,N_9091,N_9010);
xor U9396 (N_9396,N_9110,N_9093);
or U9397 (N_9397,N_9115,N_9234);
nand U9398 (N_9398,N_8798,N_9086);
nor U9399 (N_9399,N_9295,N_8936);
nor U9400 (N_9400,N_9005,N_8791);
nor U9401 (N_9401,N_9312,N_8897);
xor U9402 (N_9402,N_9152,N_9156);
xnor U9403 (N_9403,N_8806,N_9138);
xor U9404 (N_9404,N_8861,N_9116);
and U9405 (N_9405,N_8884,N_9037);
nor U9406 (N_9406,N_8995,N_8844);
nand U9407 (N_9407,N_9064,N_9215);
or U9408 (N_9408,N_9246,N_8901);
xnor U9409 (N_9409,N_8804,N_9236);
or U9410 (N_9410,N_9192,N_9291);
nor U9411 (N_9411,N_9300,N_9284);
or U9412 (N_9412,N_9032,N_8951);
or U9413 (N_9413,N_9073,N_9229);
nand U9414 (N_9414,N_9095,N_8824);
or U9415 (N_9415,N_9023,N_8870);
xor U9416 (N_9416,N_9193,N_9287);
or U9417 (N_9417,N_9173,N_9094);
nor U9418 (N_9418,N_8978,N_9230);
nand U9419 (N_9419,N_8838,N_9348);
and U9420 (N_9420,N_8922,N_8776);
nor U9421 (N_9421,N_8882,N_9290);
nor U9422 (N_9422,N_9191,N_8930);
xor U9423 (N_9423,N_8893,N_9084);
or U9424 (N_9424,N_9280,N_9273);
xnor U9425 (N_9425,N_9369,N_9004);
nand U9426 (N_9426,N_8865,N_9218);
nor U9427 (N_9427,N_8815,N_9220);
nand U9428 (N_9428,N_8900,N_9167);
xnor U9429 (N_9429,N_9195,N_9185);
or U9430 (N_9430,N_9219,N_8820);
nand U9431 (N_9431,N_9157,N_9321);
or U9432 (N_9432,N_8841,N_8881);
nand U9433 (N_9433,N_9241,N_8871);
or U9434 (N_9434,N_9140,N_8894);
xnor U9435 (N_9435,N_8760,N_9052);
nand U9436 (N_9436,N_9081,N_8810);
nor U9437 (N_9437,N_9117,N_9170);
or U9438 (N_9438,N_9360,N_8799);
nor U9439 (N_9439,N_8942,N_8949);
or U9440 (N_9440,N_9318,N_8831);
and U9441 (N_9441,N_9337,N_8879);
xnor U9442 (N_9442,N_8965,N_8864);
or U9443 (N_9443,N_9343,N_8797);
nor U9444 (N_9444,N_9024,N_8966);
nor U9445 (N_9445,N_8947,N_9145);
xnor U9446 (N_9446,N_9301,N_8913);
or U9447 (N_9447,N_9200,N_9040);
or U9448 (N_9448,N_8880,N_9126);
or U9449 (N_9449,N_8985,N_8770);
and U9450 (N_9450,N_9161,N_8967);
and U9451 (N_9451,N_9119,N_9089);
or U9452 (N_9452,N_8896,N_9262);
nand U9453 (N_9453,N_9069,N_9154);
nor U9454 (N_9454,N_9212,N_8800);
or U9455 (N_9455,N_9189,N_9031);
and U9456 (N_9456,N_8963,N_8835);
and U9457 (N_9457,N_9045,N_9068);
nor U9458 (N_9458,N_8817,N_9139);
or U9459 (N_9459,N_9351,N_9313);
or U9460 (N_9460,N_8924,N_8925);
xnor U9461 (N_9461,N_8920,N_8857);
xnor U9462 (N_9462,N_9186,N_9374);
nor U9463 (N_9463,N_9281,N_9327);
xnor U9464 (N_9464,N_9171,N_9121);
or U9465 (N_9465,N_8753,N_8998);
or U9466 (N_9466,N_8991,N_8869);
nand U9467 (N_9467,N_9108,N_8766);
and U9468 (N_9468,N_8826,N_9092);
or U9469 (N_9469,N_9225,N_9299);
and U9470 (N_9470,N_8816,N_8763);
or U9471 (N_9471,N_9277,N_9289);
nor U9472 (N_9472,N_8874,N_9151);
nor U9473 (N_9473,N_9335,N_9344);
xor U9474 (N_9474,N_8918,N_8751);
or U9475 (N_9475,N_9309,N_9254);
xor U9476 (N_9476,N_8856,N_9260);
and U9477 (N_9477,N_9333,N_9003);
nand U9478 (N_9478,N_9146,N_8773);
or U9479 (N_9479,N_9100,N_9083);
xor U9480 (N_9480,N_9322,N_9082);
nor U9481 (N_9481,N_8858,N_9067);
and U9482 (N_9482,N_8910,N_8915);
or U9483 (N_9483,N_9224,N_8796);
nor U9484 (N_9484,N_8825,N_8750);
nor U9485 (N_9485,N_8761,N_9261);
and U9486 (N_9486,N_9175,N_8958);
nand U9487 (N_9487,N_8765,N_9270);
and U9488 (N_9488,N_9199,N_9187);
nor U9489 (N_9489,N_8907,N_8916);
or U9490 (N_9490,N_8938,N_9317);
nand U9491 (N_9491,N_9362,N_9012);
nand U9492 (N_9492,N_9060,N_9223);
or U9493 (N_9493,N_9307,N_9283);
nand U9494 (N_9494,N_8756,N_8788);
and U9495 (N_9495,N_9041,N_9373);
xnor U9496 (N_9496,N_9282,N_9368);
nand U9497 (N_9497,N_8781,N_9164);
nand U9498 (N_9498,N_9129,N_8923);
nor U9499 (N_9499,N_9271,N_8828);
xnor U9500 (N_9500,N_8850,N_9204);
nor U9501 (N_9501,N_9341,N_9105);
xor U9502 (N_9502,N_9006,N_9276);
xnor U9503 (N_9503,N_8866,N_8822);
nor U9504 (N_9504,N_9345,N_9206);
or U9505 (N_9505,N_9288,N_9180);
xnor U9506 (N_9506,N_9308,N_9231);
or U9507 (N_9507,N_9063,N_9104);
xnor U9508 (N_9508,N_8886,N_9311);
nor U9509 (N_9509,N_9334,N_9051);
nor U9510 (N_9510,N_9085,N_9044);
nor U9511 (N_9511,N_8987,N_8940);
xnor U9512 (N_9512,N_9314,N_8989);
nor U9513 (N_9513,N_8859,N_9214);
xnor U9514 (N_9514,N_8769,N_8892);
xnor U9515 (N_9515,N_8843,N_8988);
or U9516 (N_9516,N_9346,N_8877);
nand U9517 (N_9517,N_9055,N_8875);
nor U9518 (N_9518,N_8876,N_8891);
nor U9519 (N_9519,N_8883,N_8908);
or U9520 (N_9520,N_9046,N_9183);
nor U9521 (N_9521,N_8846,N_8830);
nor U9522 (N_9522,N_9210,N_9017);
and U9523 (N_9523,N_9118,N_8868);
nor U9524 (N_9524,N_9015,N_9016);
and U9525 (N_9525,N_8842,N_8812);
or U9526 (N_9526,N_8853,N_9326);
and U9527 (N_9527,N_8976,N_9233);
xor U9528 (N_9528,N_9030,N_8778);
or U9529 (N_9529,N_9336,N_9319);
nand U9530 (N_9530,N_9293,N_8762);
nor U9531 (N_9531,N_9266,N_8771);
or U9532 (N_9532,N_9248,N_8974);
nand U9533 (N_9533,N_9370,N_9366);
xnor U9534 (N_9534,N_9315,N_8814);
and U9535 (N_9535,N_9097,N_8755);
nand U9536 (N_9536,N_9099,N_9257);
and U9537 (N_9537,N_9342,N_9147);
xnor U9538 (N_9538,N_8889,N_8937);
xnor U9539 (N_9539,N_9182,N_9286);
nand U9540 (N_9540,N_9077,N_8912);
and U9541 (N_9541,N_9208,N_8961);
and U9542 (N_9542,N_9196,N_9263);
nand U9543 (N_9543,N_9244,N_8809);
nand U9544 (N_9544,N_9194,N_8764);
and U9545 (N_9545,N_9338,N_9159);
and U9546 (N_9546,N_8983,N_9242);
nor U9547 (N_9547,N_9002,N_9127);
xor U9548 (N_9548,N_9324,N_8990);
or U9549 (N_9549,N_8833,N_8803);
nor U9550 (N_9550,N_8909,N_9203);
nor U9551 (N_9551,N_9359,N_9213);
xnor U9552 (N_9552,N_9298,N_9166);
or U9553 (N_9553,N_8899,N_8964);
nor U9554 (N_9554,N_9232,N_8957);
and U9555 (N_9555,N_9172,N_9162);
and U9556 (N_9556,N_9198,N_8954);
nor U9557 (N_9557,N_9240,N_9027);
and U9558 (N_9558,N_9014,N_9259);
nor U9559 (N_9559,N_8847,N_9061);
xnor U9560 (N_9560,N_8849,N_8840);
nor U9561 (N_9561,N_8848,N_9310);
or U9562 (N_9562,N_9128,N_9330);
nand U9563 (N_9563,N_8873,N_9227);
xnor U9564 (N_9564,N_8999,N_9256);
xnor U9565 (N_9565,N_8784,N_9174);
nor U9566 (N_9566,N_8802,N_8981);
or U9567 (N_9567,N_9361,N_8953);
xor U9568 (N_9568,N_8906,N_8813);
nor U9569 (N_9569,N_9120,N_8759);
nor U9570 (N_9570,N_9029,N_9352);
and U9571 (N_9571,N_9053,N_8890);
nor U9572 (N_9572,N_9228,N_9325);
nand U9573 (N_9573,N_9114,N_9305);
and U9574 (N_9574,N_9009,N_8775);
nand U9575 (N_9575,N_9274,N_8888);
xnor U9576 (N_9576,N_9323,N_9150);
or U9577 (N_9577,N_9357,N_8945);
nand U9578 (N_9578,N_9255,N_8905);
nor U9579 (N_9579,N_9306,N_9222);
nor U9580 (N_9580,N_8783,N_9144);
xor U9581 (N_9581,N_9285,N_8903);
and U9582 (N_9582,N_9178,N_9072);
nand U9583 (N_9583,N_9247,N_9316);
xor U9584 (N_9584,N_9339,N_9350);
xor U9585 (N_9585,N_9364,N_8789);
or U9586 (N_9586,N_9303,N_9137);
or U9587 (N_9587,N_9062,N_8933);
xnor U9588 (N_9588,N_8855,N_8948);
or U9589 (N_9589,N_8790,N_9007);
xnor U9590 (N_9590,N_9168,N_8768);
or U9591 (N_9591,N_8782,N_9111);
and U9592 (N_9592,N_8992,N_9155);
or U9593 (N_9593,N_9205,N_9332);
and U9594 (N_9594,N_9272,N_8867);
and U9595 (N_9595,N_8860,N_8960);
xnor U9596 (N_9596,N_8980,N_9080);
or U9597 (N_9597,N_9367,N_9142);
and U9598 (N_9598,N_9304,N_8821);
and U9599 (N_9599,N_9363,N_8950);
or U9600 (N_9600,N_8851,N_8777);
nor U9601 (N_9601,N_8795,N_9226);
xnor U9602 (N_9602,N_9297,N_8801);
or U9603 (N_9603,N_9179,N_8904);
nand U9604 (N_9604,N_9292,N_9113);
xnor U9605 (N_9605,N_8827,N_8752);
nor U9606 (N_9606,N_8996,N_9347);
and U9607 (N_9607,N_9133,N_8972);
xor U9608 (N_9608,N_8962,N_8811);
xnor U9609 (N_9609,N_9264,N_9209);
or U9610 (N_9610,N_8887,N_9028);
nand U9611 (N_9611,N_8917,N_9087);
and U9612 (N_9612,N_8994,N_8939);
nand U9613 (N_9613,N_8786,N_9036);
nand U9614 (N_9614,N_9098,N_9019);
or U9615 (N_9615,N_9071,N_9057);
nand U9616 (N_9616,N_9340,N_9021);
or U9617 (N_9617,N_8829,N_9078);
nor U9618 (N_9618,N_9124,N_8895);
nand U9619 (N_9619,N_8931,N_9216);
nor U9620 (N_9620,N_8982,N_8959);
nor U9621 (N_9621,N_8984,N_9043);
nor U9622 (N_9622,N_9328,N_8971);
and U9623 (N_9623,N_8969,N_9239);
xnor U9624 (N_9624,N_8975,N_9331);
or U9625 (N_9625,N_8818,N_9070);
nand U9626 (N_9626,N_9267,N_8852);
or U9627 (N_9627,N_9122,N_9160);
nor U9628 (N_9628,N_9048,N_9279);
xnor U9629 (N_9629,N_9011,N_9090);
nor U9630 (N_9630,N_9278,N_9106);
xnor U9631 (N_9631,N_8805,N_9197);
nand U9632 (N_9632,N_8839,N_9221);
and U9633 (N_9633,N_8819,N_9371);
or U9634 (N_9634,N_9258,N_9353);
xnor U9635 (N_9635,N_8946,N_8977);
nand U9636 (N_9636,N_8902,N_8898);
nand U9637 (N_9637,N_8832,N_8793);
nand U9638 (N_9638,N_9249,N_9349);
xor U9639 (N_9639,N_9265,N_9354);
xor U9640 (N_9640,N_9365,N_8862);
nor U9641 (N_9641,N_8935,N_9131);
or U9642 (N_9642,N_8767,N_9008);
nor U9643 (N_9643,N_8878,N_9243);
or U9644 (N_9644,N_9075,N_8932);
and U9645 (N_9645,N_9269,N_9018);
or U9646 (N_9646,N_8911,N_9109);
nor U9647 (N_9647,N_9135,N_8997);
or U9648 (N_9648,N_8807,N_9056);
xnor U9649 (N_9649,N_8993,N_8955);
or U9650 (N_9650,N_8754,N_8970);
and U9651 (N_9651,N_9035,N_9356);
or U9652 (N_9652,N_9177,N_8837);
nand U9653 (N_9653,N_8772,N_9296);
xnor U9654 (N_9654,N_9125,N_9079);
nand U9655 (N_9655,N_8928,N_8914);
and U9656 (N_9656,N_9026,N_9207);
nor U9657 (N_9657,N_9217,N_9275);
xor U9658 (N_9658,N_8872,N_8979);
or U9659 (N_9659,N_9165,N_8968);
nor U9660 (N_9660,N_8808,N_9020);
nor U9661 (N_9661,N_9112,N_9096);
or U9662 (N_9662,N_8927,N_9132);
nor U9663 (N_9663,N_9013,N_9237);
or U9664 (N_9664,N_8854,N_8934);
nor U9665 (N_9665,N_8926,N_8758);
nor U9666 (N_9666,N_9169,N_8941);
or U9667 (N_9667,N_9268,N_9329);
nand U9668 (N_9668,N_8943,N_9074);
nand U9669 (N_9669,N_9251,N_8780);
nor U9670 (N_9670,N_9050,N_9034);
nand U9671 (N_9671,N_9022,N_8952);
xor U9672 (N_9672,N_9107,N_9066);
or U9673 (N_9673,N_9054,N_9253);
and U9674 (N_9674,N_9188,N_9320);
nor U9675 (N_9675,N_9358,N_8834);
and U9676 (N_9676,N_8774,N_8785);
and U9677 (N_9677,N_9211,N_9153);
nand U9678 (N_9678,N_8779,N_9130);
nand U9679 (N_9679,N_9181,N_8885);
or U9680 (N_9680,N_9294,N_8823);
or U9681 (N_9681,N_8845,N_9163);
nor U9682 (N_9682,N_8921,N_9201);
nor U9683 (N_9683,N_8929,N_9049);
or U9684 (N_9684,N_9202,N_8986);
nand U9685 (N_9685,N_9123,N_9158);
nor U9686 (N_9686,N_9235,N_8794);
and U9687 (N_9687,N_9372,N_9306);
and U9688 (N_9688,N_9314,N_9331);
nand U9689 (N_9689,N_8970,N_9139);
nand U9690 (N_9690,N_8897,N_8904);
nand U9691 (N_9691,N_9247,N_9331);
nand U9692 (N_9692,N_9317,N_9229);
and U9693 (N_9693,N_8979,N_8770);
nor U9694 (N_9694,N_8784,N_9335);
nor U9695 (N_9695,N_9338,N_8807);
xor U9696 (N_9696,N_9044,N_8950);
nand U9697 (N_9697,N_9208,N_9243);
or U9698 (N_9698,N_8848,N_8944);
or U9699 (N_9699,N_9014,N_8876);
or U9700 (N_9700,N_8872,N_9194);
and U9701 (N_9701,N_9294,N_8751);
nand U9702 (N_9702,N_8829,N_9265);
nand U9703 (N_9703,N_9154,N_8788);
xnor U9704 (N_9704,N_9361,N_9070);
nor U9705 (N_9705,N_9006,N_8759);
xnor U9706 (N_9706,N_8806,N_9251);
and U9707 (N_9707,N_9067,N_9060);
nor U9708 (N_9708,N_9308,N_9099);
or U9709 (N_9709,N_8875,N_9036);
and U9710 (N_9710,N_8975,N_9318);
or U9711 (N_9711,N_9143,N_8821);
nand U9712 (N_9712,N_8935,N_9000);
or U9713 (N_9713,N_8829,N_8869);
xor U9714 (N_9714,N_8838,N_8888);
nor U9715 (N_9715,N_8839,N_8986);
nand U9716 (N_9716,N_9068,N_9059);
and U9717 (N_9717,N_8979,N_9308);
xor U9718 (N_9718,N_9215,N_8948);
nand U9719 (N_9719,N_9171,N_9374);
nand U9720 (N_9720,N_9165,N_9257);
and U9721 (N_9721,N_9044,N_8982);
nor U9722 (N_9722,N_9360,N_9073);
or U9723 (N_9723,N_9060,N_8849);
xor U9724 (N_9724,N_8930,N_9259);
or U9725 (N_9725,N_9255,N_9027);
nand U9726 (N_9726,N_8842,N_8895);
or U9727 (N_9727,N_9209,N_9002);
nor U9728 (N_9728,N_9227,N_9028);
xor U9729 (N_9729,N_8950,N_9271);
xnor U9730 (N_9730,N_8845,N_9025);
nor U9731 (N_9731,N_9210,N_9285);
and U9732 (N_9732,N_9108,N_9085);
nor U9733 (N_9733,N_9071,N_8944);
nor U9734 (N_9734,N_8816,N_9374);
and U9735 (N_9735,N_9086,N_9363);
and U9736 (N_9736,N_9305,N_9058);
xor U9737 (N_9737,N_9073,N_8952);
or U9738 (N_9738,N_8865,N_9175);
or U9739 (N_9739,N_9322,N_9257);
and U9740 (N_9740,N_9342,N_9195);
nor U9741 (N_9741,N_8943,N_9105);
nor U9742 (N_9742,N_9068,N_8860);
or U9743 (N_9743,N_8992,N_8801);
xnor U9744 (N_9744,N_9029,N_9142);
and U9745 (N_9745,N_9034,N_9210);
and U9746 (N_9746,N_8885,N_8799);
and U9747 (N_9747,N_8985,N_9049);
and U9748 (N_9748,N_9316,N_9234);
nor U9749 (N_9749,N_9341,N_9004);
nand U9750 (N_9750,N_9309,N_8893);
or U9751 (N_9751,N_8993,N_8775);
and U9752 (N_9752,N_8906,N_9361);
and U9753 (N_9753,N_9327,N_9082);
and U9754 (N_9754,N_9044,N_8815);
xor U9755 (N_9755,N_9071,N_9314);
nand U9756 (N_9756,N_9061,N_9361);
and U9757 (N_9757,N_8836,N_9016);
and U9758 (N_9758,N_9114,N_9060);
nor U9759 (N_9759,N_9106,N_9123);
or U9760 (N_9760,N_9210,N_9127);
nor U9761 (N_9761,N_9270,N_9112);
nor U9762 (N_9762,N_9209,N_9340);
xor U9763 (N_9763,N_9130,N_8893);
and U9764 (N_9764,N_9309,N_9080);
nor U9765 (N_9765,N_9079,N_9190);
and U9766 (N_9766,N_9217,N_8769);
xor U9767 (N_9767,N_8988,N_8875);
and U9768 (N_9768,N_8762,N_9132);
nor U9769 (N_9769,N_9283,N_9256);
nand U9770 (N_9770,N_8879,N_8881);
nand U9771 (N_9771,N_9245,N_8994);
nor U9772 (N_9772,N_8776,N_9300);
nor U9773 (N_9773,N_9041,N_8810);
xor U9774 (N_9774,N_8800,N_8807);
nor U9775 (N_9775,N_9027,N_9281);
and U9776 (N_9776,N_8897,N_9328);
or U9777 (N_9777,N_9105,N_9276);
nand U9778 (N_9778,N_9335,N_9369);
nand U9779 (N_9779,N_9039,N_9136);
nand U9780 (N_9780,N_9028,N_9334);
and U9781 (N_9781,N_8924,N_9283);
nand U9782 (N_9782,N_9168,N_9283);
nand U9783 (N_9783,N_9157,N_8921);
nor U9784 (N_9784,N_9319,N_9213);
nor U9785 (N_9785,N_9304,N_9028);
nor U9786 (N_9786,N_9187,N_8803);
or U9787 (N_9787,N_9057,N_8798);
nand U9788 (N_9788,N_8902,N_9243);
nor U9789 (N_9789,N_9273,N_9162);
xnor U9790 (N_9790,N_8856,N_8953);
nand U9791 (N_9791,N_9245,N_8956);
nand U9792 (N_9792,N_9149,N_9035);
xor U9793 (N_9793,N_8825,N_9361);
or U9794 (N_9794,N_9259,N_8760);
nor U9795 (N_9795,N_8975,N_8983);
xnor U9796 (N_9796,N_9143,N_9141);
and U9797 (N_9797,N_9331,N_8854);
nand U9798 (N_9798,N_9205,N_9054);
or U9799 (N_9799,N_8998,N_8887);
and U9800 (N_9800,N_8752,N_8814);
xnor U9801 (N_9801,N_9351,N_9028);
xnor U9802 (N_9802,N_8905,N_8966);
xor U9803 (N_9803,N_8822,N_8938);
or U9804 (N_9804,N_8929,N_9107);
and U9805 (N_9805,N_8819,N_8929);
or U9806 (N_9806,N_9207,N_9204);
nand U9807 (N_9807,N_9042,N_9212);
nor U9808 (N_9808,N_9076,N_9009);
nand U9809 (N_9809,N_9107,N_8996);
nor U9810 (N_9810,N_8892,N_8973);
nand U9811 (N_9811,N_9373,N_8933);
xor U9812 (N_9812,N_9345,N_9031);
xor U9813 (N_9813,N_9071,N_9141);
and U9814 (N_9814,N_8943,N_9229);
nand U9815 (N_9815,N_8990,N_9357);
nand U9816 (N_9816,N_9065,N_8939);
nand U9817 (N_9817,N_8793,N_9085);
or U9818 (N_9818,N_8926,N_9238);
nand U9819 (N_9819,N_8893,N_9200);
nand U9820 (N_9820,N_9038,N_9146);
and U9821 (N_9821,N_8941,N_8836);
nand U9822 (N_9822,N_8760,N_9357);
or U9823 (N_9823,N_9162,N_8862);
or U9824 (N_9824,N_8894,N_9334);
nand U9825 (N_9825,N_9109,N_8927);
or U9826 (N_9826,N_8869,N_9318);
xor U9827 (N_9827,N_9026,N_8954);
and U9828 (N_9828,N_9172,N_9148);
nand U9829 (N_9829,N_9087,N_9276);
nor U9830 (N_9830,N_9039,N_8988);
nor U9831 (N_9831,N_8766,N_9204);
nor U9832 (N_9832,N_9294,N_9028);
and U9833 (N_9833,N_8779,N_9315);
or U9834 (N_9834,N_8868,N_8943);
or U9835 (N_9835,N_8994,N_8781);
nor U9836 (N_9836,N_9194,N_9356);
or U9837 (N_9837,N_9365,N_9155);
nand U9838 (N_9838,N_9303,N_9007);
nor U9839 (N_9839,N_9063,N_9195);
nor U9840 (N_9840,N_8831,N_9213);
or U9841 (N_9841,N_9073,N_8972);
xnor U9842 (N_9842,N_8754,N_9276);
nand U9843 (N_9843,N_8921,N_8950);
xor U9844 (N_9844,N_8922,N_8882);
xor U9845 (N_9845,N_8828,N_8816);
or U9846 (N_9846,N_9173,N_9044);
nand U9847 (N_9847,N_8959,N_8895);
or U9848 (N_9848,N_8840,N_8997);
xnor U9849 (N_9849,N_9152,N_8893);
nor U9850 (N_9850,N_9248,N_9077);
xnor U9851 (N_9851,N_9234,N_8771);
nand U9852 (N_9852,N_9090,N_8832);
and U9853 (N_9853,N_8843,N_8765);
xor U9854 (N_9854,N_9311,N_9110);
or U9855 (N_9855,N_9334,N_8819);
nand U9856 (N_9856,N_9055,N_8989);
nor U9857 (N_9857,N_9147,N_8758);
or U9858 (N_9858,N_9212,N_9136);
nand U9859 (N_9859,N_9337,N_9157);
or U9860 (N_9860,N_8862,N_9176);
or U9861 (N_9861,N_9206,N_9314);
and U9862 (N_9862,N_9350,N_9323);
xor U9863 (N_9863,N_8862,N_8854);
and U9864 (N_9864,N_8920,N_8861);
nand U9865 (N_9865,N_8935,N_8930);
or U9866 (N_9866,N_8828,N_8919);
nor U9867 (N_9867,N_9252,N_9349);
nor U9868 (N_9868,N_8862,N_9089);
nand U9869 (N_9869,N_9341,N_9026);
xnor U9870 (N_9870,N_9107,N_9276);
nand U9871 (N_9871,N_9027,N_9083);
and U9872 (N_9872,N_9094,N_8991);
nor U9873 (N_9873,N_9317,N_9189);
nand U9874 (N_9874,N_9272,N_9000);
nand U9875 (N_9875,N_8979,N_9001);
nor U9876 (N_9876,N_9022,N_9273);
or U9877 (N_9877,N_8751,N_9164);
nor U9878 (N_9878,N_9109,N_9029);
nor U9879 (N_9879,N_8916,N_9368);
and U9880 (N_9880,N_9187,N_8815);
xnor U9881 (N_9881,N_9177,N_8898);
and U9882 (N_9882,N_9341,N_9049);
and U9883 (N_9883,N_8973,N_9078);
and U9884 (N_9884,N_8835,N_8792);
nor U9885 (N_9885,N_9045,N_9042);
xor U9886 (N_9886,N_9258,N_8869);
or U9887 (N_9887,N_8862,N_9345);
and U9888 (N_9888,N_8980,N_8890);
xor U9889 (N_9889,N_8952,N_9335);
nor U9890 (N_9890,N_9297,N_9157);
nor U9891 (N_9891,N_9034,N_9336);
and U9892 (N_9892,N_9307,N_9168);
and U9893 (N_9893,N_8827,N_9229);
or U9894 (N_9894,N_8997,N_8852);
nand U9895 (N_9895,N_9363,N_8907);
nand U9896 (N_9896,N_9370,N_8929);
nand U9897 (N_9897,N_9037,N_9268);
or U9898 (N_9898,N_8877,N_8855);
or U9899 (N_9899,N_9313,N_8813);
nor U9900 (N_9900,N_9280,N_9319);
xnor U9901 (N_9901,N_9154,N_9208);
and U9902 (N_9902,N_9200,N_8909);
and U9903 (N_9903,N_8839,N_8962);
nand U9904 (N_9904,N_8858,N_9301);
or U9905 (N_9905,N_8821,N_9100);
xor U9906 (N_9906,N_8928,N_9200);
nor U9907 (N_9907,N_9102,N_8839);
or U9908 (N_9908,N_9152,N_9002);
or U9909 (N_9909,N_9195,N_8884);
and U9910 (N_9910,N_9316,N_9132);
or U9911 (N_9911,N_8906,N_8805);
nor U9912 (N_9912,N_8865,N_9090);
nand U9913 (N_9913,N_8882,N_9335);
and U9914 (N_9914,N_9072,N_8997);
or U9915 (N_9915,N_9098,N_8855);
or U9916 (N_9916,N_9173,N_9348);
or U9917 (N_9917,N_8827,N_8824);
nand U9918 (N_9918,N_9294,N_8925);
or U9919 (N_9919,N_9297,N_8924);
and U9920 (N_9920,N_9352,N_8822);
xnor U9921 (N_9921,N_9262,N_8844);
nand U9922 (N_9922,N_8982,N_8784);
xor U9923 (N_9923,N_9230,N_9204);
or U9924 (N_9924,N_9128,N_8814);
nor U9925 (N_9925,N_8780,N_9027);
or U9926 (N_9926,N_9321,N_8991);
and U9927 (N_9927,N_8869,N_8938);
or U9928 (N_9928,N_8834,N_9207);
or U9929 (N_9929,N_8905,N_8818);
xnor U9930 (N_9930,N_8888,N_9008);
or U9931 (N_9931,N_9224,N_9205);
or U9932 (N_9932,N_9076,N_8944);
nor U9933 (N_9933,N_8867,N_8992);
nor U9934 (N_9934,N_9211,N_9001);
or U9935 (N_9935,N_9058,N_9230);
nand U9936 (N_9936,N_9193,N_9304);
and U9937 (N_9937,N_9256,N_9051);
and U9938 (N_9938,N_8802,N_8812);
or U9939 (N_9939,N_9060,N_9233);
xor U9940 (N_9940,N_9279,N_9160);
nand U9941 (N_9941,N_9114,N_8905);
nand U9942 (N_9942,N_9113,N_8906);
or U9943 (N_9943,N_8992,N_8764);
or U9944 (N_9944,N_8995,N_9066);
xor U9945 (N_9945,N_9286,N_9049);
or U9946 (N_9946,N_9177,N_9217);
or U9947 (N_9947,N_8780,N_9345);
and U9948 (N_9948,N_9231,N_8927);
xnor U9949 (N_9949,N_9182,N_9241);
nor U9950 (N_9950,N_9237,N_9037);
and U9951 (N_9951,N_9216,N_9127);
and U9952 (N_9952,N_9165,N_8754);
or U9953 (N_9953,N_8837,N_8779);
nand U9954 (N_9954,N_8813,N_9334);
or U9955 (N_9955,N_9134,N_8809);
xnor U9956 (N_9956,N_8803,N_9350);
xor U9957 (N_9957,N_9293,N_9175);
and U9958 (N_9958,N_8854,N_9136);
nor U9959 (N_9959,N_9292,N_8805);
or U9960 (N_9960,N_9000,N_8834);
and U9961 (N_9961,N_9159,N_9068);
or U9962 (N_9962,N_9271,N_9047);
nor U9963 (N_9963,N_9368,N_9012);
or U9964 (N_9964,N_8941,N_9320);
nor U9965 (N_9965,N_9161,N_8861);
nand U9966 (N_9966,N_9361,N_9141);
nand U9967 (N_9967,N_9359,N_8872);
xnor U9968 (N_9968,N_9076,N_9108);
and U9969 (N_9969,N_8782,N_9228);
nand U9970 (N_9970,N_8797,N_9189);
xnor U9971 (N_9971,N_9031,N_9293);
or U9972 (N_9972,N_8766,N_9122);
and U9973 (N_9973,N_9168,N_9240);
nor U9974 (N_9974,N_8840,N_8803);
nand U9975 (N_9975,N_9034,N_8837);
and U9976 (N_9976,N_8779,N_8750);
and U9977 (N_9977,N_9175,N_8803);
nand U9978 (N_9978,N_8842,N_8788);
xnor U9979 (N_9979,N_8827,N_9315);
nand U9980 (N_9980,N_9178,N_8904);
nor U9981 (N_9981,N_8791,N_8888);
nand U9982 (N_9982,N_9103,N_9116);
or U9983 (N_9983,N_9171,N_9118);
or U9984 (N_9984,N_9363,N_9092);
nand U9985 (N_9985,N_9274,N_9252);
xnor U9986 (N_9986,N_9204,N_9258);
nor U9987 (N_9987,N_9223,N_9161);
and U9988 (N_9988,N_8940,N_8829);
nand U9989 (N_9989,N_8826,N_9159);
and U9990 (N_9990,N_8888,N_9200);
or U9991 (N_9991,N_8755,N_9032);
nand U9992 (N_9992,N_8803,N_9263);
nor U9993 (N_9993,N_8899,N_9093);
and U9994 (N_9994,N_8780,N_9307);
or U9995 (N_9995,N_9295,N_8854);
and U9996 (N_9996,N_8994,N_8789);
nor U9997 (N_9997,N_9037,N_8866);
and U9998 (N_9998,N_8783,N_8897);
xnor U9999 (N_9999,N_9258,N_9218);
and U10000 (N_10000,N_9888,N_9394);
or U10001 (N_10001,N_9560,N_9674);
nand U10002 (N_10002,N_9598,N_9833);
or U10003 (N_10003,N_9995,N_9490);
xnor U10004 (N_10004,N_9879,N_9788);
or U10005 (N_10005,N_9476,N_9387);
and U10006 (N_10006,N_9969,N_9766);
nor U10007 (N_10007,N_9439,N_9672);
or U10008 (N_10008,N_9472,N_9911);
xor U10009 (N_10009,N_9548,N_9675);
or U10010 (N_10010,N_9994,N_9782);
nand U10011 (N_10011,N_9586,N_9498);
xor U10012 (N_10012,N_9558,N_9912);
xor U10013 (N_10013,N_9778,N_9650);
and U10014 (N_10014,N_9799,N_9802);
or U10015 (N_10015,N_9602,N_9666);
and U10016 (N_10016,N_9976,N_9735);
or U10017 (N_10017,N_9803,N_9577);
nand U10018 (N_10018,N_9798,N_9436);
nor U10019 (N_10019,N_9863,N_9856);
xnor U10020 (N_10020,N_9392,N_9448);
nor U10021 (N_10021,N_9730,N_9660);
xor U10022 (N_10022,N_9567,N_9382);
xnor U10023 (N_10023,N_9551,N_9688);
nand U10024 (N_10024,N_9478,N_9477);
xnor U10025 (N_10025,N_9920,N_9603);
nor U10026 (N_10026,N_9707,N_9491);
and U10027 (N_10027,N_9406,N_9703);
nand U10028 (N_10028,N_9885,N_9457);
nor U10029 (N_10029,N_9823,N_9963);
or U10030 (N_10030,N_9729,N_9752);
nand U10031 (N_10031,N_9935,N_9658);
nor U10032 (N_10032,N_9618,N_9668);
nand U10033 (N_10033,N_9619,N_9525);
or U10034 (N_10034,N_9463,N_9687);
nand U10035 (N_10035,N_9588,N_9717);
nor U10036 (N_10036,N_9846,N_9763);
and U10037 (N_10037,N_9653,N_9874);
or U10038 (N_10038,N_9924,N_9445);
xor U10039 (N_10039,N_9851,N_9795);
nor U10040 (N_10040,N_9950,N_9726);
and U10041 (N_10041,N_9840,N_9634);
nor U10042 (N_10042,N_9520,N_9628);
nor U10043 (N_10043,N_9971,N_9614);
xor U10044 (N_10044,N_9836,N_9903);
xor U10045 (N_10045,N_9739,N_9404);
and U10046 (N_10046,N_9776,N_9972);
nand U10047 (N_10047,N_9649,N_9473);
xor U10048 (N_10048,N_9461,N_9553);
and U10049 (N_10049,N_9504,N_9403);
or U10050 (N_10050,N_9640,N_9824);
or U10051 (N_10051,N_9609,N_9984);
nand U10052 (N_10052,N_9923,N_9422);
xnor U10053 (N_10053,N_9973,N_9761);
nand U10054 (N_10054,N_9952,N_9714);
and U10055 (N_10055,N_9847,N_9751);
nor U10056 (N_10056,N_9443,N_9641);
or U10057 (N_10057,N_9697,N_9512);
or U10058 (N_10058,N_9725,N_9870);
or U10059 (N_10059,N_9617,N_9575);
nor U10060 (N_10060,N_9749,N_9919);
or U10061 (N_10061,N_9953,N_9554);
or U10062 (N_10062,N_9861,N_9764);
nor U10063 (N_10063,N_9845,N_9616);
nand U10064 (N_10064,N_9775,N_9813);
nor U10065 (N_10065,N_9626,N_9702);
or U10066 (N_10066,N_9632,N_9945);
nand U10067 (N_10067,N_9471,N_9708);
nand U10068 (N_10068,N_9580,N_9837);
and U10069 (N_10069,N_9664,N_9937);
nand U10070 (N_10070,N_9777,N_9936);
nand U10071 (N_10071,N_9493,N_9916);
nor U10072 (N_10072,N_9526,N_9635);
nand U10073 (N_10073,N_9427,N_9860);
nor U10074 (N_10074,N_9850,N_9682);
or U10075 (N_10075,N_9947,N_9878);
nand U10076 (N_10076,N_9515,N_9955);
and U10077 (N_10077,N_9420,N_9556);
xor U10078 (N_10078,N_9906,N_9881);
and U10079 (N_10079,N_9582,N_9429);
nand U10080 (N_10080,N_9921,N_9931);
xor U10081 (N_10081,N_9639,N_9388);
xnor U10082 (N_10082,N_9692,N_9662);
nand U10083 (N_10083,N_9760,N_9691);
nand U10084 (N_10084,N_9742,N_9985);
xor U10085 (N_10085,N_9882,N_9944);
and U10086 (N_10086,N_9780,N_9741);
or U10087 (N_10087,N_9900,N_9711);
and U10088 (N_10088,N_9822,N_9411);
nand U10089 (N_10089,N_9982,N_9713);
nand U10090 (N_10090,N_9852,N_9880);
xor U10091 (N_10091,N_9510,N_9440);
nor U10092 (N_10092,N_9928,N_9561);
and U10093 (N_10093,N_9865,N_9968);
and U10094 (N_10094,N_9452,N_9986);
nor U10095 (N_10095,N_9670,N_9768);
and U10096 (N_10096,N_9869,N_9636);
xor U10097 (N_10097,N_9734,N_9539);
or U10098 (N_10098,N_9530,N_9622);
xnor U10099 (N_10099,N_9395,N_9638);
xor U10100 (N_10100,N_9468,N_9611);
nand U10101 (N_10101,N_9643,N_9926);
and U10102 (N_10102,N_9932,N_9594);
nor U10103 (N_10103,N_9533,N_9627);
nand U10104 (N_10104,N_9380,N_9954);
xor U10105 (N_10105,N_9946,N_9434);
and U10106 (N_10106,N_9699,N_9483);
nand U10107 (N_10107,N_9785,N_9651);
nand U10108 (N_10108,N_9905,N_9781);
nand U10109 (N_10109,N_9683,N_9818);
xor U10110 (N_10110,N_9499,N_9508);
nor U10111 (N_10111,N_9759,N_9830);
nor U10112 (N_10112,N_9466,N_9592);
nand U10113 (N_10113,N_9779,N_9571);
nand U10114 (N_10114,N_9872,N_9514);
or U10115 (N_10115,N_9416,N_9956);
nor U10116 (N_10116,N_9513,N_9893);
nor U10117 (N_10117,N_9569,N_9654);
and U10118 (N_10118,N_9549,N_9506);
nor U10119 (N_10119,N_9601,N_9964);
and U10120 (N_10120,N_9787,N_9728);
or U10121 (N_10121,N_9531,N_9769);
or U10122 (N_10122,N_9494,N_9858);
and U10123 (N_10123,N_9756,N_9610);
and U10124 (N_10124,N_9607,N_9873);
and U10125 (N_10125,N_9907,N_9480);
and U10126 (N_10126,N_9537,N_9974);
nor U10127 (N_10127,N_9705,N_9828);
or U10128 (N_10128,N_9831,N_9983);
and U10129 (N_10129,N_9421,N_9811);
xor U10130 (N_10130,N_9574,N_9904);
and U10131 (N_10131,N_9564,N_9747);
and U10132 (N_10132,N_9389,N_9940);
or U10133 (N_10133,N_9686,N_9423);
nor U10134 (N_10134,N_9736,N_9939);
nand U10135 (N_10135,N_9458,N_9765);
nand U10136 (N_10136,N_9536,N_9442);
xor U10137 (N_10137,N_9385,N_9876);
nor U10138 (N_10138,N_9678,N_9378);
xnor U10139 (N_10139,N_9857,N_9843);
nand U10140 (N_10140,N_9910,N_9731);
or U10141 (N_10141,N_9629,N_9659);
nand U10142 (N_10142,N_9425,N_9521);
and U10143 (N_10143,N_9482,N_9913);
or U10144 (N_10144,N_9993,N_9848);
nand U10145 (N_10145,N_9829,N_9431);
nor U10146 (N_10146,N_9435,N_9894);
nand U10147 (N_10147,N_9732,N_9975);
nor U10148 (N_10148,N_9897,N_9583);
nand U10149 (N_10149,N_9693,N_9767);
or U10150 (N_10150,N_9849,N_9433);
xor U10151 (N_10151,N_9698,N_9929);
and U10152 (N_10152,N_9424,N_9637);
xnor U10153 (N_10153,N_9596,N_9854);
nor U10154 (N_10154,N_9901,N_9806);
xnor U10155 (N_10155,N_9773,N_9853);
nand U10156 (N_10156,N_9718,N_9943);
xor U10157 (N_10157,N_9623,N_9656);
nand U10158 (N_10158,N_9992,N_9820);
or U10159 (N_10159,N_9685,N_9398);
nand U10160 (N_10160,N_9500,N_9488);
and U10161 (N_10161,N_9608,N_9474);
and U10162 (N_10162,N_9546,N_9645);
nor U10163 (N_10163,N_9426,N_9704);
nor U10164 (N_10164,N_9563,N_9814);
nor U10165 (N_10165,N_9565,N_9690);
or U10166 (N_10166,N_9450,N_9712);
nand U10167 (N_10167,N_9587,N_9797);
xnor U10168 (N_10168,N_9505,N_9597);
or U10169 (N_10169,N_9405,N_9784);
or U10170 (N_10170,N_9511,N_9562);
xnor U10171 (N_10171,N_9757,N_9796);
xor U10172 (N_10172,N_9838,N_9834);
nand U10173 (N_10173,N_9740,N_9459);
nand U10174 (N_10174,N_9579,N_9573);
xor U10175 (N_10175,N_9438,N_9807);
nor U10176 (N_10176,N_9475,N_9677);
and U10177 (N_10177,N_9557,N_9612);
nand U10178 (N_10178,N_9642,N_9646);
and U10179 (N_10179,N_9967,N_9960);
or U10180 (N_10180,N_9680,N_9529);
or U10181 (N_10181,N_9671,N_9655);
and U10182 (N_10182,N_9884,N_9419);
nand U10183 (N_10183,N_9615,N_9783);
and U10184 (N_10184,N_9977,N_9733);
nand U10185 (N_10185,N_9484,N_9821);
and U10186 (N_10186,N_9987,N_9408);
xnor U10187 (N_10187,N_9613,N_9750);
nor U10188 (N_10188,N_9430,N_9379);
xnor U10189 (N_10189,N_9397,N_9962);
or U10190 (N_10190,N_9891,N_9812);
nor U10191 (N_10191,N_9815,N_9770);
xor U10192 (N_10192,N_9700,N_9545);
xnor U10193 (N_10193,N_9451,N_9620);
nor U10194 (N_10194,N_9914,N_9523);
nand U10195 (N_10195,N_9844,N_9754);
xor U10196 (N_10196,N_9669,N_9927);
or U10197 (N_10197,N_9578,N_9859);
or U10198 (N_10198,N_9599,N_9661);
and U10199 (N_10199,N_9925,N_9710);
nand U10200 (N_10200,N_9386,N_9990);
nor U10201 (N_10201,N_9441,N_9786);
and U10202 (N_10202,N_9400,N_9552);
nor U10203 (N_10203,N_9867,N_9721);
and U10204 (N_10204,N_9720,N_9715);
and U10205 (N_10205,N_9809,N_9393);
and U10206 (N_10206,N_9410,N_9486);
nand U10207 (N_10207,N_9509,N_9942);
nand U10208 (N_10208,N_9444,N_9391);
nor U10209 (N_10209,N_9489,N_9568);
nand U10210 (N_10210,N_9501,N_9755);
nor U10211 (N_10211,N_9572,N_9970);
nor U10212 (N_10212,N_9738,N_9590);
nor U10213 (N_10213,N_9496,N_9892);
nor U10214 (N_10214,N_9909,N_9934);
xnor U10215 (N_10215,N_9998,N_9647);
and U10216 (N_10216,N_9566,N_9415);
or U10217 (N_10217,N_9600,N_9522);
nor U10218 (N_10218,N_9447,N_9948);
or U10219 (N_10219,N_9817,N_9502);
xor U10220 (N_10220,N_9991,N_9414);
and U10221 (N_10221,N_9538,N_9915);
nand U10222 (N_10222,N_9465,N_9542);
xnor U10223 (N_10223,N_9723,N_9673);
or U10224 (N_10224,N_9746,N_9957);
xor U10225 (N_10225,N_9396,N_9709);
and U10226 (N_10226,N_9581,N_9771);
nor U10227 (N_10227,N_9743,N_9428);
and U10228 (N_10228,N_9625,N_9469);
and U10229 (N_10229,N_9604,N_9996);
nand U10230 (N_10230,N_9933,N_9958);
nor U10231 (N_10231,N_9930,N_9497);
or U10232 (N_10232,N_9988,N_9652);
or U10233 (N_10233,N_9528,N_9722);
xnor U10234 (N_10234,N_9832,N_9657);
and U10235 (N_10235,N_9895,N_9593);
xnor U10236 (N_10236,N_9667,N_9890);
or U10237 (N_10237,N_9621,N_9432);
nor U10238 (N_10238,N_9676,N_9999);
or U10239 (N_10239,N_9997,N_9455);
or U10240 (N_10240,N_9877,N_9989);
nor U10241 (N_10241,N_9544,N_9981);
or U10242 (N_10242,N_9794,N_9527);
nor U10243 (N_10243,N_9437,N_9898);
and U10244 (N_10244,N_9390,N_9381);
xnor U10245 (N_10245,N_9835,N_9744);
and U10246 (N_10246,N_9470,N_9449);
xor U10247 (N_10247,N_9547,N_9941);
xor U10248 (N_10248,N_9978,N_9748);
and U10249 (N_10249,N_9631,N_9516);
nor U10250 (N_10250,N_9716,N_9789);
xor U10251 (N_10251,N_9805,N_9980);
xor U10252 (N_10252,N_9827,N_9816);
nor U10253 (N_10253,N_9532,N_9868);
nor U10254 (N_10254,N_9495,N_9462);
nand U10255 (N_10255,N_9464,N_9790);
or U10256 (N_10256,N_9866,N_9663);
and U10257 (N_10257,N_9961,N_9899);
xor U10258 (N_10258,N_9485,N_9375);
nand U10259 (N_10259,N_9413,N_9922);
nor U10260 (N_10260,N_9862,N_9585);
nor U10261 (N_10261,N_9684,N_9503);
nand U10262 (N_10262,N_9456,N_9519);
nand U10263 (N_10263,N_9801,N_9706);
and U10264 (N_10264,N_9605,N_9409);
and U10265 (N_10265,N_9467,N_9535);
and U10266 (N_10266,N_9804,N_9479);
xnor U10267 (N_10267,N_9772,N_9648);
or U10268 (N_10268,N_9446,N_9758);
nor U10269 (N_10269,N_9606,N_9959);
xor U10270 (N_10270,N_9384,N_9917);
or U10271 (N_10271,N_9896,N_9417);
nor U10272 (N_10272,N_9460,N_9689);
nand U10273 (N_10273,N_9595,N_9402);
xnor U10274 (N_10274,N_9633,N_9412);
or U10275 (N_10275,N_9696,N_9745);
nand U10276 (N_10276,N_9694,N_9871);
nor U10277 (N_10277,N_9454,N_9679);
nor U10278 (N_10278,N_9819,N_9918);
nor U10279 (N_10279,N_9543,N_9951);
nand U10280 (N_10280,N_9517,N_9695);
and U10281 (N_10281,N_9701,N_9518);
xnor U10282 (N_10282,N_9979,N_9541);
or U10283 (N_10283,N_9902,N_9762);
or U10284 (N_10284,N_9887,N_9570);
xor U10285 (N_10285,N_9753,N_9841);
nand U10286 (N_10286,N_9453,N_9376);
xor U10287 (N_10287,N_9883,N_9377);
and U10288 (N_10288,N_9727,N_9793);
and U10289 (N_10289,N_9576,N_9889);
and U10290 (N_10290,N_9584,N_9908);
nor U10291 (N_10291,N_9383,N_9825);
nand U10292 (N_10292,N_9589,N_9966);
nor U10293 (N_10293,N_9492,N_9524);
or U10294 (N_10294,N_9886,N_9842);
nor U10295 (N_10295,N_9418,N_9399);
nand U10296 (N_10296,N_9826,N_9737);
and U10297 (N_10297,N_9681,N_9800);
nand U10298 (N_10298,N_9559,N_9665);
nand U10299 (N_10299,N_9791,N_9401);
or U10300 (N_10300,N_9719,N_9481);
xor U10301 (N_10301,N_9407,N_9630);
xnor U10302 (N_10302,N_9864,N_9540);
and U10303 (N_10303,N_9855,N_9550);
and U10304 (N_10304,N_9507,N_9875);
or U10305 (N_10305,N_9965,N_9810);
or U10306 (N_10306,N_9724,N_9555);
nand U10307 (N_10307,N_9949,N_9534);
nand U10308 (N_10308,N_9624,N_9938);
or U10309 (N_10309,N_9774,N_9644);
or U10310 (N_10310,N_9487,N_9792);
nor U10311 (N_10311,N_9591,N_9808);
nor U10312 (N_10312,N_9839,N_9630);
or U10313 (N_10313,N_9376,N_9526);
xor U10314 (N_10314,N_9810,N_9770);
xnor U10315 (N_10315,N_9566,N_9967);
nor U10316 (N_10316,N_9634,N_9640);
and U10317 (N_10317,N_9926,N_9680);
or U10318 (N_10318,N_9961,N_9456);
nand U10319 (N_10319,N_9950,N_9378);
and U10320 (N_10320,N_9713,N_9931);
nand U10321 (N_10321,N_9868,N_9904);
and U10322 (N_10322,N_9690,N_9499);
xor U10323 (N_10323,N_9420,N_9966);
nor U10324 (N_10324,N_9831,N_9921);
and U10325 (N_10325,N_9628,N_9836);
nor U10326 (N_10326,N_9410,N_9446);
nand U10327 (N_10327,N_9749,N_9517);
or U10328 (N_10328,N_9931,N_9646);
or U10329 (N_10329,N_9904,N_9392);
nand U10330 (N_10330,N_9798,N_9566);
and U10331 (N_10331,N_9468,N_9477);
nand U10332 (N_10332,N_9778,N_9787);
and U10333 (N_10333,N_9481,N_9464);
xnor U10334 (N_10334,N_9927,N_9647);
and U10335 (N_10335,N_9980,N_9747);
nand U10336 (N_10336,N_9557,N_9696);
nand U10337 (N_10337,N_9588,N_9624);
nand U10338 (N_10338,N_9662,N_9476);
and U10339 (N_10339,N_9619,N_9997);
or U10340 (N_10340,N_9864,N_9432);
and U10341 (N_10341,N_9583,N_9968);
or U10342 (N_10342,N_9572,N_9408);
xnor U10343 (N_10343,N_9936,N_9987);
or U10344 (N_10344,N_9473,N_9574);
or U10345 (N_10345,N_9980,N_9575);
and U10346 (N_10346,N_9603,N_9411);
or U10347 (N_10347,N_9580,N_9442);
nor U10348 (N_10348,N_9768,N_9609);
xor U10349 (N_10349,N_9692,N_9656);
nor U10350 (N_10350,N_9537,N_9857);
or U10351 (N_10351,N_9674,N_9921);
or U10352 (N_10352,N_9609,N_9475);
xor U10353 (N_10353,N_9774,N_9676);
nor U10354 (N_10354,N_9866,N_9989);
nor U10355 (N_10355,N_9980,N_9399);
and U10356 (N_10356,N_9920,N_9538);
and U10357 (N_10357,N_9408,N_9653);
and U10358 (N_10358,N_9584,N_9460);
nand U10359 (N_10359,N_9918,N_9980);
or U10360 (N_10360,N_9629,N_9845);
xnor U10361 (N_10361,N_9390,N_9932);
xnor U10362 (N_10362,N_9460,N_9917);
xor U10363 (N_10363,N_9781,N_9615);
and U10364 (N_10364,N_9453,N_9978);
nor U10365 (N_10365,N_9640,N_9974);
xnor U10366 (N_10366,N_9623,N_9758);
nor U10367 (N_10367,N_9438,N_9459);
nand U10368 (N_10368,N_9848,N_9406);
nor U10369 (N_10369,N_9788,N_9795);
nor U10370 (N_10370,N_9648,N_9473);
nand U10371 (N_10371,N_9697,N_9877);
nand U10372 (N_10372,N_9714,N_9463);
nor U10373 (N_10373,N_9469,N_9808);
nor U10374 (N_10374,N_9999,N_9657);
or U10375 (N_10375,N_9438,N_9622);
or U10376 (N_10376,N_9909,N_9581);
or U10377 (N_10377,N_9605,N_9535);
or U10378 (N_10378,N_9951,N_9523);
xor U10379 (N_10379,N_9960,N_9745);
or U10380 (N_10380,N_9809,N_9940);
xnor U10381 (N_10381,N_9758,N_9518);
and U10382 (N_10382,N_9924,N_9759);
nand U10383 (N_10383,N_9706,N_9469);
xor U10384 (N_10384,N_9502,N_9946);
and U10385 (N_10385,N_9766,N_9897);
nand U10386 (N_10386,N_9843,N_9420);
or U10387 (N_10387,N_9738,N_9631);
or U10388 (N_10388,N_9864,N_9420);
or U10389 (N_10389,N_9810,N_9589);
xnor U10390 (N_10390,N_9852,N_9517);
xnor U10391 (N_10391,N_9797,N_9492);
and U10392 (N_10392,N_9765,N_9646);
xor U10393 (N_10393,N_9937,N_9383);
nor U10394 (N_10394,N_9385,N_9923);
nor U10395 (N_10395,N_9432,N_9715);
or U10396 (N_10396,N_9654,N_9607);
or U10397 (N_10397,N_9498,N_9991);
and U10398 (N_10398,N_9389,N_9804);
and U10399 (N_10399,N_9839,N_9810);
nand U10400 (N_10400,N_9867,N_9658);
nand U10401 (N_10401,N_9985,N_9830);
xor U10402 (N_10402,N_9397,N_9498);
or U10403 (N_10403,N_9527,N_9632);
nand U10404 (N_10404,N_9797,N_9622);
xnor U10405 (N_10405,N_9663,N_9736);
nand U10406 (N_10406,N_9803,N_9491);
or U10407 (N_10407,N_9525,N_9975);
or U10408 (N_10408,N_9759,N_9951);
nand U10409 (N_10409,N_9548,N_9723);
nor U10410 (N_10410,N_9401,N_9982);
xor U10411 (N_10411,N_9624,N_9947);
nand U10412 (N_10412,N_9988,N_9788);
nand U10413 (N_10413,N_9599,N_9621);
nor U10414 (N_10414,N_9624,N_9714);
nor U10415 (N_10415,N_9715,N_9843);
xor U10416 (N_10416,N_9801,N_9866);
nand U10417 (N_10417,N_9901,N_9649);
nand U10418 (N_10418,N_9637,N_9958);
nand U10419 (N_10419,N_9480,N_9582);
or U10420 (N_10420,N_9732,N_9629);
and U10421 (N_10421,N_9470,N_9581);
xor U10422 (N_10422,N_9919,N_9929);
nor U10423 (N_10423,N_9642,N_9679);
or U10424 (N_10424,N_9803,N_9854);
nand U10425 (N_10425,N_9983,N_9571);
and U10426 (N_10426,N_9647,N_9715);
xnor U10427 (N_10427,N_9752,N_9781);
and U10428 (N_10428,N_9939,N_9513);
xnor U10429 (N_10429,N_9958,N_9706);
or U10430 (N_10430,N_9632,N_9525);
or U10431 (N_10431,N_9751,N_9661);
xor U10432 (N_10432,N_9916,N_9582);
or U10433 (N_10433,N_9483,N_9986);
nor U10434 (N_10434,N_9671,N_9825);
nand U10435 (N_10435,N_9662,N_9470);
nor U10436 (N_10436,N_9811,N_9896);
xor U10437 (N_10437,N_9582,N_9566);
or U10438 (N_10438,N_9556,N_9613);
nand U10439 (N_10439,N_9997,N_9827);
or U10440 (N_10440,N_9510,N_9533);
nand U10441 (N_10441,N_9909,N_9759);
nor U10442 (N_10442,N_9616,N_9610);
or U10443 (N_10443,N_9916,N_9615);
xnor U10444 (N_10444,N_9882,N_9713);
nor U10445 (N_10445,N_9707,N_9474);
and U10446 (N_10446,N_9659,N_9532);
and U10447 (N_10447,N_9563,N_9790);
nand U10448 (N_10448,N_9980,N_9540);
and U10449 (N_10449,N_9382,N_9759);
or U10450 (N_10450,N_9799,N_9563);
or U10451 (N_10451,N_9831,N_9591);
or U10452 (N_10452,N_9815,N_9656);
xor U10453 (N_10453,N_9989,N_9593);
and U10454 (N_10454,N_9515,N_9915);
and U10455 (N_10455,N_9640,N_9509);
and U10456 (N_10456,N_9644,N_9498);
nor U10457 (N_10457,N_9934,N_9941);
and U10458 (N_10458,N_9705,N_9856);
nand U10459 (N_10459,N_9718,N_9475);
or U10460 (N_10460,N_9789,N_9982);
xnor U10461 (N_10461,N_9424,N_9635);
and U10462 (N_10462,N_9832,N_9874);
and U10463 (N_10463,N_9978,N_9645);
nand U10464 (N_10464,N_9545,N_9591);
or U10465 (N_10465,N_9419,N_9744);
or U10466 (N_10466,N_9428,N_9719);
nor U10467 (N_10467,N_9719,N_9798);
nand U10468 (N_10468,N_9873,N_9528);
xor U10469 (N_10469,N_9657,N_9497);
xor U10470 (N_10470,N_9450,N_9790);
nand U10471 (N_10471,N_9437,N_9702);
nor U10472 (N_10472,N_9500,N_9904);
or U10473 (N_10473,N_9904,N_9713);
nor U10474 (N_10474,N_9381,N_9574);
nor U10475 (N_10475,N_9912,N_9920);
and U10476 (N_10476,N_9807,N_9738);
nand U10477 (N_10477,N_9459,N_9885);
xnor U10478 (N_10478,N_9751,N_9892);
or U10479 (N_10479,N_9942,N_9730);
or U10480 (N_10480,N_9948,N_9429);
nor U10481 (N_10481,N_9634,N_9841);
xnor U10482 (N_10482,N_9387,N_9471);
nor U10483 (N_10483,N_9493,N_9411);
and U10484 (N_10484,N_9531,N_9505);
and U10485 (N_10485,N_9978,N_9440);
or U10486 (N_10486,N_9706,N_9624);
nor U10487 (N_10487,N_9891,N_9490);
nand U10488 (N_10488,N_9787,N_9471);
or U10489 (N_10489,N_9762,N_9463);
xor U10490 (N_10490,N_9960,N_9378);
and U10491 (N_10491,N_9580,N_9759);
and U10492 (N_10492,N_9957,N_9742);
or U10493 (N_10493,N_9634,N_9495);
nand U10494 (N_10494,N_9629,N_9804);
nand U10495 (N_10495,N_9437,N_9893);
nand U10496 (N_10496,N_9939,N_9483);
and U10497 (N_10497,N_9468,N_9584);
and U10498 (N_10498,N_9401,N_9445);
xnor U10499 (N_10499,N_9964,N_9589);
and U10500 (N_10500,N_9968,N_9465);
xnor U10501 (N_10501,N_9773,N_9406);
nor U10502 (N_10502,N_9482,N_9449);
and U10503 (N_10503,N_9645,N_9743);
nand U10504 (N_10504,N_9891,N_9486);
or U10505 (N_10505,N_9551,N_9813);
xnor U10506 (N_10506,N_9452,N_9597);
xor U10507 (N_10507,N_9527,N_9683);
xnor U10508 (N_10508,N_9559,N_9946);
xnor U10509 (N_10509,N_9902,N_9614);
nor U10510 (N_10510,N_9729,N_9698);
or U10511 (N_10511,N_9778,N_9380);
nor U10512 (N_10512,N_9417,N_9853);
xnor U10513 (N_10513,N_9674,N_9535);
xnor U10514 (N_10514,N_9787,N_9701);
and U10515 (N_10515,N_9448,N_9945);
and U10516 (N_10516,N_9686,N_9908);
or U10517 (N_10517,N_9602,N_9672);
and U10518 (N_10518,N_9559,N_9961);
or U10519 (N_10519,N_9976,N_9769);
or U10520 (N_10520,N_9696,N_9855);
xor U10521 (N_10521,N_9833,N_9682);
and U10522 (N_10522,N_9789,N_9823);
nand U10523 (N_10523,N_9829,N_9471);
xnor U10524 (N_10524,N_9582,N_9629);
nand U10525 (N_10525,N_9977,N_9998);
or U10526 (N_10526,N_9455,N_9906);
or U10527 (N_10527,N_9882,N_9618);
and U10528 (N_10528,N_9716,N_9409);
nand U10529 (N_10529,N_9809,N_9464);
nand U10530 (N_10530,N_9702,N_9529);
nand U10531 (N_10531,N_9589,N_9460);
nand U10532 (N_10532,N_9701,N_9411);
nand U10533 (N_10533,N_9496,N_9538);
xnor U10534 (N_10534,N_9550,N_9849);
xor U10535 (N_10535,N_9590,N_9516);
nand U10536 (N_10536,N_9475,N_9497);
xor U10537 (N_10537,N_9762,N_9418);
or U10538 (N_10538,N_9801,N_9777);
nand U10539 (N_10539,N_9422,N_9650);
or U10540 (N_10540,N_9787,N_9676);
or U10541 (N_10541,N_9604,N_9522);
nand U10542 (N_10542,N_9424,N_9409);
nor U10543 (N_10543,N_9930,N_9567);
and U10544 (N_10544,N_9950,N_9954);
and U10545 (N_10545,N_9786,N_9914);
xnor U10546 (N_10546,N_9732,N_9460);
xnor U10547 (N_10547,N_9500,N_9477);
nor U10548 (N_10548,N_9470,N_9412);
nor U10549 (N_10549,N_9692,N_9438);
nand U10550 (N_10550,N_9783,N_9710);
xnor U10551 (N_10551,N_9515,N_9741);
and U10552 (N_10552,N_9978,N_9505);
and U10553 (N_10553,N_9993,N_9563);
nand U10554 (N_10554,N_9705,N_9669);
xor U10555 (N_10555,N_9865,N_9601);
xor U10556 (N_10556,N_9669,N_9752);
nor U10557 (N_10557,N_9523,N_9615);
nor U10558 (N_10558,N_9977,N_9595);
or U10559 (N_10559,N_9884,N_9523);
nor U10560 (N_10560,N_9530,N_9597);
nand U10561 (N_10561,N_9917,N_9467);
xor U10562 (N_10562,N_9673,N_9477);
and U10563 (N_10563,N_9998,N_9424);
or U10564 (N_10564,N_9928,N_9631);
and U10565 (N_10565,N_9858,N_9603);
nand U10566 (N_10566,N_9802,N_9631);
or U10567 (N_10567,N_9447,N_9465);
nand U10568 (N_10568,N_9425,N_9641);
and U10569 (N_10569,N_9650,N_9670);
or U10570 (N_10570,N_9725,N_9782);
nand U10571 (N_10571,N_9473,N_9449);
nand U10572 (N_10572,N_9987,N_9780);
nor U10573 (N_10573,N_9874,N_9446);
nand U10574 (N_10574,N_9679,N_9770);
nor U10575 (N_10575,N_9539,N_9841);
nor U10576 (N_10576,N_9588,N_9809);
nand U10577 (N_10577,N_9496,N_9564);
xor U10578 (N_10578,N_9427,N_9705);
nand U10579 (N_10579,N_9935,N_9820);
nand U10580 (N_10580,N_9611,N_9559);
and U10581 (N_10581,N_9454,N_9678);
xor U10582 (N_10582,N_9506,N_9762);
nor U10583 (N_10583,N_9787,N_9983);
or U10584 (N_10584,N_9790,N_9713);
xnor U10585 (N_10585,N_9423,N_9862);
and U10586 (N_10586,N_9593,N_9821);
nor U10587 (N_10587,N_9561,N_9626);
or U10588 (N_10588,N_9696,N_9414);
xor U10589 (N_10589,N_9599,N_9465);
nor U10590 (N_10590,N_9769,N_9756);
or U10591 (N_10591,N_9510,N_9517);
nand U10592 (N_10592,N_9750,N_9913);
nand U10593 (N_10593,N_9782,N_9944);
or U10594 (N_10594,N_9921,N_9687);
nand U10595 (N_10595,N_9803,N_9951);
nor U10596 (N_10596,N_9915,N_9954);
nor U10597 (N_10597,N_9770,N_9417);
xnor U10598 (N_10598,N_9487,N_9645);
nand U10599 (N_10599,N_9917,N_9604);
and U10600 (N_10600,N_9439,N_9802);
nor U10601 (N_10601,N_9654,N_9891);
and U10602 (N_10602,N_9468,N_9993);
nand U10603 (N_10603,N_9959,N_9803);
nor U10604 (N_10604,N_9393,N_9782);
and U10605 (N_10605,N_9760,N_9803);
and U10606 (N_10606,N_9638,N_9424);
nand U10607 (N_10607,N_9565,N_9923);
or U10608 (N_10608,N_9542,N_9571);
nand U10609 (N_10609,N_9603,N_9802);
and U10610 (N_10610,N_9375,N_9556);
and U10611 (N_10611,N_9649,N_9965);
or U10612 (N_10612,N_9618,N_9904);
and U10613 (N_10613,N_9417,N_9533);
or U10614 (N_10614,N_9729,N_9541);
xnor U10615 (N_10615,N_9473,N_9959);
or U10616 (N_10616,N_9611,N_9709);
and U10617 (N_10617,N_9535,N_9581);
nor U10618 (N_10618,N_9468,N_9471);
or U10619 (N_10619,N_9745,N_9412);
nor U10620 (N_10620,N_9389,N_9851);
or U10621 (N_10621,N_9617,N_9479);
xor U10622 (N_10622,N_9955,N_9531);
or U10623 (N_10623,N_9596,N_9974);
xnor U10624 (N_10624,N_9435,N_9921);
nand U10625 (N_10625,N_10138,N_10359);
or U10626 (N_10626,N_10458,N_10485);
or U10627 (N_10627,N_10291,N_10373);
or U10628 (N_10628,N_10294,N_10025);
or U10629 (N_10629,N_10205,N_10327);
xnor U10630 (N_10630,N_10398,N_10571);
xor U10631 (N_10631,N_10277,N_10570);
and U10632 (N_10632,N_10079,N_10427);
or U10633 (N_10633,N_10507,N_10584);
nand U10634 (N_10634,N_10070,N_10578);
nor U10635 (N_10635,N_10032,N_10200);
and U10636 (N_10636,N_10337,N_10292);
or U10637 (N_10637,N_10434,N_10262);
nand U10638 (N_10638,N_10375,N_10467);
nand U10639 (N_10639,N_10394,N_10051);
nand U10640 (N_10640,N_10322,N_10590);
nand U10641 (N_10641,N_10141,N_10214);
and U10642 (N_10642,N_10031,N_10055);
and U10643 (N_10643,N_10133,N_10300);
nor U10644 (N_10644,N_10401,N_10391);
or U10645 (N_10645,N_10023,N_10093);
xnor U10646 (N_10646,N_10203,N_10370);
or U10647 (N_10647,N_10576,N_10046);
or U10648 (N_10648,N_10224,N_10270);
xor U10649 (N_10649,N_10037,N_10465);
and U10650 (N_10650,N_10082,N_10364);
xnor U10651 (N_10651,N_10157,N_10003);
nand U10652 (N_10652,N_10017,N_10117);
xnor U10653 (N_10653,N_10350,N_10173);
or U10654 (N_10654,N_10556,N_10144);
or U10655 (N_10655,N_10230,N_10110);
nand U10656 (N_10656,N_10457,N_10537);
nor U10657 (N_10657,N_10426,N_10605);
and U10658 (N_10658,N_10143,N_10620);
xor U10659 (N_10659,N_10125,N_10420);
nand U10660 (N_10660,N_10152,N_10387);
nor U10661 (N_10661,N_10199,N_10343);
nor U10662 (N_10662,N_10513,N_10215);
nor U10663 (N_10663,N_10073,N_10269);
nor U10664 (N_10664,N_10140,N_10357);
or U10665 (N_10665,N_10555,N_10272);
nand U10666 (N_10666,N_10597,N_10328);
or U10667 (N_10667,N_10425,N_10611);
or U10668 (N_10668,N_10080,N_10516);
nor U10669 (N_10669,N_10487,N_10542);
nand U10670 (N_10670,N_10573,N_10153);
nor U10671 (N_10671,N_10372,N_10482);
nand U10672 (N_10672,N_10547,N_10107);
or U10673 (N_10673,N_10175,N_10455);
xor U10674 (N_10674,N_10559,N_10558);
nand U10675 (N_10675,N_10560,N_10124);
nor U10676 (N_10676,N_10332,N_10338);
and U10677 (N_10677,N_10126,N_10081);
nor U10678 (N_10678,N_10354,N_10243);
and U10679 (N_10679,N_10491,N_10497);
nor U10680 (N_10680,N_10266,N_10281);
nor U10681 (N_10681,N_10399,N_10174);
xor U10682 (N_10682,N_10410,N_10260);
and U10683 (N_10683,N_10128,N_10461);
and U10684 (N_10684,N_10402,N_10217);
xor U10685 (N_10685,N_10036,N_10116);
or U10686 (N_10686,N_10526,N_10182);
nor U10687 (N_10687,N_10106,N_10474);
nor U10688 (N_10688,N_10599,N_10251);
xnor U10689 (N_10689,N_10591,N_10592);
nand U10690 (N_10690,N_10309,N_10259);
xor U10691 (N_10691,N_10183,N_10232);
nand U10692 (N_10692,N_10581,N_10532);
and U10693 (N_10693,N_10165,N_10024);
nand U10694 (N_10694,N_10225,N_10067);
or U10695 (N_10695,N_10122,N_10569);
nor U10696 (N_10696,N_10529,N_10496);
nand U10697 (N_10697,N_10154,N_10076);
nor U10698 (N_10698,N_10594,N_10190);
nor U10699 (N_10699,N_10065,N_10119);
xor U10700 (N_10700,N_10286,N_10178);
or U10701 (N_10701,N_10317,N_10180);
and U10702 (N_10702,N_10085,N_10275);
or U10703 (N_10703,N_10271,N_10472);
nand U10704 (N_10704,N_10530,N_10256);
xor U10705 (N_10705,N_10392,N_10276);
or U10706 (N_10706,N_10349,N_10617);
nand U10707 (N_10707,N_10540,N_10267);
nor U10708 (N_10708,N_10136,N_10495);
xnor U10709 (N_10709,N_10222,N_10445);
and U10710 (N_10710,N_10562,N_10273);
xnor U10711 (N_10711,N_10283,N_10139);
and U10712 (N_10712,N_10602,N_10088);
and U10713 (N_10713,N_10170,N_10518);
and U10714 (N_10714,N_10381,N_10447);
nand U10715 (N_10715,N_10614,N_10324);
nor U10716 (N_10716,N_10600,N_10428);
xnor U10717 (N_10717,N_10179,N_10563);
or U10718 (N_10718,N_10358,N_10297);
nor U10719 (N_10719,N_10534,N_10305);
or U10720 (N_10720,N_10195,N_10552);
or U10721 (N_10721,N_10198,N_10027);
nand U10722 (N_10722,N_10432,N_10288);
and U10723 (N_10723,N_10004,N_10263);
or U10724 (N_10724,N_10580,N_10466);
nor U10725 (N_10725,N_10228,N_10546);
or U10726 (N_10726,N_10607,N_10418);
or U10727 (N_10727,N_10363,N_10528);
and U10728 (N_10728,N_10500,N_10090);
nor U10729 (N_10729,N_10523,N_10084);
and U10730 (N_10730,N_10388,N_10164);
nor U10731 (N_10731,N_10265,N_10212);
and U10732 (N_10732,N_10429,N_10369);
and U10733 (N_10733,N_10544,N_10344);
xnor U10734 (N_10734,N_10331,N_10250);
xnor U10735 (N_10735,N_10621,N_10533);
nor U10736 (N_10736,N_10603,N_10156);
or U10737 (N_10737,N_10595,N_10459);
and U10738 (N_10738,N_10306,N_10210);
nor U10739 (N_10739,N_10374,N_10022);
or U10740 (N_10740,N_10083,N_10016);
or U10741 (N_10741,N_10382,N_10451);
xor U10742 (N_10742,N_10227,N_10531);
xor U10743 (N_10743,N_10041,N_10204);
nand U10744 (N_10744,N_10240,N_10226);
nor U10745 (N_10745,N_10345,N_10159);
nor U10746 (N_10746,N_10561,N_10196);
xnor U10747 (N_10747,N_10253,N_10390);
and U10748 (N_10748,N_10147,N_10335);
or U10749 (N_10749,N_10326,N_10623);
or U10750 (N_10750,N_10424,N_10453);
and U10751 (N_10751,N_10014,N_10419);
and U10752 (N_10752,N_10333,N_10450);
xnor U10753 (N_10753,N_10285,N_10356);
and U10754 (N_10754,N_10437,N_10013);
or U10755 (N_10755,N_10011,N_10411);
or U10756 (N_10756,N_10018,N_10066);
or U10757 (N_10757,N_10166,N_10063);
and U10758 (N_10758,N_10365,N_10568);
xnor U10759 (N_10759,N_10103,N_10231);
xor U10760 (N_10760,N_10545,N_10520);
nor U10761 (N_10761,N_10470,N_10118);
nand U10762 (N_10762,N_10587,N_10423);
nor U10763 (N_10763,N_10378,N_10446);
and U10764 (N_10764,N_10376,N_10311);
nand U10765 (N_10765,N_10135,N_10610);
xnor U10766 (N_10766,N_10064,N_10494);
nand U10767 (N_10767,N_10527,N_10351);
nand U10768 (N_10768,N_10238,N_10444);
and U10769 (N_10769,N_10206,N_10284);
xor U10770 (N_10770,N_10352,N_10396);
or U10771 (N_10771,N_10541,N_10188);
and U10772 (N_10772,N_10454,N_10233);
nand U10773 (N_10773,N_10463,N_10379);
and U10774 (N_10774,N_10384,N_10295);
xnor U10775 (N_10775,N_10342,N_10521);
xnor U10776 (N_10776,N_10241,N_10320);
and U10777 (N_10777,N_10104,N_10223);
nor U10778 (N_10778,N_10246,N_10236);
xor U10779 (N_10779,N_10244,N_10268);
nand U10780 (N_10780,N_10316,N_10549);
nand U10781 (N_10781,N_10468,N_10443);
nor U10782 (N_10782,N_10150,N_10339);
or U10783 (N_10783,N_10054,N_10371);
xor U10784 (N_10784,N_10535,N_10056);
and U10785 (N_10785,N_10475,N_10565);
nor U10786 (N_10786,N_10499,N_10087);
nor U10787 (N_10787,N_10334,N_10609);
xnor U10788 (N_10788,N_10367,N_10282);
xor U10789 (N_10789,N_10341,N_10476);
nor U10790 (N_10790,N_10010,N_10235);
nor U10791 (N_10791,N_10321,N_10069);
and U10792 (N_10792,N_10043,N_10261);
nand U10793 (N_10793,N_10435,N_10028);
and U10794 (N_10794,N_10194,N_10469);
nand U10795 (N_10795,N_10197,N_10131);
nor U10796 (N_10796,N_10220,N_10579);
xor U10797 (N_10797,N_10089,N_10492);
nand U10798 (N_10798,N_10422,N_10471);
or U10799 (N_10799,N_10501,N_10102);
xor U10800 (N_10800,N_10002,N_10040);
nor U10801 (N_10801,N_10514,N_10347);
nand U10802 (N_10802,N_10218,N_10008);
and U10803 (N_10803,N_10604,N_10078);
xnor U10804 (N_10804,N_10213,N_10506);
and U10805 (N_10805,N_10308,N_10524);
nand U10806 (N_10806,N_10310,N_10557);
xor U10807 (N_10807,N_10301,N_10211);
nor U10808 (N_10808,N_10409,N_10433);
or U10809 (N_10809,N_10421,N_10386);
xor U10810 (N_10810,N_10142,N_10624);
xor U10811 (N_10811,N_10302,N_10075);
nor U10812 (N_10812,N_10616,N_10299);
and U10813 (N_10813,N_10072,N_10038);
xnor U10814 (N_10814,N_10585,N_10613);
nand U10815 (N_10815,N_10313,N_10456);
or U10816 (N_10816,N_10101,N_10254);
or U10817 (N_10817,N_10171,N_10044);
or U10818 (N_10818,N_10510,N_10406);
and U10819 (N_10819,N_10130,N_10221);
and U10820 (N_10820,N_10318,N_10113);
xor U10821 (N_10821,N_10290,N_10293);
or U10822 (N_10822,N_10155,N_10033);
nand U10823 (N_10823,N_10412,N_10047);
and U10824 (N_10824,N_10052,N_10247);
and U10825 (N_10825,N_10505,N_10319);
xor U10826 (N_10826,N_10115,N_10296);
or U10827 (N_10827,N_10035,N_10449);
nor U10828 (N_10828,N_10111,N_10589);
or U10829 (N_10829,N_10020,N_10430);
and U10830 (N_10830,N_10053,N_10005);
xor U10831 (N_10831,N_10050,N_10519);
or U10832 (N_10832,N_10007,N_10478);
nor U10833 (N_10833,N_10586,N_10114);
xnor U10834 (N_10834,N_10006,N_10161);
xnor U10835 (N_10835,N_10512,N_10493);
nor U10836 (N_10836,N_10192,N_10504);
or U10837 (N_10837,N_10015,N_10353);
nand U10838 (N_10838,N_10436,N_10091);
nand U10839 (N_10839,N_10588,N_10312);
nor U10840 (N_10840,N_10538,N_10030);
xor U10841 (N_10841,N_10160,N_10149);
nor U10842 (N_10842,N_10042,N_10525);
xor U10843 (N_10843,N_10062,N_10258);
and U10844 (N_10844,N_10303,N_10314);
or U10845 (N_10845,N_10522,N_10566);
nor U10846 (N_10846,N_10034,N_10298);
nor U10847 (N_10847,N_10362,N_10105);
and U10848 (N_10848,N_10176,N_10029);
nand U10849 (N_10849,N_10554,N_10092);
xor U10850 (N_10850,N_10596,N_10257);
and U10851 (N_10851,N_10121,N_10123);
nand U10852 (N_10852,N_10209,N_10517);
or U10853 (N_10853,N_10202,N_10360);
nand U10854 (N_10854,N_10515,N_10440);
nand U10855 (N_10855,N_10278,N_10177);
or U10856 (N_10856,N_10201,N_10346);
nand U10857 (N_10857,N_10097,N_10086);
nor U10858 (N_10858,N_10404,N_10127);
nor U10859 (N_10859,N_10393,N_10577);
and U10860 (N_10860,N_10151,N_10593);
and U10861 (N_10861,N_10615,N_10408);
or U10862 (N_10862,N_10400,N_10001);
nand U10863 (N_10863,N_10168,N_10551);
and U10864 (N_10864,N_10601,N_10606);
and U10865 (N_10865,N_10255,N_10068);
nand U10866 (N_10866,N_10361,N_10488);
and U10867 (N_10867,N_10279,N_10383);
and U10868 (N_10868,N_10307,N_10059);
nand U10869 (N_10869,N_10330,N_10098);
or U10870 (N_10870,N_10368,N_10622);
or U10871 (N_10871,N_10389,N_10377);
nand U10872 (N_10872,N_10094,N_10608);
nand U10873 (N_10873,N_10489,N_10486);
xnor U10874 (N_10874,N_10567,N_10181);
nor U10875 (N_10875,N_10460,N_10574);
nand U10876 (N_10876,N_10187,N_10431);
nand U10877 (N_10877,N_10325,N_10413);
xnor U10878 (N_10878,N_10340,N_10509);
xnor U10879 (N_10879,N_10508,N_10239);
nor U10880 (N_10880,N_10264,N_10185);
and U10881 (N_10881,N_10163,N_10502);
nor U10882 (N_10882,N_10134,N_10619);
xor U10883 (N_10883,N_10287,N_10189);
xor U10884 (N_10884,N_10048,N_10323);
and U10885 (N_10885,N_10417,N_10148);
and U10886 (N_10886,N_10395,N_10120);
nand U10887 (N_10887,N_10462,N_10186);
or U10888 (N_10888,N_10039,N_10403);
nor U10889 (N_10889,N_10234,N_10405);
xnor U10890 (N_10890,N_10464,N_10045);
nand U10891 (N_10891,N_10473,N_10216);
or U10892 (N_10892,N_10503,N_10169);
xnor U10893 (N_10893,N_10100,N_10049);
nor U10894 (N_10894,N_10572,N_10193);
or U10895 (N_10895,N_10612,N_10061);
or U10896 (N_10896,N_10229,N_10553);
nand U10897 (N_10897,N_10057,N_10012);
nor U10898 (N_10898,N_10484,N_10074);
nand U10899 (N_10899,N_10490,N_10385);
nor U10900 (N_10900,N_10539,N_10129);
xor U10901 (N_10901,N_10146,N_10598);
xnor U10902 (N_10902,N_10355,N_10618);
xnor U10903 (N_10903,N_10536,N_10348);
xnor U10904 (N_10904,N_10479,N_10237);
or U10905 (N_10905,N_10366,N_10498);
or U10906 (N_10906,N_10582,N_10575);
nand U10907 (N_10907,N_10416,N_10252);
xnor U10908 (N_10908,N_10207,N_10137);
xnor U10909 (N_10909,N_10060,N_10274);
or U10910 (N_10910,N_10441,N_10280);
and U10911 (N_10911,N_10009,N_10058);
and U10912 (N_10912,N_10172,N_10249);
or U10913 (N_10913,N_10077,N_10096);
xor U10914 (N_10914,N_10315,N_10108);
xor U10915 (N_10915,N_10019,N_10336);
nand U10916 (N_10916,N_10191,N_10477);
nor U10917 (N_10917,N_10095,N_10112);
or U10918 (N_10918,N_10407,N_10242);
xnor U10919 (N_10919,N_10415,N_10304);
xor U10920 (N_10920,N_10158,N_10564);
xor U10921 (N_10921,N_10145,N_10109);
xor U10922 (N_10922,N_10162,N_10438);
xor U10923 (N_10923,N_10132,N_10219);
nor U10924 (N_10924,N_10380,N_10414);
xor U10925 (N_10925,N_10397,N_10439);
or U10926 (N_10926,N_10099,N_10511);
and U10927 (N_10927,N_10021,N_10480);
or U10928 (N_10928,N_10448,N_10184);
nor U10929 (N_10929,N_10026,N_10329);
xor U10930 (N_10930,N_10543,N_10442);
and U10931 (N_10931,N_10245,N_10071);
xnor U10932 (N_10932,N_10481,N_10167);
and U10933 (N_10933,N_10248,N_10483);
xor U10934 (N_10934,N_10289,N_10000);
nor U10935 (N_10935,N_10550,N_10208);
nor U10936 (N_10936,N_10583,N_10452);
xnor U10937 (N_10937,N_10548,N_10370);
xor U10938 (N_10938,N_10471,N_10032);
xor U10939 (N_10939,N_10594,N_10003);
nor U10940 (N_10940,N_10115,N_10095);
nor U10941 (N_10941,N_10411,N_10199);
or U10942 (N_10942,N_10505,N_10455);
xor U10943 (N_10943,N_10101,N_10438);
and U10944 (N_10944,N_10269,N_10194);
or U10945 (N_10945,N_10308,N_10154);
nor U10946 (N_10946,N_10048,N_10303);
or U10947 (N_10947,N_10334,N_10210);
or U10948 (N_10948,N_10611,N_10446);
and U10949 (N_10949,N_10176,N_10235);
or U10950 (N_10950,N_10249,N_10424);
xor U10951 (N_10951,N_10257,N_10448);
nor U10952 (N_10952,N_10235,N_10356);
xor U10953 (N_10953,N_10186,N_10396);
xnor U10954 (N_10954,N_10325,N_10361);
nand U10955 (N_10955,N_10347,N_10420);
xnor U10956 (N_10956,N_10433,N_10205);
or U10957 (N_10957,N_10452,N_10056);
xor U10958 (N_10958,N_10243,N_10413);
and U10959 (N_10959,N_10568,N_10093);
nor U10960 (N_10960,N_10374,N_10329);
and U10961 (N_10961,N_10620,N_10272);
xor U10962 (N_10962,N_10431,N_10496);
and U10963 (N_10963,N_10532,N_10539);
and U10964 (N_10964,N_10169,N_10584);
nand U10965 (N_10965,N_10624,N_10366);
nand U10966 (N_10966,N_10484,N_10506);
xor U10967 (N_10967,N_10551,N_10152);
xor U10968 (N_10968,N_10410,N_10549);
xor U10969 (N_10969,N_10220,N_10238);
nor U10970 (N_10970,N_10169,N_10332);
or U10971 (N_10971,N_10151,N_10580);
nor U10972 (N_10972,N_10475,N_10572);
or U10973 (N_10973,N_10019,N_10622);
or U10974 (N_10974,N_10442,N_10012);
nor U10975 (N_10975,N_10346,N_10273);
nand U10976 (N_10976,N_10454,N_10431);
xor U10977 (N_10977,N_10359,N_10518);
xnor U10978 (N_10978,N_10204,N_10462);
or U10979 (N_10979,N_10571,N_10093);
xor U10980 (N_10980,N_10312,N_10242);
nand U10981 (N_10981,N_10540,N_10494);
and U10982 (N_10982,N_10597,N_10054);
or U10983 (N_10983,N_10381,N_10489);
and U10984 (N_10984,N_10169,N_10571);
nand U10985 (N_10985,N_10589,N_10120);
nor U10986 (N_10986,N_10500,N_10474);
nand U10987 (N_10987,N_10401,N_10248);
and U10988 (N_10988,N_10518,N_10544);
nand U10989 (N_10989,N_10201,N_10046);
or U10990 (N_10990,N_10187,N_10454);
nor U10991 (N_10991,N_10558,N_10072);
xor U10992 (N_10992,N_10301,N_10453);
nor U10993 (N_10993,N_10096,N_10587);
nand U10994 (N_10994,N_10418,N_10438);
nand U10995 (N_10995,N_10001,N_10121);
xor U10996 (N_10996,N_10193,N_10469);
and U10997 (N_10997,N_10177,N_10285);
or U10998 (N_10998,N_10529,N_10084);
nor U10999 (N_10999,N_10033,N_10542);
and U11000 (N_11000,N_10277,N_10430);
or U11001 (N_11001,N_10424,N_10406);
or U11002 (N_11002,N_10171,N_10007);
or U11003 (N_11003,N_10556,N_10362);
xor U11004 (N_11004,N_10145,N_10593);
xnor U11005 (N_11005,N_10422,N_10415);
nor U11006 (N_11006,N_10123,N_10587);
xor U11007 (N_11007,N_10099,N_10541);
and U11008 (N_11008,N_10410,N_10452);
xnor U11009 (N_11009,N_10502,N_10291);
or U11010 (N_11010,N_10557,N_10555);
or U11011 (N_11011,N_10050,N_10575);
and U11012 (N_11012,N_10423,N_10237);
and U11013 (N_11013,N_10248,N_10085);
and U11014 (N_11014,N_10191,N_10575);
nor U11015 (N_11015,N_10348,N_10304);
nand U11016 (N_11016,N_10198,N_10320);
nor U11017 (N_11017,N_10503,N_10162);
or U11018 (N_11018,N_10232,N_10611);
nand U11019 (N_11019,N_10499,N_10067);
and U11020 (N_11020,N_10406,N_10053);
and U11021 (N_11021,N_10396,N_10624);
and U11022 (N_11022,N_10619,N_10582);
or U11023 (N_11023,N_10394,N_10244);
nor U11024 (N_11024,N_10201,N_10033);
nand U11025 (N_11025,N_10612,N_10040);
nand U11026 (N_11026,N_10339,N_10407);
nand U11027 (N_11027,N_10073,N_10230);
nand U11028 (N_11028,N_10344,N_10232);
or U11029 (N_11029,N_10577,N_10217);
xnor U11030 (N_11030,N_10457,N_10334);
nor U11031 (N_11031,N_10054,N_10220);
nor U11032 (N_11032,N_10052,N_10067);
nor U11033 (N_11033,N_10400,N_10551);
and U11034 (N_11034,N_10236,N_10135);
nand U11035 (N_11035,N_10347,N_10090);
or U11036 (N_11036,N_10149,N_10136);
xnor U11037 (N_11037,N_10422,N_10559);
nor U11038 (N_11038,N_10448,N_10375);
or U11039 (N_11039,N_10152,N_10248);
nand U11040 (N_11040,N_10037,N_10429);
nor U11041 (N_11041,N_10118,N_10104);
and U11042 (N_11042,N_10463,N_10109);
xor U11043 (N_11043,N_10237,N_10508);
xnor U11044 (N_11044,N_10506,N_10003);
or U11045 (N_11045,N_10056,N_10470);
nand U11046 (N_11046,N_10520,N_10445);
xnor U11047 (N_11047,N_10623,N_10019);
and U11048 (N_11048,N_10000,N_10126);
nor U11049 (N_11049,N_10500,N_10369);
and U11050 (N_11050,N_10208,N_10254);
nor U11051 (N_11051,N_10437,N_10271);
and U11052 (N_11052,N_10011,N_10550);
nand U11053 (N_11053,N_10009,N_10065);
nor U11054 (N_11054,N_10523,N_10043);
and U11055 (N_11055,N_10211,N_10571);
xnor U11056 (N_11056,N_10425,N_10017);
xor U11057 (N_11057,N_10238,N_10377);
and U11058 (N_11058,N_10345,N_10405);
nor U11059 (N_11059,N_10296,N_10125);
nand U11060 (N_11060,N_10071,N_10420);
or U11061 (N_11061,N_10491,N_10334);
and U11062 (N_11062,N_10414,N_10396);
and U11063 (N_11063,N_10492,N_10114);
and U11064 (N_11064,N_10552,N_10144);
nand U11065 (N_11065,N_10376,N_10390);
xor U11066 (N_11066,N_10454,N_10181);
nand U11067 (N_11067,N_10358,N_10466);
or U11068 (N_11068,N_10527,N_10606);
xnor U11069 (N_11069,N_10614,N_10166);
and U11070 (N_11070,N_10544,N_10334);
or U11071 (N_11071,N_10399,N_10556);
and U11072 (N_11072,N_10234,N_10605);
nand U11073 (N_11073,N_10187,N_10170);
nand U11074 (N_11074,N_10582,N_10287);
xor U11075 (N_11075,N_10466,N_10341);
nor U11076 (N_11076,N_10076,N_10624);
or U11077 (N_11077,N_10374,N_10320);
nor U11078 (N_11078,N_10006,N_10280);
or U11079 (N_11079,N_10126,N_10216);
nand U11080 (N_11080,N_10033,N_10524);
or U11081 (N_11081,N_10138,N_10197);
and U11082 (N_11082,N_10270,N_10328);
xor U11083 (N_11083,N_10588,N_10035);
xor U11084 (N_11084,N_10168,N_10516);
and U11085 (N_11085,N_10146,N_10079);
xnor U11086 (N_11086,N_10397,N_10069);
and U11087 (N_11087,N_10290,N_10189);
nor U11088 (N_11088,N_10557,N_10440);
xnor U11089 (N_11089,N_10511,N_10086);
and U11090 (N_11090,N_10307,N_10455);
nand U11091 (N_11091,N_10475,N_10022);
and U11092 (N_11092,N_10084,N_10241);
nand U11093 (N_11093,N_10377,N_10597);
nor U11094 (N_11094,N_10337,N_10489);
or U11095 (N_11095,N_10318,N_10244);
nor U11096 (N_11096,N_10087,N_10127);
xnor U11097 (N_11097,N_10094,N_10071);
nor U11098 (N_11098,N_10515,N_10270);
xor U11099 (N_11099,N_10293,N_10286);
nor U11100 (N_11100,N_10248,N_10279);
or U11101 (N_11101,N_10381,N_10410);
and U11102 (N_11102,N_10380,N_10479);
or U11103 (N_11103,N_10193,N_10100);
or U11104 (N_11104,N_10001,N_10382);
nand U11105 (N_11105,N_10508,N_10413);
xor U11106 (N_11106,N_10583,N_10146);
or U11107 (N_11107,N_10017,N_10291);
xor U11108 (N_11108,N_10170,N_10563);
and U11109 (N_11109,N_10121,N_10300);
or U11110 (N_11110,N_10220,N_10021);
xor U11111 (N_11111,N_10124,N_10295);
nand U11112 (N_11112,N_10056,N_10050);
nor U11113 (N_11113,N_10302,N_10217);
xnor U11114 (N_11114,N_10065,N_10057);
nand U11115 (N_11115,N_10133,N_10473);
nand U11116 (N_11116,N_10523,N_10461);
nor U11117 (N_11117,N_10359,N_10390);
xnor U11118 (N_11118,N_10506,N_10459);
nor U11119 (N_11119,N_10182,N_10349);
nor U11120 (N_11120,N_10177,N_10575);
xnor U11121 (N_11121,N_10154,N_10578);
or U11122 (N_11122,N_10098,N_10239);
or U11123 (N_11123,N_10026,N_10085);
and U11124 (N_11124,N_10049,N_10333);
nand U11125 (N_11125,N_10128,N_10412);
or U11126 (N_11126,N_10357,N_10201);
nor U11127 (N_11127,N_10525,N_10030);
xnor U11128 (N_11128,N_10116,N_10379);
and U11129 (N_11129,N_10615,N_10393);
and U11130 (N_11130,N_10347,N_10012);
or U11131 (N_11131,N_10040,N_10482);
xnor U11132 (N_11132,N_10363,N_10150);
or U11133 (N_11133,N_10308,N_10406);
or U11134 (N_11134,N_10427,N_10321);
nand U11135 (N_11135,N_10396,N_10555);
xor U11136 (N_11136,N_10415,N_10309);
and U11137 (N_11137,N_10487,N_10396);
and U11138 (N_11138,N_10391,N_10113);
or U11139 (N_11139,N_10245,N_10268);
xnor U11140 (N_11140,N_10137,N_10267);
and U11141 (N_11141,N_10216,N_10109);
nor U11142 (N_11142,N_10120,N_10262);
and U11143 (N_11143,N_10029,N_10303);
and U11144 (N_11144,N_10393,N_10160);
nor U11145 (N_11145,N_10596,N_10359);
and U11146 (N_11146,N_10535,N_10217);
and U11147 (N_11147,N_10452,N_10352);
xor U11148 (N_11148,N_10038,N_10407);
or U11149 (N_11149,N_10447,N_10362);
nand U11150 (N_11150,N_10039,N_10356);
or U11151 (N_11151,N_10134,N_10550);
nand U11152 (N_11152,N_10423,N_10310);
nor U11153 (N_11153,N_10294,N_10590);
nor U11154 (N_11154,N_10496,N_10239);
or U11155 (N_11155,N_10570,N_10599);
nor U11156 (N_11156,N_10562,N_10618);
and U11157 (N_11157,N_10470,N_10402);
nand U11158 (N_11158,N_10093,N_10603);
nor U11159 (N_11159,N_10614,N_10237);
xor U11160 (N_11160,N_10209,N_10176);
or U11161 (N_11161,N_10562,N_10420);
nand U11162 (N_11162,N_10511,N_10327);
xnor U11163 (N_11163,N_10560,N_10080);
nor U11164 (N_11164,N_10047,N_10043);
or U11165 (N_11165,N_10479,N_10467);
xnor U11166 (N_11166,N_10462,N_10166);
xnor U11167 (N_11167,N_10435,N_10391);
and U11168 (N_11168,N_10308,N_10610);
nand U11169 (N_11169,N_10070,N_10288);
and U11170 (N_11170,N_10225,N_10098);
nor U11171 (N_11171,N_10327,N_10176);
nand U11172 (N_11172,N_10296,N_10384);
or U11173 (N_11173,N_10288,N_10623);
nor U11174 (N_11174,N_10381,N_10188);
nor U11175 (N_11175,N_10362,N_10000);
and U11176 (N_11176,N_10204,N_10247);
and U11177 (N_11177,N_10019,N_10349);
nand U11178 (N_11178,N_10472,N_10120);
nor U11179 (N_11179,N_10412,N_10605);
or U11180 (N_11180,N_10368,N_10491);
and U11181 (N_11181,N_10495,N_10410);
or U11182 (N_11182,N_10500,N_10493);
xnor U11183 (N_11183,N_10509,N_10226);
nand U11184 (N_11184,N_10227,N_10261);
or U11185 (N_11185,N_10332,N_10386);
or U11186 (N_11186,N_10142,N_10090);
nand U11187 (N_11187,N_10572,N_10621);
or U11188 (N_11188,N_10596,N_10351);
and U11189 (N_11189,N_10021,N_10022);
or U11190 (N_11190,N_10144,N_10255);
xor U11191 (N_11191,N_10556,N_10264);
nor U11192 (N_11192,N_10050,N_10104);
and U11193 (N_11193,N_10557,N_10485);
nor U11194 (N_11194,N_10427,N_10086);
and U11195 (N_11195,N_10150,N_10503);
and U11196 (N_11196,N_10070,N_10427);
or U11197 (N_11197,N_10464,N_10323);
xor U11198 (N_11198,N_10534,N_10321);
xor U11199 (N_11199,N_10060,N_10009);
or U11200 (N_11200,N_10353,N_10581);
and U11201 (N_11201,N_10184,N_10296);
nor U11202 (N_11202,N_10406,N_10242);
and U11203 (N_11203,N_10476,N_10288);
or U11204 (N_11204,N_10068,N_10257);
and U11205 (N_11205,N_10224,N_10283);
nand U11206 (N_11206,N_10283,N_10325);
or U11207 (N_11207,N_10441,N_10418);
and U11208 (N_11208,N_10589,N_10030);
nand U11209 (N_11209,N_10569,N_10399);
or U11210 (N_11210,N_10197,N_10067);
nor U11211 (N_11211,N_10203,N_10150);
or U11212 (N_11212,N_10360,N_10045);
nand U11213 (N_11213,N_10260,N_10104);
nand U11214 (N_11214,N_10013,N_10587);
nor U11215 (N_11215,N_10339,N_10233);
nand U11216 (N_11216,N_10042,N_10173);
nand U11217 (N_11217,N_10596,N_10210);
and U11218 (N_11218,N_10494,N_10032);
and U11219 (N_11219,N_10609,N_10061);
and U11220 (N_11220,N_10174,N_10356);
and U11221 (N_11221,N_10180,N_10576);
nand U11222 (N_11222,N_10183,N_10615);
nor U11223 (N_11223,N_10327,N_10015);
nor U11224 (N_11224,N_10296,N_10484);
and U11225 (N_11225,N_10046,N_10393);
or U11226 (N_11226,N_10231,N_10354);
or U11227 (N_11227,N_10384,N_10287);
and U11228 (N_11228,N_10012,N_10231);
nand U11229 (N_11229,N_10400,N_10487);
nor U11230 (N_11230,N_10479,N_10445);
nor U11231 (N_11231,N_10322,N_10031);
and U11232 (N_11232,N_10189,N_10178);
and U11233 (N_11233,N_10414,N_10021);
nor U11234 (N_11234,N_10139,N_10566);
nand U11235 (N_11235,N_10435,N_10229);
or U11236 (N_11236,N_10517,N_10096);
nand U11237 (N_11237,N_10299,N_10456);
nand U11238 (N_11238,N_10507,N_10135);
nor U11239 (N_11239,N_10398,N_10412);
nand U11240 (N_11240,N_10308,N_10321);
nand U11241 (N_11241,N_10488,N_10038);
nand U11242 (N_11242,N_10288,N_10117);
nand U11243 (N_11243,N_10131,N_10172);
or U11244 (N_11244,N_10325,N_10603);
and U11245 (N_11245,N_10123,N_10441);
nand U11246 (N_11246,N_10415,N_10575);
xnor U11247 (N_11247,N_10144,N_10214);
or U11248 (N_11248,N_10273,N_10149);
nand U11249 (N_11249,N_10295,N_10460);
or U11250 (N_11250,N_11188,N_10856);
xor U11251 (N_11251,N_10663,N_10922);
xnor U11252 (N_11252,N_10918,N_10980);
nor U11253 (N_11253,N_11025,N_10944);
or U11254 (N_11254,N_10822,N_11097);
nor U11255 (N_11255,N_10758,N_11099);
nand U11256 (N_11256,N_10643,N_11110);
nor U11257 (N_11257,N_10733,N_10642);
or U11258 (N_11258,N_11135,N_10798);
xnor U11259 (N_11259,N_10973,N_11202);
nand U11260 (N_11260,N_10915,N_11201);
nand U11261 (N_11261,N_10993,N_11065);
or U11262 (N_11262,N_10636,N_10847);
nand U11263 (N_11263,N_10755,N_10893);
nand U11264 (N_11264,N_10888,N_10930);
xnor U11265 (N_11265,N_11054,N_10675);
or U11266 (N_11266,N_10705,N_11217);
xnor U11267 (N_11267,N_10778,N_10972);
nor U11268 (N_11268,N_10690,N_10630);
and U11269 (N_11269,N_10999,N_11043);
nand U11270 (N_11270,N_11011,N_10725);
xor U11271 (N_11271,N_10830,N_11209);
nand U11272 (N_11272,N_11245,N_11024);
nand U11273 (N_11273,N_10985,N_10939);
and U11274 (N_11274,N_10669,N_10754);
xnor U11275 (N_11275,N_11145,N_10760);
nand U11276 (N_11276,N_11242,N_11170);
nor U11277 (N_11277,N_10729,N_10874);
or U11278 (N_11278,N_11225,N_11111);
xor U11279 (N_11279,N_11056,N_10748);
nor U11280 (N_11280,N_11138,N_10794);
xnor U11281 (N_11281,N_11048,N_11147);
or U11282 (N_11282,N_11093,N_10841);
and U11283 (N_11283,N_11162,N_10717);
or U11284 (N_11284,N_10708,N_11222);
nor U11285 (N_11285,N_10774,N_10911);
xor U11286 (N_11286,N_11243,N_11184);
nand U11287 (N_11287,N_11075,N_10765);
nand U11288 (N_11288,N_10635,N_10728);
or U11289 (N_11289,N_10923,N_10989);
and U11290 (N_11290,N_11030,N_11109);
nand U11291 (N_11291,N_10880,N_10685);
xnor U11292 (N_11292,N_11010,N_10773);
and U11293 (N_11293,N_10682,N_10892);
nor U11294 (N_11294,N_10793,N_10819);
or U11295 (N_11295,N_10843,N_11226);
nor U11296 (N_11296,N_10820,N_11079);
xnor U11297 (N_11297,N_11151,N_11122);
and U11298 (N_11298,N_11081,N_10965);
and U11299 (N_11299,N_11073,N_11244);
nand U11300 (N_11300,N_10872,N_10861);
nor U11301 (N_11301,N_11103,N_10704);
xor U11302 (N_11302,N_10987,N_11215);
nand U11303 (N_11303,N_10837,N_10964);
nand U11304 (N_11304,N_10886,N_11029);
and U11305 (N_11305,N_11080,N_10813);
and U11306 (N_11306,N_10916,N_10720);
or U11307 (N_11307,N_10898,N_11041);
nand U11308 (N_11308,N_10736,N_11022);
xnor U11309 (N_11309,N_11241,N_11091);
nand U11310 (N_11310,N_10796,N_10829);
nand U11311 (N_11311,N_11036,N_11074);
xor U11312 (N_11312,N_10637,N_10711);
nand U11313 (N_11313,N_10741,N_10900);
and U11314 (N_11314,N_11161,N_10994);
xnor U11315 (N_11315,N_10929,N_10633);
xnor U11316 (N_11316,N_10827,N_11013);
or U11317 (N_11317,N_11064,N_10681);
xnor U11318 (N_11318,N_10718,N_11142);
xnor U11319 (N_11319,N_10785,N_10657);
nor U11320 (N_11320,N_10730,N_10802);
xnor U11321 (N_11321,N_10775,N_10815);
xnor U11322 (N_11322,N_10885,N_11211);
and U11323 (N_11323,N_11114,N_10851);
nand U11324 (N_11324,N_11026,N_11078);
xnor U11325 (N_11325,N_11157,N_11045);
or U11326 (N_11326,N_11062,N_10701);
nand U11327 (N_11327,N_10875,N_11001);
and U11328 (N_11328,N_11132,N_10865);
and U11329 (N_11329,N_11082,N_10659);
nor U11330 (N_11330,N_10654,N_11148);
and U11331 (N_11331,N_10768,N_11218);
xnor U11332 (N_11332,N_10703,N_11120);
and U11333 (N_11333,N_11016,N_11169);
and U11334 (N_11334,N_10716,N_10629);
nor U11335 (N_11335,N_10848,N_11186);
nor U11336 (N_11336,N_10897,N_11171);
nand U11337 (N_11337,N_10766,N_11067);
and U11338 (N_11338,N_10828,N_10871);
and U11339 (N_11339,N_11233,N_10684);
or U11340 (N_11340,N_11200,N_11131);
xor U11341 (N_11341,N_10818,N_11140);
xor U11342 (N_11342,N_10974,N_11107);
and U11343 (N_11343,N_10791,N_10671);
nor U11344 (N_11344,N_11037,N_11046);
xnor U11345 (N_11345,N_10839,N_11006);
nand U11346 (N_11346,N_11027,N_10960);
nor U11347 (N_11347,N_11129,N_11072);
and U11348 (N_11348,N_10638,N_10783);
nand U11349 (N_11349,N_10978,N_10801);
and U11350 (N_11350,N_10662,N_11003);
nand U11351 (N_11351,N_11127,N_11015);
and U11352 (N_11352,N_11137,N_11070);
or U11353 (N_11353,N_10832,N_11071);
or U11354 (N_11354,N_10764,N_10655);
xor U11355 (N_11355,N_11168,N_10938);
or U11356 (N_11356,N_11197,N_11032);
and U11357 (N_11357,N_10749,N_10772);
nand U11358 (N_11358,N_11207,N_11042);
xor U11359 (N_11359,N_10756,N_10723);
nor U11360 (N_11360,N_11194,N_10855);
and U11361 (N_11361,N_10628,N_10850);
or U11362 (N_11362,N_10858,N_11237);
and U11363 (N_11363,N_10714,N_11094);
nand U11364 (N_11364,N_11180,N_11153);
xnor U11365 (N_11365,N_10650,N_10644);
nor U11366 (N_11366,N_11149,N_10984);
nor U11367 (N_11367,N_11087,N_10761);
and U11368 (N_11368,N_11182,N_10645);
or U11369 (N_11369,N_10735,N_11066);
and U11370 (N_11370,N_11058,N_10873);
nand U11371 (N_11371,N_11177,N_11141);
and U11372 (N_11372,N_10626,N_10879);
and U11373 (N_11373,N_11038,N_10975);
xor U11374 (N_11374,N_10894,N_10920);
and U11375 (N_11375,N_11192,N_11158);
nand U11376 (N_11376,N_11223,N_11101);
nand U11377 (N_11377,N_10835,N_10710);
nand U11378 (N_11378,N_11133,N_10899);
nand U11379 (N_11379,N_11235,N_10912);
nor U11380 (N_11380,N_10821,N_11152);
nand U11381 (N_11381,N_10670,N_11166);
xnor U11382 (N_11382,N_11176,N_10936);
nor U11383 (N_11383,N_11203,N_10838);
or U11384 (N_11384,N_10666,N_10658);
or U11385 (N_11385,N_10906,N_11144);
nand U11386 (N_11386,N_10932,N_10763);
nand U11387 (N_11387,N_11155,N_10870);
xnor U11388 (N_11388,N_10933,N_10876);
or U11389 (N_11389,N_10997,N_11118);
nor U11390 (N_11390,N_10660,N_10868);
xor U11391 (N_11391,N_10686,N_10940);
nor U11392 (N_11392,N_11221,N_11165);
or U11393 (N_11393,N_11249,N_10988);
nand U11394 (N_11394,N_10625,N_11076);
and U11395 (N_11395,N_10726,N_11047);
and U11396 (N_11396,N_10895,N_10823);
nand U11397 (N_11397,N_11102,N_10786);
and U11398 (N_11398,N_11181,N_11017);
nand U11399 (N_11399,N_11130,N_10904);
xnor U11400 (N_11400,N_10910,N_10928);
and U11401 (N_11401,N_10889,N_11100);
nor U11402 (N_11402,N_10652,N_10805);
xor U11403 (N_11403,N_10840,N_11159);
nor U11404 (N_11404,N_11219,N_11061);
and U11405 (N_11405,N_10712,N_10992);
nor U11406 (N_11406,N_10687,N_11035);
and U11407 (N_11407,N_10734,N_10653);
and U11408 (N_11408,N_10702,N_11113);
xnor U11409 (N_11409,N_11123,N_10713);
and U11410 (N_11410,N_10862,N_11204);
or U11411 (N_11411,N_11183,N_10715);
xnor U11412 (N_11412,N_10807,N_10700);
nand U11413 (N_11413,N_10676,N_10824);
xor U11414 (N_11414,N_10942,N_11005);
nor U11415 (N_11415,N_10903,N_11049);
nor U11416 (N_11416,N_11063,N_10753);
nand U11417 (N_11417,N_10864,N_11224);
xnor U11418 (N_11418,N_10639,N_10699);
xor U11419 (N_11419,N_10665,N_10640);
nor U11420 (N_11420,N_10995,N_11086);
or U11421 (N_11421,N_10863,N_11214);
and U11422 (N_11422,N_10921,N_11057);
nor U11423 (N_11423,N_11034,N_10648);
nor U11424 (N_11424,N_10935,N_10831);
nor U11425 (N_11425,N_10731,N_10694);
or U11426 (N_11426,N_10747,N_10806);
xnor U11427 (N_11427,N_10692,N_11179);
and U11428 (N_11428,N_10762,N_11033);
and U11429 (N_11429,N_11228,N_10803);
nand U11430 (N_11430,N_10634,N_11238);
nor U11431 (N_11431,N_10746,N_10991);
and U11432 (N_11432,N_10673,N_10890);
or U11433 (N_11433,N_10649,N_11106);
or U11434 (N_11434,N_10963,N_10695);
xor U11435 (N_11435,N_11227,N_11189);
nor U11436 (N_11436,N_10981,N_11172);
nand U11437 (N_11437,N_11187,N_10808);
nand U11438 (N_11438,N_10790,N_10924);
nor U11439 (N_11439,N_10891,N_10743);
xor U11440 (N_11440,N_10852,N_10941);
and U11441 (N_11441,N_11231,N_11083);
and U11442 (N_11442,N_10950,N_11096);
xor U11443 (N_11443,N_10954,N_11089);
and U11444 (N_11444,N_10709,N_10949);
xor U11445 (N_11445,N_11002,N_10919);
xor U11446 (N_11446,N_11044,N_10943);
and U11447 (N_11447,N_10719,N_11178);
and U11448 (N_11448,N_11248,N_11028);
xnor U11449 (N_11449,N_11234,N_11098);
or U11450 (N_11450,N_10784,N_11164);
and U11451 (N_11451,N_10826,N_11175);
and U11452 (N_11452,N_10842,N_11007);
nor U11453 (N_11453,N_11090,N_10816);
xnor U11454 (N_11454,N_11206,N_11050);
and U11455 (N_11455,N_11167,N_11150);
or U11456 (N_11456,N_11156,N_10752);
nand U11457 (N_11457,N_10983,N_11134);
nand U11458 (N_11458,N_10846,N_10744);
nand U11459 (N_11459,N_10905,N_10721);
nor U11460 (N_11460,N_11163,N_10647);
or U11461 (N_11461,N_10811,N_11216);
xor U11462 (N_11462,N_11051,N_10792);
nor U11463 (N_11463,N_10966,N_11205);
and U11464 (N_11464,N_10641,N_10958);
xnor U11465 (N_11465,N_11108,N_10740);
xnor U11466 (N_11466,N_11240,N_10800);
and U11467 (N_11467,N_10896,N_10745);
and U11468 (N_11468,N_10779,N_10854);
and U11469 (N_11469,N_10750,N_11069);
nor U11470 (N_11470,N_10934,N_11023);
xor U11471 (N_11471,N_10878,N_10902);
and U11472 (N_11472,N_11146,N_10881);
xor U11473 (N_11473,N_10759,N_10913);
xnor U11474 (N_11474,N_10857,N_10672);
xnor U11475 (N_11475,N_11229,N_10698);
xnor U11476 (N_11476,N_10887,N_10697);
nor U11477 (N_11477,N_10707,N_10706);
xnor U11478 (N_11478,N_10967,N_10844);
or U11479 (N_11479,N_11236,N_10834);
or U11480 (N_11480,N_11191,N_10849);
and U11481 (N_11481,N_11239,N_11213);
nand U11482 (N_11482,N_10945,N_10656);
or U11483 (N_11483,N_11190,N_11210);
or U11484 (N_11484,N_10782,N_10948);
nor U11485 (N_11485,N_10925,N_10957);
nor U11486 (N_11486,N_10877,N_10696);
nand U11487 (N_11487,N_10998,N_11126);
xnor U11488 (N_11488,N_11019,N_10688);
or U11489 (N_11489,N_10727,N_11008);
or U11490 (N_11490,N_11125,N_10795);
nor U11491 (N_11491,N_10979,N_11128);
or U11492 (N_11492,N_10969,N_11020);
and U11493 (N_11493,N_10677,N_10959);
and U11494 (N_11494,N_10787,N_10953);
and U11495 (N_11495,N_11230,N_10901);
or U11496 (N_11496,N_11198,N_11139);
or U11497 (N_11497,N_11018,N_10836);
nor U11498 (N_11498,N_10908,N_10971);
or U11499 (N_11499,N_11117,N_11000);
xor U11500 (N_11500,N_10869,N_11092);
nand U11501 (N_11501,N_10661,N_10693);
and U11502 (N_11502,N_10738,N_11232);
or U11503 (N_11503,N_11185,N_10951);
and U11504 (N_11504,N_10691,N_10799);
xnor U11505 (N_11505,N_10739,N_10679);
and U11506 (N_11506,N_10757,N_10884);
nor U11507 (N_11507,N_10627,N_10825);
nand U11508 (N_11508,N_10977,N_11124);
nand U11509 (N_11509,N_11039,N_11220);
nand U11510 (N_11510,N_10777,N_10814);
xor U11511 (N_11511,N_10742,N_11055);
and U11512 (N_11512,N_10917,N_10770);
or U11513 (N_11513,N_11012,N_10859);
xor U11514 (N_11514,N_10781,N_10809);
or U11515 (N_11515,N_11009,N_11077);
nand U11516 (N_11516,N_10937,N_11014);
nand U11517 (N_11517,N_10962,N_11119);
xnor U11518 (N_11518,N_11095,N_10631);
nand U11519 (N_11519,N_10689,N_10646);
nor U11520 (N_11520,N_10683,N_11068);
nor U11521 (N_11521,N_10678,N_10664);
nand U11522 (N_11522,N_10952,N_11121);
xnor U11523 (N_11523,N_10946,N_11246);
xor U11524 (N_11524,N_11085,N_11115);
and U11525 (N_11525,N_11193,N_10955);
nand U11526 (N_11526,N_10812,N_11173);
nor U11527 (N_11527,N_11021,N_10996);
nand U11528 (N_11528,N_10927,N_11212);
nand U11529 (N_11529,N_11136,N_10833);
nor U11530 (N_11530,N_10724,N_10776);
and U11531 (N_11531,N_10845,N_10926);
nor U11532 (N_11532,N_10722,N_10732);
nand U11533 (N_11533,N_10982,N_10797);
nor U11534 (N_11534,N_11004,N_10986);
nand U11535 (N_11535,N_11116,N_11059);
nand U11536 (N_11536,N_11105,N_10668);
or U11537 (N_11537,N_10632,N_11053);
or U11538 (N_11538,N_10853,N_10769);
nor U11539 (N_11539,N_11195,N_10947);
nor U11540 (N_11540,N_11143,N_10767);
or U11541 (N_11541,N_10804,N_10914);
nand U11542 (N_11542,N_10970,N_11174);
nand U11543 (N_11543,N_11031,N_10990);
nor U11544 (N_11544,N_10817,N_11199);
nand U11545 (N_11545,N_10651,N_11160);
nor U11546 (N_11546,N_10976,N_11247);
and U11547 (N_11547,N_10961,N_11112);
nor U11548 (N_11548,N_10907,N_10882);
or U11549 (N_11549,N_10788,N_10931);
nand U11550 (N_11550,N_10674,N_10789);
and U11551 (N_11551,N_10771,N_10968);
or U11552 (N_11552,N_10867,N_10667);
or U11553 (N_11553,N_11196,N_10866);
nor U11554 (N_11554,N_11154,N_11208);
and U11555 (N_11555,N_10680,N_11088);
and U11556 (N_11556,N_10751,N_11084);
nor U11557 (N_11557,N_10860,N_10956);
nor U11558 (N_11558,N_10883,N_11040);
nand U11559 (N_11559,N_10909,N_11052);
and U11560 (N_11560,N_11104,N_10780);
xnor U11561 (N_11561,N_10810,N_10737);
and U11562 (N_11562,N_11060,N_10889);
xnor U11563 (N_11563,N_10755,N_10933);
xnor U11564 (N_11564,N_10997,N_10639);
xor U11565 (N_11565,N_10939,N_10987);
nor U11566 (N_11566,N_10812,N_10854);
and U11567 (N_11567,N_10906,N_10805);
and U11568 (N_11568,N_11101,N_10871);
xnor U11569 (N_11569,N_11233,N_10836);
and U11570 (N_11570,N_10636,N_10813);
nand U11571 (N_11571,N_11103,N_10963);
and U11572 (N_11572,N_10699,N_11009);
nor U11573 (N_11573,N_11191,N_10986);
or U11574 (N_11574,N_10716,N_11109);
or U11575 (N_11575,N_10674,N_10983);
nand U11576 (N_11576,N_10955,N_11035);
or U11577 (N_11577,N_11182,N_10726);
nand U11578 (N_11578,N_10936,N_11024);
or U11579 (N_11579,N_11126,N_11121);
and U11580 (N_11580,N_10631,N_10890);
nand U11581 (N_11581,N_11200,N_10716);
nand U11582 (N_11582,N_10651,N_11146);
and U11583 (N_11583,N_11190,N_10695);
or U11584 (N_11584,N_10882,N_11042);
xnor U11585 (N_11585,N_11110,N_10670);
or U11586 (N_11586,N_11111,N_10711);
and U11587 (N_11587,N_11135,N_10981);
or U11588 (N_11588,N_10916,N_11243);
nand U11589 (N_11589,N_11220,N_10763);
nand U11590 (N_11590,N_10699,N_10691);
xor U11591 (N_11591,N_11003,N_11218);
nor U11592 (N_11592,N_11125,N_10750);
xnor U11593 (N_11593,N_10940,N_11042);
nor U11594 (N_11594,N_10878,N_10656);
and U11595 (N_11595,N_10693,N_11193);
and U11596 (N_11596,N_11158,N_11173);
xnor U11597 (N_11597,N_11237,N_10823);
xnor U11598 (N_11598,N_10694,N_11107);
nand U11599 (N_11599,N_10820,N_11225);
nand U11600 (N_11600,N_10686,N_10830);
and U11601 (N_11601,N_10842,N_11121);
or U11602 (N_11602,N_11027,N_10738);
nand U11603 (N_11603,N_11106,N_10830);
and U11604 (N_11604,N_11193,N_10998);
xor U11605 (N_11605,N_10848,N_11168);
nor U11606 (N_11606,N_11065,N_11141);
or U11607 (N_11607,N_11056,N_10979);
nor U11608 (N_11608,N_11049,N_11140);
nand U11609 (N_11609,N_11001,N_10628);
or U11610 (N_11610,N_10658,N_10678);
xnor U11611 (N_11611,N_10694,N_11134);
nand U11612 (N_11612,N_10739,N_10847);
and U11613 (N_11613,N_10747,N_11160);
or U11614 (N_11614,N_10763,N_11063);
nor U11615 (N_11615,N_11043,N_10679);
xor U11616 (N_11616,N_11217,N_10998);
nand U11617 (N_11617,N_10922,N_10873);
nor U11618 (N_11618,N_11236,N_10638);
nor U11619 (N_11619,N_11043,N_11045);
or U11620 (N_11620,N_10806,N_10649);
and U11621 (N_11621,N_10876,N_11180);
and U11622 (N_11622,N_11031,N_11042);
or U11623 (N_11623,N_10829,N_10785);
nor U11624 (N_11624,N_11084,N_10946);
nor U11625 (N_11625,N_10633,N_10693);
nand U11626 (N_11626,N_10855,N_10644);
nand U11627 (N_11627,N_10934,N_10690);
nor U11628 (N_11628,N_11191,N_11131);
and U11629 (N_11629,N_11079,N_11052);
and U11630 (N_11630,N_11014,N_10982);
xor U11631 (N_11631,N_10885,N_10659);
nand U11632 (N_11632,N_10817,N_11104);
and U11633 (N_11633,N_11203,N_10656);
or U11634 (N_11634,N_10744,N_11204);
nand U11635 (N_11635,N_10723,N_11149);
and U11636 (N_11636,N_11214,N_10648);
nor U11637 (N_11637,N_10716,N_10684);
nand U11638 (N_11638,N_10774,N_11237);
nand U11639 (N_11639,N_10637,N_10885);
or U11640 (N_11640,N_11247,N_10854);
and U11641 (N_11641,N_10985,N_10924);
or U11642 (N_11642,N_10925,N_11074);
nand U11643 (N_11643,N_10720,N_11106);
nand U11644 (N_11644,N_11068,N_10801);
or U11645 (N_11645,N_10973,N_10770);
xor U11646 (N_11646,N_10932,N_11015);
nand U11647 (N_11647,N_10743,N_10745);
and U11648 (N_11648,N_11095,N_11004);
xor U11649 (N_11649,N_10669,N_11133);
or U11650 (N_11650,N_11054,N_11196);
or U11651 (N_11651,N_11038,N_11169);
or U11652 (N_11652,N_10681,N_11028);
and U11653 (N_11653,N_10672,N_11153);
nor U11654 (N_11654,N_11182,N_10662);
and U11655 (N_11655,N_11172,N_11036);
xor U11656 (N_11656,N_10885,N_11049);
nor U11657 (N_11657,N_10984,N_10800);
xnor U11658 (N_11658,N_11044,N_10880);
xor U11659 (N_11659,N_10919,N_10941);
or U11660 (N_11660,N_10843,N_10773);
nor U11661 (N_11661,N_10924,N_10975);
or U11662 (N_11662,N_10709,N_11185);
xor U11663 (N_11663,N_10859,N_10811);
nand U11664 (N_11664,N_10749,N_10968);
or U11665 (N_11665,N_10647,N_10674);
xnor U11666 (N_11666,N_10936,N_10827);
nor U11667 (N_11667,N_11151,N_10886);
nor U11668 (N_11668,N_11047,N_10962);
xnor U11669 (N_11669,N_10723,N_10630);
or U11670 (N_11670,N_10983,N_11225);
xnor U11671 (N_11671,N_10903,N_11122);
and U11672 (N_11672,N_11041,N_10862);
or U11673 (N_11673,N_10986,N_10712);
xor U11674 (N_11674,N_10640,N_10777);
nor U11675 (N_11675,N_11110,N_11175);
nor U11676 (N_11676,N_11219,N_11205);
or U11677 (N_11677,N_10972,N_11060);
xnor U11678 (N_11678,N_10939,N_11159);
and U11679 (N_11679,N_11065,N_10974);
xnor U11680 (N_11680,N_11102,N_10938);
nor U11681 (N_11681,N_10845,N_11050);
and U11682 (N_11682,N_10924,N_11207);
and U11683 (N_11683,N_10759,N_10867);
nor U11684 (N_11684,N_10744,N_11175);
and U11685 (N_11685,N_10706,N_10838);
xnor U11686 (N_11686,N_10675,N_10969);
nand U11687 (N_11687,N_10860,N_11192);
nand U11688 (N_11688,N_11046,N_10887);
nand U11689 (N_11689,N_10721,N_11163);
xnor U11690 (N_11690,N_10849,N_10894);
nor U11691 (N_11691,N_11191,N_11217);
or U11692 (N_11692,N_10732,N_11247);
nor U11693 (N_11693,N_11237,N_11163);
nand U11694 (N_11694,N_11125,N_11002);
nor U11695 (N_11695,N_10875,N_11123);
or U11696 (N_11696,N_10985,N_10846);
xnor U11697 (N_11697,N_10916,N_10805);
nand U11698 (N_11698,N_10650,N_10764);
or U11699 (N_11699,N_10915,N_10647);
or U11700 (N_11700,N_10686,N_11156);
or U11701 (N_11701,N_10940,N_10738);
nor U11702 (N_11702,N_11061,N_10655);
and U11703 (N_11703,N_10979,N_10637);
xor U11704 (N_11704,N_11031,N_10745);
and U11705 (N_11705,N_11102,N_11200);
nand U11706 (N_11706,N_11140,N_11035);
or U11707 (N_11707,N_11036,N_10902);
and U11708 (N_11708,N_10979,N_10664);
or U11709 (N_11709,N_11222,N_11059);
nor U11710 (N_11710,N_11201,N_11192);
or U11711 (N_11711,N_10788,N_10669);
nor U11712 (N_11712,N_11064,N_10923);
nor U11713 (N_11713,N_10962,N_11165);
nor U11714 (N_11714,N_10637,N_11081);
and U11715 (N_11715,N_11190,N_11003);
nand U11716 (N_11716,N_10806,N_11109);
xor U11717 (N_11717,N_10994,N_11221);
and U11718 (N_11718,N_11062,N_10713);
and U11719 (N_11719,N_10811,N_11217);
nand U11720 (N_11720,N_10802,N_10833);
and U11721 (N_11721,N_11075,N_10647);
and U11722 (N_11722,N_11115,N_10998);
or U11723 (N_11723,N_10903,N_10967);
nand U11724 (N_11724,N_10933,N_10968);
nand U11725 (N_11725,N_11208,N_11076);
xnor U11726 (N_11726,N_10803,N_10839);
nand U11727 (N_11727,N_10914,N_10668);
or U11728 (N_11728,N_10644,N_11152);
xnor U11729 (N_11729,N_10951,N_10743);
nand U11730 (N_11730,N_10948,N_11122);
or U11731 (N_11731,N_10689,N_10921);
or U11732 (N_11732,N_10812,N_10953);
and U11733 (N_11733,N_10925,N_10963);
or U11734 (N_11734,N_11104,N_10924);
or U11735 (N_11735,N_10916,N_10692);
or U11736 (N_11736,N_11143,N_10759);
xor U11737 (N_11737,N_11053,N_10962);
nor U11738 (N_11738,N_10904,N_10787);
nor U11739 (N_11739,N_10908,N_10898);
nor U11740 (N_11740,N_11157,N_11069);
and U11741 (N_11741,N_10725,N_11031);
nand U11742 (N_11742,N_10838,N_10829);
nor U11743 (N_11743,N_10935,N_10644);
nand U11744 (N_11744,N_11197,N_11200);
or U11745 (N_11745,N_11192,N_11096);
nand U11746 (N_11746,N_10961,N_10843);
or U11747 (N_11747,N_10715,N_10989);
xor U11748 (N_11748,N_10984,N_11216);
nand U11749 (N_11749,N_10804,N_11045);
or U11750 (N_11750,N_11235,N_11076);
xnor U11751 (N_11751,N_10883,N_11191);
xor U11752 (N_11752,N_10632,N_11242);
nor U11753 (N_11753,N_10663,N_10852);
and U11754 (N_11754,N_10662,N_10944);
nand U11755 (N_11755,N_11214,N_10745);
xnor U11756 (N_11756,N_11039,N_11082);
and U11757 (N_11757,N_10759,N_11185);
or U11758 (N_11758,N_11036,N_11024);
nand U11759 (N_11759,N_10905,N_11008);
and U11760 (N_11760,N_10996,N_10973);
xor U11761 (N_11761,N_10995,N_10647);
nor U11762 (N_11762,N_10939,N_10806);
nand U11763 (N_11763,N_10654,N_10673);
nor U11764 (N_11764,N_10636,N_10726);
nor U11765 (N_11765,N_10969,N_11241);
or U11766 (N_11766,N_11193,N_10891);
nor U11767 (N_11767,N_10952,N_10946);
nor U11768 (N_11768,N_11217,N_10903);
and U11769 (N_11769,N_11109,N_11147);
nor U11770 (N_11770,N_10892,N_10819);
or U11771 (N_11771,N_10849,N_10825);
and U11772 (N_11772,N_11078,N_11062);
nor U11773 (N_11773,N_11114,N_10691);
and U11774 (N_11774,N_11176,N_10806);
nand U11775 (N_11775,N_10718,N_10667);
and U11776 (N_11776,N_11241,N_11236);
xnor U11777 (N_11777,N_10863,N_11200);
xnor U11778 (N_11778,N_10673,N_11077);
xor U11779 (N_11779,N_10923,N_10759);
nor U11780 (N_11780,N_10844,N_10654);
nand U11781 (N_11781,N_10698,N_11144);
and U11782 (N_11782,N_11181,N_10976);
or U11783 (N_11783,N_10947,N_10998);
or U11784 (N_11784,N_11068,N_10888);
or U11785 (N_11785,N_10880,N_11200);
and U11786 (N_11786,N_10781,N_11052);
and U11787 (N_11787,N_11016,N_11101);
xor U11788 (N_11788,N_11040,N_10648);
nor U11789 (N_11789,N_10695,N_11100);
xor U11790 (N_11790,N_11189,N_11174);
xnor U11791 (N_11791,N_10740,N_11097);
and U11792 (N_11792,N_11123,N_10677);
xor U11793 (N_11793,N_10681,N_11212);
and U11794 (N_11794,N_10983,N_10919);
nor U11795 (N_11795,N_10841,N_10702);
xor U11796 (N_11796,N_10768,N_11071);
or U11797 (N_11797,N_11003,N_11159);
or U11798 (N_11798,N_10826,N_11217);
nor U11799 (N_11799,N_10684,N_10947);
nor U11800 (N_11800,N_11033,N_10651);
xnor U11801 (N_11801,N_10935,N_10873);
nor U11802 (N_11802,N_10656,N_11007);
and U11803 (N_11803,N_10795,N_10934);
and U11804 (N_11804,N_11034,N_10870);
and U11805 (N_11805,N_10767,N_10817);
xnor U11806 (N_11806,N_10710,N_10636);
nor U11807 (N_11807,N_10880,N_10722);
nand U11808 (N_11808,N_10956,N_10787);
or U11809 (N_11809,N_11039,N_11068);
nor U11810 (N_11810,N_10980,N_10763);
nor U11811 (N_11811,N_10999,N_10975);
or U11812 (N_11812,N_10795,N_10723);
and U11813 (N_11813,N_10726,N_10818);
nor U11814 (N_11814,N_11236,N_10670);
nor U11815 (N_11815,N_10631,N_10950);
and U11816 (N_11816,N_10813,N_10958);
and U11817 (N_11817,N_10831,N_11118);
nand U11818 (N_11818,N_10899,N_10974);
or U11819 (N_11819,N_10691,N_10982);
nor U11820 (N_11820,N_10685,N_11048);
nor U11821 (N_11821,N_10849,N_10800);
nor U11822 (N_11822,N_10632,N_11016);
or U11823 (N_11823,N_11158,N_10725);
and U11824 (N_11824,N_11187,N_10764);
nor U11825 (N_11825,N_11064,N_11226);
nand U11826 (N_11826,N_10899,N_10756);
or U11827 (N_11827,N_11103,N_11153);
or U11828 (N_11828,N_10925,N_10938);
nand U11829 (N_11829,N_11235,N_11092);
nand U11830 (N_11830,N_10801,N_10652);
or U11831 (N_11831,N_10647,N_10862);
nor U11832 (N_11832,N_11117,N_10765);
nor U11833 (N_11833,N_11226,N_10837);
nand U11834 (N_11834,N_11034,N_10709);
and U11835 (N_11835,N_11068,N_10700);
and U11836 (N_11836,N_10941,N_11075);
xor U11837 (N_11837,N_11037,N_10838);
or U11838 (N_11838,N_11212,N_10656);
or U11839 (N_11839,N_11197,N_10666);
nor U11840 (N_11840,N_11186,N_11108);
or U11841 (N_11841,N_10627,N_11132);
nor U11842 (N_11842,N_10816,N_11139);
nor U11843 (N_11843,N_10722,N_10657);
xor U11844 (N_11844,N_10679,N_11153);
or U11845 (N_11845,N_11022,N_11157);
nand U11846 (N_11846,N_11126,N_11123);
nor U11847 (N_11847,N_10880,N_11051);
nor U11848 (N_11848,N_11210,N_11079);
xor U11849 (N_11849,N_10981,N_10892);
xor U11850 (N_11850,N_10662,N_10630);
and U11851 (N_11851,N_11080,N_10658);
nand U11852 (N_11852,N_11157,N_11096);
nor U11853 (N_11853,N_11117,N_11149);
xnor U11854 (N_11854,N_10988,N_11081);
or U11855 (N_11855,N_10824,N_10745);
nor U11856 (N_11856,N_10834,N_11079);
nand U11857 (N_11857,N_11190,N_10931);
nand U11858 (N_11858,N_10645,N_11220);
nor U11859 (N_11859,N_11060,N_11030);
nand U11860 (N_11860,N_10892,N_11127);
nand U11861 (N_11861,N_10862,N_10651);
or U11862 (N_11862,N_10815,N_11012);
nor U11863 (N_11863,N_10803,N_10933);
nor U11864 (N_11864,N_10639,N_10664);
or U11865 (N_11865,N_10919,N_11117);
nor U11866 (N_11866,N_10841,N_11136);
or U11867 (N_11867,N_11021,N_10947);
or U11868 (N_11868,N_11167,N_10704);
nand U11869 (N_11869,N_11154,N_10748);
xor U11870 (N_11870,N_11099,N_10743);
nand U11871 (N_11871,N_11247,N_10968);
nand U11872 (N_11872,N_10775,N_11006);
nor U11873 (N_11873,N_11036,N_10890);
nand U11874 (N_11874,N_10708,N_11117);
or U11875 (N_11875,N_11593,N_11541);
nand U11876 (N_11876,N_11835,N_11274);
nor U11877 (N_11877,N_11337,N_11414);
xnor U11878 (N_11878,N_11436,N_11317);
or U11879 (N_11879,N_11527,N_11851);
nor U11880 (N_11880,N_11759,N_11347);
nand U11881 (N_11881,N_11309,N_11356);
nand U11882 (N_11882,N_11656,N_11754);
xor U11883 (N_11883,N_11498,N_11558);
nand U11884 (N_11884,N_11269,N_11318);
xnor U11885 (N_11885,N_11836,N_11769);
nand U11886 (N_11886,N_11789,N_11502);
xor U11887 (N_11887,N_11720,N_11506);
nor U11888 (N_11888,N_11731,N_11590);
or U11889 (N_11889,N_11391,N_11440);
xor U11890 (N_11890,N_11516,N_11804);
or U11891 (N_11891,N_11536,N_11788);
nand U11892 (N_11892,N_11409,N_11618);
nand U11893 (N_11893,N_11297,N_11487);
nand U11894 (N_11894,N_11844,N_11796);
nand U11895 (N_11895,N_11744,N_11296);
nor U11896 (N_11896,N_11629,N_11730);
xor U11897 (N_11897,N_11524,N_11698);
and U11898 (N_11898,N_11304,N_11323);
nand U11899 (N_11899,N_11480,N_11494);
xor U11900 (N_11900,N_11329,N_11684);
xor U11901 (N_11901,N_11483,N_11375);
or U11902 (N_11902,N_11282,N_11529);
nand U11903 (N_11903,N_11530,N_11484);
nand U11904 (N_11904,N_11660,N_11363);
nand U11905 (N_11905,N_11532,N_11547);
and U11906 (N_11906,N_11841,N_11373);
and U11907 (N_11907,N_11777,N_11735);
nor U11908 (N_11908,N_11517,N_11652);
nor U11909 (N_11909,N_11685,N_11848);
xnor U11910 (N_11910,N_11458,N_11668);
nor U11911 (N_11911,N_11772,N_11340);
nor U11912 (N_11912,N_11383,N_11467);
and U11913 (N_11913,N_11559,N_11411);
xor U11914 (N_11914,N_11461,N_11543);
and U11915 (N_11915,N_11605,N_11650);
xor U11916 (N_11916,N_11473,N_11679);
and U11917 (N_11917,N_11299,N_11768);
or U11918 (N_11918,N_11315,N_11589);
nand U11919 (N_11919,N_11291,N_11349);
or U11920 (N_11920,N_11840,N_11654);
nor U11921 (N_11921,N_11594,N_11621);
nor U11922 (N_11922,N_11466,N_11533);
and U11923 (N_11923,N_11424,N_11397);
xnor U11924 (N_11924,N_11393,N_11403);
or U11925 (N_11925,N_11686,N_11272);
nor U11926 (N_11926,N_11724,N_11265);
nor U11927 (N_11927,N_11402,N_11722);
nor U11928 (N_11928,N_11812,N_11413);
nor U11929 (N_11929,N_11587,N_11710);
xor U11930 (N_11930,N_11763,N_11301);
and U11931 (N_11931,N_11806,N_11277);
xor U11932 (N_11932,N_11279,N_11616);
or U11933 (N_11933,N_11603,N_11354);
nand U11934 (N_11934,N_11770,N_11408);
nor U11935 (N_11935,N_11258,N_11577);
and U11936 (N_11936,N_11442,N_11697);
xnor U11937 (N_11937,N_11750,N_11764);
and U11938 (N_11938,N_11569,N_11737);
nor U11939 (N_11939,N_11694,N_11361);
or U11940 (N_11940,N_11701,N_11575);
nand U11941 (N_11941,N_11302,N_11747);
and U11942 (N_11942,N_11452,N_11479);
nand U11943 (N_11943,N_11713,N_11678);
or U11944 (N_11944,N_11465,N_11670);
and U11945 (N_11945,N_11776,N_11597);
nand U11946 (N_11946,N_11264,N_11644);
and U11947 (N_11947,N_11649,N_11734);
nand U11948 (N_11948,N_11716,N_11578);
nor U11949 (N_11949,N_11853,N_11427);
nand U11950 (N_11950,N_11374,N_11481);
and U11951 (N_11951,N_11420,N_11485);
or U11952 (N_11952,N_11858,N_11787);
nand U11953 (N_11953,N_11680,N_11625);
and U11954 (N_11954,N_11740,N_11672);
nor U11955 (N_11955,N_11478,N_11666);
xnor U11956 (N_11956,N_11310,N_11288);
and U11957 (N_11957,N_11511,N_11350);
and U11958 (N_11958,N_11434,N_11749);
xnor U11959 (N_11959,N_11389,N_11614);
and U11960 (N_11960,N_11663,N_11266);
nand U11961 (N_11961,N_11606,N_11544);
and U11962 (N_11962,N_11596,N_11570);
nand U11963 (N_11963,N_11433,N_11542);
nor U11964 (N_11964,N_11795,N_11676);
nor U11965 (N_11965,N_11286,N_11378);
or U11966 (N_11966,N_11718,N_11800);
xnor U11967 (N_11967,N_11564,N_11460);
nor U11968 (N_11968,N_11861,N_11627);
xor U11969 (N_11969,N_11583,N_11552);
xor U11970 (N_11970,N_11617,N_11774);
nand U11971 (N_11971,N_11445,N_11691);
or U11972 (N_11972,N_11430,N_11534);
and U11973 (N_11973,N_11550,N_11438);
or U11974 (N_11974,N_11364,N_11521);
and U11975 (N_11975,N_11406,N_11692);
nand U11976 (N_11976,N_11820,N_11312);
nor U11977 (N_11977,N_11798,N_11637);
nand U11978 (N_11978,N_11439,N_11762);
and U11979 (N_11979,N_11548,N_11448);
nand U11980 (N_11980,N_11803,N_11275);
nand U11981 (N_11981,N_11797,N_11689);
or U11982 (N_11982,N_11289,N_11818);
and U11983 (N_11983,N_11615,N_11845);
nor U11984 (N_11984,N_11872,N_11492);
nand U11985 (N_11985,N_11659,N_11281);
xnor U11986 (N_11986,N_11786,N_11566);
nor U11987 (N_11987,N_11690,N_11355);
or U11988 (N_11988,N_11251,N_11854);
nand U11989 (N_11989,N_11733,N_11714);
nor U11990 (N_11990,N_11280,N_11715);
or U11991 (N_11991,N_11599,N_11306);
and U11992 (N_11992,N_11647,N_11554);
and U11993 (N_11993,N_11802,N_11608);
and U11994 (N_11994,N_11539,N_11719);
and U11995 (N_11995,N_11741,N_11344);
xor U11996 (N_11996,N_11324,N_11600);
nand U11997 (N_11997,N_11334,N_11869);
or U11998 (N_11998,N_11295,N_11419);
nand U11999 (N_11999,N_11362,N_11790);
or U12000 (N_12000,N_11586,N_11783);
nand U12001 (N_12001,N_11610,N_11874);
xnor U12002 (N_12002,N_11751,N_11518);
nor U12003 (N_12003,N_11252,N_11842);
xnor U12004 (N_12004,N_11695,N_11346);
nor U12005 (N_12005,N_11681,N_11815);
nor U12006 (N_12006,N_11867,N_11462);
and U12007 (N_12007,N_11386,N_11773);
nand U12008 (N_12008,N_11784,N_11646);
or U12009 (N_12009,N_11450,N_11416);
or U12010 (N_12010,N_11817,N_11256);
or U12011 (N_12011,N_11604,N_11658);
nor U12012 (N_12012,N_11285,N_11400);
or U12013 (N_12013,N_11418,N_11551);
nand U12014 (N_12014,N_11838,N_11863);
nor U12015 (N_12015,N_11794,N_11417);
and U12016 (N_12016,N_11866,N_11602);
and U12017 (N_12017,N_11669,N_11619);
nand U12018 (N_12018,N_11855,N_11753);
and U12019 (N_12019,N_11331,N_11488);
nor U12020 (N_12020,N_11415,N_11468);
nor U12021 (N_12021,N_11368,N_11808);
and U12022 (N_12022,N_11307,N_11320);
xor U12023 (N_12023,N_11809,N_11702);
nand U12024 (N_12024,N_11476,N_11852);
nand U12025 (N_12025,N_11816,N_11860);
xnor U12026 (N_12026,N_11345,N_11497);
nand U12027 (N_12027,N_11847,N_11477);
xnor U12028 (N_12028,N_11352,N_11626);
nand U12029 (N_12029,N_11699,N_11765);
or U12030 (N_12030,N_11563,N_11636);
and U12031 (N_12031,N_11336,N_11292);
nor U12032 (N_12032,N_11531,N_11683);
nor U12033 (N_12033,N_11831,N_11696);
or U12034 (N_12034,N_11263,N_11755);
nand U12035 (N_12035,N_11523,N_11367);
nor U12036 (N_12036,N_11574,N_11642);
nand U12037 (N_12037,N_11513,N_11509);
nand U12038 (N_12038,N_11333,N_11833);
xnor U12039 (N_12039,N_11819,N_11585);
and U12040 (N_12040,N_11813,N_11454);
nor U12041 (N_12041,N_11451,N_11567);
nor U12042 (N_12042,N_11711,N_11839);
nand U12043 (N_12043,N_11412,N_11556);
or U12044 (N_12044,N_11426,N_11515);
or U12045 (N_12045,N_11598,N_11328);
xnor U12046 (N_12046,N_11388,N_11657);
and U12047 (N_12047,N_11671,N_11261);
nand U12048 (N_12048,N_11490,N_11782);
nand U12049 (N_12049,N_11736,N_11775);
and U12050 (N_12050,N_11834,N_11634);
or U12051 (N_12051,N_11827,N_11607);
nor U12052 (N_12052,N_11553,N_11661);
or U12053 (N_12053,N_11538,N_11377);
nor U12054 (N_12054,N_11298,N_11394);
or U12055 (N_12055,N_11864,N_11766);
nor U12056 (N_12056,N_11581,N_11365);
xnor U12057 (N_12057,N_11253,N_11767);
or U12058 (N_12058,N_11601,N_11528);
or U12059 (N_12059,N_11405,N_11793);
nor U12060 (N_12060,N_11837,N_11358);
or U12061 (N_12061,N_11821,N_11846);
or U12062 (N_12062,N_11540,N_11791);
nor U12063 (N_12063,N_11276,N_11360);
or U12064 (N_12064,N_11822,N_11771);
nand U12065 (N_12065,N_11464,N_11641);
nor U12066 (N_12066,N_11571,N_11469);
nand U12067 (N_12067,N_11395,N_11475);
and U12068 (N_12068,N_11392,N_11379);
nand U12069 (N_12069,N_11341,N_11327);
nand U12070 (N_12070,N_11510,N_11491);
nand U12071 (N_12071,N_11868,N_11700);
nand U12072 (N_12072,N_11756,N_11675);
nand U12073 (N_12073,N_11457,N_11259);
nor U12074 (N_12074,N_11313,N_11332);
nand U12075 (N_12075,N_11287,N_11828);
xnor U12076 (N_12076,N_11537,N_11682);
nand U12077 (N_12077,N_11584,N_11503);
nor U12078 (N_12078,N_11508,N_11568);
nand U12079 (N_12079,N_11351,N_11260);
nor U12080 (N_12080,N_11723,N_11343);
or U12081 (N_12081,N_11664,N_11645);
nand U12082 (N_12082,N_11823,N_11499);
and U12083 (N_12083,N_11739,N_11330);
and U12084 (N_12084,N_11612,N_11255);
nand U12085 (N_12085,N_11832,N_11278);
and U12086 (N_12086,N_11425,N_11482);
nor U12087 (N_12087,N_11294,N_11579);
nand U12088 (N_12088,N_11522,N_11717);
nor U12089 (N_12089,N_11549,N_11758);
and U12090 (N_12090,N_11453,N_11335);
nand U12091 (N_12091,N_11369,N_11339);
or U12092 (N_12092,N_11742,N_11807);
xnor U12093 (N_12093,N_11843,N_11385);
or U12094 (N_12094,N_11592,N_11325);
nor U12095 (N_12095,N_11792,N_11825);
and U12096 (N_12096,N_11293,N_11609);
and U12097 (N_12097,N_11372,N_11435);
nand U12098 (N_12098,N_11613,N_11257);
and U12099 (N_12099,N_11655,N_11428);
and U12100 (N_12100,N_11449,N_11801);
and U12101 (N_12101,N_11631,N_11582);
xor U12102 (N_12102,N_11849,N_11673);
xnor U12103 (N_12103,N_11624,N_11588);
and U12104 (N_12104,N_11546,N_11580);
or U12105 (N_12105,N_11651,N_11338);
and U12106 (N_12106,N_11489,N_11665);
xnor U12107 (N_12107,N_11779,N_11371);
and U12108 (N_12108,N_11305,N_11705);
nand U12109 (N_12109,N_11757,N_11396);
nand U12110 (N_12110,N_11496,N_11830);
nor U12111 (N_12111,N_11727,N_11519);
xor U12112 (N_12112,N_11726,N_11353);
nand U12113 (N_12113,N_11729,N_11611);
and U12114 (N_12114,N_11814,N_11507);
xnor U12115 (N_12115,N_11623,N_11545);
xnor U12116 (N_12116,N_11688,N_11643);
nand U12117 (N_12117,N_11423,N_11562);
and U12118 (N_12118,N_11778,N_11250);
or U12119 (N_12119,N_11525,N_11576);
and U12120 (N_12120,N_11662,N_11640);
xnor U12121 (N_12121,N_11850,N_11653);
nand U12122 (N_12122,N_11382,N_11270);
nand U12123 (N_12123,N_11455,N_11471);
and U12124 (N_12124,N_11314,N_11704);
xor U12125 (N_12125,N_11348,N_11622);
or U12126 (N_12126,N_11573,N_11459);
and U12127 (N_12127,N_11639,N_11780);
or U12128 (N_12128,N_11535,N_11474);
and U12129 (N_12129,N_11284,N_11514);
nor U12130 (N_12130,N_11752,N_11572);
and U12131 (N_12131,N_11446,N_11321);
and U12132 (N_12132,N_11667,N_11384);
xnor U12133 (N_12133,N_11303,N_11493);
and U12134 (N_12134,N_11504,N_11632);
nand U12135 (N_12135,N_11707,N_11381);
or U12136 (N_12136,N_11591,N_11512);
and U12137 (N_12137,N_11404,N_11745);
xor U12138 (N_12138,N_11677,N_11370);
or U12139 (N_12139,N_11501,N_11322);
nor U12140 (N_12140,N_11871,N_11709);
or U12141 (N_12141,N_11811,N_11859);
or U12142 (N_12142,N_11376,N_11273);
or U12143 (N_12143,N_11638,N_11805);
or U12144 (N_12144,N_11421,N_11380);
and U12145 (N_12145,N_11443,N_11633);
or U12146 (N_12146,N_11262,N_11500);
and U12147 (N_12147,N_11781,N_11635);
and U12148 (N_12148,N_11555,N_11271);
nand U12149 (N_12149,N_11743,N_11398);
nor U12150 (N_12150,N_11456,N_11268);
and U12151 (N_12151,N_11721,N_11620);
and U12152 (N_12152,N_11437,N_11873);
nand U12153 (N_12153,N_11432,N_11748);
and U12154 (N_12154,N_11390,N_11687);
and U12155 (N_12155,N_11799,N_11422);
or U12156 (N_12156,N_11495,N_11746);
nand U12157 (N_12157,N_11674,N_11387);
nand U12158 (N_12158,N_11824,N_11520);
or U12159 (N_12159,N_11444,N_11254);
xor U12160 (N_12160,N_11441,N_11319);
xor U12161 (N_12161,N_11357,N_11708);
nor U12162 (N_12162,N_11732,N_11447);
nand U12163 (N_12163,N_11267,N_11486);
and U12164 (N_12164,N_11470,N_11401);
and U12165 (N_12165,N_11862,N_11316);
and U12166 (N_12166,N_11300,N_11725);
or U12167 (N_12167,N_11761,N_11630);
and U12168 (N_12168,N_11505,N_11785);
nor U12169 (N_12169,N_11410,N_11628);
nand U12170 (N_12170,N_11565,N_11829);
nor U12171 (N_12171,N_11311,N_11366);
nor U12172 (N_12172,N_11290,N_11308);
xor U12173 (N_12173,N_11359,N_11407);
or U12174 (N_12174,N_11557,N_11856);
or U12175 (N_12175,N_11826,N_11560);
and U12176 (N_12176,N_11648,N_11399);
nand U12177 (N_12177,N_11712,N_11429);
or U12178 (N_12178,N_11728,N_11595);
nand U12179 (N_12179,N_11431,N_11561);
nand U12180 (N_12180,N_11760,N_11857);
xor U12181 (N_12181,N_11472,N_11703);
xor U12182 (N_12182,N_11326,N_11738);
and U12183 (N_12183,N_11463,N_11706);
or U12184 (N_12184,N_11810,N_11526);
xnor U12185 (N_12185,N_11693,N_11870);
nor U12186 (N_12186,N_11342,N_11865);
and U12187 (N_12187,N_11283,N_11637);
and U12188 (N_12188,N_11447,N_11495);
and U12189 (N_12189,N_11648,N_11768);
and U12190 (N_12190,N_11400,N_11255);
nand U12191 (N_12191,N_11341,N_11616);
or U12192 (N_12192,N_11300,N_11723);
nor U12193 (N_12193,N_11551,N_11797);
nor U12194 (N_12194,N_11802,N_11541);
xor U12195 (N_12195,N_11503,N_11751);
and U12196 (N_12196,N_11645,N_11595);
nand U12197 (N_12197,N_11819,N_11509);
nor U12198 (N_12198,N_11551,N_11765);
xor U12199 (N_12199,N_11300,N_11686);
xor U12200 (N_12200,N_11455,N_11830);
nor U12201 (N_12201,N_11688,N_11759);
or U12202 (N_12202,N_11616,N_11524);
xor U12203 (N_12203,N_11371,N_11761);
xor U12204 (N_12204,N_11567,N_11361);
xnor U12205 (N_12205,N_11606,N_11853);
nand U12206 (N_12206,N_11561,N_11517);
nor U12207 (N_12207,N_11601,N_11558);
and U12208 (N_12208,N_11292,N_11467);
or U12209 (N_12209,N_11751,N_11579);
xor U12210 (N_12210,N_11830,N_11502);
xnor U12211 (N_12211,N_11785,N_11350);
nor U12212 (N_12212,N_11836,N_11609);
or U12213 (N_12213,N_11319,N_11345);
xnor U12214 (N_12214,N_11580,N_11619);
nor U12215 (N_12215,N_11448,N_11589);
or U12216 (N_12216,N_11432,N_11334);
xor U12217 (N_12217,N_11492,N_11708);
nand U12218 (N_12218,N_11357,N_11664);
or U12219 (N_12219,N_11394,N_11710);
nor U12220 (N_12220,N_11338,N_11636);
or U12221 (N_12221,N_11571,N_11484);
and U12222 (N_12222,N_11532,N_11684);
or U12223 (N_12223,N_11483,N_11756);
nand U12224 (N_12224,N_11870,N_11319);
xor U12225 (N_12225,N_11263,N_11488);
or U12226 (N_12226,N_11310,N_11279);
and U12227 (N_12227,N_11276,N_11739);
nor U12228 (N_12228,N_11394,N_11345);
xor U12229 (N_12229,N_11419,N_11372);
xor U12230 (N_12230,N_11654,N_11455);
or U12231 (N_12231,N_11735,N_11765);
or U12232 (N_12232,N_11695,N_11868);
nand U12233 (N_12233,N_11749,N_11353);
xnor U12234 (N_12234,N_11526,N_11749);
nor U12235 (N_12235,N_11696,N_11808);
xor U12236 (N_12236,N_11428,N_11307);
xor U12237 (N_12237,N_11269,N_11320);
nand U12238 (N_12238,N_11655,N_11538);
and U12239 (N_12239,N_11617,N_11301);
nand U12240 (N_12240,N_11668,N_11585);
xnor U12241 (N_12241,N_11838,N_11777);
or U12242 (N_12242,N_11538,N_11806);
and U12243 (N_12243,N_11274,N_11411);
and U12244 (N_12244,N_11670,N_11357);
or U12245 (N_12245,N_11802,N_11466);
and U12246 (N_12246,N_11709,N_11792);
or U12247 (N_12247,N_11843,N_11752);
or U12248 (N_12248,N_11659,N_11424);
or U12249 (N_12249,N_11765,N_11255);
nand U12250 (N_12250,N_11452,N_11496);
nand U12251 (N_12251,N_11826,N_11480);
nor U12252 (N_12252,N_11637,N_11469);
nand U12253 (N_12253,N_11251,N_11827);
nand U12254 (N_12254,N_11694,N_11343);
or U12255 (N_12255,N_11493,N_11278);
nor U12256 (N_12256,N_11279,N_11792);
nor U12257 (N_12257,N_11352,N_11360);
or U12258 (N_12258,N_11579,N_11347);
nor U12259 (N_12259,N_11304,N_11712);
nand U12260 (N_12260,N_11436,N_11747);
nand U12261 (N_12261,N_11726,N_11301);
xor U12262 (N_12262,N_11273,N_11806);
nor U12263 (N_12263,N_11778,N_11446);
nand U12264 (N_12264,N_11604,N_11332);
nand U12265 (N_12265,N_11336,N_11318);
xnor U12266 (N_12266,N_11298,N_11462);
and U12267 (N_12267,N_11554,N_11532);
xnor U12268 (N_12268,N_11665,N_11349);
xor U12269 (N_12269,N_11822,N_11453);
nand U12270 (N_12270,N_11558,N_11571);
nand U12271 (N_12271,N_11734,N_11659);
nand U12272 (N_12272,N_11824,N_11581);
and U12273 (N_12273,N_11321,N_11835);
xnor U12274 (N_12274,N_11418,N_11270);
or U12275 (N_12275,N_11834,N_11719);
and U12276 (N_12276,N_11417,N_11255);
nor U12277 (N_12277,N_11253,N_11467);
nand U12278 (N_12278,N_11620,N_11322);
or U12279 (N_12279,N_11843,N_11433);
nand U12280 (N_12280,N_11842,N_11380);
and U12281 (N_12281,N_11683,N_11439);
nand U12282 (N_12282,N_11554,N_11617);
nand U12283 (N_12283,N_11562,N_11364);
or U12284 (N_12284,N_11381,N_11501);
xor U12285 (N_12285,N_11711,N_11784);
nor U12286 (N_12286,N_11611,N_11517);
xnor U12287 (N_12287,N_11516,N_11852);
xnor U12288 (N_12288,N_11720,N_11600);
nor U12289 (N_12289,N_11583,N_11378);
nor U12290 (N_12290,N_11279,N_11402);
nor U12291 (N_12291,N_11790,N_11407);
and U12292 (N_12292,N_11354,N_11411);
xor U12293 (N_12293,N_11847,N_11680);
or U12294 (N_12294,N_11718,N_11761);
xnor U12295 (N_12295,N_11520,N_11657);
or U12296 (N_12296,N_11374,N_11778);
nor U12297 (N_12297,N_11259,N_11332);
and U12298 (N_12298,N_11340,N_11625);
or U12299 (N_12299,N_11355,N_11867);
xor U12300 (N_12300,N_11716,N_11354);
xnor U12301 (N_12301,N_11289,N_11368);
and U12302 (N_12302,N_11720,N_11427);
and U12303 (N_12303,N_11291,N_11815);
nand U12304 (N_12304,N_11659,N_11354);
and U12305 (N_12305,N_11616,N_11778);
xnor U12306 (N_12306,N_11342,N_11378);
or U12307 (N_12307,N_11301,N_11557);
nor U12308 (N_12308,N_11399,N_11374);
nor U12309 (N_12309,N_11730,N_11551);
and U12310 (N_12310,N_11592,N_11479);
nor U12311 (N_12311,N_11465,N_11497);
nor U12312 (N_12312,N_11544,N_11607);
and U12313 (N_12313,N_11532,N_11314);
nor U12314 (N_12314,N_11420,N_11490);
xnor U12315 (N_12315,N_11273,N_11769);
or U12316 (N_12316,N_11648,N_11794);
and U12317 (N_12317,N_11342,N_11461);
or U12318 (N_12318,N_11561,N_11745);
or U12319 (N_12319,N_11811,N_11611);
xnor U12320 (N_12320,N_11622,N_11604);
nand U12321 (N_12321,N_11705,N_11506);
or U12322 (N_12322,N_11556,N_11780);
nand U12323 (N_12323,N_11663,N_11573);
xnor U12324 (N_12324,N_11711,N_11517);
nand U12325 (N_12325,N_11830,N_11444);
nand U12326 (N_12326,N_11383,N_11844);
xor U12327 (N_12327,N_11413,N_11706);
nor U12328 (N_12328,N_11388,N_11636);
nand U12329 (N_12329,N_11592,N_11303);
and U12330 (N_12330,N_11873,N_11258);
xnor U12331 (N_12331,N_11692,N_11495);
xor U12332 (N_12332,N_11327,N_11742);
nor U12333 (N_12333,N_11791,N_11400);
nor U12334 (N_12334,N_11511,N_11459);
nor U12335 (N_12335,N_11404,N_11816);
nor U12336 (N_12336,N_11647,N_11843);
and U12337 (N_12337,N_11561,N_11647);
or U12338 (N_12338,N_11543,N_11352);
and U12339 (N_12339,N_11449,N_11414);
or U12340 (N_12340,N_11283,N_11302);
nor U12341 (N_12341,N_11675,N_11374);
xor U12342 (N_12342,N_11502,N_11410);
xnor U12343 (N_12343,N_11253,N_11724);
and U12344 (N_12344,N_11402,N_11855);
nand U12345 (N_12345,N_11607,N_11528);
and U12346 (N_12346,N_11535,N_11663);
nor U12347 (N_12347,N_11706,N_11313);
or U12348 (N_12348,N_11315,N_11678);
nand U12349 (N_12349,N_11836,N_11668);
nand U12350 (N_12350,N_11754,N_11858);
or U12351 (N_12351,N_11451,N_11300);
and U12352 (N_12352,N_11651,N_11601);
nor U12353 (N_12353,N_11673,N_11601);
nor U12354 (N_12354,N_11781,N_11459);
and U12355 (N_12355,N_11528,N_11595);
and U12356 (N_12356,N_11592,N_11475);
or U12357 (N_12357,N_11859,N_11576);
xnor U12358 (N_12358,N_11714,N_11723);
and U12359 (N_12359,N_11842,N_11535);
and U12360 (N_12360,N_11756,N_11753);
or U12361 (N_12361,N_11855,N_11435);
xnor U12362 (N_12362,N_11376,N_11430);
nor U12363 (N_12363,N_11675,N_11730);
nor U12364 (N_12364,N_11414,N_11277);
and U12365 (N_12365,N_11829,N_11706);
nand U12366 (N_12366,N_11259,N_11363);
and U12367 (N_12367,N_11290,N_11747);
and U12368 (N_12368,N_11713,N_11348);
xnor U12369 (N_12369,N_11724,N_11367);
nand U12370 (N_12370,N_11808,N_11754);
xor U12371 (N_12371,N_11650,N_11280);
xor U12372 (N_12372,N_11600,N_11510);
nand U12373 (N_12373,N_11686,N_11389);
nor U12374 (N_12374,N_11835,N_11350);
and U12375 (N_12375,N_11479,N_11565);
and U12376 (N_12376,N_11652,N_11393);
nor U12377 (N_12377,N_11382,N_11359);
and U12378 (N_12378,N_11466,N_11591);
or U12379 (N_12379,N_11812,N_11852);
or U12380 (N_12380,N_11617,N_11702);
or U12381 (N_12381,N_11845,N_11837);
or U12382 (N_12382,N_11809,N_11361);
and U12383 (N_12383,N_11695,N_11257);
or U12384 (N_12384,N_11720,N_11363);
nor U12385 (N_12385,N_11346,N_11484);
and U12386 (N_12386,N_11712,N_11790);
xor U12387 (N_12387,N_11270,N_11748);
or U12388 (N_12388,N_11703,N_11856);
xor U12389 (N_12389,N_11831,N_11656);
or U12390 (N_12390,N_11868,N_11353);
xor U12391 (N_12391,N_11707,N_11610);
nor U12392 (N_12392,N_11371,N_11690);
xnor U12393 (N_12393,N_11343,N_11490);
and U12394 (N_12394,N_11270,N_11433);
and U12395 (N_12395,N_11688,N_11619);
nor U12396 (N_12396,N_11535,N_11493);
or U12397 (N_12397,N_11790,N_11748);
xnor U12398 (N_12398,N_11326,N_11511);
nand U12399 (N_12399,N_11317,N_11318);
and U12400 (N_12400,N_11726,N_11473);
or U12401 (N_12401,N_11533,N_11813);
xnor U12402 (N_12402,N_11567,N_11430);
nor U12403 (N_12403,N_11826,N_11844);
and U12404 (N_12404,N_11577,N_11666);
xnor U12405 (N_12405,N_11364,N_11860);
or U12406 (N_12406,N_11679,N_11658);
nor U12407 (N_12407,N_11316,N_11648);
xor U12408 (N_12408,N_11823,N_11368);
and U12409 (N_12409,N_11703,N_11604);
xnor U12410 (N_12410,N_11626,N_11519);
and U12411 (N_12411,N_11828,N_11674);
nand U12412 (N_12412,N_11501,N_11741);
nand U12413 (N_12413,N_11484,N_11297);
and U12414 (N_12414,N_11442,N_11687);
xnor U12415 (N_12415,N_11865,N_11364);
nor U12416 (N_12416,N_11538,N_11539);
nor U12417 (N_12417,N_11647,N_11459);
nor U12418 (N_12418,N_11503,N_11664);
and U12419 (N_12419,N_11809,N_11634);
and U12420 (N_12420,N_11487,N_11869);
nor U12421 (N_12421,N_11662,N_11341);
nand U12422 (N_12422,N_11552,N_11506);
nand U12423 (N_12423,N_11470,N_11595);
nand U12424 (N_12424,N_11402,N_11371);
or U12425 (N_12425,N_11716,N_11332);
nor U12426 (N_12426,N_11612,N_11337);
nor U12427 (N_12427,N_11548,N_11345);
nor U12428 (N_12428,N_11304,N_11361);
and U12429 (N_12429,N_11333,N_11461);
nand U12430 (N_12430,N_11820,N_11554);
and U12431 (N_12431,N_11532,N_11323);
or U12432 (N_12432,N_11522,N_11599);
or U12433 (N_12433,N_11326,N_11586);
and U12434 (N_12434,N_11506,N_11824);
nand U12435 (N_12435,N_11442,N_11829);
xor U12436 (N_12436,N_11810,N_11595);
or U12437 (N_12437,N_11803,N_11542);
or U12438 (N_12438,N_11336,N_11531);
nor U12439 (N_12439,N_11871,N_11632);
nor U12440 (N_12440,N_11693,N_11464);
xnor U12441 (N_12441,N_11677,N_11357);
xor U12442 (N_12442,N_11258,N_11833);
or U12443 (N_12443,N_11704,N_11441);
nor U12444 (N_12444,N_11253,N_11408);
and U12445 (N_12445,N_11857,N_11842);
nor U12446 (N_12446,N_11773,N_11810);
xnor U12447 (N_12447,N_11358,N_11288);
xnor U12448 (N_12448,N_11767,N_11758);
nand U12449 (N_12449,N_11310,N_11282);
xnor U12450 (N_12450,N_11722,N_11467);
and U12451 (N_12451,N_11533,N_11763);
xnor U12452 (N_12452,N_11423,N_11396);
xor U12453 (N_12453,N_11485,N_11591);
and U12454 (N_12454,N_11380,N_11736);
xnor U12455 (N_12455,N_11831,N_11828);
nor U12456 (N_12456,N_11459,N_11794);
nor U12457 (N_12457,N_11792,N_11312);
and U12458 (N_12458,N_11305,N_11787);
nor U12459 (N_12459,N_11527,N_11251);
nor U12460 (N_12460,N_11347,N_11833);
nor U12461 (N_12461,N_11518,N_11617);
nand U12462 (N_12462,N_11440,N_11872);
or U12463 (N_12463,N_11661,N_11370);
or U12464 (N_12464,N_11562,N_11753);
and U12465 (N_12465,N_11829,N_11424);
nand U12466 (N_12466,N_11565,N_11377);
xor U12467 (N_12467,N_11836,N_11482);
nand U12468 (N_12468,N_11587,N_11381);
or U12469 (N_12469,N_11370,N_11669);
xor U12470 (N_12470,N_11497,N_11604);
or U12471 (N_12471,N_11424,N_11338);
nand U12472 (N_12472,N_11292,N_11331);
nand U12473 (N_12473,N_11466,N_11534);
nand U12474 (N_12474,N_11768,N_11774);
xor U12475 (N_12475,N_11381,N_11446);
and U12476 (N_12476,N_11302,N_11284);
or U12477 (N_12477,N_11372,N_11278);
or U12478 (N_12478,N_11744,N_11709);
xnor U12479 (N_12479,N_11866,N_11712);
and U12480 (N_12480,N_11814,N_11490);
nor U12481 (N_12481,N_11318,N_11456);
xor U12482 (N_12482,N_11571,N_11349);
xnor U12483 (N_12483,N_11365,N_11776);
or U12484 (N_12484,N_11328,N_11678);
nand U12485 (N_12485,N_11562,N_11798);
nor U12486 (N_12486,N_11574,N_11644);
nand U12487 (N_12487,N_11286,N_11510);
or U12488 (N_12488,N_11458,N_11853);
nor U12489 (N_12489,N_11290,N_11836);
nor U12490 (N_12490,N_11809,N_11727);
xor U12491 (N_12491,N_11817,N_11267);
and U12492 (N_12492,N_11664,N_11826);
or U12493 (N_12493,N_11601,N_11498);
nor U12494 (N_12494,N_11376,N_11587);
and U12495 (N_12495,N_11711,N_11807);
nand U12496 (N_12496,N_11790,N_11730);
or U12497 (N_12497,N_11423,N_11542);
or U12498 (N_12498,N_11444,N_11313);
nor U12499 (N_12499,N_11774,N_11846);
or U12500 (N_12500,N_12499,N_12358);
nor U12501 (N_12501,N_12019,N_12395);
nand U12502 (N_12502,N_12181,N_12281);
nand U12503 (N_12503,N_12208,N_12115);
nor U12504 (N_12504,N_12299,N_11876);
nand U12505 (N_12505,N_11927,N_12165);
and U12506 (N_12506,N_12390,N_12069);
nand U12507 (N_12507,N_12397,N_12369);
nand U12508 (N_12508,N_12394,N_12344);
nand U12509 (N_12509,N_12391,N_12347);
and U12510 (N_12510,N_12139,N_12210);
and U12511 (N_12511,N_12207,N_11966);
nand U12512 (N_12512,N_12310,N_12434);
nor U12513 (N_12513,N_11963,N_12167);
nand U12514 (N_12514,N_12349,N_12444);
or U12515 (N_12515,N_12414,N_12017);
xor U12516 (N_12516,N_12380,N_12376);
or U12517 (N_12517,N_12042,N_12327);
and U12518 (N_12518,N_12236,N_11923);
xor U12519 (N_12519,N_12011,N_11891);
nor U12520 (N_12520,N_12475,N_12476);
nand U12521 (N_12521,N_12145,N_11917);
nand U12522 (N_12522,N_11916,N_11895);
xor U12523 (N_12523,N_12201,N_12126);
or U12524 (N_12524,N_11987,N_12151);
xnor U12525 (N_12525,N_12421,N_12137);
nand U12526 (N_12526,N_12027,N_12152);
nand U12527 (N_12527,N_12399,N_12334);
and U12528 (N_12528,N_12100,N_12315);
nand U12529 (N_12529,N_12332,N_12097);
xnor U12530 (N_12530,N_12345,N_12287);
and U12531 (N_12531,N_12498,N_12381);
xnor U12532 (N_12532,N_12452,N_12050);
nor U12533 (N_12533,N_12193,N_12166);
xor U12534 (N_12534,N_11933,N_12229);
nand U12535 (N_12535,N_12138,N_12159);
nand U12536 (N_12536,N_12295,N_11905);
nand U12537 (N_12537,N_12328,N_12062);
and U12538 (N_12538,N_12464,N_12238);
nand U12539 (N_12539,N_11886,N_12075);
xor U12540 (N_12540,N_12154,N_12186);
xnor U12541 (N_12541,N_12226,N_12018);
nor U12542 (N_12542,N_11990,N_12418);
and U12543 (N_12543,N_12179,N_12259);
nor U12544 (N_12544,N_12492,N_12266);
xor U12545 (N_12545,N_12455,N_12090);
xnor U12546 (N_12546,N_12038,N_12083);
nand U12547 (N_12547,N_11913,N_12180);
and U12548 (N_12548,N_12121,N_12023);
or U12549 (N_12549,N_12463,N_12483);
or U12550 (N_12550,N_11964,N_11888);
xnor U12551 (N_12551,N_12346,N_12077);
or U12552 (N_12552,N_12136,N_11984);
xnor U12553 (N_12553,N_12454,N_12158);
nand U12554 (N_12554,N_12248,N_11911);
nor U12555 (N_12555,N_12211,N_12339);
nor U12556 (N_12556,N_12191,N_12085);
or U12557 (N_12557,N_12044,N_12348);
nand U12558 (N_12558,N_12196,N_12417);
nand U12559 (N_12559,N_12387,N_12477);
and U12560 (N_12560,N_12024,N_12053);
nor U12561 (N_12561,N_11968,N_12441);
or U12562 (N_12562,N_12330,N_12448);
and U12563 (N_12563,N_12322,N_12325);
xnor U12564 (N_12564,N_12192,N_12060);
nor U12565 (N_12565,N_12102,N_12013);
or U12566 (N_12566,N_12222,N_12131);
and U12567 (N_12567,N_12362,N_11887);
nand U12568 (N_12568,N_12064,N_12220);
and U12569 (N_12569,N_12480,N_12262);
xnor U12570 (N_12570,N_11962,N_12146);
or U12571 (N_12571,N_12081,N_11985);
nand U12572 (N_12572,N_12438,N_12244);
nand U12573 (N_12573,N_11920,N_12405);
xnor U12574 (N_12574,N_11953,N_12355);
nor U12575 (N_12575,N_12103,N_12482);
and U12576 (N_12576,N_12401,N_12384);
and U12577 (N_12577,N_11991,N_12089);
nor U12578 (N_12578,N_11909,N_12361);
nor U12579 (N_12579,N_12304,N_12489);
nand U12580 (N_12580,N_12134,N_12486);
and U12581 (N_12581,N_12016,N_11881);
nand U12582 (N_12582,N_12010,N_12288);
nand U12583 (N_12583,N_12432,N_12487);
and U12584 (N_12584,N_12471,N_12264);
nand U12585 (N_12585,N_12459,N_12130);
nand U12586 (N_12586,N_12247,N_12243);
xnor U12587 (N_12587,N_12224,N_12048);
nor U12588 (N_12588,N_11918,N_12305);
or U12589 (N_12589,N_11976,N_12172);
or U12590 (N_12590,N_11978,N_12034);
and U12591 (N_12591,N_12485,N_11974);
and U12592 (N_12592,N_11970,N_12363);
xor U12593 (N_12593,N_12123,N_12317);
nand U12594 (N_12594,N_12200,N_12422);
nor U12595 (N_12595,N_12036,N_12292);
nor U12596 (N_12596,N_12311,N_12231);
and U12597 (N_12597,N_12219,N_12338);
nor U12598 (N_12598,N_12319,N_12007);
and U12599 (N_12599,N_11982,N_11921);
nand U12600 (N_12600,N_12240,N_12080);
nor U12601 (N_12601,N_12020,N_11961);
nand U12602 (N_12602,N_12415,N_12357);
nand U12603 (N_12603,N_12368,N_11906);
and U12604 (N_12604,N_11935,N_11930);
nand U12605 (N_12605,N_12284,N_12261);
and U12606 (N_12606,N_11983,N_11879);
nand U12607 (N_12607,N_12120,N_12199);
xor U12608 (N_12608,N_12300,N_12128);
xor U12609 (N_12609,N_12353,N_12169);
and U12610 (N_12610,N_12105,N_11952);
and U12611 (N_12611,N_12478,N_12263);
nor U12612 (N_12612,N_12116,N_12450);
or U12613 (N_12613,N_12155,N_11892);
and U12614 (N_12614,N_12407,N_12323);
nand U12615 (N_12615,N_12135,N_12253);
xor U12616 (N_12616,N_12141,N_12076);
or U12617 (N_12617,N_12337,N_12271);
xor U12618 (N_12618,N_12379,N_12051);
nor U12619 (N_12619,N_12096,N_12178);
nand U12620 (N_12620,N_12117,N_12443);
and U12621 (N_12621,N_12177,N_12230);
nand U12622 (N_12622,N_12213,N_12067);
or U12623 (N_12623,N_11902,N_12406);
xor U12624 (N_12624,N_12043,N_11986);
xor U12625 (N_12625,N_11956,N_12101);
nor U12626 (N_12626,N_11955,N_12484);
or U12627 (N_12627,N_12298,N_12351);
and U12628 (N_12628,N_11925,N_12065);
nand U12629 (N_12629,N_12112,N_11960);
nand U12630 (N_12630,N_12082,N_12119);
xor U12631 (N_12631,N_11979,N_12419);
and U12632 (N_12632,N_12257,N_12205);
nand U12633 (N_12633,N_12092,N_12110);
or U12634 (N_12634,N_12129,N_12197);
or U12635 (N_12635,N_12184,N_12140);
nor U12636 (N_12636,N_12424,N_12250);
nor U12637 (N_12637,N_12233,N_12153);
nor U12638 (N_12638,N_12469,N_12370);
nand U12639 (N_12639,N_12467,N_12458);
or U12640 (N_12640,N_12033,N_12055);
nand U12641 (N_12641,N_12239,N_12289);
xnor U12642 (N_12642,N_12326,N_12286);
and U12643 (N_12643,N_12331,N_12133);
nand U12644 (N_12644,N_12256,N_12160);
xor U12645 (N_12645,N_12147,N_12277);
nand U12646 (N_12646,N_12366,N_11877);
nor U12647 (N_12647,N_11882,N_11901);
nand U12648 (N_12648,N_11999,N_12021);
or U12649 (N_12649,N_12070,N_12296);
nor U12650 (N_12650,N_11893,N_12161);
or U12651 (N_12651,N_12047,N_12314);
or U12652 (N_12652,N_12308,N_12212);
and U12653 (N_12653,N_12113,N_11958);
nor U12654 (N_12654,N_11915,N_12496);
nor U12655 (N_12655,N_12061,N_11939);
xor U12656 (N_12656,N_12462,N_12378);
or U12657 (N_12657,N_12079,N_12371);
nor U12658 (N_12658,N_12254,N_12383);
nand U12659 (N_12659,N_12290,N_11994);
and U12660 (N_12660,N_12251,N_12106);
nand U12661 (N_12661,N_11929,N_12400);
xnor U12662 (N_12662,N_12218,N_11965);
nor U12663 (N_12663,N_12059,N_11972);
nor U12664 (N_12664,N_12031,N_12143);
xnor U12665 (N_12665,N_11938,N_12427);
or U12666 (N_12666,N_12258,N_12375);
and U12667 (N_12667,N_12148,N_12402);
and U12668 (N_12668,N_12012,N_12303);
and U12669 (N_12669,N_12189,N_11880);
or U12670 (N_12670,N_12056,N_12360);
nand U12671 (N_12671,N_12388,N_12194);
nor U12672 (N_12672,N_11949,N_12009);
nor U12673 (N_12673,N_12037,N_12445);
or U12674 (N_12674,N_12490,N_12282);
nor U12675 (N_12675,N_11971,N_12086);
or U12676 (N_12676,N_12260,N_12124);
nand U12677 (N_12677,N_12202,N_11885);
or U12678 (N_12678,N_12472,N_11910);
nor U12679 (N_12679,N_12175,N_12431);
or U12680 (N_12680,N_11937,N_12150);
and U12681 (N_12681,N_12227,N_11948);
xnor U12682 (N_12682,N_11980,N_11977);
nor U12683 (N_12683,N_11907,N_12393);
nand U12684 (N_12684,N_12108,N_11903);
nand U12685 (N_12685,N_12000,N_12099);
nor U12686 (N_12686,N_12412,N_12029);
nand U12687 (N_12687,N_12275,N_12032);
or U12688 (N_12688,N_12234,N_11969);
nor U12689 (N_12689,N_12392,N_12232);
and U12690 (N_12690,N_11878,N_12035);
xor U12691 (N_12691,N_12267,N_11889);
nand U12692 (N_12692,N_12206,N_11973);
or U12693 (N_12693,N_12335,N_12365);
or U12694 (N_12694,N_11942,N_12474);
nor U12695 (N_12695,N_12372,N_12001);
or U12696 (N_12696,N_12428,N_12408);
or U12697 (N_12697,N_11950,N_12276);
or U12698 (N_12698,N_12409,N_12359);
or U12699 (N_12699,N_11941,N_12190);
nand U12700 (N_12700,N_12057,N_12403);
xnor U12701 (N_12701,N_12203,N_12309);
nor U12702 (N_12702,N_12350,N_12214);
xnor U12703 (N_12703,N_12066,N_12249);
and U12704 (N_12704,N_12336,N_11912);
nor U12705 (N_12705,N_12285,N_12301);
or U12706 (N_12706,N_12235,N_12142);
xnor U12707 (N_12707,N_12283,N_12374);
or U12708 (N_12708,N_12026,N_11997);
or U12709 (N_12709,N_11940,N_12488);
or U12710 (N_12710,N_11975,N_12280);
nor U12711 (N_12711,N_11992,N_11995);
nor U12712 (N_12712,N_12164,N_11936);
nor U12713 (N_12713,N_12479,N_12246);
nand U12714 (N_12714,N_12420,N_12041);
nor U12715 (N_12715,N_12265,N_12003);
xnor U12716 (N_12716,N_12342,N_12429);
and U12717 (N_12717,N_12049,N_11928);
or U12718 (N_12718,N_12094,N_12430);
xor U12719 (N_12719,N_12436,N_12063);
nor U12720 (N_12720,N_12216,N_12447);
nor U12721 (N_12721,N_12198,N_12377);
and U12722 (N_12722,N_11988,N_12183);
or U12723 (N_12723,N_12343,N_11900);
nand U12724 (N_12724,N_12188,N_12095);
and U12725 (N_12725,N_12302,N_12237);
and U12726 (N_12726,N_11943,N_12209);
nor U12727 (N_12727,N_12457,N_12114);
nor U12728 (N_12728,N_12078,N_12093);
and U12729 (N_12729,N_11926,N_12015);
nor U12730 (N_12730,N_12386,N_12473);
or U12731 (N_12731,N_11946,N_12127);
or U12732 (N_12732,N_12091,N_12320);
nor U12733 (N_12733,N_12149,N_12088);
xor U12734 (N_12734,N_12118,N_12404);
nand U12735 (N_12735,N_12030,N_12045);
and U12736 (N_12736,N_12341,N_12410);
nor U12737 (N_12737,N_12221,N_12252);
and U12738 (N_12738,N_12312,N_11947);
nand U12739 (N_12739,N_12170,N_12187);
nor U12740 (N_12740,N_11924,N_12456);
or U12741 (N_12741,N_11908,N_12356);
nor U12742 (N_12742,N_12125,N_12435);
nor U12743 (N_12743,N_12052,N_12451);
or U12744 (N_12744,N_11897,N_12367);
nor U12745 (N_12745,N_12382,N_11934);
xor U12746 (N_12746,N_12316,N_11884);
and U12747 (N_12747,N_12468,N_12493);
nand U12748 (N_12748,N_12109,N_12497);
nor U12749 (N_12749,N_12002,N_12228);
xnor U12750 (N_12750,N_12278,N_11914);
xnor U12751 (N_12751,N_12491,N_12040);
xor U12752 (N_12752,N_11959,N_12306);
and U12753 (N_12753,N_12416,N_12460);
nor U12754 (N_12754,N_11945,N_12297);
and U12755 (N_12755,N_12269,N_12425);
and U12756 (N_12756,N_12398,N_12274);
or U12757 (N_12757,N_11899,N_12225);
nand U12758 (N_12758,N_12072,N_12074);
nand U12759 (N_12759,N_12071,N_12329);
and U12760 (N_12760,N_12279,N_11898);
nand U12761 (N_12761,N_11875,N_12058);
nand U12762 (N_12762,N_12433,N_11989);
nand U12763 (N_12763,N_12204,N_12272);
and U12764 (N_12764,N_12162,N_11996);
xnor U12765 (N_12765,N_12087,N_12122);
or U12766 (N_12766,N_12255,N_12446);
and U12767 (N_12767,N_11967,N_12163);
or U12768 (N_12768,N_12453,N_11932);
xnor U12769 (N_12769,N_12268,N_12111);
xor U12770 (N_12770,N_12084,N_12270);
xnor U12771 (N_12771,N_12157,N_11954);
and U12772 (N_12772,N_12465,N_12364);
xnor U12773 (N_12773,N_12006,N_11922);
nor U12774 (N_12774,N_12294,N_12132);
and U12775 (N_12775,N_12470,N_12440);
nand U12776 (N_12776,N_12004,N_12413);
nor U12777 (N_12777,N_12173,N_11944);
and U12778 (N_12778,N_12046,N_12340);
nand U12779 (N_12779,N_12373,N_12307);
xnor U12780 (N_12780,N_12008,N_12068);
and U12781 (N_12781,N_12171,N_12494);
or U12782 (N_12782,N_11998,N_12324);
and U12783 (N_12783,N_12442,N_12423);
nor U12784 (N_12784,N_12466,N_12182);
nor U12785 (N_12785,N_12449,N_12385);
or U12786 (N_12786,N_12025,N_11993);
and U12787 (N_12787,N_12005,N_12333);
nor U12788 (N_12788,N_12437,N_12411);
nand U12789 (N_12789,N_12176,N_12389);
and U12790 (N_12790,N_12273,N_12215);
nor U12791 (N_12791,N_12321,N_12104);
nand U12792 (N_12792,N_12481,N_11883);
and U12793 (N_12793,N_12242,N_11951);
nand U12794 (N_12794,N_12014,N_11904);
or U12795 (N_12795,N_12426,N_12168);
xnor U12796 (N_12796,N_12241,N_12291);
nand U12797 (N_12797,N_12293,N_12028);
or U12798 (N_12798,N_12223,N_12174);
nand U12799 (N_12799,N_11896,N_12054);
nand U12800 (N_12800,N_12073,N_12245);
nand U12801 (N_12801,N_12107,N_11957);
and U12802 (N_12802,N_12495,N_12185);
nand U12803 (N_12803,N_12039,N_12318);
nor U12804 (N_12804,N_12156,N_11894);
nor U12805 (N_12805,N_12217,N_11981);
or U12806 (N_12806,N_12313,N_11919);
nor U12807 (N_12807,N_11890,N_12098);
or U12808 (N_12808,N_12195,N_12352);
or U12809 (N_12809,N_11931,N_12396);
nand U12810 (N_12810,N_12439,N_12022);
xnor U12811 (N_12811,N_12354,N_12461);
nor U12812 (N_12812,N_12144,N_12057);
nor U12813 (N_12813,N_12325,N_12370);
or U12814 (N_12814,N_12439,N_11892);
nand U12815 (N_12815,N_12423,N_12013);
nor U12816 (N_12816,N_12031,N_12331);
nand U12817 (N_12817,N_12232,N_12349);
or U12818 (N_12818,N_11926,N_11969);
xor U12819 (N_12819,N_12215,N_12307);
nor U12820 (N_12820,N_12488,N_12286);
and U12821 (N_12821,N_12177,N_12223);
nor U12822 (N_12822,N_12317,N_12239);
and U12823 (N_12823,N_12251,N_12151);
nor U12824 (N_12824,N_12339,N_12497);
nor U12825 (N_12825,N_12193,N_11884);
or U12826 (N_12826,N_11987,N_12458);
nor U12827 (N_12827,N_11926,N_12277);
or U12828 (N_12828,N_12059,N_12369);
nand U12829 (N_12829,N_11987,N_12329);
and U12830 (N_12830,N_11925,N_12307);
and U12831 (N_12831,N_12088,N_11963);
xnor U12832 (N_12832,N_12243,N_12439);
and U12833 (N_12833,N_12491,N_11959);
or U12834 (N_12834,N_12067,N_12376);
and U12835 (N_12835,N_12275,N_12481);
xnor U12836 (N_12836,N_12266,N_12023);
xnor U12837 (N_12837,N_11989,N_12020);
nor U12838 (N_12838,N_12394,N_12427);
nand U12839 (N_12839,N_12346,N_11967);
and U12840 (N_12840,N_11999,N_12397);
xnor U12841 (N_12841,N_11994,N_12339);
nand U12842 (N_12842,N_12019,N_11933);
xor U12843 (N_12843,N_12008,N_11965);
or U12844 (N_12844,N_12487,N_12365);
and U12845 (N_12845,N_12082,N_11897);
nand U12846 (N_12846,N_11987,N_12208);
and U12847 (N_12847,N_12256,N_12194);
nor U12848 (N_12848,N_12170,N_12165);
nor U12849 (N_12849,N_11932,N_12308);
and U12850 (N_12850,N_12477,N_12479);
and U12851 (N_12851,N_12169,N_12419);
nand U12852 (N_12852,N_12417,N_12118);
nand U12853 (N_12853,N_12474,N_12162);
and U12854 (N_12854,N_12242,N_12104);
and U12855 (N_12855,N_12249,N_12161);
nor U12856 (N_12856,N_12303,N_12341);
nand U12857 (N_12857,N_12327,N_12431);
or U12858 (N_12858,N_12109,N_11977);
and U12859 (N_12859,N_12046,N_12222);
xnor U12860 (N_12860,N_12346,N_12037);
nor U12861 (N_12861,N_12180,N_12075);
or U12862 (N_12862,N_12133,N_12309);
nand U12863 (N_12863,N_11950,N_12434);
xor U12864 (N_12864,N_12003,N_12206);
xnor U12865 (N_12865,N_12175,N_12203);
and U12866 (N_12866,N_12479,N_12393);
or U12867 (N_12867,N_12025,N_11954);
and U12868 (N_12868,N_12090,N_12141);
or U12869 (N_12869,N_11919,N_12190);
nor U12870 (N_12870,N_12316,N_12346);
nor U12871 (N_12871,N_12498,N_11988);
nor U12872 (N_12872,N_12348,N_12060);
xnor U12873 (N_12873,N_12489,N_12384);
or U12874 (N_12874,N_12091,N_12156);
and U12875 (N_12875,N_11922,N_12416);
nand U12876 (N_12876,N_12449,N_12452);
xnor U12877 (N_12877,N_12015,N_11977);
xor U12878 (N_12878,N_12440,N_12412);
nor U12879 (N_12879,N_11955,N_12005);
and U12880 (N_12880,N_12159,N_12178);
or U12881 (N_12881,N_12300,N_12108);
and U12882 (N_12882,N_12107,N_12282);
nor U12883 (N_12883,N_12089,N_12266);
nand U12884 (N_12884,N_12258,N_12230);
nor U12885 (N_12885,N_11964,N_12225);
and U12886 (N_12886,N_11941,N_12335);
nand U12887 (N_12887,N_11930,N_12383);
and U12888 (N_12888,N_12492,N_12454);
nand U12889 (N_12889,N_12348,N_12143);
and U12890 (N_12890,N_12065,N_12009);
or U12891 (N_12891,N_12199,N_12214);
xnor U12892 (N_12892,N_12336,N_12270);
nor U12893 (N_12893,N_12451,N_12414);
nand U12894 (N_12894,N_12022,N_12476);
nand U12895 (N_12895,N_12039,N_12082);
and U12896 (N_12896,N_12338,N_12185);
and U12897 (N_12897,N_12378,N_12329);
nor U12898 (N_12898,N_12417,N_12119);
xnor U12899 (N_12899,N_12026,N_12022);
nand U12900 (N_12900,N_12334,N_11886);
and U12901 (N_12901,N_11910,N_12370);
and U12902 (N_12902,N_12257,N_12131);
nor U12903 (N_12903,N_12169,N_12162);
nor U12904 (N_12904,N_12206,N_11948);
nor U12905 (N_12905,N_12425,N_12006);
or U12906 (N_12906,N_12162,N_12282);
or U12907 (N_12907,N_12086,N_12425);
and U12908 (N_12908,N_12167,N_11903);
xor U12909 (N_12909,N_11929,N_12301);
nor U12910 (N_12910,N_12001,N_12082);
or U12911 (N_12911,N_12126,N_11877);
nor U12912 (N_12912,N_12469,N_12018);
nor U12913 (N_12913,N_12166,N_11948);
nor U12914 (N_12914,N_12185,N_12018);
and U12915 (N_12915,N_12062,N_12150);
or U12916 (N_12916,N_12427,N_12151);
or U12917 (N_12917,N_12475,N_11931);
nor U12918 (N_12918,N_12090,N_12148);
nand U12919 (N_12919,N_12473,N_12450);
nor U12920 (N_12920,N_12036,N_12104);
nor U12921 (N_12921,N_12187,N_12138);
and U12922 (N_12922,N_12143,N_11953);
xor U12923 (N_12923,N_11911,N_11907);
nor U12924 (N_12924,N_12144,N_12383);
nor U12925 (N_12925,N_12418,N_12314);
and U12926 (N_12926,N_12225,N_12294);
or U12927 (N_12927,N_12127,N_11933);
xnor U12928 (N_12928,N_12288,N_11908);
or U12929 (N_12929,N_11949,N_11957);
and U12930 (N_12930,N_12168,N_11985);
nor U12931 (N_12931,N_12004,N_12015);
or U12932 (N_12932,N_12277,N_12091);
nand U12933 (N_12933,N_12178,N_11921);
nor U12934 (N_12934,N_12072,N_11947);
nand U12935 (N_12935,N_12205,N_12480);
and U12936 (N_12936,N_12319,N_12090);
nand U12937 (N_12937,N_12040,N_12150);
and U12938 (N_12938,N_12241,N_12429);
and U12939 (N_12939,N_12398,N_12486);
nor U12940 (N_12940,N_12319,N_12428);
and U12941 (N_12941,N_12147,N_12258);
nand U12942 (N_12942,N_12042,N_12209);
or U12943 (N_12943,N_12424,N_11896);
and U12944 (N_12944,N_12287,N_12478);
xnor U12945 (N_12945,N_12085,N_11929);
or U12946 (N_12946,N_12020,N_12072);
xor U12947 (N_12947,N_12043,N_12246);
xnor U12948 (N_12948,N_12378,N_12464);
and U12949 (N_12949,N_12048,N_12307);
and U12950 (N_12950,N_12203,N_12188);
xnor U12951 (N_12951,N_12084,N_12332);
nor U12952 (N_12952,N_11894,N_12497);
xnor U12953 (N_12953,N_11917,N_12347);
nand U12954 (N_12954,N_11997,N_11947);
or U12955 (N_12955,N_12045,N_12410);
or U12956 (N_12956,N_12244,N_12414);
and U12957 (N_12957,N_12073,N_12236);
nand U12958 (N_12958,N_12183,N_12492);
nand U12959 (N_12959,N_12195,N_12444);
nand U12960 (N_12960,N_12215,N_12368);
and U12961 (N_12961,N_11989,N_11935);
or U12962 (N_12962,N_12278,N_12218);
xnor U12963 (N_12963,N_12325,N_12051);
nand U12964 (N_12964,N_11994,N_12424);
xnor U12965 (N_12965,N_12194,N_12125);
nand U12966 (N_12966,N_12045,N_12492);
nor U12967 (N_12967,N_12049,N_12418);
or U12968 (N_12968,N_12074,N_12491);
nand U12969 (N_12969,N_12229,N_12322);
xnor U12970 (N_12970,N_11976,N_12262);
nor U12971 (N_12971,N_12378,N_11955);
nand U12972 (N_12972,N_11940,N_12079);
nor U12973 (N_12973,N_12238,N_12298);
or U12974 (N_12974,N_12231,N_12422);
nand U12975 (N_12975,N_12011,N_12289);
nor U12976 (N_12976,N_12251,N_11899);
and U12977 (N_12977,N_12227,N_12425);
and U12978 (N_12978,N_12342,N_12305);
nor U12979 (N_12979,N_11937,N_12060);
xor U12980 (N_12980,N_12085,N_12230);
xnor U12981 (N_12981,N_12078,N_12124);
and U12982 (N_12982,N_12401,N_12406);
nor U12983 (N_12983,N_12332,N_12306);
nand U12984 (N_12984,N_12247,N_11893);
or U12985 (N_12985,N_11943,N_12072);
nand U12986 (N_12986,N_11883,N_12350);
nor U12987 (N_12987,N_12490,N_12474);
xnor U12988 (N_12988,N_12395,N_11962);
or U12989 (N_12989,N_12474,N_11965);
and U12990 (N_12990,N_12155,N_12274);
nor U12991 (N_12991,N_12430,N_12458);
or U12992 (N_12992,N_11881,N_12105);
and U12993 (N_12993,N_11987,N_12301);
nand U12994 (N_12994,N_11926,N_11978);
xnor U12995 (N_12995,N_12210,N_11914);
nor U12996 (N_12996,N_12234,N_11994);
xnor U12997 (N_12997,N_11887,N_12401);
or U12998 (N_12998,N_12129,N_12188);
nor U12999 (N_12999,N_12241,N_12243);
and U13000 (N_13000,N_12089,N_12038);
and U13001 (N_13001,N_12429,N_11899);
or U13002 (N_13002,N_12317,N_11925);
or U13003 (N_13003,N_12146,N_12124);
xnor U13004 (N_13004,N_12330,N_12135);
xor U13005 (N_13005,N_12188,N_12349);
and U13006 (N_13006,N_12482,N_11929);
nor U13007 (N_13007,N_12166,N_12065);
or U13008 (N_13008,N_11913,N_12347);
nor U13009 (N_13009,N_12343,N_12479);
xnor U13010 (N_13010,N_11891,N_12016);
xor U13011 (N_13011,N_12399,N_11895);
nand U13012 (N_13012,N_12350,N_12102);
nor U13013 (N_13013,N_12290,N_12131);
nand U13014 (N_13014,N_12128,N_12022);
and U13015 (N_13015,N_12225,N_11995);
nor U13016 (N_13016,N_11937,N_12429);
and U13017 (N_13017,N_11980,N_12438);
xnor U13018 (N_13018,N_12494,N_12435);
and U13019 (N_13019,N_12095,N_12435);
xor U13020 (N_13020,N_12273,N_12475);
or U13021 (N_13021,N_12165,N_12348);
xor U13022 (N_13022,N_12392,N_11954);
nand U13023 (N_13023,N_12401,N_11951);
xnor U13024 (N_13024,N_12113,N_12394);
nor U13025 (N_13025,N_12254,N_12311);
nand U13026 (N_13026,N_12053,N_12224);
or U13027 (N_13027,N_12021,N_12150);
nand U13028 (N_13028,N_12429,N_12075);
nor U13029 (N_13029,N_11895,N_12327);
nor U13030 (N_13030,N_12342,N_12134);
nand U13031 (N_13031,N_11924,N_12439);
nand U13032 (N_13032,N_12487,N_12206);
and U13033 (N_13033,N_12439,N_11950);
and U13034 (N_13034,N_12196,N_12262);
and U13035 (N_13035,N_12274,N_12130);
or U13036 (N_13036,N_12412,N_11880);
xnor U13037 (N_13037,N_12222,N_12302);
or U13038 (N_13038,N_11953,N_11884);
and U13039 (N_13039,N_11946,N_12256);
nand U13040 (N_13040,N_12420,N_11883);
xor U13041 (N_13041,N_12345,N_12397);
or U13042 (N_13042,N_12245,N_12107);
or U13043 (N_13043,N_12375,N_12273);
nand U13044 (N_13044,N_12225,N_12163);
or U13045 (N_13045,N_12407,N_12395);
or U13046 (N_13046,N_12434,N_12098);
nand U13047 (N_13047,N_11983,N_12222);
or U13048 (N_13048,N_12040,N_12003);
xnor U13049 (N_13049,N_11929,N_11902);
and U13050 (N_13050,N_12497,N_12066);
or U13051 (N_13051,N_12414,N_12331);
or U13052 (N_13052,N_12019,N_12288);
and U13053 (N_13053,N_12025,N_12410);
nor U13054 (N_13054,N_12327,N_12290);
nand U13055 (N_13055,N_12130,N_12286);
nand U13056 (N_13056,N_12190,N_12104);
nand U13057 (N_13057,N_12083,N_12223);
xor U13058 (N_13058,N_12419,N_12015);
and U13059 (N_13059,N_12117,N_12468);
xnor U13060 (N_13060,N_12380,N_12437);
or U13061 (N_13061,N_12214,N_11875);
and U13062 (N_13062,N_12238,N_12478);
nor U13063 (N_13063,N_11974,N_12328);
or U13064 (N_13064,N_12325,N_12213);
nand U13065 (N_13065,N_12196,N_12015);
nand U13066 (N_13066,N_11908,N_12289);
and U13067 (N_13067,N_12388,N_12176);
xnor U13068 (N_13068,N_11934,N_12042);
or U13069 (N_13069,N_12100,N_12205);
and U13070 (N_13070,N_12286,N_12368);
nand U13071 (N_13071,N_12480,N_11957);
and U13072 (N_13072,N_12487,N_12372);
xor U13073 (N_13073,N_11962,N_12176);
xnor U13074 (N_13074,N_12249,N_12376);
xor U13075 (N_13075,N_11921,N_12372);
nor U13076 (N_13076,N_12130,N_12023);
nand U13077 (N_13077,N_12062,N_11926);
xnor U13078 (N_13078,N_12474,N_12478);
and U13079 (N_13079,N_11967,N_12303);
xnor U13080 (N_13080,N_12363,N_12152);
nor U13081 (N_13081,N_12266,N_12002);
nor U13082 (N_13082,N_12392,N_12464);
nor U13083 (N_13083,N_12399,N_12488);
xnor U13084 (N_13084,N_12087,N_12050);
nor U13085 (N_13085,N_12284,N_12165);
or U13086 (N_13086,N_12199,N_12337);
nand U13087 (N_13087,N_12205,N_12145);
nor U13088 (N_13088,N_12437,N_12485);
nand U13089 (N_13089,N_12348,N_12031);
nand U13090 (N_13090,N_11912,N_11916);
nor U13091 (N_13091,N_12393,N_12406);
xnor U13092 (N_13092,N_12000,N_12491);
or U13093 (N_13093,N_12236,N_12254);
or U13094 (N_13094,N_12031,N_12476);
nor U13095 (N_13095,N_12185,N_12216);
nand U13096 (N_13096,N_12475,N_12299);
and U13097 (N_13097,N_12035,N_11940);
xnor U13098 (N_13098,N_12358,N_12121);
and U13099 (N_13099,N_12025,N_12499);
xnor U13100 (N_13100,N_12170,N_12271);
and U13101 (N_13101,N_12252,N_12427);
nand U13102 (N_13102,N_12337,N_12235);
nand U13103 (N_13103,N_12161,N_12443);
nor U13104 (N_13104,N_12204,N_12293);
or U13105 (N_13105,N_12473,N_12128);
and U13106 (N_13106,N_12129,N_12432);
or U13107 (N_13107,N_11953,N_12206);
nand U13108 (N_13108,N_12333,N_12099);
nand U13109 (N_13109,N_11883,N_12218);
and U13110 (N_13110,N_12292,N_12390);
nor U13111 (N_13111,N_12293,N_12363);
and U13112 (N_13112,N_12151,N_12083);
or U13113 (N_13113,N_11928,N_11910);
nor U13114 (N_13114,N_12039,N_12116);
or U13115 (N_13115,N_12492,N_12408);
and U13116 (N_13116,N_12452,N_11884);
nand U13117 (N_13117,N_12368,N_12389);
xor U13118 (N_13118,N_12435,N_11893);
or U13119 (N_13119,N_11883,N_11901);
nand U13120 (N_13120,N_12305,N_12085);
nand U13121 (N_13121,N_12076,N_12365);
or U13122 (N_13122,N_12379,N_12080);
nor U13123 (N_13123,N_12182,N_11903);
xor U13124 (N_13124,N_12379,N_12068);
and U13125 (N_13125,N_12996,N_12647);
xnor U13126 (N_13126,N_13060,N_12706);
nor U13127 (N_13127,N_12838,N_12762);
nor U13128 (N_13128,N_12746,N_12726);
and U13129 (N_13129,N_12504,N_12569);
or U13130 (N_13130,N_12781,N_12829);
and U13131 (N_13131,N_12512,N_12533);
nand U13132 (N_13132,N_13048,N_12947);
nand U13133 (N_13133,N_12670,N_12946);
xor U13134 (N_13134,N_12652,N_13067);
or U13135 (N_13135,N_13062,N_13011);
nand U13136 (N_13136,N_13002,N_13025);
nand U13137 (N_13137,N_12925,N_12978);
or U13138 (N_13138,N_13096,N_12803);
nor U13139 (N_13139,N_13109,N_12683);
or U13140 (N_13140,N_13049,N_12539);
or U13141 (N_13141,N_12842,N_12780);
and U13142 (N_13142,N_12753,N_12974);
xor U13143 (N_13143,N_12547,N_12676);
xor U13144 (N_13144,N_12735,N_12855);
and U13145 (N_13145,N_12963,N_12743);
nor U13146 (N_13146,N_12699,N_12568);
xnor U13147 (N_13147,N_12987,N_13115);
xnor U13148 (N_13148,N_12961,N_13070);
nand U13149 (N_13149,N_12942,N_12562);
xor U13150 (N_13150,N_12542,N_12815);
nand U13151 (N_13151,N_12975,N_12894);
and U13152 (N_13152,N_12649,N_12601);
nor U13153 (N_13153,N_12953,N_12864);
or U13154 (N_13154,N_13009,N_12638);
nand U13155 (N_13155,N_12993,N_12981);
nor U13156 (N_13156,N_13050,N_13086);
nand U13157 (N_13157,N_12879,N_12725);
or U13158 (N_13158,N_12596,N_12966);
nor U13159 (N_13159,N_12761,N_12692);
nor U13160 (N_13160,N_12721,N_12710);
and U13161 (N_13161,N_12916,N_13065);
nand U13162 (N_13162,N_12932,N_12639);
and U13163 (N_13163,N_12679,N_12592);
nor U13164 (N_13164,N_12962,N_12728);
nor U13165 (N_13165,N_12874,N_13039);
xnor U13166 (N_13166,N_12723,N_13121);
or U13167 (N_13167,N_12612,N_12671);
or U13168 (N_13168,N_12703,N_13092);
nand U13169 (N_13169,N_12826,N_12570);
xor U13170 (N_13170,N_12605,N_13089);
and U13171 (N_13171,N_12702,N_12905);
nand U13172 (N_13172,N_12816,N_12663);
and U13173 (N_13173,N_12715,N_12920);
nor U13174 (N_13174,N_12989,N_12903);
nand U13175 (N_13175,N_12907,N_13035);
and U13176 (N_13176,N_12790,N_12621);
and U13177 (N_13177,N_12581,N_12675);
or U13178 (N_13178,N_12766,N_12866);
nand U13179 (N_13179,N_12640,N_12751);
and U13180 (N_13180,N_12629,N_13090);
xor U13181 (N_13181,N_12731,N_12552);
nor U13182 (N_13182,N_12856,N_12834);
and U13183 (N_13183,N_12757,N_12736);
nand U13184 (N_13184,N_12549,N_12811);
or U13185 (N_13185,N_12930,N_12954);
nand U13186 (N_13186,N_13017,N_12783);
and U13187 (N_13187,N_13029,N_12602);
and U13188 (N_13188,N_13008,N_12580);
nor U13189 (N_13189,N_12599,N_12887);
and U13190 (N_13190,N_12984,N_12525);
nor U13191 (N_13191,N_12796,N_13069);
nor U13192 (N_13192,N_12818,N_12955);
nand U13193 (N_13193,N_13117,N_12660);
nand U13194 (N_13194,N_12899,N_13031);
or U13195 (N_13195,N_12538,N_12734);
nor U13196 (N_13196,N_12840,N_13053);
nand U13197 (N_13197,N_12574,N_13122);
nor U13198 (N_13198,N_12886,N_12729);
xor U13199 (N_13199,N_13023,N_12997);
nor U13200 (N_13200,N_13010,N_12541);
and U13201 (N_13201,N_12852,N_13005);
xor U13202 (N_13202,N_12982,N_12802);
or U13203 (N_13203,N_12686,N_12906);
and U13204 (N_13204,N_12998,N_12794);
or U13205 (N_13205,N_13123,N_12738);
xnor U13206 (N_13206,N_12784,N_12832);
and U13207 (N_13207,N_12850,N_12551);
nand U13208 (N_13208,N_12940,N_13093);
xor U13209 (N_13209,N_12884,N_13038);
and U13210 (N_13210,N_12511,N_13037);
nand U13211 (N_13211,N_12559,N_13058);
nor U13212 (N_13212,N_12968,N_12651);
nand U13213 (N_13213,N_12583,N_12587);
and U13214 (N_13214,N_12824,N_12633);
xnor U13215 (N_13215,N_12666,N_12988);
xnor U13216 (N_13216,N_13059,N_12754);
nor U13217 (N_13217,N_12617,N_12804);
nor U13218 (N_13218,N_12656,N_13064);
nand U13219 (N_13219,N_12584,N_12682);
xor U13220 (N_13220,N_13057,N_13105);
or U13221 (N_13221,N_12926,N_13052);
xnor U13222 (N_13222,N_13013,N_12880);
or U13223 (N_13223,N_12892,N_12820);
nor U13224 (N_13224,N_12724,N_12708);
xor U13225 (N_13225,N_12582,N_12673);
nor U13226 (N_13226,N_12876,N_12586);
and U13227 (N_13227,N_12748,N_12716);
nor U13228 (N_13228,N_12898,N_12520);
nor U13229 (N_13229,N_13019,N_12878);
or U13230 (N_13230,N_12732,N_12752);
nor U13231 (N_13231,N_12608,N_12910);
nor U13232 (N_13232,N_13006,N_12756);
and U13233 (N_13233,N_12566,N_12628);
and U13234 (N_13234,N_13055,N_12972);
xnor U13235 (N_13235,N_12677,N_12604);
or U13236 (N_13236,N_12741,N_13020);
or U13237 (N_13237,N_12807,N_13102);
and U13238 (N_13238,N_12700,N_12970);
and U13239 (N_13239,N_12529,N_12672);
and U13240 (N_13240,N_12645,N_12825);
xor U13241 (N_13241,N_12923,N_13026);
and U13242 (N_13242,N_12623,N_12994);
nor U13243 (N_13243,N_12918,N_13012);
and U13244 (N_13244,N_12848,N_12661);
nor U13245 (N_13245,N_12875,N_12691);
nand U13246 (N_13246,N_13077,N_12607);
nor U13247 (N_13247,N_12793,N_12759);
nand U13248 (N_13248,N_12517,N_12833);
or U13249 (N_13249,N_13108,N_12775);
and U13250 (N_13250,N_12631,N_12870);
and U13251 (N_13251,N_12610,N_12507);
nand U13252 (N_13252,N_12544,N_12615);
nand U13253 (N_13253,N_12573,N_12701);
xor U13254 (N_13254,N_12619,N_12983);
xor U13255 (N_13255,N_12977,N_12719);
nor U13256 (N_13256,N_12814,N_12801);
nor U13257 (N_13257,N_12618,N_12653);
and U13258 (N_13258,N_12915,N_12969);
xnor U13259 (N_13259,N_13097,N_13068);
or U13260 (N_13260,N_12516,N_12554);
nor U13261 (N_13261,N_12534,N_12792);
xor U13262 (N_13262,N_12717,N_12749);
and U13263 (N_13263,N_12755,N_12556);
nor U13264 (N_13264,N_12819,N_12873);
xnor U13265 (N_13265,N_12821,N_12854);
xnor U13266 (N_13266,N_12967,N_12900);
or U13267 (N_13267,N_13061,N_12658);
xor U13268 (N_13268,N_12822,N_12914);
or U13269 (N_13269,N_12847,N_12561);
or U13270 (N_13270,N_13094,N_12941);
nand U13271 (N_13271,N_13083,N_12800);
nor U13272 (N_13272,N_12540,N_13000);
nand U13273 (N_13273,N_13074,N_13099);
nor U13274 (N_13274,N_12797,N_12558);
or U13275 (N_13275,N_12785,N_12613);
nand U13276 (N_13276,N_12659,N_12768);
or U13277 (N_13277,N_12908,N_12902);
and U13278 (N_13278,N_12722,N_13032);
nand U13279 (N_13279,N_12585,N_12509);
nor U13280 (N_13280,N_12626,N_12789);
and U13281 (N_13281,N_13040,N_12883);
nand U13282 (N_13282,N_12553,N_12503);
xnor U13283 (N_13283,N_12634,N_12944);
nor U13284 (N_13284,N_13041,N_13043);
xnor U13285 (N_13285,N_12861,N_12571);
nand U13286 (N_13286,N_13116,N_12664);
and U13287 (N_13287,N_12519,N_12575);
xor U13288 (N_13288,N_12560,N_12705);
and U13289 (N_13289,N_12846,N_12857);
and U13290 (N_13290,N_12805,N_12830);
and U13291 (N_13291,N_12839,N_12665);
nor U13292 (N_13292,N_12745,N_12841);
and U13293 (N_13293,N_12588,N_13001);
xnor U13294 (N_13294,N_12537,N_12893);
or U13295 (N_13295,N_12860,N_12550);
nor U13296 (N_13296,N_12798,N_12808);
or U13297 (N_13297,N_12648,N_12545);
or U13298 (N_13298,N_12791,N_12636);
xnor U13299 (N_13299,N_12637,N_12685);
or U13300 (N_13300,N_12885,N_12505);
or U13301 (N_13301,N_13075,N_12718);
and U13302 (N_13302,N_12952,N_13046);
and U13303 (N_13303,N_13007,N_12630);
xnor U13304 (N_13304,N_12526,N_12956);
or U13305 (N_13305,N_12865,N_13063);
and U13306 (N_13306,N_12991,N_13016);
and U13307 (N_13307,N_12933,N_12971);
and U13308 (N_13308,N_12597,N_12712);
xor U13309 (N_13309,N_12868,N_12888);
xnor U13310 (N_13310,N_12958,N_12578);
nand U13311 (N_13311,N_12711,N_13051);
xnor U13312 (N_13312,N_13054,N_12555);
or U13313 (N_13313,N_12843,N_12845);
or U13314 (N_13314,N_12782,N_12622);
nor U13315 (N_13315,N_12823,N_12591);
xor U13316 (N_13316,N_12849,N_12973);
and U13317 (N_13317,N_12799,N_13022);
xor U13318 (N_13318,N_12787,N_13024);
nor U13319 (N_13319,N_12546,N_12641);
or U13320 (N_13320,N_12646,N_12851);
nor U13321 (N_13321,N_12837,N_12684);
xor U13322 (N_13322,N_12606,N_12779);
or U13323 (N_13323,N_12502,N_12901);
and U13324 (N_13324,N_13106,N_13066);
nand U13325 (N_13325,N_12867,N_12812);
xor U13326 (N_13326,N_12891,N_12727);
nor U13327 (N_13327,N_12620,N_12853);
xor U13328 (N_13328,N_12928,N_12935);
nor U13329 (N_13329,N_12943,N_13095);
and U13330 (N_13330,N_12871,N_12770);
nand U13331 (N_13331,N_12750,N_13056);
and U13332 (N_13332,N_12657,N_12508);
xnor U13333 (N_13333,N_12668,N_12603);
xor U13334 (N_13334,N_12938,N_12609);
xnor U13335 (N_13335,N_12774,N_12600);
or U13336 (N_13336,N_12698,N_12862);
nand U13337 (N_13337,N_12614,N_12616);
or U13338 (N_13338,N_13047,N_12939);
and U13339 (N_13339,N_12523,N_12912);
and U13340 (N_13340,N_12598,N_12536);
nor U13341 (N_13341,N_12521,N_12522);
nor U13342 (N_13342,N_12742,N_12689);
nand U13343 (N_13343,N_12627,N_13045);
xnor U13344 (N_13344,N_12828,N_12709);
xor U13345 (N_13345,N_12650,N_12590);
nand U13346 (N_13346,N_12810,N_12773);
nor U13347 (N_13347,N_12931,N_12913);
and U13348 (N_13348,N_12949,N_12758);
nor U13349 (N_13349,N_12909,N_12514);
xnor U13350 (N_13350,N_13044,N_12524);
nand U13351 (N_13351,N_12662,N_13103);
nor U13352 (N_13352,N_12795,N_12625);
nor U13353 (N_13353,N_12957,N_12872);
nor U13354 (N_13354,N_13027,N_12714);
nand U13355 (N_13355,N_12747,N_12720);
nor U13356 (N_13356,N_12593,N_13104);
and U13357 (N_13357,N_12567,N_12895);
nand U13358 (N_13358,N_12869,N_12889);
or U13359 (N_13359,N_12506,N_12979);
nor U13360 (N_13360,N_13003,N_13073);
or U13361 (N_13361,N_12632,N_12681);
or U13362 (N_13362,N_12786,N_12528);
nor U13363 (N_13363,N_12986,N_12992);
nand U13364 (N_13364,N_12817,N_12595);
nand U13365 (N_13365,N_12548,N_12744);
nor U13366 (N_13366,N_12579,N_13124);
and U13367 (N_13367,N_12730,N_13004);
and U13368 (N_13368,N_13112,N_12896);
and U13369 (N_13369,N_12919,N_12576);
or U13370 (N_13370,N_12844,N_12788);
nor U13371 (N_13371,N_13113,N_13091);
xnor U13372 (N_13372,N_12642,N_13080);
or U13373 (N_13373,N_12929,N_12624);
or U13374 (N_13374,N_12733,N_12964);
xnor U13375 (N_13375,N_12927,N_13018);
and U13376 (N_13376,N_12863,N_12543);
nor U13377 (N_13377,N_12767,N_12501);
xnor U13378 (N_13378,N_12980,N_12688);
and U13379 (N_13379,N_12760,N_12960);
nor U13380 (N_13380,N_12881,N_13111);
nor U13381 (N_13381,N_13082,N_13101);
nand U13382 (N_13382,N_12577,N_13072);
nand U13383 (N_13383,N_12531,N_12589);
and U13384 (N_13384,N_13098,N_12937);
nand U13385 (N_13385,N_12674,N_12687);
nand U13386 (N_13386,N_12765,N_12999);
xnor U13387 (N_13387,N_12917,N_13015);
or U13388 (N_13388,N_12936,N_12835);
nand U13389 (N_13389,N_12611,N_12769);
or U13390 (N_13390,N_12518,N_12704);
xnor U13391 (N_13391,N_12667,N_12776);
xnor U13392 (N_13392,N_13120,N_12921);
and U13393 (N_13393,N_12763,N_12922);
nor U13394 (N_13394,N_13036,N_12530);
xor U13395 (N_13395,N_12959,N_12680);
and U13396 (N_13396,N_12924,N_13085);
and U13397 (N_13397,N_12911,N_12965);
xnor U13398 (N_13398,N_12945,N_13078);
xnor U13399 (N_13399,N_12513,N_12563);
and U13400 (N_13400,N_12693,N_12890);
xnor U13401 (N_13401,N_13100,N_12515);
xnor U13402 (N_13402,N_13028,N_12655);
nand U13403 (N_13403,N_12565,N_12713);
and U13404 (N_13404,N_12535,N_12644);
and U13405 (N_13405,N_12806,N_12985);
nor U13406 (N_13406,N_13087,N_12897);
or U13407 (N_13407,N_13076,N_12831);
nand U13408 (N_13408,N_12500,N_12696);
nand U13409 (N_13409,N_12904,N_12859);
or U13410 (N_13410,N_13030,N_12778);
and U13411 (N_13411,N_12695,N_12527);
and U13412 (N_13412,N_12557,N_12858);
xor U13413 (N_13413,N_12532,N_12690);
xor U13414 (N_13414,N_12740,N_12697);
nand U13415 (N_13415,N_12813,N_13079);
nand U13416 (N_13416,N_13071,N_13107);
xnor U13417 (N_13417,N_12882,N_12877);
nand U13418 (N_13418,N_13021,N_12771);
nand U13419 (N_13419,N_13110,N_12995);
nor U13420 (N_13420,N_12654,N_13042);
and U13421 (N_13421,N_13119,N_13084);
and U13422 (N_13422,N_12951,N_12739);
and U13423 (N_13423,N_12934,N_12572);
and U13424 (N_13424,N_13114,N_12827);
and U13425 (N_13425,N_12948,N_13014);
nor U13426 (N_13426,N_13088,N_12737);
and U13427 (N_13427,N_12772,N_13118);
nor U13428 (N_13428,N_12564,N_12694);
or U13429 (N_13429,N_12809,N_12777);
nand U13430 (N_13430,N_12643,N_12678);
nand U13431 (N_13431,N_12510,N_12950);
nand U13432 (N_13432,N_12976,N_12635);
and U13433 (N_13433,N_13081,N_13034);
xnor U13434 (N_13434,N_12836,N_12594);
or U13435 (N_13435,N_13033,N_12990);
and U13436 (N_13436,N_12669,N_12707);
xnor U13437 (N_13437,N_12764,N_12622);
nand U13438 (N_13438,N_12574,N_12920);
or U13439 (N_13439,N_12898,N_12654);
and U13440 (N_13440,N_12911,N_12758);
nand U13441 (N_13441,N_12977,N_12765);
xor U13442 (N_13442,N_13030,N_12669);
nand U13443 (N_13443,N_12759,N_13111);
or U13444 (N_13444,N_12934,N_12721);
nor U13445 (N_13445,N_12933,N_12934);
nor U13446 (N_13446,N_12680,N_12757);
and U13447 (N_13447,N_12810,N_12893);
nand U13448 (N_13448,N_12826,N_12934);
or U13449 (N_13449,N_12901,N_12643);
nor U13450 (N_13450,N_12747,N_12699);
and U13451 (N_13451,N_12588,N_13050);
nor U13452 (N_13452,N_12990,N_13094);
nor U13453 (N_13453,N_12810,N_12520);
xnor U13454 (N_13454,N_12541,N_12869);
nor U13455 (N_13455,N_13006,N_12828);
nor U13456 (N_13456,N_12844,N_12968);
xor U13457 (N_13457,N_13059,N_12610);
or U13458 (N_13458,N_13011,N_12830);
nor U13459 (N_13459,N_12537,N_13016);
nand U13460 (N_13460,N_12623,N_12983);
and U13461 (N_13461,N_12599,N_12831);
nand U13462 (N_13462,N_12701,N_12923);
nand U13463 (N_13463,N_13042,N_12596);
nand U13464 (N_13464,N_13014,N_12558);
or U13465 (N_13465,N_12910,N_13083);
or U13466 (N_13466,N_12707,N_12686);
and U13467 (N_13467,N_12596,N_13047);
xnor U13468 (N_13468,N_12766,N_12847);
nand U13469 (N_13469,N_12649,N_12550);
xor U13470 (N_13470,N_12888,N_12595);
nor U13471 (N_13471,N_13088,N_13122);
or U13472 (N_13472,N_12656,N_12627);
or U13473 (N_13473,N_12730,N_12687);
nor U13474 (N_13474,N_12620,N_13072);
or U13475 (N_13475,N_12775,N_13030);
and U13476 (N_13476,N_12667,N_12635);
or U13477 (N_13477,N_12766,N_12765);
xor U13478 (N_13478,N_12800,N_12767);
nand U13479 (N_13479,N_12818,N_12561);
xnor U13480 (N_13480,N_12612,N_12501);
nor U13481 (N_13481,N_12990,N_12911);
nor U13482 (N_13482,N_12666,N_13070);
nor U13483 (N_13483,N_12709,N_12576);
xor U13484 (N_13484,N_12856,N_12840);
xnor U13485 (N_13485,N_12626,N_12991);
nand U13486 (N_13486,N_13065,N_12828);
nand U13487 (N_13487,N_12911,N_12519);
or U13488 (N_13488,N_12687,N_13072);
or U13489 (N_13489,N_12706,N_12606);
nor U13490 (N_13490,N_12869,N_12815);
nand U13491 (N_13491,N_12656,N_12605);
nor U13492 (N_13492,N_13040,N_12915);
xnor U13493 (N_13493,N_13110,N_12730);
or U13494 (N_13494,N_12690,N_12708);
nand U13495 (N_13495,N_12738,N_13019);
nand U13496 (N_13496,N_12528,N_13050);
or U13497 (N_13497,N_12958,N_12830);
nor U13498 (N_13498,N_12547,N_13085);
nand U13499 (N_13499,N_12785,N_13059);
xnor U13500 (N_13500,N_12794,N_12771);
or U13501 (N_13501,N_13080,N_12506);
and U13502 (N_13502,N_12823,N_12875);
nor U13503 (N_13503,N_12876,N_12822);
xor U13504 (N_13504,N_12645,N_12507);
and U13505 (N_13505,N_12971,N_13063);
or U13506 (N_13506,N_12782,N_12718);
xor U13507 (N_13507,N_12819,N_12955);
nor U13508 (N_13508,N_12505,N_13007);
nor U13509 (N_13509,N_12620,N_12696);
xor U13510 (N_13510,N_12921,N_13002);
or U13511 (N_13511,N_12640,N_13013);
nor U13512 (N_13512,N_12924,N_12952);
xnor U13513 (N_13513,N_12961,N_12655);
nand U13514 (N_13514,N_13020,N_13009);
xnor U13515 (N_13515,N_12917,N_13062);
and U13516 (N_13516,N_13044,N_12734);
and U13517 (N_13517,N_13091,N_12530);
nor U13518 (N_13518,N_12774,N_12520);
nor U13519 (N_13519,N_12904,N_13124);
or U13520 (N_13520,N_12834,N_12832);
nor U13521 (N_13521,N_13090,N_13124);
xor U13522 (N_13522,N_12915,N_12896);
nand U13523 (N_13523,N_12919,N_12835);
xnor U13524 (N_13524,N_13006,N_12819);
nor U13525 (N_13525,N_12607,N_12761);
nor U13526 (N_13526,N_13023,N_12543);
nor U13527 (N_13527,N_12502,N_12516);
and U13528 (N_13528,N_12670,N_12970);
and U13529 (N_13529,N_12682,N_12962);
and U13530 (N_13530,N_12579,N_13069);
nor U13531 (N_13531,N_12735,N_12960);
xor U13532 (N_13532,N_12815,N_12602);
nand U13533 (N_13533,N_12562,N_12539);
nand U13534 (N_13534,N_13113,N_12865);
nand U13535 (N_13535,N_12889,N_12921);
and U13536 (N_13536,N_12519,N_12760);
and U13537 (N_13537,N_12701,N_12700);
xnor U13538 (N_13538,N_13075,N_12881);
and U13539 (N_13539,N_12565,N_12582);
xnor U13540 (N_13540,N_12656,N_12898);
or U13541 (N_13541,N_12887,N_12575);
nor U13542 (N_13542,N_12615,N_12529);
or U13543 (N_13543,N_12658,N_12955);
and U13544 (N_13544,N_12908,N_12927);
and U13545 (N_13545,N_12505,N_12834);
xnor U13546 (N_13546,N_12578,N_12740);
or U13547 (N_13547,N_12705,N_12916);
and U13548 (N_13548,N_12942,N_12916);
and U13549 (N_13549,N_13069,N_12765);
nand U13550 (N_13550,N_13075,N_13017);
nor U13551 (N_13551,N_13123,N_13122);
and U13552 (N_13552,N_12954,N_12723);
nor U13553 (N_13553,N_13041,N_13048);
nor U13554 (N_13554,N_12854,N_12901);
xor U13555 (N_13555,N_12777,N_12989);
and U13556 (N_13556,N_13101,N_12730);
nor U13557 (N_13557,N_12724,N_13064);
xnor U13558 (N_13558,N_12637,N_13067);
nor U13559 (N_13559,N_12779,N_13053);
or U13560 (N_13560,N_13051,N_13104);
xor U13561 (N_13561,N_12793,N_12944);
or U13562 (N_13562,N_12792,N_12972);
xor U13563 (N_13563,N_12876,N_12710);
xnor U13564 (N_13564,N_12871,N_12743);
nand U13565 (N_13565,N_12759,N_12504);
nor U13566 (N_13566,N_13116,N_12797);
and U13567 (N_13567,N_13113,N_12665);
or U13568 (N_13568,N_12997,N_13091);
and U13569 (N_13569,N_12552,N_12874);
nor U13570 (N_13570,N_12746,N_12704);
or U13571 (N_13571,N_12897,N_12998);
nand U13572 (N_13572,N_12739,N_12864);
nand U13573 (N_13573,N_12508,N_12785);
nand U13574 (N_13574,N_12995,N_12535);
and U13575 (N_13575,N_12954,N_12603);
nor U13576 (N_13576,N_13038,N_12535);
and U13577 (N_13577,N_13123,N_12923);
nand U13578 (N_13578,N_13026,N_12603);
or U13579 (N_13579,N_13041,N_13046);
or U13580 (N_13580,N_12579,N_12556);
xor U13581 (N_13581,N_12532,N_12941);
or U13582 (N_13582,N_12577,N_12601);
or U13583 (N_13583,N_12867,N_13073);
and U13584 (N_13584,N_13052,N_12951);
nor U13585 (N_13585,N_12523,N_12539);
and U13586 (N_13586,N_12894,N_12974);
or U13587 (N_13587,N_13062,N_12807);
and U13588 (N_13588,N_13109,N_12621);
nor U13589 (N_13589,N_12693,N_12613);
and U13590 (N_13590,N_12518,N_12732);
and U13591 (N_13591,N_13103,N_12504);
nor U13592 (N_13592,N_12740,N_12897);
and U13593 (N_13593,N_13099,N_12502);
nand U13594 (N_13594,N_12837,N_13020);
nor U13595 (N_13595,N_12939,N_13088);
nor U13596 (N_13596,N_12802,N_12667);
and U13597 (N_13597,N_13032,N_13073);
nand U13598 (N_13598,N_12804,N_12815);
or U13599 (N_13599,N_12616,N_12856);
or U13600 (N_13600,N_12938,N_12759);
or U13601 (N_13601,N_12652,N_12814);
nor U13602 (N_13602,N_12984,N_12996);
and U13603 (N_13603,N_12739,N_12907);
or U13604 (N_13604,N_13019,N_12766);
and U13605 (N_13605,N_12865,N_12759);
xnor U13606 (N_13606,N_12614,N_12619);
nor U13607 (N_13607,N_12748,N_13049);
nor U13608 (N_13608,N_12595,N_12799);
nand U13609 (N_13609,N_12524,N_12761);
nand U13610 (N_13610,N_12740,N_12743);
xor U13611 (N_13611,N_12720,N_12614);
nand U13612 (N_13612,N_12513,N_12841);
and U13613 (N_13613,N_12795,N_13123);
or U13614 (N_13614,N_12887,N_12510);
xnor U13615 (N_13615,N_12968,N_13061);
nor U13616 (N_13616,N_12683,N_12698);
or U13617 (N_13617,N_12999,N_12525);
or U13618 (N_13618,N_12850,N_12669);
or U13619 (N_13619,N_12819,N_12910);
or U13620 (N_13620,N_12820,N_12540);
and U13621 (N_13621,N_12800,N_13009);
nor U13622 (N_13622,N_13095,N_12694);
and U13623 (N_13623,N_12810,N_12626);
xnor U13624 (N_13624,N_12956,N_12651);
and U13625 (N_13625,N_12831,N_13067);
or U13626 (N_13626,N_12652,N_13084);
xnor U13627 (N_13627,N_12944,N_12838);
or U13628 (N_13628,N_12905,N_12543);
xor U13629 (N_13629,N_12842,N_12985);
or U13630 (N_13630,N_12562,N_12535);
or U13631 (N_13631,N_12826,N_12552);
nor U13632 (N_13632,N_13106,N_12756);
and U13633 (N_13633,N_12802,N_12920);
xnor U13634 (N_13634,N_13114,N_12878);
xor U13635 (N_13635,N_12787,N_12628);
xnor U13636 (N_13636,N_12543,N_12592);
xnor U13637 (N_13637,N_12774,N_12832);
nor U13638 (N_13638,N_12855,N_12552);
or U13639 (N_13639,N_12549,N_12574);
nor U13640 (N_13640,N_12723,N_12702);
or U13641 (N_13641,N_12732,N_12991);
and U13642 (N_13642,N_12924,N_12731);
xor U13643 (N_13643,N_12862,N_12932);
xnor U13644 (N_13644,N_12861,N_12505);
nor U13645 (N_13645,N_12554,N_12511);
nor U13646 (N_13646,N_12637,N_12734);
and U13647 (N_13647,N_12543,N_12797);
or U13648 (N_13648,N_12588,N_12990);
nor U13649 (N_13649,N_13081,N_13076);
or U13650 (N_13650,N_12513,N_12537);
nor U13651 (N_13651,N_12589,N_12567);
nand U13652 (N_13652,N_12586,N_12833);
xor U13653 (N_13653,N_12591,N_12951);
or U13654 (N_13654,N_12882,N_13083);
nor U13655 (N_13655,N_12834,N_12879);
xor U13656 (N_13656,N_13059,N_12717);
nand U13657 (N_13657,N_12930,N_12960);
nand U13658 (N_13658,N_12596,N_12895);
nand U13659 (N_13659,N_12828,N_12624);
and U13660 (N_13660,N_12838,N_13124);
nor U13661 (N_13661,N_12636,N_12533);
nand U13662 (N_13662,N_12696,N_12788);
nor U13663 (N_13663,N_12694,N_12820);
xnor U13664 (N_13664,N_12848,N_12517);
xor U13665 (N_13665,N_13037,N_12662);
or U13666 (N_13666,N_12735,N_12796);
or U13667 (N_13667,N_12561,N_12539);
nand U13668 (N_13668,N_12632,N_12706);
nand U13669 (N_13669,N_13116,N_13107);
nand U13670 (N_13670,N_12650,N_12527);
or U13671 (N_13671,N_12569,N_12752);
nor U13672 (N_13672,N_12835,N_12826);
xnor U13673 (N_13673,N_12825,N_12906);
nand U13674 (N_13674,N_12710,N_13118);
xor U13675 (N_13675,N_12716,N_12732);
nor U13676 (N_13676,N_12830,N_12712);
or U13677 (N_13677,N_12918,N_12765);
and U13678 (N_13678,N_12803,N_12881);
nand U13679 (N_13679,N_12781,N_13060);
nand U13680 (N_13680,N_12681,N_12601);
nand U13681 (N_13681,N_12729,N_12995);
xnor U13682 (N_13682,N_12978,N_12591);
nor U13683 (N_13683,N_13073,N_12903);
nand U13684 (N_13684,N_12559,N_12840);
xor U13685 (N_13685,N_12865,N_12524);
nor U13686 (N_13686,N_12634,N_12751);
xnor U13687 (N_13687,N_12979,N_12958);
and U13688 (N_13688,N_12767,N_13074);
or U13689 (N_13689,N_12985,N_12536);
xor U13690 (N_13690,N_12839,N_13075);
nor U13691 (N_13691,N_12953,N_12628);
or U13692 (N_13692,N_12566,N_12956);
and U13693 (N_13693,N_12742,N_12569);
nor U13694 (N_13694,N_12936,N_12880);
or U13695 (N_13695,N_13118,N_12844);
or U13696 (N_13696,N_12937,N_12737);
or U13697 (N_13697,N_12781,N_12789);
or U13698 (N_13698,N_12565,N_12721);
or U13699 (N_13699,N_12719,N_13060);
nor U13700 (N_13700,N_13048,N_12928);
and U13701 (N_13701,N_12835,N_12650);
nor U13702 (N_13702,N_12873,N_12642);
xor U13703 (N_13703,N_12810,N_13053);
xnor U13704 (N_13704,N_12871,N_12648);
nor U13705 (N_13705,N_12773,N_12925);
and U13706 (N_13706,N_12686,N_12895);
or U13707 (N_13707,N_12607,N_12941);
or U13708 (N_13708,N_12737,N_13026);
nand U13709 (N_13709,N_12500,N_13030);
nand U13710 (N_13710,N_12604,N_13012);
and U13711 (N_13711,N_12555,N_12651);
or U13712 (N_13712,N_12624,N_12714);
xnor U13713 (N_13713,N_12584,N_12837);
and U13714 (N_13714,N_12664,N_13041);
nand U13715 (N_13715,N_12905,N_12642);
nor U13716 (N_13716,N_12948,N_12753);
or U13717 (N_13717,N_12505,N_12868);
and U13718 (N_13718,N_12865,N_12632);
and U13719 (N_13719,N_12882,N_12961);
nor U13720 (N_13720,N_13039,N_12640);
nand U13721 (N_13721,N_12977,N_12907);
and U13722 (N_13722,N_12588,N_12552);
or U13723 (N_13723,N_12739,N_12576);
xnor U13724 (N_13724,N_12790,N_12716);
nand U13725 (N_13725,N_12787,N_12647);
xnor U13726 (N_13726,N_12701,N_12865);
or U13727 (N_13727,N_13017,N_13046);
nand U13728 (N_13728,N_12811,N_12832);
and U13729 (N_13729,N_12936,N_12875);
and U13730 (N_13730,N_12985,N_12742);
nor U13731 (N_13731,N_12680,N_12835);
xor U13732 (N_13732,N_12947,N_12505);
xor U13733 (N_13733,N_12807,N_12969);
and U13734 (N_13734,N_12750,N_12839);
or U13735 (N_13735,N_12612,N_12993);
nand U13736 (N_13736,N_12685,N_13094);
xor U13737 (N_13737,N_12802,N_13047);
or U13738 (N_13738,N_12726,N_12799);
nand U13739 (N_13739,N_12758,N_13117);
and U13740 (N_13740,N_12604,N_12949);
xor U13741 (N_13741,N_12970,N_12829);
nand U13742 (N_13742,N_13025,N_12970);
nand U13743 (N_13743,N_12730,N_12858);
and U13744 (N_13744,N_12664,N_12657);
and U13745 (N_13745,N_12902,N_12895);
nor U13746 (N_13746,N_12998,N_12712);
nand U13747 (N_13747,N_12810,N_13068);
nor U13748 (N_13748,N_13087,N_12918);
xor U13749 (N_13749,N_12552,N_13034);
and U13750 (N_13750,N_13606,N_13273);
or U13751 (N_13751,N_13535,N_13743);
nand U13752 (N_13752,N_13192,N_13169);
nand U13753 (N_13753,N_13187,N_13496);
xor U13754 (N_13754,N_13504,N_13387);
nand U13755 (N_13755,N_13695,N_13141);
and U13756 (N_13756,N_13623,N_13545);
nand U13757 (N_13757,N_13225,N_13585);
xnor U13758 (N_13758,N_13488,N_13170);
xnor U13759 (N_13759,N_13566,N_13221);
nand U13760 (N_13760,N_13349,N_13228);
xor U13761 (N_13761,N_13309,N_13322);
nor U13762 (N_13762,N_13211,N_13474);
and U13763 (N_13763,N_13492,N_13138);
nor U13764 (N_13764,N_13625,N_13583);
and U13765 (N_13765,N_13346,N_13411);
xor U13766 (N_13766,N_13718,N_13588);
xnor U13767 (N_13767,N_13604,N_13708);
nor U13768 (N_13768,N_13540,N_13638);
nor U13769 (N_13769,N_13136,N_13125);
and U13770 (N_13770,N_13392,N_13373);
xor U13771 (N_13771,N_13272,N_13716);
nand U13772 (N_13772,N_13577,N_13439);
or U13773 (N_13773,N_13325,N_13723);
or U13774 (N_13774,N_13151,N_13436);
nor U13775 (N_13775,N_13455,N_13527);
nor U13776 (N_13776,N_13135,N_13269);
nor U13777 (N_13777,N_13683,N_13520);
and U13778 (N_13778,N_13641,N_13271);
nand U13779 (N_13779,N_13429,N_13354);
or U13780 (N_13780,N_13658,N_13579);
or U13781 (N_13781,N_13596,N_13480);
and U13782 (N_13782,N_13290,N_13654);
or U13783 (N_13783,N_13155,N_13469);
and U13784 (N_13784,N_13539,N_13476);
and U13785 (N_13785,N_13149,N_13453);
or U13786 (N_13786,N_13414,N_13637);
and U13787 (N_13787,N_13157,N_13681);
or U13788 (N_13788,N_13674,N_13191);
or U13789 (N_13789,N_13531,N_13489);
nor U13790 (N_13790,N_13701,N_13340);
or U13791 (N_13791,N_13445,N_13441);
nand U13792 (N_13792,N_13407,N_13163);
and U13793 (N_13793,N_13569,N_13460);
nand U13794 (N_13794,N_13288,N_13655);
xnor U13795 (N_13795,N_13334,N_13398);
and U13796 (N_13796,N_13481,N_13224);
or U13797 (N_13797,N_13458,N_13289);
nand U13798 (N_13798,N_13247,N_13675);
nand U13799 (N_13799,N_13516,N_13150);
nand U13800 (N_13800,N_13512,N_13602);
nor U13801 (N_13801,N_13353,N_13307);
xor U13802 (N_13802,N_13194,N_13131);
or U13803 (N_13803,N_13692,N_13295);
or U13804 (N_13804,N_13217,N_13287);
or U13805 (N_13805,N_13555,N_13282);
nand U13806 (N_13806,N_13222,N_13600);
xor U13807 (N_13807,N_13215,N_13470);
xor U13808 (N_13808,N_13345,N_13365);
or U13809 (N_13809,N_13649,N_13721);
and U13810 (N_13810,N_13327,N_13359);
nand U13811 (N_13811,N_13567,N_13454);
nand U13812 (N_13812,N_13375,N_13632);
and U13813 (N_13813,N_13261,N_13212);
xnor U13814 (N_13814,N_13680,N_13337);
nor U13815 (N_13815,N_13475,N_13582);
xor U13816 (N_13816,N_13145,N_13742);
and U13817 (N_13817,N_13616,N_13142);
and U13818 (N_13818,N_13580,N_13661);
and U13819 (N_13819,N_13530,N_13199);
nor U13820 (N_13820,N_13497,N_13595);
or U13821 (N_13821,N_13313,N_13293);
nor U13822 (N_13822,N_13733,N_13564);
xnor U13823 (N_13823,N_13646,N_13719);
and U13824 (N_13824,N_13171,N_13185);
or U13825 (N_13825,N_13491,N_13328);
nand U13826 (N_13826,N_13578,N_13154);
nand U13827 (N_13827,N_13350,N_13635);
nand U13828 (N_13828,N_13697,N_13296);
xor U13829 (N_13829,N_13158,N_13134);
or U13830 (N_13830,N_13343,N_13438);
xnor U13831 (N_13831,N_13368,N_13576);
and U13832 (N_13832,N_13371,N_13533);
and U13833 (N_13833,N_13312,N_13613);
nor U13834 (N_13834,N_13226,N_13372);
nand U13835 (N_13835,N_13419,N_13402);
nand U13836 (N_13836,N_13541,N_13597);
nor U13837 (N_13837,N_13227,N_13746);
or U13838 (N_13838,N_13418,N_13745);
or U13839 (N_13839,N_13729,N_13378);
and U13840 (N_13840,N_13216,N_13709);
nor U13841 (N_13841,N_13736,N_13202);
nand U13842 (N_13842,N_13669,N_13725);
nor U13843 (N_13843,N_13711,N_13198);
xor U13844 (N_13844,N_13361,N_13687);
or U13845 (N_13845,N_13690,N_13234);
nand U13846 (N_13846,N_13663,N_13315);
nand U13847 (N_13847,N_13208,N_13406);
nor U13848 (N_13848,N_13724,N_13240);
nor U13849 (N_13849,N_13720,N_13627);
nor U13850 (N_13850,N_13586,N_13332);
xnor U13851 (N_13851,N_13292,N_13570);
and U13852 (N_13852,N_13451,N_13220);
and U13853 (N_13853,N_13647,N_13223);
or U13854 (N_13854,N_13331,N_13153);
nand U13855 (N_13855,N_13508,N_13173);
nor U13856 (N_13856,N_13560,N_13703);
and U13857 (N_13857,N_13415,N_13642);
xor U13858 (N_13858,N_13236,N_13548);
xor U13859 (N_13859,N_13446,N_13473);
nand U13860 (N_13860,N_13213,N_13525);
nand U13861 (N_13861,N_13645,N_13706);
nor U13862 (N_13862,N_13147,N_13524);
nor U13863 (N_13863,N_13182,N_13630);
and U13864 (N_13864,N_13274,N_13132);
and U13865 (N_13865,N_13667,N_13197);
nand U13866 (N_13866,N_13682,N_13693);
nor U13867 (N_13867,N_13726,N_13139);
or U13868 (N_13868,N_13360,N_13214);
nand U13869 (N_13869,N_13389,N_13400);
or U13870 (N_13870,N_13507,N_13270);
xnor U13871 (N_13871,N_13152,N_13188);
nand U13872 (N_13872,N_13739,N_13463);
and U13873 (N_13873,N_13503,N_13558);
xor U13874 (N_13874,N_13688,N_13561);
nor U13875 (N_13875,N_13133,N_13741);
or U13876 (N_13876,N_13559,N_13517);
nand U13877 (N_13877,N_13390,N_13614);
and U13878 (N_13878,N_13342,N_13624);
nor U13879 (N_13879,N_13549,N_13676);
and U13880 (N_13880,N_13581,N_13383);
or U13881 (N_13881,N_13622,N_13668);
and U13882 (N_13882,N_13506,N_13643);
or U13883 (N_13883,N_13461,N_13382);
nand U13884 (N_13884,N_13529,N_13665);
nand U13885 (N_13885,N_13210,N_13483);
nand U13886 (N_13886,N_13266,N_13657);
and U13887 (N_13887,N_13466,N_13421);
and U13888 (N_13888,N_13189,N_13707);
and U13889 (N_13889,N_13388,N_13568);
nand U13890 (N_13890,N_13543,N_13652);
or U13891 (N_13891,N_13490,N_13615);
and U13892 (N_13892,N_13294,N_13352);
nor U13893 (N_13893,N_13493,N_13256);
xor U13894 (N_13894,N_13732,N_13651);
and U13895 (N_13895,N_13181,N_13485);
nor U13896 (N_13896,N_13403,N_13174);
xnor U13897 (N_13897,N_13457,N_13162);
nor U13898 (N_13898,N_13547,N_13513);
and U13899 (N_13899,N_13143,N_13633);
nand U13900 (N_13900,N_13209,N_13509);
or U13901 (N_13901,N_13422,N_13691);
and U13902 (N_13902,N_13207,N_13357);
xnor U13903 (N_13903,N_13737,N_13175);
nor U13904 (N_13904,N_13195,N_13394);
and U13905 (N_13905,N_13740,N_13333);
nor U13906 (N_13906,N_13341,N_13329);
and U13907 (N_13907,N_13502,N_13629);
nand U13908 (N_13908,N_13268,N_13728);
or U13909 (N_13909,N_13444,N_13511);
xor U13910 (N_13910,N_13621,N_13593);
xnor U13911 (N_13911,N_13714,N_13704);
nor U13912 (N_13912,N_13601,N_13374);
and U13913 (N_13913,N_13320,N_13250);
nand U13914 (N_13914,N_13205,N_13631);
nor U13915 (N_13915,N_13130,N_13204);
xor U13916 (N_13916,N_13563,N_13698);
nor U13917 (N_13917,N_13308,N_13554);
nand U13918 (N_13918,N_13467,N_13717);
xor U13919 (N_13919,N_13424,N_13144);
and U13920 (N_13920,N_13370,N_13286);
or U13921 (N_13921,N_13184,N_13159);
nor U13922 (N_13922,N_13542,N_13246);
nor U13923 (N_13923,N_13310,N_13727);
nor U13924 (N_13924,N_13664,N_13434);
nor U13925 (N_13925,N_13620,N_13298);
xnor U13926 (N_13926,N_13355,N_13348);
xnor U13927 (N_13927,N_13526,N_13285);
xor U13928 (N_13928,N_13326,N_13584);
and U13929 (N_13929,N_13306,N_13433);
xnor U13930 (N_13930,N_13180,N_13267);
or U13931 (N_13931,N_13238,N_13347);
nor U13932 (N_13932,N_13249,N_13515);
xor U13933 (N_13933,N_13425,N_13660);
nand U13934 (N_13934,N_13607,N_13605);
and U13935 (N_13935,N_13409,N_13413);
and U13936 (N_13936,N_13468,N_13744);
nand U13937 (N_13937,N_13248,N_13514);
nand U13938 (N_13938,N_13203,N_13678);
and U13939 (N_13939,N_13479,N_13505);
and U13940 (N_13940,N_13659,N_13364);
or U13941 (N_13941,N_13459,N_13335);
xor U13942 (N_13942,N_13730,N_13177);
or U13943 (N_13943,N_13283,N_13280);
nand U13944 (N_13944,N_13423,N_13275);
nand U13945 (N_13945,N_13735,N_13747);
and U13946 (N_13946,N_13702,N_13471);
and U13947 (N_13947,N_13166,N_13462);
xnor U13948 (N_13948,N_13219,N_13685);
xor U13949 (N_13949,N_13608,N_13302);
nor U13950 (N_13950,N_13500,N_13305);
and U13951 (N_13951,N_13450,N_13179);
xnor U13952 (N_13952,N_13279,N_13722);
and U13953 (N_13953,N_13447,N_13519);
or U13954 (N_13954,N_13129,N_13127);
or U13955 (N_13955,N_13257,N_13395);
xor U13956 (N_13956,N_13628,N_13694);
xor U13957 (N_13957,N_13550,N_13190);
xor U13958 (N_13958,N_13229,N_13178);
nand U13959 (N_13959,N_13265,N_13231);
and U13960 (N_13960,N_13393,N_13677);
or U13961 (N_13961,N_13551,N_13599);
nor U13962 (N_13962,N_13532,N_13253);
nor U13963 (N_13963,N_13437,N_13431);
nand U13964 (N_13964,N_13258,N_13399);
and U13965 (N_13965,N_13319,N_13594);
or U13966 (N_13966,N_13230,N_13501);
nor U13967 (N_13967,N_13260,N_13731);
nand U13968 (N_13968,N_13160,N_13358);
xnor U13969 (N_13969,N_13408,N_13672);
or U13970 (N_13970,N_13617,N_13715);
and U13971 (N_13971,N_13465,N_13251);
or U13972 (N_13972,N_13478,N_13321);
nor U13973 (N_13973,N_13510,N_13684);
or U13974 (N_13974,N_13264,N_13573);
and U13975 (N_13975,N_13610,N_13299);
nor U13976 (N_13976,N_13410,N_13700);
nor U13977 (N_13977,N_13262,N_13571);
and U13978 (N_13978,N_13304,N_13379);
or U13979 (N_13979,N_13653,N_13553);
xor U13980 (N_13980,N_13435,N_13536);
and U13981 (N_13981,N_13591,N_13330);
xor U13982 (N_13982,N_13278,N_13277);
or U13983 (N_13983,N_13301,N_13405);
nor U13984 (N_13984,N_13430,N_13362);
nand U13985 (N_13985,N_13156,N_13689);
nor U13986 (N_13986,N_13537,N_13252);
xor U13987 (N_13987,N_13412,N_13148);
nand U13988 (N_13988,N_13670,N_13748);
nor U13989 (N_13989,N_13734,N_13486);
or U13990 (N_13990,N_13546,N_13538);
nand U13991 (N_13991,N_13432,N_13218);
xor U13992 (N_13992,N_13477,N_13167);
or U13993 (N_13993,N_13126,N_13464);
xor U13994 (N_13994,N_13200,N_13164);
and U13995 (N_13995,N_13523,N_13233);
xor U13996 (N_13996,N_13245,N_13448);
nor U13997 (N_13997,N_13534,N_13259);
xnor U13998 (N_13998,N_13656,N_13589);
and U13999 (N_13999,N_13416,N_13235);
and U14000 (N_14000,N_13255,N_13562);
and U14001 (N_14001,N_13172,N_13618);
nor U14002 (N_14002,N_13140,N_13699);
nand U14003 (N_14003,N_13254,N_13452);
or U14004 (N_14004,N_13603,N_13574);
or U14005 (N_14005,N_13612,N_13544);
nor U14006 (N_14006,N_13161,N_13239);
and U14007 (N_14007,N_13644,N_13317);
nand U14008 (N_14008,N_13487,N_13590);
or U14009 (N_14009,N_13324,N_13376);
and U14010 (N_14010,N_13377,N_13611);
or U14011 (N_14011,N_13738,N_13356);
nor U14012 (N_14012,N_13587,N_13232);
nand U14013 (N_14013,N_13640,N_13671);
xnor U14014 (N_14014,N_13183,N_13565);
nand U14015 (N_14015,N_13557,N_13165);
nor U14016 (N_14016,N_13201,N_13206);
or U14017 (N_14017,N_13339,N_13498);
and U14018 (N_14018,N_13679,N_13440);
nor U14019 (N_14019,N_13648,N_13186);
nand U14020 (N_14020,N_13385,N_13673);
nand U14021 (N_14021,N_13713,N_13363);
nor U14022 (N_14022,N_13241,N_13401);
nor U14023 (N_14023,N_13314,N_13442);
and U14024 (N_14024,N_13193,N_13381);
nand U14025 (N_14025,N_13495,N_13336);
or U14026 (N_14026,N_13284,N_13367);
or U14027 (N_14027,N_13619,N_13176);
and U14028 (N_14028,N_13297,N_13420);
nand U14029 (N_14029,N_13316,N_13344);
xnor U14030 (N_14030,N_13311,N_13300);
nand U14031 (N_14031,N_13291,N_13662);
nor U14032 (N_14032,N_13243,N_13705);
and U14033 (N_14033,N_13318,N_13168);
and U14034 (N_14034,N_13518,N_13443);
nand U14035 (N_14035,N_13634,N_13696);
nor U14036 (N_14036,N_13196,N_13276);
and U14037 (N_14037,N_13499,N_13380);
xnor U14038 (N_14038,N_13396,N_13449);
and U14039 (N_14039,N_13639,N_13397);
and U14040 (N_14040,N_13386,N_13472);
nand U14041 (N_14041,N_13242,N_13427);
xor U14042 (N_14042,N_13426,N_13636);
nand U14043 (N_14043,N_13391,N_13556);
and U14044 (N_14044,N_13666,N_13137);
nor U14045 (N_14045,N_13686,N_13303);
nor U14046 (N_14046,N_13650,N_13626);
or U14047 (N_14047,N_13244,N_13575);
and U14048 (N_14048,N_13609,N_13598);
or U14049 (N_14049,N_13281,N_13528);
and U14050 (N_14050,N_13351,N_13749);
nor U14051 (N_14051,N_13146,N_13712);
xnor U14052 (N_14052,N_13552,N_13482);
or U14053 (N_14053,N_13263,N_13417);
and U14054 (N_14054,N_13456,N_13366);
nor U14055 (N_14055,N_13592,N_13521);
nand U14056 (N_14056,N_13494,N_13338);
nor U14057 (N_14057,N_13404,N_13128);
nor U14058 (N_14058,N_13384,N_13428);
or U14059 (N_14059,N_13522,N_13484);
nand U14060 (N_14060,N_13323,N_13572);
nor U14061 (N_14061,N_13237,N_13710);
xnor U14062 (N_14062,N_13369,N_13255);
nor U14063 (N_14063,N_13508,N_13461);
or U14064 (N_14064,N_13639,N_13385);
or U14065 (N_14065,N_13286,N_13395);
nor U14066 (N_14066,N_13653,N_13516);
xor U14067 (N_14067,N_13451,N_13377);
nor U14068 (N_14068,N_13303,N_13554);
xor U14069 (N_14069,N_13184,N_13372);
or U14070 (N_14070,N_13658,N_13445);
xnor U14071 (N_14071,N_13556,N_13269);
or U14072 (N_14072,N_13179,N_13644);
nor U14073 (N_14073,N_13199,N_13314);
nor U14074 (N_14074,N_13496,N_13210);
xnor U14075 (N_14075,N_13325,N_13578);
or U14076 (N_14076,N_13550,N_13389);
xor U14077 (N_14077,N_13285,N_13474);
xor U14078 (N_14078,N_13581,N_13159);
xor U14079 (N_14079,N_13202,N_13416);
or U14080 (N_14080,N_13699,N_13285);
and U14081 (N_14081,N_13400,N_13738);
nor U14082 (N_14082,N_13281,N_13496);
and U14083 (N_14083,N_13137,N_13541);
nor U14084 (N_14084,N_13305,N_13142);
nand U14085 (N_14085,N_13288,N_13183);
or U14086 (N_14086,N_13420,N_13647);
xnor U14087 (N_14087,N_13608,N_13648);
nor U14088 (N_14088,N_13445,N_13673);
or U14089 (N_14089,N_13511,N_13303);
or U14090 (N_14090,N_13250,N_13389);
nor U14091 (N_14091,N_13515,N_13325);
and U14092 (N_14092,N_13338,N_13500);
xor U14093 (N_14093,N_13336,N_13126);
xor U14094 (N_14094,N_13664,N_13285);
or U14095 (N_14095,N_13163,N_13351);
nor U14096 (N_14096,N_13727,N_13741);
and U14097 (N_14097,N_13591,N_13277);
nand U14098 (N_14098,N_13468,N_13403);
and U14099 (N_14099,N_13408,N_13222);
xor U14100 (N_14100,N_13477,N_13656);
xnor U14101 (N_14101,N_13547,N_13167);
xnor U14102 (N_14102,N_13607,N_13139);
nand U14103 (N_14103,N_13155,N_13160);
nor U14104 (N_14104,N_13609,N_13606);
or U14105 (N_14105,N_13244,N_13637);
nand U14106 (N_14106,N_13417,N_13730);
and U14107 (N_14107,N_13259,N_13435);
and U14108 (N_14108,N_13284,N_13652);
or U14109 (N_14109,N_13161,N_13427);
nor U14110 (N_14110,N_13653,N_13673);
nor U14111 (N_14111,N_13575,N_13204);
nand U14112 (N_14112,N_13165,N_13648);
or U14113 (N_14113,N_13371,N_13262);
or U14114 (N_14114,N_13582,N_13371);
xor U14115 (N_14115,N_13225,N_13434);
or U14116 (N_14116,N_13230,N_13710);
and U14117 (N_14117,N_13742,N_13675);
nor U14118 (N_14118,N_13286,N_13315);
and U14119 (N_14119,N_13488,N_13356);
nand U14120 (N_14120,N_13662,N_13443);
xor U14121 (N_14121,N_13226,N_13219);
or U14122 (N_14122,N_13337,N_13547);
nand U14123 (N_14123,N_13327,N_13610);
nand U14124 (N_14124,N_13325,N_13511);
and U14125 (N_14125,N_13348,N_13326);
xnor U14126 (N_14126,N_13255,N_13174);
nand U14127 (N_14127,N_13686,N_13530);
or U14128 (N_14128,N_13532,N_13190);
nand U14129 (N_14129,N_13567,N_13528);
or U14130 (N_14130,N_13624,N_13156);
xor U14131 (N_14131,N_13279,N_13361);
xnor U14132 (N_14132,N_13333,N_13157);
and U14133 (N_14133,N_13605,N_13139);
xnor U14134 (N_14134,N_13244,N_13175);
or U14135 (N_14135,N_13422,N_13475);
xor U14136 (N_14136,N_13364,N_13676);
nor U14137 (N_14137,N_13501,N_13697);
or U14138 (N_14138,N_13429,N_13545);
and U14139 (N_14139,N_13391,N_13699);
nand U14140 (N_14140,N_13686,N_13358);
nor U14141 (N_14141,N_13741,N_13486);
or U14142 (N_14142,N_13533,N_13583);
nand U14143 (N_14143,N_13423,N_13431);
nor U14144 (N_14144,N_13238,N_13209);
xor U14145 (N_14145,N_13643,N_13142);
nor U14146 (N_14146,N_13290,N_13528);
or U14147 (N_14147,N_13723,N_13571);
and U14148 (N_14148,N_13559,N_13401);
and U14149 (N_14149,N_13292,N_13296);
xnor U14150 (N_14150,N_13247,N_13158);
nor U14151 (N_14151,N_13230,N_13343);
nand U14152 (N_14152,N_13646,N_13337);
nand U14153 (N_14153,N_13341,N_13720);
or U14154 (N_14154,N_13417,N_13231);
xor U14155 (N_14155,N_13316,N_13204);
xnor U14156 (N_14156,N_13184,N_13425);
nand U14157 (N_14157,N_13698,N_13442);
nor U14158 (N_14158,N_13428,N_13659);
and U14159 (N_14159,N_13738,N_13601);
or U14160 (N_14160,N_13651,N_13502);
or U14161 (N_14161,N_13614,N_13192);
and U14162 (N_14162,N_13610,N_13389);
nand U14163 (N_14163,N_13125,N_13586);
xor U14164 (N_14164,N_13610,N_13407);
nor U14165 (N_14165,N_13438,N_13346);
or U14166 (N_14166,N_13274,N_13238);
nor U14167 (N_14167,N_13335,N_13195);
or U14168 (N_14168,N_13283,N_13213);
and U14169 (N_14169,N_13294,N_13689);
xor U14170 (N_14170,N_13295,N_13554);
or U14171 (N_14171,N_13580,N_13601);
and U14172 (N_14172,N_13400,N_13151);
xor U14173 (N_14173,N_13159,N_13298);
and U14174 (N_14174,N_13140,N_13580);
nor U14175 (N_14175,N_13206,N_13512);
xnor U14176 (N_14176,N_13377,N_13408);
nor U14177 (N_14177,N_13352,N_13342);
or U14178 (N_14178,N_13174,N_13239);
xnor U14179 (N_14179,N_13656,N_13440);
and U14180 (N_14180,N_13637,N_13727);
or U14181 (N_14181,N_13640,N_13354);
nand U14182 (N_14182,N_13411,N_13688);
and U14183 (N_14183,N_13233,N_13360);
nand U14184 (N_14184,N_13579,N_13572);
nand U14185 (N_14185,N_13353,N_13673);
nand U14186 (N_14186,N_13158,N_13548);
xor U14187 (N_14187,N_13532,N_13407);
and U14188 (N_14188,N_13443,N_13342);
and U14189 (N_14189,N_13723,N_13548);
nor U14190 (N_14190,N_13149,N_13205);
and U14191 (N_14191,N_13678,N_13285);
xnor U14192 (N_14192,N_13207,N_13527);
nand U14193 (N_14193,N_13256,N_13139);
nand U14194 (N_14194,N_13319,N_13181);
nor U14195 (N_14195,N_13253,N_13713);
xnor U14196 (N_14196,N_13126,N_13583);
and U14197 (N_14197,N_13567,N_13312);
nor U14198 (N_14198,N_13477,N_13138);
or U14199 (N_14199,N_13483,N_13173);
nand U14200 (N_14200,N_13300,N_13196);
or U14201 (N_14201,N_13493,N_13496);
xor U14202 (N_14202,N_13438,N_13381);
nor U14203 (N_14203,N_13340,N_13599);
and U14204 (N_14204,N_13326,N_13430);
nor U14205 (N_14205,N_13532,N_13674);
xnor U14206 (N_14206,N_13267,N_13168);
xnor U14207 (N_14207,N_13625,N_13515);
xor U14208 (N_14208,N_13365,N_13718);
nand U14209 (N_14209,N_13640,N_13482);
nand U14210 (N_14210,N_13458,N_13631);
xor U14211 (N_14211,N_13141,N_13701);
or U14212 (N_14212,N_13150,N_13176);
or U14213 (N_14213,N_13187,N_13406);
nand U14214 (N_14214,N_13396,N_13339);
nor U14215 (N_14215,N_13691,N_13500);
nand U14216 (N_14216,N_13417,N_13601);
nor U14217 (N_14217,N_13143,N_13293);
and U14218 (N_14218,N_13696,N_13548);
xor U14219 (N_14219,N_13395,N_13670);
nand U14220 (N_14220,N_13673,N_13714);
nand U14221 (N_14221,N_13240,N_13348);
xor U14222 (N_14222,N_13703,N_13387);
nand U14223 (N_14223,N_13721,N_13561);
nor U14224 (N_14224,N_13199,N_13333);
nor U14225 (N_14225,N_13434,N_13234);
nand U14226 (N_14226,N_13607,N_13581);
nor U14227 (N_14227,N_13530,N_13186);
nand U14228 (N_14228,N_13289,N_13627);
xnor U14229 (N_14229,N_13141,N_13315);
nand U14230 (N_14230,N_13622,N_13287);
and U14231 (N_14231,N_13379,N_13154);
or U14232 (N_14232,N_13501,N_13669);
or U14233 (N_14233,N_13462,N_13583);
nor U14234 (N_14234,N_13666,N_13133);
nand U14235 (N_14235,N_13552,N_13462);
and U14236 (N_14236,N_13272,N_13145);
xnor U14237 (N_14237,N_13641,N_13424);
nand U14238 (N_14238,N_13183,N_13648);
nor U14239 (N_14239,N_13627,N_13172);
nand U14240 (N_14240,N_13598,N_13155);
and U14241 (N_14241,N_13488,N_13299);
nor U14242 (N_14242,N_13243,N_13129);
or U14243 (N_14243,N_13451,N_13743);
and U14244 (N_14244,N_13406,N_13376);
or U14245 (N_14245,N_13687,N_13421);
and U14246 (N_14246,N_13614,N_13675);
and U14247 (N_14247,N_13652,N_13481);
and U14248 (N_14248,N_13386,N_13691);
xor U14249 (N_14249,N_13424,N_13232);
xnor U14250 (N_14250,N_13197,N_13476);
nand U14251 (N_14251,N_13587,N_13656);
or U14252 (N_14252,N_13700,N_13271);
and U14253 (N_14253,N_13146,N_13342);
or U14254 (N_14254,N_13390,N_13346);
or U14255 (N_14255,N_13429,N_13473);
and U14256 (N_14256,N_13170,N_13706);
nand U14257 (N_14257,N_13694,N_13278);
nor U14258 (N_14258,N_13448,N_13281);
and U14259 (N_14259,N_13247,N_13356);
and U14260 (N_14260,N_13581,N_13176);
xor U14261 (N_14261,N_13389,N_13247);
xnor U14262 (N_14262,N_13596,N_13684);
xnor U14263 (N_14263,N_13296,N_13537);
or U14264 (N_14264,N_13413,N_13589);
and U14265 (N_14265,N_13328,N_13243);
nor U14266 (N_14266,N_13172,N_13643);
and U14267 (N_14267,N_13372,N_13525);
or U14268 (N_14268,N_13156,N_13716);
and U14269 (N_14269,N_13442,N_13241);
or U14270 (N_14270,N_13635,N_13628);
nor U14271 (N_14271,N_13492,N_13523);
or U14272 (N_14272,N_13387,N_13210);
nor U14273 (N_14273,N_13628,N_13322);
xnor U14274 (N_14274,N_13436,N_13577);
xor U14275 (N_14275,N_13160,N_13376);
and U14276 (N_14276,N_13557,N_13161);
xor U14277 (N_14277,N_13595,N_13605);
nand U14278 (N_14278,N_13644,N_13461);
xnor U14279 (N_14279,N_13176,N_13466);
or U14280 (N_14280,N_13155,N_13555);
xor U14281 (N_14281,N_13158,N_13620);
or U14282 (N_14282,N_13741,N_13491);
and U14283 (N_14283,N_13385,N_13643);
or U14284 (N_14284,N_13249,N_13220);
nand U14285 (N_14285,N_13395,N_13547);
nor U14286 (N_14286,N_13433,N_13397);
and U14287 (N_14287,N_13354,N_13672);
xnor U14288 (N_14288,N_13673,N_13434);
nor U14289 (N_14289,N_13645,N_13287);
and U14290 (N_14290,N_13310,N_13630);
and U14291 (N_14291,N_13469,N_13239);
or U14292 (N_14292,N_13150,N_13210);
or U14293 (N_14293,N_13388,N_13394);
or U14294 (N_14294,N_13270,N_13681);
nor U14295 (N_14295,N_13417,N_13469);
and U14296 (N_14296,N_13563,N_13514);
nand U14297 (N_14297,N_13386,N_13545);
nor U14298 (N_14298,N_13686,N_13692);
xor U14299 (N_14299,N_13418,N_13319);
or U14300 (N_14300,N_13137,N_13745);
and U14301 (N_14301,N_13689,N_13537);
nand U14302 (N_14302,N_13372,N_13695);
nand U14303 (N_14303,N_13277,N_13715);
xor U14304 (N_14304,N_13187,N_13292);
xor U14305 (N_14305,N_13260,N_13453);
xnor U14306 (N_14306,N_13252,N_13264);
nand U14307 (N_14307,N_13346,N_13243);
xor U14308 (N_14308,N_13664,N_13425);
and U14309 (N_14309,N_13212,N_13349);
and U14310 (N_14310,N_13374,N_13570);
nor U14311 (N_14311,N_13150,N_13441);
nand U14312 (N_14312,N_13203,N_13398);
nand U14313 (N_14313,N_13378,N_13736);
or U14314 (N_14314,N_13168,N_13137);
and U14315 (N_14315,N_13444,N_13309);
nor U14316 (N_14316,N_13628,N_13315);
and U14317 (N_14317,N_13680,N_13405);
nor U14318 (N_14318,N_13527,N_13370);
and U14319 (N_14319,N_13265,N_13533);
xnor U14320 (N_14320,N_13658,N_13499);
xor U14321 (N_14321,N_13396,N_13473);
nor U14322 (N_14322,N_13349,N_13323);
and U14323 (N_14323,N_13256,N_13708);
nand U14324 (N_14324,N_13162,N_13481);
xnor U14325 (N_14325,N_13559,N_13384);
or U14326 (N_14326,N_13142,N_13514);
and U14327 (N_14327,N_13687,N_13416);
nor U14328 (N_14328,N_13400,N_13683);
xnor U14329 (N_14329,N_13661,N_13551);
nor U14330 (N_14330,N_13494,N_13671);
or U14331 (N_14331,N_13417,N_13270);
or U14332 (N_14332,N_13387,N_13159);
and U14333 (N_14333,N_13217,N_13444);
nand U14334 (N_14334,N_13363,N_13658);
nor U14335 (N_14335,N_13302,N_13636);
and U14336 (N_14336,N_13394,N_13680);
nand U14337 (N_14337,N_13632,N_13298);
nor U14338 (N_14338,N_13327,N_13740);
nand U14339 (N_14339,N_13446,N_13401);
nor U14340 (N_14340,N_13150,N_13539);
nor U14341 (N_14341,N_13427,N_13202);
or U14342 (N_14342,N_13281,N_13381);
or U14343 (N_14343,N_13587,N_13373);
nor U14344 (N_14344,N_13680,N_13139);
and U14345 (N_14345,N_13259,N_13183);
xor U14346 (N_14346,N_13361,N_13612);
nand U14347 (N_14347,N_13405,N_13717);
xnor U14348 (N_14348,N_13542,N_13594);
nand U14349 (N_14349,N_13250,N_13406);
and U14350 (N_14350,N_13455,N_13146);
nand U14351 (N_14351,N_13742,N_13489);
xnor U14352 (N_14352,N_13214,N_13479);
or U14353 (N_14353,N_13302,N_13337);
or U14354 (N_14354,N_13424,N_13324);
or U14355 (N_14355,N_13163,N_13621);
or U14356 (N_14356,N_13130,N_13161);
nor U14357 (N_14357,N_13282,N_13210);
xor U14358 (N_14358,N_13477,N_13719);
nor U14359 (N_14359,N_13499,N_13506);
nand U14360 (N_14360,N_13536,N_13343);
or U14361 (N_14361,N_13291,N_13482);
and U14362 (N_14362,N_13603,N_13529);
or U14363 (N_14363,N_13506,N_13135);
and U14364 (N_14364,N_13639,N_13200);
and U14365 (N_14365,N_13214,N_13340);
or U14366 (N_14366,N_13505,N_13739);
nand U14367 (N_14367,N_13620,N_13465);
nor U14368 (N_14368,N_13585,N_13403);
or U14369 (N_14369,N_13611,N_13226);
xor U14370 (N_14370,N_13147,N_13715);
and U14371 (N_14371,N_13734,N_13587);
nor U14372 (N_14372,N_13452,N_13400);
nand U14373 (N_14373,N_13749,N_13154);
nor U14374 (N_14374,N_13168,N_13294);
nor U14375 (N_14375,N_14106,N_14325);
and U14376 (N_14376,N_14128,N_13818);
xor U14377 (N_14377,N_13857,N_13921);
xnor U14378 (N_14378,N_14109,N_13762);
and U14379 (N_14379,N_13946,N_14118);
nor U14380 (N_14380,N_13897,N_13759);
or U14381 (N_14381,N_13884,N_13779);
xor U14382 (N_14382,N_13766,N_13951);
and U14383 (N_14383,N_13904,N_13957);
xor U14384 (N_14384,N_14161,N_13767);
xnor U14385 (N_14385,N_13819,N_14186);
nand U14386 (N_14386,N_13781,N_14262);
nand U14387 (N_14387,N_14143,N_13913);
or U14388 (N_14388,N_13796,N_13961);
or U14389 (N_14389,N_14367,N_14238);
or U14390 (N_14390,N_14196,N_14122);
xnor U14391 (N_14391,N_14111,N_14212);
nand U14392 (N_14392,N_13987,N_13863);
or U14393 (N_14393,N_13976,N_14183);
and U14394 (N_14394,N_14064,N_13886);
nor U14395 (N_14395,N_13812,N_13825);
xnor U14396 (N_14396,N_14038,N_13873);
nor U14397 (N_14397,N_13864,N_14136);
xor U14398 (N_14398,N_13968,N_13817);
xnor U14399 (N_14399,N_13808,N_14032);
xor U14400 (N_14400,N_14241,N_13983);
nor U14401 (N_14401,N_14301,N_13772);
and U14402 (N_14402,N_14160,N_14075);
or U14403 (N_14403,N_13794,N_14069);
nor U14404 (N_14404,N_14133,N_14104);
xnor U14405 (N_14405,N_14170,N_14073);
nand U14406 (N_14406,N_13756,N_14278);
or U14407 (N_14407,N_14013,N_13908);
nand U14408 (N_14408,N_13947,N_14276);
and U14409 (N_14409,N_14326,N_14090);
nor U14410 (N_14410,N_13958,N_14313);
xor U14411 (N_14411,N_14357,N_14131);
xor U14412 (N_14412,N_14072,N_13815);
and U14413 (N_14413,N_13888,N_13950);
or U14414 (N_14414,N_14173,N_14284);
nand U14415 (N_14415,N_14221,N_14211);
and U14416 (N_14416,N_13985,N_13805);
nand U14417 (N_14417,N_14201,N_14327);
and U14418 (N_14418,N_13820,N_14004);
xor U14419 (N_14419,N_14076,N_13835);
nor U14420 (N_14420,N_14029,N_14156);
nand U14421 (N_14421,N_14268,N_14034);
and U14422 (N_14422,N_14130,N_13850);
nand U14423 (N_14423,N_13870,N_14341);
and U14424 (N_14424,N_13934,N_14081);
or U14425 (N_14425,N_14297,N_13930);
nand U14426 (N_14426,N_14062,N_14292);
nand U14427 (N_14427,N_13937,N_14263);
nor U14428 (N_14428,N_14197,N_13885);
xnor U14429 (N_14429,N_14203,N_14324);
xor U14430 (N_14430,N_14174,N_13956);
nand U14431 (N_14431,N_14120,N_14189);
nand U14432 (N_14432,N_13901,N_13875);
xor U14433 (N_14433,N_13970,N_14152);
xnor U14434 (N_14434,N_13971,N_13973);
nor U14435 (N_14435,N_13920,N_14222);
or U14436 (N_14436,N_14051,N_13892);
and U14437 (N_14437,N_13940,N_14220);
or U14438 (N_14438,N_14010,N_14359);
or U14439 (N_14439,N_14307,N_13926);
xor U14440 (N_14440,N_14146,N_14151);
nor U14441 (N_14441,N_13752,N_14138);
and U14442 (N_14442,N_13997,N_13963);
and U14443 (N_14443,N_13878,N_14372);
nor U14444 (N_14444,N_13979,N_14056);
xor U14445 (N_14445,N_14205,N_13755);
nand U14446 (N_14446,N_14250,N_13959);
and U14447 (N_14447,N_14270,N_14192);
nand U14448 (N_14448,N_13999,N_14112);
xor U14449 (N_14449,N_13900,N_14187);
nor U14450 (N_14450,N_14330,N_14286);
and U14451 (N_14451,N_13758,N_14225);
nor U14452 (N_14452,N_14157,N_13816);
or U14453 (N_14453,N_13811,N_13977);
nor U14454 (N_14454,N_14349,N_14318);
xnor U14455 (N_14455,N_13866,N_14177);
nor U14456 (N_14456,N_14331,N_14235);
or U14457 (N_14457,N_13949,N_14208);
and U14458 (N_14458,N_14098,N_14281);
nor U14459 (N_14459,N_14336,N_14125);
xnor U14460 (N_14460,N_14345,N_13865);
or U14461 (N_14461,N_13790,N_14181);
xnor U14462 (N_14462,N_13822,N_14167);
or U14463 (N_14463,N_13799,N_13981);
or U14464 (N_14464,N_14310,N_14265);
nand U14465 (N_14465,N_14258,N_13938);
and U14466 (N_14466,N_14371,N_14364);
and U14467 (N_14467,N_14351,N_13982);
and U14468 (N_14468,N_14057,N_14074);
nor U14469 (N_14469,N_14145,N_13778);
nand U14470 (N_14470,N_14086,N_13750);
and U14471 (N_14471,N_13757,N_13909);
nor U14472 (N_14472,N_14119,N_14030);
nor U14473 (N_14473,N_13876,N_13975);
xor U14474 (N_14474,N_14103,N_14300);
xor U14475 (N_14475,N_13771,N_14308);
nor U14476 (N_14476,N_13889,N_14155);
nand U14477 (N_14477,N_13830,N_14148);
or U14478 (N_14478,N_14317,N_14094);
xor U14479 (N_14479,N_14025,N_13782);
xnor U14480 (N_14480,N_13916,N_13896);
or U14481 (N_14481,N_14059,N_14287);
or U14482 (N_14482,N_14343,N_13753);
or U14483 (N_14483,N_14328,N_13871);
nand U14484 (N_14484,N_14003,N_14141);
or U14485 (N_14485,N_13774,N_14063);
nand U14486 (N_14486,N_13824,N_14065);
and U14487 (N_14487,N_14215,N_14066);
nand U14488 (N_14488,N_14117,N_14037);
xnor U14489 (N_14489,N_14009,N_14243);
xor U14490 (N_14490,N_13927,N_13823);
nor U14491 (N_14491,N_14071,N_13907);
or U14492 (N_14492,N_14289,N_13854);
or U14493 (N_14493,N_14230,N_14001);
or U14494 (N_14494,N_13905,N_14044);
nor U14495 (N_14495,N_14045,N_14269);
or U14496 (N_14496,N_14362,N_13841);
nor U14497 (N_14497,N_14061,N_14022);
nor U14498 (N_14498,N_14279,N_14231);
nand U14499 (N_14499,N_14288,N_13809);
xor U14500 (N_14500,N_14067,N_14018);
xor U14501 (N_14501,N_13986,N_14035);
nand U14502 (N_14502,N_14312,N_13802);
xnor U14503 (N_14503,N_14114,N_14095);
xor U14504 (N_14504,N_14058,N_13960);
xor U14505 (N_14505,N_14368,N_13763);
nand U14506 (N_14506,N_14246,N_13972);
or U14507 (N_14507,N_14194,N_13966);
xor U14508 (N_14508,N_14190,N_13821);
and U14509 (N_14509,N_13845,N_14015);
nor U14510 (N_14510,N_13860,N_14153);
or U14511 (N_14511,N_13989,N_13915);
nor U14512 (N_14512,N_13839,N_13784);
or U14513 (N_14513,N_13906,N_14089);
nand U14514 (N_14514,N_13847,N_13846);
nand U14515 (N_14515,N_14020,N_14280);
or U14516 (N_14516,N_13929,N_14031);
or U14517 (N_14517,N_13840,N_14242);
nand U14518 (N_14518,N_13978,N_13848);
or U14519 (N_14519,N_14115,N_14294);
or U14520 (N_14520,N_14232,N_14171);
nor U14521 (N_14521,N_14274,N_14169);
nor U14522 (N_14522,N_14185,N_14100);
xnor U14523 (N_14523,N_14337,N_13806);
nor U14524 (N_14524,N_13980,N_14110);
nand U14525 (N_14525,N_14333,N_14306);
nor U14526 (N_14526,N_14296,N_13941);
nand U14527 (N_14527,N_13944,N_13931);
xnor U14528 (N_14528,N_13932,N_13935);
and U14529 (N_14529,N_14226,N_14369);
and U14530 (N_14530,N_13945,N_13964);
or U14531 (N_14531,N_14097,N_13836);
xnor U14532 (N_14532,N_13785,N_13895);
or U14533 (N_14533,N_13786,N_14224);
nor U14534 (N_14534,N_14135,N_14162);
xnor U14535 (N_14535,N_14079,N_14083);
xnor U14536 (N_14536,N_14244,N_13899);
nand U14537 (N_14537,N_14251,N_14093);
or U14538 (N_14538,N_13925,N_14043);
xnor U14539 (N_14539,N_13891,N_14356);
xor U14540 (N_14540,N_13874,N_14210);
and U14541 (N_14541,N_14322,N_13974);
and U14542 (N_14542,N_14339,N_13902);
and U14543 (N_14543,N_14099,N_14055);
nand U14544 (N_14544,N_14291,N_14245);
xnor U14545 (N_14545,N_14199,N_14040);
and U14546 (N_14546,N_14223,N_13800);
nor U14547 (N_14547,N_14159,N_14091);
xnor U14548 (N_14548,N_13793,N_14373);
nor U14549 (N_14549,N_13832,N_14023);
nand U14550 (N_14550,N_14033,N_14374);
xnor U14551 (N_14551,N_13912,N_14188);
xnor U14552 (N_14552,N_14275,N_14149);
nor U14553 (N_14553,N_13965,N_14234);
nand U14554 (N_14554,N_14012,N_14361);
or U14555 (N_14555,N_13862,N_13883);
or U14556 (N_14556,N_13910,N_13914);
or U14557 (N_14557,N_14264,N_13898);
nor U14558 (N_14558,N_14132,N_14116);
xor U14559 (N_14559,N_14008,N_14080);
nand U14560 (N_14560,N_14311,N_14158);
or U14561 (N_14561,N_14028,N_13969);
and U14562 (N_14562,N_13911,N_14365);
and U14563 (N_14563,N_13761,N_13924);
nand U14564 (N_14564,N_13787,N_13780);
nand U14565 (N_14565,N_13887,N_14358);
xnor U14566 (N_14566,N_13813,N_14126);
and U14567 (N_14567,N_14124,N_13988);
nor U14568 (N_14568,N_14253,N_14366);
and U14569 (N_14569,N_14085,N_13826);
xor U14570 (N_14570,N_13953,N_13844);
and U14571 (N_14571,N_14127,N_13998);
or U14572 (N_14572,N_13807,N_13996);
or U14573 (N_14573,N_14218,N_13992);
nor U14574 (N_14574,N_14178,N_14323);
or U14575 (N_14575,N_14048,N_14207);
and U14576 (N_14576,N_14191,N_14180);
nor U14577 (N_14577,N_14248,N_13955);
nor U14578 (N_14578,N_14283,N_13804);
and U14579 (N_14579,N_14216,N_13872);
nand U14580 (N_14580,N_14236,N_13797);
xnor U14581 (N_14581,N_13837,N_13827);
nand U14582 (N_14582,N_14202,N_14219);
or U14583 (N_14583,N_14140,N_14233);
and U14584 (N_14584,N_14154,N_14092);
nor U14585 (N_14585,N_14036,N_13834);
nor U14586 (N_14586,N_13993,N_14305);
and U14587 (N_14587,N_14321,N_14184);
nor U14588 (N_14588,N_14053,N_14249);
xnor U14589 (N_14589,N_13942,N_14350);
nand U14590 (N_14590,N_14261,N_14087);
or U14591 (N_14591,N_13893,N_14237);
or U14592 (N_14592,N_14206,N_14335);
xor U14593 (N_14593,N_13881,N_13754);
and U14594 (N_14594,N_13984,N_14193);
and U14595 (N_14595,N_13798,N_14285);
nor U14596 (N_14596,N_13922,N_13879);
xnor U14597 (N_14597,N_14000,N_13928);
nor U14598 (N_14598,N_14355,N_13810);
nand U14599 (N_14599,N_13855,N_14163);
nor U14600 (N_14600,N_13990,N_14121);
nand U14601 (N_14601,N_14200,N_13919);
nand U14602 (N_14602,N_14314,N_14047);
nand U14603 (N_14603,N_14239,N_14198);
nand U14604 (N_14604,N_14182,N_14272);
or U14605 (N_14605,N_13903,N_14217);
or U14606 (N_14606,N_13918,N_14293);
nor U14607 (N_14607,N_14108,N_14077);
nand U14608 (N_14608,N_13995,N_14266);
xnor U14609 (N_14609,N_14113,N_14303);
xor U14610 (N_14610,N_14332,N_14024);
and U14611 (N_14611,N_13952,N_14107);
nor U14612 (N_14612,N_14102,N_13765);
and U14613 (N_14613,N_14084,N_14016);
or U14614 (N_14614,N_14070,N_14214);
and U14615 (N_14615,N_14176,N_14342);
nand U14616 (N_14616,N_14166,N_14046);
or U14617 (N_14617,N_13751,N_14348);
nand U14618 (N_14618,N_14354,N_14257);
xnor U14619 (N_14619,N_14137,N_14011);
nand U14620 (N_14620,N_14340,N_14172);
nor U14621 (N_14621,N_14299,N_14088);
and U14622 (N_14622,N_13788,N_14360);
nor U14623 (N_14623,N_14255,N_13861);
or U14624 (N_14624,N_13776,N_13843);
xor U14625 (N_14625,N_14282,N_14240);
nand U14626 (N_14626,N_13933,N_14319);
and U14627 (N_14627,N_13877,N_13948);
and U14628 (N_14628,N_13939,N_13856);
or U14629 (N_14629,N_14309,N_13894);
xor U14630 (N_14630,N_14134,N_14054);
or U14631 (N_14631,N_13954,N_14259);
or U14632 (N_14632,N_13882,N_13789);
nor U14633 (N_14633,N_13775,N_14247);
or U14634 (N_14634,N_14363,N_13859);
nand U14635 (N_14635,N_13994,N_13783);
nor U14636 (N_14636,N_13852,N_14168);
and U14637 (N_14637,N_13768,N_14123);
nand U14638 (N_14638,N_13801,N_14267);
xnor U14639 (N_14639,N_14179,N_14175);
or U14640 (N_14640,N_14019,N_13880);
xnor U14641 (N_14641,N_14142,N_14370);
xnor U14642 (N_14642,N_14352,N_14213);
and U14643 (N_14643,N_14039,N_14105);
nor U14644 (N_14644,N_13769,N_14147);
or U14645 (N_14645,N_13858,N_14344);
xnor U14646 (N_14646,N_14026,N_13814);
nand U14647 (N_14647,N_13770,N_14052);
and U14648 (N_14648,N_14334,N_13890);
nand U14649 (N_14649,N_13849,N_14329);
nor U14650 (N_14650,N_14068,N_13842);
or U14651 (N_14651,N_14227,N_13923);
nand U14652 (N_14652,N_13868,N_14347);
xnor U14653 (N_14653,N_14165,N_14298);
and U14654 (N_14654,N_13838,N_14320);
and U14655 (N_14655,N_14295,N_13760);
nor U14656 (N_14656,N_14050,N_14256);
xor U14657 (N_14657,N_13795,N_14260);
xnor U14658 (N_14658,N_14082,N_14273);
nand U14659 (N_14659,N_13773,N_14271);
and U14660 (N_14660,N_13791,N_14049);
or U14661 (N_14661,N_14007,N_14150);
and U14662 (N_14662,N_14078,N_14096);
and U14663 (N_14663,N_14353,N_14129);
or U14664 (N_14664,N_14002,N_14021);
or U14665 (N_14665,N_14228,N_14315);
nor U14666 (N_14666,N_13829,N_14164);
nor U14667 (N_14667,N_14195,N_14060);
nand U14668 (N_14668,N_14229,N_14139);
nand U14669 (N_14669,N_13991,N_13792);
nor U14670 (N_14670,N_13967,N_13777);
nor U14671 (N_14671,N_14005,N_14316);
xor U14672 (N_14672,N_14302,N_13867);
or U14673 (N_14673,N_14277,N_14101);
nand U14674 (N_14674,N_14027,N_13803);
xor U14675 (N_14675,N_14252,N_14144);
nand U14676 (N_14676,N_14041,N_13917);
or U14677 (N_14677,N_13943,N_13831);
and U14678 (N_14678,N_14014,N_13833);
or U14679 (N_14679,N_13764,N_14304);
or U14680 (N_14680,N_14254,N_14338);
nand U14681 (N_14681,N_14290,N_13828);
and U14682 (N_14682,N_13851,N_14006);
and U14683 (N_14683,N_14017,N_13962);
or U14684 (N_14684,N_13936,N_13853);
nor U14685 (N_14685,N_13869,N_14346);
nor U14686 (N_14686,N_14209,N_14204);
nand U14687 (N_14687,N_14042,N_14299);
and U14688 (N_14688,N_13834,N_14345);
and U14689 (N_14689,N_13901,N_14102);
or U14690 (N_14690,N_13966,N_14307);
xnor U14691 (N_14691,N_13983,N_14005);
nand U14692 (N_14692,N_13813,N_14076);
nor U14693 (N_14693,N_13762,N_14327);
and U14694 (N_14694,N_14167,N_13831);
nor U14695 (N_14695,N_14008,N_14233);
nand U14696 (N_14696,N_14025,N_13882);
xnor U14697 (N_14697,N_13786,N_13944);
or U14698 (N_14698,N_14031,N_14032);
or U14699 (N_14699,N_13916,N_14097);
nand U14700 (N_14700,N_14187,N_14314);
xnor U14701 (N_14701,N_14218,N_13757);
xnor U14702 (N_14702,N_13849,N_13830);
or U14703 (N_14703,N_14034,N_14211);
or U14704 (N_14704,N_13770,N_14174);
and U14705 (N_14705,N_13996,N_14229);
and U14706 (N_14706,N_14058,N_13782);
nor U14707 (N_14707,N_14243,N_14186);
nand U14708 (N_14708,N_14191,N_14102);
nor U14709 (N_14709,N_13764,N_14273);
nor U14710 (N_14710,N_14238,N_14105);
nand U14711 (N_14711,N_13821,N_14254);
nand U14712 (N_14712,N_13959,N_14348);
and U14713 (N_14713,N_14302,N_13869);
nor U14714 (N_14714,N_13904,N_14078);
nor U14715 (N_14715,N_14200,N_14203);
xor U14716 (N_14716,N_14229,N_13869);
and U14717 (N_14717,N_13868,N_14308);
xor U14718 (N_14718,N_14372,N_13973);
or U14719 (N_14719,N_14040,N_14000);
nor U14720 (N_14720,N_13976,N_13789);
and U14721 (N_14721,N_14224,N_13940);
and U14722 (N_14722,N_13851,N_13893);
nand U14723 (N_14723,N_13984,N_13924);
nor U14724 (N_14724,N_13985,N_13821);
and U14725 (N_14725,N_13804,N_14311);
xor U14726 (N_14726,N_13799,N_13775);
nand U14727 (N_14727,N_13978,N_13920);
xor U14728 (N_14728,N_14122,N_14036);
nand U14729 (N_14729,N_14284,N_14071);
and U14730 (N_14730,N_13868,N_13902);
nor U14731 (N_14731,N_14035,N_14020);
and U14732 (N_14732,N_14045,N_13795);
or U14733 (N_14733,N_14142,N_13911);
and U14734 (N_14734,N_14196,N_14329);
xnor U14735 (N_14735,N_14163,N_14134);
nand U14736 (N_14736,N_13789,N_14192);
and U14737 (N_14737,N_13834,N_14173);
xor U14738 (N_14738,N_14091,N_14212);
and U14739 (N_14739,N_13925,N_13761);
and U14740 (N_14740,N_13872,N_14293);
and U14741 (N_14741,N_14098,N_14126);
nor U14742 (N_14742,N_14317,N_14229);
nand U14743 (N_14743,N_14138,N_14003);
and U14744 (N_14744,N_14004,N_14117);
nor U14745 (N_14745,N_14180,N_14302);
nor U14746 (N_14746,N_14081,N_14353);
and U14747 (N_14747,N_13767,N_13828);
or U14748 (N_14748,N_14267,N_13750);
xnor U14749 (N_14749,N_14360,N_14225);
xor U14750 (N_14750,N_14068,N_14097);
xor U14751 (N_14751,N_13819,N_14058);
and U14752 (N_14752,N_13877,N_14122);
nand U14753 (N_14753,N_14351,N_14171);
xnor U14754 (N_14754,N_13941,N_14199);
or U14755 (N_14755,N_13752,N_14253);
or U14756 (N_14756,N_13944,N_13856);
nand U14757 (N_14757,N_14327,N_13938);
nor U14758 (N_14758,N_13751,N_14330);
or U14759 (N_14759,N_13918,N_14298);
xor U14760 (N_14760,N_14120,N_13964);
and U14761 (N_14761,N_14200,N_14139);
and U14762 (N_14762,N_14213,N_14333);
and U14763 (N_14763,N_14032,N_14209);
nor U14764 (N_14764,N_14354,N_14117);
xnor U14765 (N_14765,N_13751,N_14034);
and U14766 (N_14766,N_14232,N_13964);
xnor U14767 (N_14767,N_14035,N_14295);
or U14768 (N_14768,N_14047,N_13842);
and U14769 (N_14769,N_13996,N_14205);
xnor U14770 (N_14770,N_14079,N_13755);
nor U14771 (N_14771,N_13862,N_14108);
nand U14772 (N_14772,N_14122,N_13873);
and U14773 (N_14773,N_13809,N_14287);
nor U14774 (N_14774,N_14202,N_14161);
and U14775 (N_14775,N_14042,N_13952);
or U14776 (N_14776,N_13855,N_14197);
nand U14777 (N_14777,N_13763,N_14227);
nand U14778 (N_14778,N_14100,N_14177);
and U14779 (N_14779,N_14196,N_14117);
and U14780 (N_14780,N_13947,N_13789);
or U14781 (N_14781,N_14352,N_14089);
and U14782 (N_14782,N_14363,N_14280);
nand U14783 (N_14783,N_13826,N_13921);
nand U14784 (N_14784,N_13964,N_14131);
or U14785 (N_14785,N_13782,N_14357);
xor U14786 (N_14786,N_13972,N_13776);
nand U14787 (N_14787,N_14010,N_13998);
or U14788 (N_14788,N_14189,N_14019);
nor U14789 (N_14789,N_13770,N_14101);
and U14790 (N_14790,N_14195,N_13765);
or U14791 (N_14791,N_14288,N_14009);
and U14792 (N_14792,N_14346,N_14177);
nand U14793 (N_14793,N_14259,N_14098);
xnor U14794 (N_14794,N_13809,N_13815);
nor U14795 (N_14795,N_14365,N_13842);
nand U14796 (N_14796,N_14202,N_14189);
or U14797 (N_14797,N_13792,N_14156);
xnor U14798 (N_14798,N_14300,N_14087);
and U14799 (N_14799,N_13750,N_14278);
nor U14800 (N_14800,N_13807,N_14359);
or U14801 (N_14801,N_14155,N_13792);
nand U14802 (N_14802,N_14353,N_14118);
nand U14803 (N_14803,N_13883,N_13992);
and U14804 (N_14804,N_14204,N_14110);
nand U14805 (N_14805,N_14084,N_14342);
nand U14806 (N_14806,N_14084,N_13941);
xnor U14807 (N_14807,N_14105,N_13768);
nand U14808 (N_14808,N_13833,N_13873);
nor U14809 (N_14809,N_14357,N_13993);
nor U14810 (N_14810,N_14126,N_14357);
xor U14811 (N_14811,N_14011,N_14343);
nand U14812 (N_14812,N_13768,N_13967);
and U14813 (N_14813,N_13866,N_13889);
xor U14814 (N_14814,N_14211,N_14111);
and U14815 (N_14815,N_14337,N_13924);
nand U14816 (N_14816,N_14263,N_13827);
xnor U14817 (N_14817,N_14305,N_14001);
and U14818 (N_14818,N_14209,N_14066);
or U14819 (N_14819,N_13986,N_13783);
and U14820 (N_14820,N_14320,N_13938);
and U14821 (N_14821,N_13973,N_14264);
nor U14822 (N_14822,N_13906,N_14121);
and U14823 (N_14823,N_14119,N_14214);
xnor U14824 (N_14824,N_13986,N_14344);
nor U14825 (N_14825,N_13976,N_14002);
nand U14826 (N_14826,N_13943,N_13981);
or U14827 (N_14827,N_13761,N_14010);
nand U14828 (N_14828,N_14205,N_14134);
and U14829 (N_14829,N_14348,N_14043);
and U14830 (N_14830,N_14187,N_13889);
nor U14831 (N_14831,N_13925,N_13835);
and U14832 (N_14832,N_13808,N_14291);
nand U14833 (N_14833,N_14150,N_14086);
and U14834 (N_14834,N_13843,N_14227);
and U14835 (N_14835,N_13884,N_13766);
nand U14836 (N_14836,N_14157,N_14155);
nand U14837 (N_14837,N_13768,N_14279);
nand U14838 (N_14838,N_14150,N_13999);
nor U14839 (N_14839,N_14273,N_13993);
xor U14840 (N_14840,N_14072,N_13887);
nor U14841 (N_14841,N_14095,N_14284);
xor U14842 (N_14842,N_13780,N_13904);
nor U14843 (N_14843,N_14369,N_13846);
or U14844 (N_14844,N_14150,N_13821);
and U14845 (N_14845,N_14168,N_13953);
nor U14846 (N_14846,N_14093,N_14123);
nand U14847 (N_14847,N_14241,N_14069);
and U14848 (N_14848,N_13928,N_14237);
or U14849 (N_14849,N_13930,N_14081);
nor U14850 (N_14850,N_14000,N_13914);
or U14851 (N_14851,N_14143,N_14205);
and U14852 (N_14852,N_14001,N_13780);
and U14853 (N_14853,N_14187,N_13783);
xnor U14854 (N_14854,N_14265,N_14101);
xor U14855 (N_14855,N_14124,N_14106);
nand U14856 (N_14856,N_14023,N_14358);
or U14857 (N_14857,N_13899,N_13873);
or U14858 (N_14858,N_13936,N_14282);
xnor U14859 (N_14859,N_13818,N_14187);
xor U14860 (N_14860,N_14138,N_14215);
xor U14861 (N_14861,N_14244,N_14251);
and U14862 (N_14862,N_14058,N_13854);
and U14863 (N_14863,N_14157,N_13901);
or U14864 (N_14864,N_13900,N_14209);
and U14865 (N_14865,N_13832,N_13794);
nand U14866 (N_14866,N_13903,N_13783);
nand U14867 (N_14867,N_13879,N_13859);
or U14868 (N_14868,N_14061,N_14174);
and U14869 (N_14869,N_14196,N_14280);
or U14870 (N_14870,N_13851,N_13860);
nand U14871 (N_14871,N_14290,N_14282);
xnor U14872 (N_14872,N_14122,N_14310);
nand U14873 (N_14873,N_13761,N_14352);
nor U14874 (N_14874,N_14080,N_13819);
nand U14875 (N_14875,N_14253,N_14167);
nand U14876 (N_14876,N_14283,N_13937);
or U14877 (N_14877,N_14102,N_14201);
nor U14878 (N_14878,N_13932,N_13769);
nor U14879 (N_14879,N_14022,N_13757);
or U14880 (N_14880,N_13875,N_13920);
or U14881 (N_14881,N_13939,N_14007);
nor U14882 (N_14882,N_13866,N_13899);
and U14883 (N_14883,N_13835,N_14092);
nor U14884 (N_14884,N_14333,N_13959);
and U14885 (N_14885,N_13973,N_14138);
and U14886 (N_14886,N_14315,N_14084);
or U14887 (N_14887,N_13800,N_14117);
or U14888 (N_14888,N_14059,N_13943);
nor U14889 (N_14889,N_13762,N_14253);
and U14890 (N_14890,N_14053,N_14013);
nor U14891 (N_14891,N_14338,N_14009);
or U14892 (N_14892,N_13938,N_13760);
and U14893 (N_14893,N_14351,N_13767);
xnor U14894 (N_14894,N_14129,N_14124);
nand U14895 (N_14895,N_14204,N_13913);
xnor U14896 (N_14896,N_14193,N_14207);
and U14897 (N_14897,N_13866,N_13909);
and U14898 (N_14898,N_14320,N_14268);
or U14899 (N_14899,N_14242,N_13928);
nor U14900 (N_14900,N_14359,N_14217);
and U14901 (N_14901,N_14368,N_14276);
and U14902 (N_14902,N_14132,N_14078);
and U14903 (N_14903,N_14355,N_14044);
and U14904 (N_14904,N_14158,N_14004);
xnor U14905 (N_14905,N_14105,N_14167);
and U14906 (N_14906,N_13916,N_13892);
xor U14907 (N_14907,N_13794,N_13761);
and U14908 (N_14908,N_14111,N_13836);
nor U14909 (N_14909,N_13980,N_14090);
and U14910 (N_14910,N_13755,N_14060);
or U14911 (N_14911,N_14166,N_13822);
xor U14912 (N_14912,N_14171,N_14033);
and U14913 (N_14913,N_13765,N_13898);
or U14914 (N_14914,N_14345,N_14323);
nand U14915 (N_14915,N_14309,N_14370);
xnor U14916 (N_14916,N_13851,N_14211);
nand U14917 (N_14917,N_13865,N_14239);
xnor U14918 (N_14918,N_13911,N_14350);
xor U14919 (N_14919,N_14337,N_14358);
nand U14920 (N_14920,N_13787,N_14241);
or U14921 (N_14921,N_13857,N_14334);
and U14922 (N_14922,N_14355,N_14321);
nor U14923 (N_14923,N_13761,N_14259);
or U14924 (N_14924,N_13968,N_13831);
nand U14925 (N_14925,N_14294,N_13941);
nand U14926 (N_14926,N_14018,N_13825);
and U14927 (N_14927,N_13751,N_13784);
xnor U14928 (N_14928,N_14305,N_14077);
and U14929 (N_14929,N_14326,N_14021);
xnor U14930 (N_14930,N_13773,N_13899);
nand U14931 (N_14931,N_14232,N_14137);
nand U14932 (N_14932,N_13785,N_14194);
xnor U14933 (N_14933,N_14338,N_13915);
nand U14934 (N_14934,N_14363,N_14119);
or U14935 (N_14935,N_14230,N_14158);
xnor U14936 (N_14936,N_14172,N_14054);
or U14937 (N_14937,N_13949,N_14272);
nand U14938 (N_14938,N_14179,N_14137);
nor U14939 (N_14939,N_14033,N_14310);
and U14940 (N_14940,N_13926,N_13885);
nor U14941 (N_14941,N_14135,N_13916);
nor U14942 (N_14942,N_14356,N_13772);
nor U14943 (N_14943,N_14308,N_14163);
xor U14944 (N_14944,N_14266,N_14045);
nor U14945 (N_14945,N_14064,N_13896);
or U14946 (N_14946,N_14131,N_13803);
or U14947 (N_14947,N_14304,N_13755);
and U14948 (N_14948,N_13995,N_14167);
nand U14949 (N_14949,N_14183,N_14059);
nand U14950 (N_14950,N_14263,N_14282);
nor U14951 (N_14951,N_14192,N_14142);
or U14952 (N_14952,N_14363,N_14178);
or U14953 (N_14953,N_13995,N_13810);
or U14954 (N_14954,N_14234,N_14271);
xor U14955 (N_14955,N_14138,N_13965);
xor U14956 (N_14956,N_14341,N_13968);
or U14957 (N_14957,N_14329,N_14066);
nor U14958 (N_14958,N_14254,N_14038);
nor U14959 (N_14959,N_14201,N_14174);
or U14960 (N_14960,N_14145,N_13928);
nand U14961 (N_14961,N_13895,N_14110);
or U14962 (N_14962,N_13900,N_14011);
nand U14963 (N_14963,N_14220,N_14184);
and U14964 (N_14964,N_13807,N_14040);
nor U14965 (N_14965,N_14224,N_14056);
or U14966 (N_14966,N_14363,N_14089);
nand U14967 (N_14967,N_13912,N_13808);
and U14968 (N_14968,N_14149,N_14225);
nor U14969 (N_14969,N_13903,N_14233);
nor U14970 (N_14970,N_14278,N_13839);
nand U14971 (N_14971,N_13880,N_13791);
and U14972 (N_14972,N_14000,N_14240);
and U14973 (N_14973,N_14042,N_14068);
nand U14974 (N_14974,N_14188,N_14006);
nor U14975 (N_14975,N_14278,N_13978);
nand U14976 (N_14976,N_13850,N_14296);
xor U14977 (N_14977,N_14044,N_14313);
nor U14978 (N_14978,N_14287,N_14262);
or U14979 (N_14979,N_14300,N_13888);
nand U14980 (N_14980,N_14261,N_14066);
xnor U14981 (N_14981,N_14165,N_14354);
or U14982 (N_14982,N_13821,N_14092);
xor U14983 (N_14983,N_14142,N_14076);
or U14984 (N_14984,N_14076,N_14081);
xnor U14985 (N_14985,N_14219,N_13894);
xnor U14986 (N_14986,N_13883,N_14068);
and U14987 (N_14987,N_13824,N_13865);
nand U14988 (N_14988,N_14085,N_13955);
and U14989 (N_14989,N_13976,N_14279);
xnor U14990 (N_14990,N_14053,N_14048);
xnor U14991 (N_14991,N_13853,N_13951);
xor U14992 (N_14992,N_14240,N_13819);
nor U14993 (N_14993,N_13984,N_14316);
xnor U14994 (N_14994,N_13801,N_14011);
and U14995 (N_14995,N_14315,N_13889);
or U14996 (N_14996,N_14299,N_13877);
xnor U14997 (N_14997,N_14300,N_13855);
xnor U14998 (N_14998,N_14178,N_14117);
nor U14999 (N_14999,N_14090,N_13906);
xnor U15000 (N_15000,N_14635,N_14995);
nand U15001 (N_15001,N_14875,N_14741);
and U15002 (N_15002,N_14726,N_14891);
xor U15003 (N_15003,N_14547,N_14833);
or U15004 (N_15004,N_14558,N_14944);
nand U15005 (N_15005,N_14950,N_14821);
or U15006 (N_15006,N_14556,N_14988);
and U15007 (N_15007,N_14610,N_14529);
xor U15008 (N_15008,N_14580,N_14502);
nand U15009 (N_15009,N_14861,N_14870);
nor U15010 (N_15010,N_14649,N_14605);
nor U15011 (N_15011,N_14800,N_14923);
xnor U15012 (N_15012,N_14485,N_14948);
xor U15013 (N_15013,N_14664,N_14389);
and U15014 (N_15014,N_14492,N_14714);
nor U15015 (N_15015,N_14673,N_14447);
nand U15016 (N_15016,N_14657,N_14983);
nor U15017 (N_15017,N_14534,N_14849);
xnor U15018 (N_15018,N_14907,N_14910);
xnor U15019 (N_15019,N_14515,N_14552);
or U15020 (N_15020,N_14382,N_14452);
xnor U15021 (N_15021,N_14810,N_14520);
xor U15022 (N_15022,N_14876,N_14507);
xor U15023 (N_15023,N_14844,N_14874);
or U15024 (N_15024,N_14450,N_14981);
and U15025 (N_15025,N_14393,N_14932);
nand U15026 (N_15026,N_14665,N_14440);
xor U15027 (N_15027,N_14648,N_14766);
or U15028 (N_15028,N_14873,N_14445);
and U15029 (N_15029,N_14390,N_14656);
nor U15030 (N_15030,N_14585,N_14544);
nand U15031 (N_15031,N_14623,N_14476);
nor U15032 (N_15032,N_14663,N_14410);
and U15033 (N_15033,N_14537,N_14750);
nand U15034 (N_15034,N_14512,N_14557);
and U15035 (N_15035,N_14900,N_14666);
or U15036 (N_15036,N_14715,N_14501);
or U15037 (N_15037,N_14942,N_14961);
and U15038 (N_15038,N_14417,N_14830);
and U15039 (N_15039,N_14574,N_14508);
xor U15040 (N_15040,N_14409,N_14818);
nand U15041 (N_15041,N_14549,N_14444);
and U15042 (N_15042,N_14438,N_14634);
and U15043 (N_15043,N_14879,N_14587);
or U15044 (N_15044,N_14839,N_14647);
nand U15045 (N_15045,N_14639,N_14397);
nand U15046 (N_15046,N_14769,N_14976);
nand U15047 (N_15047,N_14560,N_14985);
nand U15048 (N_15048,N_14434,N_14436);
or U15049 (N_15049,N_14866,N_14676);
and U15050 (N_15050,N_14624,N_14783);
xor U15051 (N_15051,N_14472,N_14883);
xor U15052 (N_15052,N_14483,N_14926);
and U15053 (N_15053,N_14375,N_14475);
nand U15054 (N_15054,N_14765,N_14841);
and U15055 (N_15055,N_14531,N_14627);
nand U15056 (N_15056,N_14572,N_14615);
and U15057 (N_15057,N_14380,N_14859);
and U15058 (N_15058,N_14947,N_14752);
or U15059 (N_15059,N_14723,N_14897);
xnor U15060 (N_15060,N_14621,N_14898);
nor U15061 (N_15061,N_14736,N_14761);
nand U15062 (N_15062,N_14743,N_14806);
xnor U15063 (N_15063,N_14809,N_14601);
xnor U15064 (N_15064,N_14376,N_14681);
and U15065 (N_15065,N_14916,N_14845);
nand U15066 (N_15066,N_14862,N_14790);
nor U15067 (N_15067,N_14396,N_14991);
nor U15068 (N_15068,N_14786,N_14685);
or U15069 (N_15069,N_14922,N_14598);
nand U15070 (N_15070,N_14645,N_14398);
and U15071 (N_15071,N_14509,N_14578);
xnor U15072 (N_15072,N_14887,N_14734);
and U15073 (N_15073,N_14513,N_14427);
or U15074 (N_15074,N_14764,N_14654);
xor U15075 (N_15075,N_14488,N_14928);
nor U15076 (N_15076,N_14545,N_14419);
nor U15077 (N_15077,N_14586,N_14962);
nor U15078 (N_15078,N_14827,N_14391);
nand U15079 (N_15079,N_14538,N_14936);
nor U15080 (N_15080,N_14933,N_14780);
nor U15081 (N_15081,N_14795,N_14503);
or U15082 (N_15082,N_14680,N_14405);
and U15083 (N_15083,N_14996,N_14459);
or U15084 (N_15084,N_14804,N_14642);
and U15085 (N_15085,N_14829,N_14671);
or U15086 (N_15086,N_14379,N_14805);
xor U15087 (N_15087,N_14994,N_14798);
nor U15088 (N_15088,N_14954,N_14668);
or U15089 (N_15089,N_14834,N_14869);
nand U15090 (N_15090,N_14978,N_14500);
nor U15091 (N_15091,N_14729,N_14628);
and U15092 (N_15092,N_14892,N_14888);
nor U15093 (N_15093,N_14791,N_14394);
or U15094 (N_15094,N_14696,N_14757);
nor U15095 (N_15095,N_14963,N_14816);
and U15096 (N_15096,N_14386,N_14902);
or U15097 (N_15097,N_14388,N_14644);
and U15098 (N_15098,N_14530,N_14630);
nor U15099 (N_15099,N_14579,N_14739);
nand U15100 (N_15100,N_14969,N_14808);
xnor U15101 (N_15101,N_14895,N_14385);
xor U15102 (N_15102,N_14433,N_14826);
nor U15103 (N_15103,N_14784,N_14911);
nor U15104 (N_15104,N_14486,N_14838);
nand U15105 (N_15105,N_14555,N_14442);
or U15106 (N_15106,N_14925,N_14774);
xnor U15107 (N_15107,N_14720,N_14918);
and U15108 (N_15108,N_14504,N_14992);
nand U15109 (N_15109,N_14421,N_14612);
xor U15110 (N_15110,N_14506,N_14480);
and U15111 (N_15111,N_14518,N_14464);
and U15112 (N_15112,N_14903,N_14675);
or U15113 (N_15113,N_14406,N_14958);
nand U15114 (N_15114,N_14904,N_14770);
xor U15115 (N_15115,N_14441,N_14446);
and U15116 (N_15116,N_14777,N_14599);
and U15117 (N_15117,N_14470,N_14987);
nor U15118 (N_15118,N_14746,N_14825);
xor U15119 (N_15119,N_14575,N_14443);
nand U15120 (N_15120,N_14835,N_14411);
and U15121 (N_15121,N_14539,N_14408);
or U15122 (N_15122,N_14738,N_14456);
nor U15123 (N_15123,N_14522,N_14425);
nor U15124 (N_15124,N_14953,N_14707);
xor U15125 (N_15125,N_14453,N_14955);
or U15126 (N_15126,N_14633,N_14940);
and U15127 (N_15127,N_14863,N_14617);
or U15128 (N_15128,N_14528,N_14758);
and U15129 (N_15129,N_14687,N_14814);
and U15130 (N_15130,N_14966,N_14751);
nor U15131 (N_15131,N_14619,N_14709);
nor U15132 (N_15132,N_14763,N_14819);
or U15133 (N_15133,N_14519,N_14993);
or U15134 (N_15134,N_14867,N_14716);
nand U15135 (N_15135,N_14677,N_14896);
and U15136 (N_15136,N_14855,N_14820);
or U15137 (N_15137,N_14889,N_14594);
or U15138 (N_15138,N_14514,N_14740);
nand U15139 (N_15139,N_14546,N_14454);
nand U15140 (N_15140,N_14971,N_14455);
or U15141 (N_15141,N_14864,N_14625);
nand U15142 (N_15142,N_14626,N_14817);
or U15143 (N_15143,N_14779,N_14510);
and U15144 (N_15144,N_14679,N_14516);
xnor U15145 (N_15145,N_14699,N_14846);
nor U15146 (N_15146,N_14517,N_14813);
nor U15147 (N_15147,N_14597,N_14583);
xnor U15148 (N_15148,N_14882,N_14384);
or U15149 (N_15149,N_14998,N_14553);
xnor U15150 (N_15150,N_14793,N_14493);
nor U15151 (N_15151,N_14692,N_14865);
and U15152 (N_15152,N_14484,N_14497);
and U15153 (N_15153,N_14400,N_14785);
nor U15154 (N_15154,N_14551,N_14850);
xor U15155 (N_15155,N_14693,N_14908);
xor U15156 (N_15156,N_14781,N_14684);
nor U15157 (N_15157,N_14979,N_14670);
and U15158 (N_15158,N_14650,N_14423);
and U15159 (N_15159,N_14886,N_14802);
and U15160 (N_15160,N_14872,N_14489);
or U15161 (N_15161,N_14689,N_14525);
or U15162 (N_15162,N_14986,N_14837);
xnor U15163 (N_15163,N_14713,N_14392);
nor U15164 (N_15164,N_14843,N_14458);
and U15165 (N_15165,N_14694,N_14956);
or U15166 (N_15166,N_14473,N_14402);
nor U15167 (N_15167,N_14468,N_14749);
nor U15168 (N_15168,N_14554,N_14768);
and U15169 (N_15169,N_14951,N_14678);
nand U15170 (N_15170,N_14964,N_14616);
nand U15171 (N_15171,N_14906,N_14611);
nand U15172 (N_15172,N_14767,N_14487);
nor U15173 (N_15173,N_14430,N_14705);
nor U15174 (N_15174,N_14762,N_14658);
xnor U15175 (N_15175,N_14852,N_14822);
and U15176 (N_15176,N_14941,N_14403);
nor U15177 (N_15177,N_14420,N_14466);
xor U15178 (N_15178,N_14478,N_14968);
or U15179 (N_15179,N_14915,N_14881);
xnor U15180 (N_15180,N_14532,N_14686);
and U15181 (N_15181,N_14660,N_14812);
or U15182 (N_15182,N_14416,N_14573);
and U15183 (N_15183,N_14935,N_14797);
and U15184 (N_15184,N_14943,N_14776);
and U15185 (N_15185,N_14383,N_14710);
nor U15186 (N_15186,N_14412,N_14989);
nand U15187 (N_15187,N_14490,N_14429);
and U15188 (N_15188,N_14931,N_14930);
or U15189 (N_15189,N_14496,N_14727);
nand U15190 (N_15190,N_14787,N_14742);
or U15191 (N_15191,N_14788,N_14701);
and U15192 (N_15192,N_14526,N_14595);
nand U15193 (N_15193,N_14600,N_14377);
or U15194 (N_15194,N_14609,N_14945);
or U15195 (N_15195,N_14494,N_14858);
xor U15196 (N_15196,N_14719,N_14772);
nand U15197 (N_15197,N_14857,N_14773);
or U15198 (N_15198,N_14655,N_14728);
nor U15199 (N_15199,N_14498,N_14744);
and U15200 (N_15200,N_14499,N_14541);
xor U15201 (N_15201,N_14414,N_14570);
or U15202 (N_15202,N_14533,N_14691);
nand U15203 (N_15203,N_14461,N_14927);
nor U15204 (N_15204,N_14880,N_14982);
nor U15205 (N_15205,N_14620,N_14702);
and U15206 (N_15206,N_14721,N_14563);
and U15207 (N_15207,N_14540,N_14973);
nand U15208 (N_15208,N_14511,N_14437);
or U15209 (N_15209,N_14878,N_14815);
and U15210 (N_15210,N_14856,N_14413);
or U15211 (N_15211,N_14637,N_14682);
nand U15212 (N_15212,N_14934,N_14536);
xnor U15213 (N_15213,N_14548,N_14792);
or U15214 (N_15214,N_14471,N_14789);
xnor U15215 (N_15215,N_14667,N_14596);
and U15216 (N_15216,N_14439,N_14724);
nand U15217 (N_15217,N_14571,N_14424);
or U15218 (N_15218,N_14703,N_14463);
and U15219 (N_15219,N_14823,N_14618);
and U15220 (N_15220,N_14604,N_14708);
xnor U15221 (N_15221,N_14460,N_14877);
nor U15222 (N_15222,N_14569,N_14733);
or U15223 (N_15223,N_14491,N_14695);
nand U15224 (N_15224,N_14426,N_14381);
xnor U15225 (N_15225,N_14836,N_14451);
nor U15226 (N_15226,N_14431,N_14568);
nand U15227 (N_15227,N_14760,N_14807);
or U15228 (N_15228,N_14975,N_14576);
xnor U15229 (N_15229,N_14632,N_14672);
nor U15230 (N_15230,N_14999,N_14588);
and U15231 (N_15231,N_14893,N_14965);
xor U15232 (N_15232,N_14775,N_14737);
nand U15233 (N_15233,N_14824,N_14730);
xnor U15234 (N_15234,N_14957,N_14567);
or U15235 (N_15235,N_14909,N_14479);
and U15236 (N_15236,N_14828,N_14755);
xor U15237 (N_15237,N_14745,N_14946);
xnor U15238 (N_15238,N_14984,N_14467);
and U15239 (N_15239,N_14854,N_14629);
nand U15240 (N_15240,N_14415,N_14495);
xnor U15241 (N_15241,N_14613,N_14832);
or U15242 (N_15242,N_14698,N_14581);
nor U15243 (N_15243,N_14614,N_14748);
and U15244 (N_15244,N_14938,N_14564);
nand U15245 (N_15245,N_14735,N_14469);
xor U15246 (N_15246,N_14462,N_14700);
nor U15247 (N_15247,N_14924,N_14477);
nor U15248 (N_15248,N_14523,N_14378);
or U15249 (N_15249,N_14646,N_14937);
or U15250 (N_15250,N_14591,N_14972);
xor U15251 (N_15251,N_14921,N_14662);
or U15252 (N_15252,N_14606,N_14917);
and U15253 (N_15253,N_14640,N_14593);
and U15254 (N_15254,N_14607,N_14725);
xor U15255 (N_15255,N_14592,N_14884);
nor U15256 (N_15256,N_14566,N_14542);
nand U15257 (N_15257,N_14997,N_14561);
nand U15258 (N_15258,N_14659,N_14717);
and U15259 (N_15259,N_14885,N_14914);
and U15260 (N_15260,N_14505,N_14527);
and U15261 (N_15261,N_14919,N_14712);
and U15262 (N_15262,N_14401,N_14688);
nand U15263 (N_15263,N_14731,N_14465);
nand U15264 (N_15264,N_14949,N_14706);
and U15265 (N_15265,N_14890,N_14894);
nor U15266 (N_15266,N_14474,N_14589);
nand U15267 (N_15267,N_14543,N_14718);
and U15268 (N_15268,N_14771,N_14481);
nand U15269 (N_15269,N_14636,N_14435);
xnor U15270 (N_15270,N_14747,N_14562);
xor U15271 (N_15271,N_14603,N_14754);
and U15272 (N_15272,N_14697,N_14550);
and U15273 (N_15273,N_14559,N_14868);
and U15274 (N_15274,N_14448,N_14722);
xor U15275 (N_15275,N_14418,N_14905);
and U15276 (N_15276,N_14799,N_14669);
and U15277 (N_15277,N_14831,N_14395);
nand U15278 (N_15278,N_14960,N_14959);
nand U15279 (N_15279,N_14848,N_14801);
xor U15280 (N_15280,N_14652,N_14977);
xnor U15281 (N_15281,N_14860,N_14428);
and U15282 (N_15282,N_14638,N_14590);
nand U15283 (N_15283,N_14952,N_14732);
nor U15284 (N_15284,N_14811,N_14967);
or U15285 (N_15285,N_14794,N_14651);
and U15286 (N_15286,N_14704,N_14577);
xor U15287 (N_15287,N_14929,N_14674);
or U15288 (N_15288,N_14399,N_14840);
nor U15289 (N_15289,N_14803,N_14387);
nand U15290 (N_15290,N_14990,N_14901);
and U15291 (N_15291,N_14683,N_14535);
and U15292 (N_15292,N_14939,N_14482);
or U15293 (N_15293,N_14602,N_14641);
nand U15294 (N_15294,N_14920,N_14404);
and U15295 (N_15295,N_14449,N_14871);
nor U15296 (N_15296,N_14753,N_14521);
xor U15297 (N_15297,N_14643,N_14653);
or U15298 (N_15298,N_14974,N_14970);
nor U15299 (N_15299,N_14912,N_14690);
nand U15300 (N_15300,N_14584,N_14759);
nand U15301 (N_15301,N_14407,N_14565);
xor U15302 (N_15302,N_14899,N_14847);
and U15303 (N_15303,N_14432,N_14796);
and U15304 (N_15304,N_14853,N_14913);
nor U15305 (N_15305,N_14711,N_14756);
nor U15306 (N_15306,N_14631,N_14457);
xnor U15307 (N_15307,N_14622,N_14842);
nand U15308 (N_15308,N_14778,N_14582);
nand U15309 (N_15309,N_14661,N_14851);
xor U15310 (N_15310,N_14422,N_14524);
nand U15311 (N_15311,N_14782,N_14608);
and U15312 (N_15312,N_14980,N_14971);
and U15313 (N_15313,N_14654,N_14975);
xor U15314 (N_15314,N_14944,N_14859);
nand U15315 (N_15315,N_14761,N_14954);
nand U15316 (N_15316,N_14615,N_14830);
xor U15317 (N_15317,N_14477,N_14576);
nor U15318 (N_15318,N_14531,N_14666);
nand U15319 (N_15319,N_14731,N_14548);
and U15320 (N_15320,N_14661,N_14830);
nor U15321 (N_15321,N_14497,N_14861);
nand U15322 (N_15322,N_14400,N_14901);
xor U15323 (N_15323,N_14395,N_14900);
nor U15324 (N_15324,N_14852,N_14779);
nor U15325 (N_15325,N_14717,N_14962);
and U15326 (N_15326,N_14758,N_14446);
nor U15327 (N_15327,N_14947,N_14823);
and U15328 (N_15328,N_14634,N_14899);
xnor U15329 (N_15329,N_14763,N_14889);
nand U15330 (N_15330,N_14573,N_14895);
or U15331 (N_15331,N_14781,N_14919);
xor U15332 (N_15332,N_14891,N_14916);
nor U15333 (N_15333,N_14602,N_14394);
xor U15334 (N_15334,N_14536,N_14390);
xor U15335 (N_15335,N_14656,N_14795);
nand U15336 (N_15336,N_14380,N_14892);
or U15337 (N_15337,N_14762,N_14404);
nor U15338 (N_15338,N_14757,N_14971);
or U15339 (N_15339,N_14814,N_14435);
nor U15340 (N_15340,N_14389,N_14848);
nor U15341 (N_15341,N_14656,N_14433);
nor U15342 (N_15342,N_14924,N_14915);
or U15343 (N_15343,N_14846,N_14955);
and U15344 (N_15344,N_14469,N_14731);
or U15345 (N_15345,N_14797,N_14696);
nor U15346 (N_15346,N_14826,N_14974);
xnor U15347 (N_15347,N_14585,N_14623);
and U15348 (N_15348,N_14572,N_14753);
or U15349 (N_15349,N_14411,N_14515);
nand U15350 (N_15350,N_14458,N_14854);
and U15351 (N_15351,N_14854,N_14517);
xor U15352 (N_15352,N_14576,N_14616);
xor U15353 (N_15353,N_14911,N_14729);
xor U15354 (N_15354,N_14498,N_14402);
and U15355 (N_15355,N_14701,N_14673);
nor U15356 (N_15356,N_14820,N_14497);
xnor U15357 (N_15357,N_14755,N_14873);
nor U15358 (N_15358,N_14749,N_14541);
and U15359 (N_15359,N_14523,N_14542);
or U15360 (N_15360,N_14723,N_14736);
nand U15361 (N_15361,N_14967,N_14669);
nand U15362 (N_15362,N_14730,N_14614);
and U15363 (N_15363,N_14902,N_14734);
or U15364 (N_15364,N_14386,N_14573);
or U15365 (N_15365,N_14904,N_14738);
nand U15366 (N_15366,N_14496,N_14638);
nand U15367 (N_15367,N_14388,N_14716);
or U15368 (N_15368,N_14876,N_14535);
and U15369 (N_15369,N_14633,N_14939);
and U15370 (N_15370,N_14421,N_14842);
nand U15371 (N_15371,N_14791,N_14387);
xor U15372 (N_15372,N_14745,N_14412);
nor U15373 (N_15373,N_14793,N_14752);
or U15374 (N_15374,N_14635,N_14387);
or U15375 (N_15375,N_14703,N_14592);
nand U15376 (N_15376,N_14919,N_14739);
nor U15377 (N_15377,N_14750,N_14820);
nor U15378 (N_15378,N_14824,N_14497);
xor U15379 (N_15379,N_14610,N_14571);
nand U15380 (N_15380,N_14606,N_14573);
xnor U15381 (N_15381,N_14660,N_14415);
nor U15382 (N_15382,N_14851,N_14722);
or U15383 (N_15383,N_14853,N_14469);
nor U15384 (N_15384,N_14963,N_14651);
and U15385 (N_15385,N_14731,N_14870);
nand U15386 (N_15386,N_14644,N_14791);
xnor U15387 (N_15387,N_14966,N_14911);
xnor U15388 (N_15388,N_14720,N_14983);
xor U15389 (N_15389,N_14722,N_14504);
and U15390 (N_15390,N_14573,N_14398);
nor U15391 (N_15391,N_14714,N_14937);
nand U15392 (N_15392,N_14970,N_14526);
nand U15393 (N_15393,N_14490,N_14491);
nor U15394 (N_15394,N_14757,N_14966);
nor U15395 (N_15395,N_14721,N_14634);
xor U15396 (N_15396,N_14586,N_14766);
xor U15397 (N_15397,N_14933,N_14801);
nor U15398 (N_15398,N_14400,N_14985);
nand U15399 (N_15399,N_14653,N_14803);
and U15400 (N_15400,N_14465,N_14930);
and U15401 (N_15401,N_14775,N_14492);
nor U15402 (N_15402,N_14701,N_14679);
or U15403 (N_15403,N_14419,N_14510);
nor U15404 (N_15404,N_14424,N_14405);
and U15405 (N_15405,N_14718,N_14606);
nand U15406 (N_15406,N_14889,N_14691);
or U15407 (N_15407,N_14927,N_14751);
xnor U15408 (N_15408,N_14860,N_14900);
nor U15409 (N_15409,N_14597,N_14761);
or U15410 (N_15410,N_14859,N_14387);
and U15411 (N_15411,N_14891,N_14485);
nor U15412 (N_15412,N_14560,N_14839);
or U15413 (N_15413,N_14450,N_14445);
or U15414 (N_15414,N_14943,N_14503);
nand U15415 (N_15415,N_14971,N_14897);
xnor U15416 (N_15416,N_14915,N_14850);
or U15417 (N_15417,N_14534,N_14639);
or U15418 (N_15418,N_14622,N_14512);
and U15419 (N_15419,N_14657,N_14976);
nand U15420 (N_15420,N_14462,N_14733);
nand U15421 (N_15421,N_14402,N_14415);
or U15422 (N_15422,N_14936,N_14937);
xor U15423 (N_15423,N_14866,N_14689);
nor U15424 (N_15424,N_14973,N_14603);
xnor U15425 (N_15425,N_14962,N_14440);
nand U15426 (N_15426,N_14791,N_14397);
xnor U15427 (N_15427,N_14673,N_14956);
xnor U15428 (N_15428,N_14950,N_14699);
nor U15429 (N_15429,N_14665,N_14625);
or U15430 (N_15430,N_14851,N_14852);
and U15431 (N_15431,N_14507,N_14791);
nor U15432 (N_15432,N_14714,N_14837);
xnor U15433 (N_15433,N_14647,N_14825);
xor U15434 (N_15434,N_14609,N_14555);
or U15435 (N_15435,N_14780,N_14549);
nand U15436 (N_15436,N_14422,N_14696);
xnor U15437 (N_15437,N_14390,N_14594);
and U15438 (N_15438,N_14639,N_14935);
nand U15439 (N_15439,N_14470,N_14423);
and U15440 (N_15440,N_14991,N_14598);
nand U15441 (N_15441,N_14411,N_14783);
and U15442 (N_15442,N_14864,N_14619);
xnor U15443 (N_15443,N_14398,N_14782);
and U15444 (N_15444,N_14740,N_14765);
and U15445 (N_15445,N_14869,N_14816);
and U15446 (N_15446,N_14479,N_14743);
xor U15447 (N_15447,N_14614,N_14975);
nand U15448 (N_15448,N_14619,N_14951);
nand U15449 (N_15449,N_14697,N_14922);
and U15450 (N_15450,N_14964,N_14958);
xor U15451 (N_15451,N_14966,N_14846);
and U15452 (N_15452,N_14978,N_14732);
nor U15453 (N_15453,N_14935,N_14832);
and U15454 (N_15454,N_14637,N_14906);
nand U15455 (N_15455,N_14733,N_14685);
xor U15456 (N_15456,N_14616,N_14851);
xor U15457 (N_15457,N_14748,N_14611);
xnor U15458 (N_15458,N_14862,N_14963);
and U15459 (N_15459,N_14655,N_14552);
or U15460 (N_15460,N_14823,N_14444);
and U15461 (N_15461,N_14565,N_14840);
or U15462 (N_15462,N_14425,N_14587);
or U15463 (N_15463,N_14694,N_14652);
xor U15464 (N_15464,N_14842,N_14711);
or U15465 (N_15465,N_14898,N_14697);
nand U15466 (N_15466,N_14431,N_14863);
or U15467 (N_15467,N_14567,N_14935);
and U15468 (N_15468,N_14561,N_14884);
nand U15469 (N_15469,N_14728,N_14726);
and U15470 (N_15470,N_14398,N_14947);
or U15471 (N_15471,N_14983,N_14607);
and U15472 (N_15472,N_14602,N_14791);
xnor U15473 (N_15473,N_14978,N_14969);
nand U15474 (N_15474,N_14477,N_14811);
xor U15475 (N_15475,N_14885,N_14810);
nor U15476 (N_15476,N_14784,N_14452);
nor U15477 (N_15477,N_14951,N_14995);
and U15478 (N_15478,N_14734,N_14830);
xnor U15479 (N_15479,N_14851,N_14797);
nand U15480 (N_15480,N_14778,N_14421);
or U15481 (N_15481,N_14870,N_14397);
nor U15482 (N_15482,N_14582,N_14683);
nand U15483 (N_15483,N_14890,N_14885);
nor U15484 (N_15484,N_14867,N_14429);
and U15485 (N_15485,N_14949,N_14538);
nand U15486 (N_15486,N_14921,N_14772);
or U15487 (N_15487,N_14978,N_14970);
or U15488 (N_15488,N_14774,N_14946);
nand U15489 (N_15489,N_14553,N_14564);
and U15490 (N_15490,N_14388,N_14847);
nor U15491 (N_15491,N_14740,N_14560);
or U15492 (N_15492,N_14815,N_14417);
nor U15493 (N_15493,N_14899,N_14844);
and U15494 (N_15494,N_14429,N_14912);
nor U15495 (N_15495,N_14685,N_14833);
and U15496 (N_15496,N_14400,N_14868);
nand U15497 (N_15497,N_14451,N_14434);
xor U15498 (N_15498,N_14471,N_14967);
xnor U15499 (N_15499,N_14735,N_14841);
or U15500 (N_15500,N_14846,N_14839);
xor U15501 (N_15501,N_14760,N_14866);
nor U15502 (N_15502,N_14799,N_14461);
nor U15503 (N_15503,N_14455,N_14988);
or U15504 (N_15504,N_14794,N_14616);
nor U15505 (N_15505,N_14765,N_14891);
nor U15506 (N_15506,N_14613,N_14979);
and U15507 (N_15507,N_14501,N_14713);
and U15508 (N_15508,N_14919,N_14813);
and U15509 (N_15509,N_14457,N_14649);
and U15510 (N_15510,N_14462,N_14408);
nor U15511 (N_15511,N_14848,N_14831);
xnor U15512 (N_15512,N_14818,N_14459);
nand U15513 (N_15513,N_14420,N_14933);
and U15514 (N_15514,N_14713,N_14482);
xor U15515 (N_15515,N_14956,N_14786);
or U15516 (N_15516,N_14817,N_14793);
or U15517 (N_15517,N_14738,N_14987);
xnor U15518 (N_15518,N_14913,N_14792);
nor U15519 (N_15519,N_14755,N_14904);
and U15520 (N_15520,N_14443,N_14461);
nor U15521 (N_15521,N_14997,N_14569);
nand U15522 (N_15522,N_14704,N_14852);
and U15523 (N_15523,N_14587,N_14719);
nor U15524 (N_15524,N_14946,N_14852);
nand U15525 (N_15525,N_14975,N_14981);
or U15526 (N_15526,N_14719,N_14488);
or U15527 (N_15527,N_14428,N_14848);
and U15528 (N_15528,N_14909,N_14994);
or U15529 (N_15529,N_14643,N_14456);
nand U15530 (N_15530,N_14688,N_14474);
nand U15531 (N_15531,N_14691,N_14666);
or U15532 (N_15532,N_14877,N_14543);
and U15533 (N_15533,N_14448,N_14411);
or U15534 (N_15534,N_14545,N_14584);
nor U15535 (N_15535,N_14686,N_14408);
nor U15536 (N_15536,N_14432,N_14910);
nor U15537 (N_15537,N_14930,N_14765);
nand U15538 (N_15538,N_14995,N_14850);
or U15539 (N_15539,N_14573,N_14553);
nor U15540 (N_15540,N_14492,N_14766);
and U15541 (N_15541,N_14772,N_14940);
nand U15542 (N_15542,N_14483,N_14663);
xor U15543 (N_15543,N_14928,N_14449);
or U15544 (N_15544,N_14809,N_14924);
nand U15545 (N_15545,N_14953,N_14517);
xnor U15546 (N_15546,N_14882,N_14922);
nand U15547 (N_15547,N_14468,N_14488);
and U15548 (N_15548,N_14873,N_14861);
nand U15549 (N_15549,N_14639,N_14540);
and U15550 (N_15550,N_14918,N_14832);
and U15551 (N_15551,N_14826,N_14569);
nor U15552 (N_15552,N_14759,N_14739);
nor U15553 (N_15553,N_14937,N_14626);
xnor U15554 (N_15554,N_14451,N_14817);
nand U15555 (N_15555,N_14684,N_14640);
xnor U15556 (N_15556,N_14801,N_14578);
xnor U15557 (N_15557,N_14872,N_14894);
or U15558 (N_15558,N_14385,N_14491);
xnor U15559 (N_15559,N_14693,N_14942);
xnor U15560 (N_15560,N_14556,N_14523);
nor U15561 (N_15561,N_14940,N_14414);
nor U15562 (N_15562,N_14640,N_14384);
nand U15563 (N_15563,N_14561,N_14413);
xor U15564 (N_15564,N_14526,N_14770);
and U15565 (N_15565,N_14517,N_14814);
and U15566 (N_15566,N_14834,N_14550);
or U15567 (N_15567,N_14689,N_14867);
or U15568 (N_15568,N_14825,N_14882);
and U15569 (N_15569,N_14531,N_14526);
and U15570 (N_15570,N_14933,N_14965);
xor U15571 (N_15571,N_14714,N_14863);
or U15572 (N_15572,N_14989,N_14623);
xor U15573 (N_15573,N_14700,N_14684);
and U15574 (N_15574,N_14735,N_14713);
nand U15575 (N_15575,N_14831,N_14946);
nand U15576 (N_15576,N_14624,N_14677);
nor U15577 (N_15577,N_14501,N_14384);
or U15578 (N_15578,N_14696,N_14521);
and U15579 (N_15579,N_14668,N_14903);
xor U15580 (N_15580,N_14422,N_14406);
xnor U15581 (N_15581,N_14980,N_14487);
or U15582 (N_15582,N_14642,N_14389);
and U15583 (N_15583,N_14472,N_14719);
and U15584 (N_15584,N_14664,N_14815);
or U15585 (N_15585,N_14420,N_14402);
nor U15586 (N_15586,N_14522,N_14408);
or U15587 (N_15587,N_14884,N_14736);
nor U15588 (N_15588,N_14643,N_14666);
xnor U15589 (N_15589,N_14719,N_14596);
nor U15590 (N_15590,N_14424,N_14533);
and U15591 (N_15591,N_14892,N_14540);
and U15592 (N_15592,N_14473,N_14852);
or U15593 (N_15593,N_14757,N_14862);
and U15594 (N_15594,N_14727,N_14693);
nor U15595 (N_15595,N_14762,N_14495);
nand U15596 (N_15596,N_14751,N_14430);
nor U15597 (N_15597,N_14825,N_14723);
nor U15598 (N_15598,N_14464,N_14945);
nor U15599 (N_15599,N_14393,N_14536);
or U15600 (N_15600,N_14910,N_14461);
nor U15601 (N_15601,N_14395,N_14398);
or U15602 (N_15602,N_14580,N_14507);
xnor U15603 (N_15603,N_14574,N_14969);
xnor U15604 (N_15604,N_14491,N_14589);
and U15605 (N_15605,N_14526,N_14626);
xnor U15606 (N_15606,N_14600,N_14484);
xnor U15607 (N_15607,N_14487,N_14486);
and U15608 (N_15608,N_14784,N_14704);
nand U15609 (N_15609,N_14580,N_14839);
or U15610 (N_15610,N_14581,N_14610);
xor U15611 (N_15611,N_14877,N_14781);
nand U15612 (N_15612,N_14586,N_14620);
or U15613 (N_15613,N_14922,N_14642);
or U15614 (N_15614,N_14603,N_14991);
nand U15615 (N_15615,N_14915,N_14422);
or U15616 (N_15616,N_14775,N_14546);
or U15617 (N_15617,N_14485,N_14651);
xnor U15618 (N_15618,N_14651,N_14755);
or U15619 (N_15619,N_14926,N_14714);
nand U15620 (N_15620,N_14808,N_14620);
xnor U15621 (N_15621,N_14916,N_14521);
nand U15622 (N_15622,N_14418,N_14532);
and U15623 (N_15623,N_14714,N_14615);
nand U15624 (N_15624,N_14672,N_14986);
or U15625 (N_15625,N_15309,N_15513);
xnor U15626 (N_15626,N_15319,N_15115);
and U15627 (N_15627,N_15540,N_15181);
nand U15628 (N_15628,N_15325,N_15246);
and U15629 (N_15629,N_15601,N_15275);
and U15630 (N_15630,N_15384,N_15088);
nand U15631 (N_15631,N_15004,N_15530);
and U15632 (N_15632,N_15476,N_15395);
xnor U15633 (N_15633,N_15251,N_15278);
nor U15634 (N_15634,N_15333,N_15177);
xor U15635 (N_15635,N_15014,N_15566);
xnor U15636 (N_15636,N_15422,N_15436);
nor U15637 (N_15637,N_15244,N_15053);
xor U15638 (N_15638,N_15287,N_15093);
nor U15639 (N_15639,N_15060,N_15425);
nand U15640 (N_15640,N_15126,N_15335);
xor U15641 (N_15641,N_15462,N_15184);
or U15642 (N_15642,N_15327,N_15102);
and U15643 (N_15643,N_15588,N_15592);
and U15644 (N_15644,N_15057,N_15344);
nor U15645 (N_15645,N_15065,N_15572);
nor U15646 (N_15646,N_15548,N_15135);
nor U15647 (N_15647,N_15405,N_15371);
or U15648 (N_15648,N_15162,N_15130);
or U15649 (N_15649,N_15310,N_15468);
nor U15650 (N_15650,N_15370,N_15170);
xnor U15651 (N_15651,N_15159,N_15147);
nor U15652 (N_15652,N_15612,N_15006);
or U15653 (N_15653,N_15536,N_15078);
xor U15654 (N_15654,N_15377,N_15291);
and U15655 (N_15655,N_15271,N_15040);
or U15656 (N_15656,N_15293,N_15461);
nor U15657 (N_15657,N_15488,N_15522);
or U15658 (N_15658,N_15492,N_15276);
or U15659 (N_15659,N_15457,N_15072);
xor U15660 (N_15660,N_15109,N_15059);
and U15661 (N_15661,N_15311,N_15264);
xor U15662 (N_15662,N_15290,N_15454);
or U15663 (N_15663,N_15401,N_15213);
or U15664 (N_15664,N_15104,N_15447);
xor U15665 (N_15665,N_15316,N_15535);
or U15666 (N_15666,N_15208,N_15336);
xor U15667 (N_15667,N_15166,N_15391);
nor U15668 (N_15668,N_15283,N_15015);
xnor U15669 (N_15669,N_15118,N_15042);
nor U15670 (N_15670,N_15367,N_15539);
nand U15671 (N_15671,N_15002,N_15498);
or U15672 (N_15672,N_15146,N_15527);
and U15673 (N_15673,N_15240,N_15201);
xnor U15674 (N_15674,N_15050,N_15107);
nor U15675 (N_15675,N_15351,N_15451);
and U15676 (N_15676,N_15397,N_15236);
xor U15677 (N_15677,N_15175,N_15314);
and U15678 (N_15678,N_15086,N_15226);
xor U15679 (N_15679,N_15589,N_15355);
nand U15680 (N_15680,N_15420,N_15494);
nor U15681 (N_15681,N_15321,N_15521);
or U15682 (N_15682,N_15400,N_15211);
nand U15683 (N_15683,N_15055,N_15474);
nand U15684 (N_15684,N_15259,N_15173);
or U15685 (N_15685,N_15149,N_15305);
and U15686 (N_15686,N_15419,N_15571);
nor U15687 (N_15687,N_15010,N_15545);
nand U15688 (N_15688,N_15153,N_15496);
and U15689 (N_15689,N_15140,N_15503);
xor U15690 (N_15690,N_15483,N_15315);
nand U15691 (N_15691,N_15207,N_15368);
nand U15692 (N_15692,N_15141,N_15339);
xor U15693 (N_15693,N_15332,N_15360);
xor U15694 (N_15694,N_15191,N_15217);
or U15695 (N_15695,N_15414,N_15594);
xor U15696 (N_15696,N_15475,N_15117);
or U15697 (N_15697,N_15373,N_15005);
nand U15698 (N_15698,N_15026,N_15445);
xnor U15699 (N_15699,N_15304,N_15206);
xor U15700 (N_15700,N_15101,N_15577);
nand U15701 (N_15701,N_15322,N_15605);
nand U15702 (N_15702,N_15575,N_15242);
xor U15703 (N_15703,N_15353,N_15134);
and U15704 (N_15704,N_15340,N_15039);
xor U15705 (N_15705,N_15453,N_15262);
or U15706 (N_15706,N_15407,N_15263);
nor U15707 (N_15707,N_15533,N_15103);
nand U15708 (N_15708,N_15379,N_15179);
nor U15709 (N_15709,N_15127,N_15615);
nand U15710 (N_15710,N_15441,N_15112);
or U15711 (N_15711,N_15218,N_15435);
or U15712 (N_15712,N_15564,N_15038);
nand U15713 (N_15713,N_15614,N_15458);
nand U15714 (N_15714,N_15035,N_15392);
or U15715 (N_15715,N_15348,N_15524);
xnor U15716 (N_15716,N_15043,N_15227);
or U15717 (N_15717,N_15215,N_15075);
or U15718 (N_15718,N_15427,N_15347);
and U15719 (N_15719,N_15220,N_15624);
and U15720 (N_15720,N_15094,N_15049);
xnor U15721 (N_15721,N_15125,N_15477);
or U15722 (N_15722,N_15029,N_15358);
nor U15723 (N_15723,N_15495,N_15460);
xor U15724 (N_15724,N_15559,N_15531);
or U15725 (N_15725,N_15168,N_15025);
nand U15726 (N_15726,N_15113,N_15001);
nand U15727 (N_15727,N_15187,N_15223);
nand U15728 (N_15728,N_15324,N_15058);
and U15729 (N_15729,N_15409,N_15408);
nor U15730 (N_15730,N_15560,N_15455);
nand U15731 (N_15731,N_15066,N_15359);
nand U15732 (N_15732,N_15144,N_15390);
nand U15733 (N_15733,N_15267,N_15183);
or U15734 (N_15734,N_15423,N_15288);
or U15735 (N_15735,N_15543,N_15511);
and U15736 (N_15736,N_15216,N_15334);
nand U15737 (N_15737,N_15501,N_15248);
xnor U15738 (N_15738,N_15580,N_15583);
xnor U15739 (N_15739,N_15538,N_15214);
nor U15740 (N_15740,N_15136,N_15192);
xor U15741 (N_15741,N_15519,N_15128);
or U15742 (N_15742,N_15547,N_15222);
xor U15743 (N_15743,N_15196,N_15526);
nand U15744 (N_15744,N_15169,N_15607);
and U15745 (N_15745,N_15027,N_15597);
xnor U15746 (N_15746,N_15361,N_15092);
nand U15747 (N_15747,N_15326,N_15330);
nand U15748 (N_15748,N_15106,N_15070);
nor U15749 (N_15749,N_15163,N_15064);
nand U15750 (N_15750,N_15398,N_15228);
nor U15751 (N_15751,N_15443,N_15329);
and U15752 (N_15752,N_15616,N_15234);
nand U15753 (N_15753,N_15020,N_15229);
and U15754 (N_15754,N_15051,N_15255);
nand U15755 (N_15755,N_15033,N_15591);
or U15756 (N_15756,N_15415,N_15489);
and U15757 (N_15757,N_15341,N_15097);
xor U15758 (N_15758,N_15481,N_15257);
xor U15759 (N_15759,N_15582,N_15487);
nand U15760 (N_15760,N_15108,N_15139);
nand U15761 (N_15761,N_15131,N_15444);
or U15762 (N_15762,N_15578,N_15525);
or U15763 (N_15763,N_15194,N_15016);
nand U15764 (N_15764,N_15551,N_15084);
and U15765 (N_15765,N_15268,N_15412);
nor U15766 (N_15766,N_15432,N_15045);
or U15767 (N_15767,N_15449,N_15343);
and U15768 (N_15768,N_15385,N_15562);
or U15769 (N_15769,N_15294,N_15478);
and U15770 (N_15770,N_15362,N_15486);
and U15771 (N_15771,N_15044,N_15479);
and U15772 (N_15772,N_15532,N_15349);
and U15773 (N_15773,N_15584,N_15600);
xnor U15774 (N_15774,N_15265,N_15138);
or U15775 (N_15775,N_15553,N_15317);
xnor U15776 (N_15776,N_15202,N_15541);
nand U15777 (N_15777,N_15151,N_15537);
and U15778 (N_15778,N_15137,N_15174);
nand U15779 (N_15779,N_15021,N_15369);
nand U15780 (N_15780,N_15429,N_15123);
and U15781 (N_15781,N_15160,N_15593);
nor U15782 (N_15782,N_15514,N_15313);
and U15783 (N_15783,N_15312,N_15260);
and U15784 (N_15784,N_15345,N_15365);
or U15785 (N_15785,N_15285,N_15561);
and U15786 (N_15786,N_15424,N_15504);
or U15787 (N_15787,N_15258,N_15007);
or U15788 (N_15788,N_15599,N_15205);
nor U15789 (N_15789,N_15523,N_15596);
nand U15790 (N_15790,N_15497,N_15609);
nor U15791 (N_15791,N_15095,N_15011);
nor U15792 (N_15792,N_15032,N_15438);
or U15793 (N_15793,N_15224,N_15402);
nand U15794 (N_15794,N_15046,N_15249);
nor U15795 (N_15795,N_15197,N_15366);
or U15796 (N_15796,N_15375,N_15142);
nor U15797 (N_15797,N_15469,N_15150);
xor U15798 (N_15798,N_15085,N_15171);
xnor U15799 (N_15799,N_15230,N_15281);
nor U15800 (N_15800,N_15133,N_15387);
nand U15801 (N_15801,N_15555,N_15354);
or U15802 (N_15802,N_15404,N_15490);
nor U15803 (N_15803,N_15235,N_15069);
or U15804 (N_15804,N_15210,N_15132);
or U15805 (N_15805,N_15156,N_15620);
and U15806 (N_15806,N_15299,N_15048);
and U15807 (N_15807,N_15546,N_15338);
or U15808 (N_15808,N_15516,N_15618);
nand U15809 (N_15809,N_15509,N_15182);
or U15810 (N_15810,N_15081,N_15037);
or U15811 (N_15811,N_15426,N_15467);
xnor U15812 (N_15812,N_15018,N_15195);
xnor U15813 (N_15813,N_15396,N_15623);
and U15814 (N_15814,N_15071,N_15382);
nor U15815 (N_15815,N_15298,N_15376);
xor U15816 (N_15816,N_15091,N_15485);
and U15817 (N_15817,N_15111,N_15000);
nand U15818 (N_15818,N_15180,N_15297);
xnor U15819 (N_15819,N_15581,N_15500);
nor U15820 (N_15820,N_15225,N_15399);
nor U15821 (N_15821,N_15129,N_15012);
nor U15822 (N_15822,N_15089,N_15212);
xnor U15823 (N_15823,N_15161,N_15269);
nor U15824 (N_15824,N_15076,N_15586);
or U15825 (N_15825,N_15052,N_15518);
nor U15826 (N_15826,N_15507,N_15472);
and U15827 (N_15827,N_15284,N_15544);
nor U15828 (N_15828,N_15074,N_15493);
xor U15829 (N_15829,N_15569,N_15254);
xor U15830 (N_15830,N_15013,N_15610);
xnor U15831 (N_15831,N_15590,N_15148);
or U15832 (N_15832,N_15252,N_15606);
xnor U15833 (N_15833,N_15352,N_15036);
nor U15834 (N_15834,N_15245,N_15250);
xor U15835 (N_15835,N_15186,N_15303);
xnor U15836 (N_15836,N_15570,N_15080);
nand U15837 (N_15837,N_15296,N_15506);
nor U15838 (N_15838,N_15009,N_15099);
xor U15839 (N_15839,N_15198,N_15617);
and U15840 (N_15840,N_15356,N_15556);
and U15841 (N_15841,N_15022,N_15534);
xor U15842 (N_15842,N_15337,N_15439);
nand U15843 (N_15843,N_15172,N_15239);
or U15844 (N_15844,N_15346,N_15003);
or U15845 (N_15845,N_15155,N_15266);
or U15846 (N_15846,N_15189,N_15122);
xnor U15847 (N_15847,N_15017,N_15034);
nor U15848 (N_15848,N_15077,N_15096);
nand U15849 (N_15849,N_15098,N_15484);
and U15850 (N_15850,N_15430,N_15433);
or U15851 (N_15851,N_15558,N_15528);
and U15852 (N_15852,N_15437,N_15190);
nand U15853 (N_15853,N_15434,N_15056);
and U15854 (N_15854,N_15219,N_15517);
and U15855 (N_15855,N_15272,N_15200);
nand U15856 (N_15856,N_15008,N_15199);
xor U15857 (N_15857,N_15167,N_15185);
nor U15858 (N_15858,N_15178,N_15466);
or U15859 (N_15859,N_15054,N_15188);
and U15860 (N_15860,N_15243,N_15090);
or U15861 (N_15861,N_15579,N_15237);
and U15862 (N_15862,N_15087,N_15381);
xor U15863 (N_15863,N_15410,N_15510);
and U15864 (N_15864,N_15473,N_15386);
nand U15865 (N_15865,N_15440,N_15100);
nand U15866 (N_15866,N_15549,N_15233);
or U15867 (N_15867,N_15068,N_15273);
or U15868 (N_15868,N_15350,N_15413);
or U15869 (N_15869,N_15231,N_15302);
xnor U15870 (N_15870,N_15030,N_15221);
xnor U15871 (N_15871,N_15550,N_15574);
nand U15872 (N_15872,N_15120,N_15418);
or U15873 (N_15873,N_15431,N_15567);
nand U15874 (N_15874,N_15411,N_15062);
or U15875 (N_15875,N_15274,N_15568);
nor U15876 (N_15876,N_15480,N_15031);
nand U15877 (N_15877,N_15595,N_15270);
xor U15878 (N_15878,N_15482,N_15318);
or U15879 (N_15879,N_15613,N_15619);
or U15880 (N_15880,N_15331,N_15116);
and U15881 (N_15881,N_15622,N_15491);
and U15882 (N_15882,N_15576,N_15552);
xnor U15883 (N_15883,N_15119,N_15383);
xor U15884 (N_15884,N_15105,N_15611);
nor U15885 (N_15885,N_15416,N_15621);
xnor U15886 (N_15886,N_15515,N_15204);
xor U15887 (N_15887,N_15028,N_15061);
nor U15888 (N_15888,N_15389,N_15520);
nor U15889 (N_15889,N_15176,N_15152);
xnor U15890 (N_15890,N_15306,N_15301);
xnor U15891 (N_15891,N_15286,N_15421);
xnor U15892 (N_15892,N_15193,N_15428);
or U15893 (N_15893,N_15024,N_15364);
nor U15894 (N_15894,N_15585,N_15463);
nor U15895 (N_15895,N_15602,N_15542);
xnor U15896 (N_15896,N_15241,N_15452);
nand U15897 (N_15897,N_15279,N_15378);
xnor U15898 (N_15898,N_15357,N_15502);
xor U15899 (N_15899,N_15456,N_15573);
nand U15900 (N_15900,N_15406,N_15063);
and U15901 (N_15901,N_15403,N_15124);
or U15902 (N_15902,N_15121,N_15470);
xnor U15903 (N_15903,N_15067,N_15529);
or U15904 (N_15904,N_15465,N_15598);
or U15905 (N_15905,N_15083,N_15393);
or U15906 (N_15906,N_15143,N_15110);
or U15907 (N_15907,N_15505,N_15459);
and U15908 (N_15908,N_15145,N_15446);
nand U15909 (N_15909,N_15388,N_15165);
or U15910 (N_15910,N_15563,N_15247);
xnor U15911 (N_15911,N_15565,N_15464);
or U15912 (N_15912,N_15256,N_15442);
nand U15913 (N_15913,N_15261,N_15342);
xor U15914 (N_15914,N_15158,N_15079);
and U15915 (N_15915,N_15450,N_15238);
xnor U15916 (N_15916,N_15073,N_15554);
nand U15917 (N_15917,N_15328,N_15019);
nand U15918 (N_15918,N_15154,N_15082);
nor U15919 (N_15919,N_15282,N_15308);
xnor U15920 (N_15920,N_15280,N_15295);
xnor U15921 (N_15921,N_15253,N_15323);
nor U15922 (N_15922,N_15603,N_15300);
nand U15923 (N_15923,N_15512,N_15372);
xor U15924 (N_15924,N_15380,N_15604);
or U15925 (N_15925,N_15232,N_15471);
xor U15926 (N_15926,N_15209,N_15114);
nand U15927 (N_15927,N_15363,N_15289);
nand U15928 (N_15928,N_15448,N_15164);
and U15929 (N_15929,N_15307,N_15374);
nand U15930 (N_15930,N_15203,N_15320);
nor U15931 (N_15931,N_15587,N_15292);
xnor U15932 (N_15932,N_15417,N_15608);
nor U15933 (N_15933,N_15394,N_15157);
or U15934 (N_15934,N_15277,N_15041);
xor U15935 (N_15935,N_15023,N_15047);
or U15936 (N_15936,N_15499,N_15557);
and U15937 (N_15937,N_15508,N_15317);
or U15938 (N_15938,N_15511,N_15299);
nand U15939 (N_15939,N_15596,N_15022);
nor U15940 (N_15940,N_15516,N_15415);
and U15941 (N_15941,N_15607,N_15101);
or U15942 (N_15942,N_15194,N_15039);
nor U15943 (N_15943,N_15528,N_15403);
nor U15944 (N_15944,N_15362,N_15415);
and U15945 (N_15945,N_15284,N_15191);
xnor U15946 (N_15946,N_15029,N_15081);
xor U15947 (N_15947,N_15606,N_15297);
and U15948 (N_15948,N_15365,N_15100);
nand U15949 (N_15949,N_15459,N_15525);
xor U15950 (N_15950,N_15292,N_15479);
and U15951 (N_15951,N_15219,N_15408);
nor U15952 (N_15952,N_15170,N_15113);
and U15953 (N_15953,N_15067,N_15362);
nand U15954 (N_15954,N_15108,N_15239);
xor U15955 (N_15955,N_15313,N_15525);
and U15956 (N_15956,N_15547,N_15374);
nand U15957 (N_15957,N_15151,N_15534);
nor U15958 (N_15958,N_15367,N_15441);
or U15959 (N_15959,N_15596,N_15126);
nor U15960 (N_15960,N_15098,N_15129);
or U15961 (N_15961,N_15405,N_15074);
nor U15962 (N_15962,N_15260,N_15599);
nand U15963 (N_15963,N_15271,N_15029);
xnor U15964 (N_15964,N_15149,N_15203);
nand U15965 (N_15965,N_15614,N_15266);
xor U15966 (N_15966,N_15595,N_15180);
or U15967 (N_15967,N_15270,N_15409);
nand U15968 (N_15968,N_15523,N_15377);
xor U15969 (N_15969,N_15522,N_15073);
and U15970 (N_15970,N_15432,N_15404);
nor U15971 (N_15971,N_15242,N_15370);
xnor U15972 (N_15972,N_15224,N_15354);
or U15973 (N_15973,N_15608,N_15506);
xor U15974 (N_15974,N_15103,N_15567);
nor U15975 (N_15975,N_15263,N_15580);
or U15976 (N_15976,N_15289,N_15242);
nor U15977 (N_15977,N_15426,N_15349);
xnor U15978 (N_15978,N_15516,N_15155);
nor U15979 (N_15979,N_15592,N_15269);
nand U15980 (N_15980,N_15366,N_15040);
nand U15981 (N_15981,N_15011,N_15126);
and U15982 (N_15982,N_15109,N_15448);
or U15983 (N_15983,N_15344,N_15523);
or U15984 (N_15984,N_15120,N_15428);
and U15985 (N_15985,N_15491,N_15476);
and U15986 (N_15986,N_15330,N_15040);
nor U15987 (N_15987,N_15280,N_15354);
nand U15988 (N_15988,N_15337,N_15160);
xnor U15989 (N_15989,N_15347,N_15358);
nand U15990 (N_15990,N_15149,N_15176);
nor U15991 (N_15991,N_15259,N_15313);
xnor U15992 (N_15992,N_15284,N_15390);
nor U15993 (N_15993,N_15062,N_15555);
and U15994 (N_15994,N_15476,N_15077);
or U15995 (N_15995,N_15196,N_15242);
or U15996 (N_15996,N_15461,N_15568);
or U15997 (N_15997,N_15126,N_15309);
nor U15998 (N_15998,N_15488,N_15102);
or U15999 (N_15999,N_15440,N_15009);
and U16000 (N_16000,N_15454,N_15307);
nor U16001 (N_16001,N_15523,N_15023);
nor U16002 (N_16002,N_15033,N_15410);
and U16003 (N_16003,N_15108,N_15288);
nand U16004 (N_16004,N_15119,N_15001);
nor U16005 (N_16005,N_15418,N_15329);
or U16006 (N_16006,N_15143,N_15016);
nor U16007 (N_16007,N_15045,N_15368);
xnor U16008 (N_16008,N_15455,N_15152);
or U16009 (N_16009,N_15623,N_15268);
or U16010 (N_16010,N_15483,N_15527);
or U16011 (N_16011,N_15535,N_15136);
nor U16012 (N_16012,N_15376,N_15249);
nand U16013 (N_16013,N_15019,N_15172);
xor U16014 (N_16014,N_15457,N_15498);
nor U16015 (N_16015,N_15554,N_15162);
or U16016 (N_16016,N_15556,N_15462);
nor U16017 (N_16017,N_15571,N_15565);
or U16018 (N_16018,N_15568,N_15088);
and U16019 (N_16019,N_15036,N_15309);
or U16020 (N_16020,N_15167,N_15401);
or U16021 (N_16021,N_15012,N_15264);
and U16022 (N_16022,N_15392,N_15115);
nor U16023 (N_16023,N_15264,N_15309);
or U16024 (N_16024,N_15025,N_15024);
nand U16025 (N_16025,N_15538,N_15585);
or U16026 (N_16026,N_15468,N_15499);
nand U16027 (N_16027,N_15073,N_15241);
or U16028 (N_16028,N_15217,N_15565);
or U16029 (N_16029,N_15574,N_15548);
nand U16030 (N_16030,N_15499,N_15046);
nor U16031 (N_16031,N_15063,N_15483);
or U16032 (N_16032,N_15397,N_15189);
and U16033 (N_16033,N_15136,N_15029);
or U16034 (N_16034,N_15344,N_15507);
nor U16035 (N_16035,N_15444,N_15151);
nand U16036 (N_16036,N_15555,N_15457);
or U16037 (N_16037,N_15226,N_15373);
nor U16038 (N_16038,N_15192,N_15191);
and U16039 (N_16039,N_15600,N_15178);
nor U16040 (N_16040,N_15403,N_15354);
and U16041 (N_16041,N_15096,N_15529);
nand U16042 (N_16042,N_15390,N_15326);
and U16043 (N_16043,N_15294,N_15268);
xnor U16044 (N_16044,N_15492,N_15042);
xnor U16045 (N_16045,N_15243,N_15155);
nor U16046 (N_16046,N_15126,N_15117);
nor U16047 (N_16047,N_15073,N_15432);
nand U16048 (N_16048,N_15505,N_15568);
nor U16049 (N_16049,N_15432,N_15486);
xor U16050 (N_16050,N_15435,N_15129);
xnor U16051 (N_16051,N_15092,N_15167);
and U16052 (N_16052,N_15207,N_15361);
and U16053 (N_16053,N_15525,N_15240);
xnor U16054 (N_16054,N_15200,N_15314);
nor U16055 (N_16055,N_15527,N_15152);
xnor U16056 (N_16056,N_15459,N_15465);
nand U16057 (N_16057,N_15392,N_15020);
xor U16058 (N_16058,N_15172,N_15040);
xnor U16059 (N_16059,N_15124,N_15548);
xnor U16060 (N_16060,N_15504,N_15313);
or U16061 (N_16061,N_15108,N_15081);
nor U16062 (N_16062,N_15127,N_15238);
nor U16063 (N_16063,N_15443,N_15515);
nor U16064 (N_16064,N_15124,N_15489);
or U16065 (N_16065,N_15459,N_15491);
xor U16066 (N_16066,N_15551,N_15358);
nor U16067 (N_16067,N_15106,N_15447);
xor U16068 (N_16068,N_15017,N_15316);
xor U16069 (N_16069,N_15341,N_15287);
and U16070 (N_16070,N_15393,N_15213);
nor U16071 (N_16071,N_15475,N_15288);
nand U16072 (N_16072,N_15196,N_15441);
nand U16073 (N_16073,N_15381,N_15402);
nor U16074 (N_16074,N_15545,N_15244);
xor U16075 (N_16075,N_15571,N_15213);
or U16076 (N_16076,N_15586,N_15513);
xnor U16077 (N_16077,N_15454,N_15432);
xnor U16078 (N_16078,N_15453,N_15268);
nor U16079 (N_16079,N_15340,N_15118);
nor U16080 (N_16080,N_15115,N_15009);
or U16081 (N_16081,N_15284,N_15593);
nand U16082 (N_16082,N_15255,N_15518);
xor U16083 (N_16083,N_15275,N_15239);
nand U16084 (N_16084,N_15506,N_15249);
nor U16085 (N_16085,N_15262,N_15611);
and U16086 (N_16086,N_15482,N_15356);
and U16087 (N_16087,N_15215,N_15357);
and U16088 (N_16088,N_15398,N_15155);
xnor U16089 (N_16089,N_15342,N_15051);
xnor U16090 (N_16090,N_15553,N_15607);
xnor U16091 (N_16091,N_15345,N_15173);
or U16092 (N_16092,N_15167,N_15062);
nand U16093 (N_16093,N_15066,N_15188);
or U16094 (N_16094,N_15285,N_15186);
and U16095 (N_16095,N_15557,N_15389);
and U16096 (N_16096,N_15384,N_15463);
nand U16097 (N_16097,N_15198,N_15335);
or U16098 (N_16098,N_15142,N_15119);
xor U16099 (N_16099,N_15597,N_15081);
or U16100 (N_16100,N_15030,N_15624);
nand U16101 (N_16101,N_15562,N_15190);
nand U16102 (N_16102,N_15196,N_15125);
xor U16103 (N_16103,N_15555,N_15147);
and U16104 (N_16104,N_15369,N_15160);
nand U16105 (N_16105,N_15208,N_15141);
nor U16106 (N_16106,N_15362,N_15412);
nor U16107 (N_16107,N_15318,N_15140);
and U16108 (N_16108,N_15070,N_15232);
nand U16109 (N_16109,N_15501,N_15223);
or U16110 (N_16110,N_15386,N_15314);
or U16111 (N_16111,N_15237,N_15209);
nand U16112 (N_16112,N_15344,N_15015);
xor U16113 (N_16113,N_15588,N_15573);
nor U16114 (N_16114,N_15374,N_15050);
or U16115 (N_16115,N_15184,N_15052);
and U16116 (N_16116,N_15160,N_15394);
nor U16117 (N_16117,N_15581,N_15536);
or U16118 (N_16118,N_15287,N_15236);
or U16119 (N_16119,N_15025,N_15188);
and U16120 (N_16120,N_15130,N_15028);
nand U16121 (N_16121,N_15163,N_15007);
nand U16122 (N_16122,N_15614,N_15178);
or U16123 (N_16123,N_15355,N_15125);
and U16124 (N_16124,N_15621,N_15440);
or U16125 (N_16125,N_15576,N_15142);
nand U16126 (N_16126,N_15017,N_15280);
or U16127 (N_16127,N_15404,N_15172);
nand U16128 (N_16128,N_15122,N_15324);
xnor U16129 (N_16129,N_15344,N_15561);
xor U16130 (N_16130,N_15616,N_15305);
and U16131 (N_16131,N_15255,N_15259);
and U16132 (N_16132,N_15460,N_15126);
xor U16133 (N_16133,N_15426,N_15046);
nand U16134 (N_16134,N_15001,N_15091);
xnor U16135 (N_16135,N_15171,N_15116);
nand U16136 (N_16136,N_15323,N_15374);
and U16137 (N_16137,N_15049,N_15311);
or U16138 (N_16138,N_15194,N_15604);
xnor U16139 (N_16139,N_15169,N_15046);
xor U16140 (N_16140,N_15060,N_15512);
xor U16141 (N_16141,N_15068,N_15161);
nand U16142 (N_16142,N_15102,N_15523);
xor U16143 (N_16143,N_15522,N_15335);
xor U16144 (N_16144,N_15307,N_15123);
nor U16145 (N_16145,N_15180,N_15415);
or U16146 (N_16146,N_15277,N_15282);
and U16147 (N_16147,N_15461,N_15476);
and U16148 (N_16148,N_15222,N_15106);
xnor U16149 (N_16149,N_15068,N_15174);
or U16150 (N_16150,N_15447,N_15289);
nand U16151 (N_16151,N_15191,N_15109);
and U16152 (N_16152,N_15202,N_15420);
nor U16153 (N_16153,N_15235,N_15420);
nand U16154 (N_16154,N_15433,N_15225);
xnor U16155 (N_16155,N_15042,N_15353);
nand U16156 (N_16156,N_15143,N_15043);
or U16157 (N_16157,N_15431,N_15494);
nand U16158 (N_16158,N_15319,N_15127);
nor U16159 (N_16159,N_15504,N_15425);
xnor U16160 (N_16160,N_15373,N_15331);
nand U16161 (N_16161,N_15369,N_15041);
xnor U16162 (N_16162,N_15000,N_15476);
xor U16163 (N_16163,N_15362,N_15065);
xor U16164 (N_16164,N_15576,N_15291);
and U16165 (N_16165,N_15022,N_15445);
nand U16166 (N_16166,N_15201,N_15520);
nand U16167 (N_16167,N_15437,N_15605);
and U16168 (N_16168,N_15467,N_15451);
nor U16169 (N_16169,N_15104,N_15174);
nor U16170 (N_16170,N_15379,N_15136);
and U16171 (N_16171,N_15147,N_15177);
xor U16172 (N_16172,N_15016,N_15411);
and U16173 (N_16173,N_15035,N_15002);
and U16174 (N_16174,N_15394,N_15540);
nand U16175 (N_16175,N_15204,N_15435);
or U16176 (N_16176,N_15016,N_15452);
and U16177 (N_16177,N_15613,N_15512);
nor U16178 (N_16178,N_15025,N_15411);
or U16179 (N_16179,N_15337,N_15050);
or U16180 (N_16180,N_15069,N_15444);
nor U16181 (N_16181,N_15223,N_15153);
nand U16182 (N_16182,N_15527,N_15101);
or U16183 (N_16183,N_15262,N_15215);
nand U16184 (N_16184,N_15599,N_15614);
nand U16185 (N_16185,N_15059,N_15064);
xor U16186 (N_16186,N_15618,N_15439);
nand U16187 (N_16187,N_15023,N_15053);
xnor U16188 (N_16188,N_15518,N_15330);
nor U16189 (N_16189,N_15350,N_15294);
or U16190 (N_16190,N_15164,N_15188);
and U16191 (N_16191,N_15388,N_15135);
xnor U16192 (N_16192,N_15489,N_15049);
nor U16193 (N_16193,N_15600,N_15612);
nand U16194 (N_16194,N_15545,N_15264);
nand U16195 (N_16195,N_15496,N_15595);
and U16196 (N_16196,N_15350,N_15326);
xnor U16197 (N_16197,N_15431,N_15409);
and U16198 (N_16198,N_15222,N_15152);
nor U16199 (N_16199,N_15189,N_15075);
nand U16200 (N_16200,N_15308,N_15423);
nand U16201 (N_16201,N_15293,N_15514);
xor U16202 (N_16202,N_15364,N_15398);
or U16203 (N_16203,N_15480,N_15120);
nor U16204 (N_16204,N_15487,N_15490);
nor U16205 (N_16205,N_15148,N_15010);
nor U16206 (N_16206,N_15099,N_15492);
xnor U16207 (N_16207,N_15607,N_15002);
nor U16208 (N_16208,N_15595,N_15304);
xor U16209 (N_16209,N_15423,N_15561);
xnor U16210 (N_16210,N_15127,N_15165);
or U16211 (N_16211,N_15614,N_15072);
nand U16212 (N_16212,N_15313,N_15444);
and U16213 (N_16213,N_15418,N_15518);
and U16214 (N_16214,N_15435,N_15157);
nand U16215 (N_16215,N_15439,N_15562);
xor U16216 (N_16216,N_15320,N_15053);
nand U16217 (N_16217,N_15043,N_15456);
nand U16218 (N_16218,N_15442,N_15620);
or U16219 (N_16219,N_15347,N_15186);
or U16220 (N_16220,N_15066,N_15431);
and U16221 (N_16221,N_15055,N_15566);
nand U16222 (N_16222,N_15095,N_15297);
nand U16223 (N_16223,N_15195,N_15359);
nand U16224 (N_16224,N_15531,N_15041);
nor U16225 (N_16225,N_15353,N_15349);
nand U16226 (N_16226,N_15523,N_15423);
xnor U16227 (N_16227,N_15558,N_15466);
and U16228 (N_16228,N_15559,N_15233);
nor U16229 (N_16229,N_15482,N_15337);
nand U16230 (N_16230,N_15222,N_15290);
nor U16231 (N_16231,N_15451,N_15504);
nand U16232 (N_16232,N_15509,N_15250);
nor U16233 (N_16233,N_15546,N_15493);
nor U16234 (N_16234,N_15420,N_15472);
nand U16235 (N_16235,N_15164,N_15192);
xnor U16236 (N_16236,N_15429,N_15481);
or U16237 (N_16237,N_15188,N_15096);
nor U16238 (N_16238,N_15354,N_15287);
and U16239 (N_16239,N_15158,N_15093);
and U16240 (N_16240,N_15263,N_15565);
nor U16241 (N_16241,N_15617,N_15211);
nand U16242 (N_16242,N_15528,N_15330);
or U16243 (N_16243,N_15133,N_15257);
xnor U16244 (N_16244,N_15220,N_15377);
xor U16245 (N_16245,N_15576,N_15222);
xnor U16246 (N_16246,N_15384,N_15558);
nor U16247 (N_16247,N_15476,N_15248);
nor U16248 (N_16248,N_15480,N_15342);
or U16249 (N_16249,N_15142,N_15392);
and U16250 (N_16250,N_16019,N_15958);
nor U16251 (N_16251,N_16072,N_15782);
or U16252 (N_16252,N_16153,N_16176);
or U16253 (N_16253,N_16136,N_15689);
nand U16254 (N_16254,N_15778,N_15976);
and U16255 (N_16255,N_16225,N_16124);
or U16256 (N_16256,N_15718,N_16249);
nor U16257 (N_16257,N_15786,N_16195);
xor U16258 (N_16258,N_15665,N_15925);
nand U16259 (N_16259,N_16146,N_16165);
or U16260 (N_16260,N_15835,N_15815);
nor U16261 (N_16261,N_15964,N_15747);
or U16262 (N_16262,N_15781,N_15967);
nor U16263 (N_16263,N_15851,N_15787);
nand U16264 (N_16264,N_15711,N_15949);
nor U16265 (N_16265,N_15807,N_15765);
nor U16266 (N_16266,N_16123,N_15779);
nand U16267 (N_16267,N_15713,N_16138);
nor U16268 (N_16268,N_15630,N_15750);
nand U16269 (N_16269,N_15784,N_15797);
or U16270 (N_16270,N_16015,N_16073);
nor U16271 (N_16271,N_15848,N_15654);
nand U16272 (N_16272,N_16111,N_15738);
or U16273 (N_16273,N_16022,N_16033);
nor U16274 (N_16274,N_15868,N_15668);
nor U16275 (N_16275,N_15725,N_16100);
xnor U16276 (N_16276,N_16235,N_15902);
xor U16277 (N_16277,N_15977,N_15938);
nand U16278 (N_16278,N_15694,N_15876);
nor U16279 (N_16279,N_16219,N_16067);
nand U16280 (N_16280,N_16117,N_16102);
nor U16281 (N_16281,N_15794,N_15777);
xnor U16282 (N_16282,N_16128,N_16240);
or U16283 (N_16283,N_16002,N_15878);
and U16284 (N_16284,N_16094,N_15972);
and U16285 (N_16285,N_15864,N_16142);
and U16286 (N_16286,N_16139,N_15648);
or U16287 (N_16287,N_16133,N_15974);
or U16288 (N_16288,N_15772,N_16004);
or U16289 (N_16289,N_15880,N_15673);
nor U16290 (N_16290,N_16049,N_16213);
xnor U16291 (N_16291,N_16129,N_15907);
nand U16292 (N_16292,N_15915,N_16242);
and U16293 (N_16293,N_16070,N_15686);
xor U16294 (N_16294,N_15803,N_16081);
xnor U16295 (N_16295,N_16125,N_15692);
nor U16296 (N_16296,N_15914,N_15773);
nor U16297 (N_16297,N_16036,N_15709);
and U16298 (N_16298,N_16104,N_15840);
and U16299 (N_16299,N_15985,N_16056);
nand U16300 (N_16300,N_15965,N_15882);
xor U16301 (N_16301,N_16144,N_15953);
and U16302 (N_16302,N_15679,N_16155);
and U16303 (N_16303,N_15946,N_15683);
nor U16304 (N_16304,N_16157,N_15741);
and U16305 (N_16305,N_16211,N_15969);
nand U16306 (N_16306,N_15687,N_16046);
and U16307 (N_16307,N_15704,N_15961);
or U16308 (N_16308,N_15829,N_15962);
xnor U16309 (N_16309,N_16044,N_15918);
and U16310 (N_16310,N_16172,N_15720);
xor U16311 (N_16311,N_15831,N_16210);
nand U16312 (N_16312,N_15879,N_15729);
or U16313 (N_16313,N_15629,N_15978);
or U16314 (N_16314,N_15955,N_16075);
xnor U16315 (N_16315,N_15724,N_16215);
nor U16316 (N_16316,N_15759,N_15853);
xor U16317 (N_16317,N_16032,N_15633);
and U16318 (N_16318,N_16188,N_15688);
nand U16319 (N_16319,N_15875,N_15798);
or U16320 (N_16320,N_16180,N_16167);
nand U16321 (N_16321,N_15641,N_16244);
or U16322 (N_16322,N_15874,N_16080);
xnor U16323 (N_16323,N_16151,N_15651);
and U16324 (N_16324,N_15952,N_15968);
or U16325 (N_16325,N_15942,N_15761);
or U16326 (N_16326,N_15793,N_15884);
nand U16327 (N_16327,N_15647,N_15762);
nand U16328 (N_16328,N_16234,N_15821);
nand U16329 (N_16329,N_15693,N_15842);
nor U16330 (N_16330,N_15987,N_15894);
and U16331 (N_16331,N_16012,N_16085);
and U16332 (N_16332,N_15963,N_15819);
xnor U16333 (N_16333,N_16190,N_16077);
or U16334 (N_16334,N_15854,N_15789);
xnor U16335 (N_16335,N_16071,N_16241);
nand U16336 (N_16336,N_15660,N_15856);
nand U16337 (N_16337,N_16184,N_15828);
nor U16338 (N_16338,N_15727,N_15810);
nor U16339 (N_16339,N_15714,N_16065);
or U16340 (N_16340,N_15684,N_15642);
or U16341 (N_16341,N_16160,N_15717);
and U16342 (N_16342,N_16107,N_15712);
nand U16343 (N_16343,N_15939,N_15674);
nor U16344 (N_16344,N_16243,N_16057);
xor U16345 (N_16345,N_16003,N_15749);
nor U16346 (N_16346,N_16039,N_15910);
xnor U16347 (N_16347,N_15986,N_15802);
nor U16348 (N_16348,N_16187,N_16137);
nand U16349 (N_16349,N_15883,N_15924);
or U16350 (N_16350,N_16086,N_16096);
or U16351 (N_16351,N_15701,N_15913);
nand U16352 (N_16352,N_15706,N_15659);
xor U16353 (N_16353,N_16202,N_15852);
and U16354 (N_16354,N_16222,N_15635);
or U16355 (N_16355,N_15752,N_16217);
nor U16356 (N_16356,N_16062,N_16200);
or U16357 (N_16357,N_16247,N_16161);
nand U16358 (N_16358,N_15678,N_16109);
xor U16359 (N_16359,N_16166,N_15935);
and U16360 (N_16360,N_15979,N_16163);
xor U16361 (N_16361,N_15945,N_16134);
or U16362 (N_16362,N_16060,N_15818);
xor U16363 (N_16363,N_15664,N_15893);
xor U16364 (N_16364,N_15824,N_15857);
and U16365 (N_16365,N_15870,N_15703);
or U16366 (N_16366,N_16236,N_16021);
and U16367 (N_16367,N_16246,N_16148);
nor U16368 (N_16368,N_16207,N_15917);
nand U16369 (N_16369,N_16145,N_15655);
and U16370 (N_16370,N_15859,N_15638);
xnor U16371 (N_16371,N_16231,N_15716);
nor U16372 (N_16372,N_16122,N_15719);
nor U16373 (N_16373,N_15626,N_15931);
or U16374 (N_16374,N_15998,N_15643);
nor U16375 (N_16375,N_16189,N_15801);
and U16376 (N_16376,N_16024,N_15943);
nand U16377 (N_16377,N_16209,N_15715);
nor U16378 (N_16378,N_15627,N_16101);
or U16379 (N_16379,N_16112,N_15912);
or U16380 (N_16380,N_15780,N_16055);
and U16381 (N_16381,N_15636,N_16181);
or U16382 (N_16382,N_15947,N_15896);
xnor U16383 (N_16383,N_15911,N_15923);
and U16384 (N_16384,N_15652,N_15930);
nor U16385 (N_16385,N_15858,N_15774);
nand U16386 (N_16386,N_15639,N_15739);
or U16387 (N_16387,N_15685,N_16226);
nor U16388 (N_16388,N_16054,N_15696);
and U16389 (N_16389,N_16179,N_15785);
and U16390 (N_16390,N_15806,N_15754);
nor U16391 (N_16391,N_15653,N_16152);
nor U16392 (N_16392,N_16011,N_15887);
xor U16393 (N_16393,N_15834,N_16061);
and U16394 (N_16394,N_15861,N_15996);
nand U16395 (N_16395,N_15649,N_16013);
or U16396 (N_16396,N_15932,N_15640);
nand U16397 (N_16397,N_15920,N_15755);
nor U16398 (N_16398,N_15690,N_15700);
or U16399 (N_16399,N_16227,N_15993);
xnor U16400 (N_16400,N_16079,N_16238);
or U16401 (N_16401,N_15885,N_15676);
and U16402 (N_16402,N_15733,N_16230);
nor U16403 (N_16403,N_16214,N_16237);
nor U16404 (N_16404,N_16232,N_15847);
nor U16405 (N_16405,N_15812,N_15743);
and U16406 (N_16406,N_15865,N_16186);
and U16407 (N_16407,N_16141,N_15916);
or U16408 (N_16408,N_15708,N_15644);
xor U16409 (N_16409,N_15988,N_15705);
or U16410 (N_16410,N_15732,N_15899);
nor U16411 (N_16411,N_16051,N_16204);
nand U16412 (N_16412,N_16088,N_15768);
and U16413 (N_16413,N_15790,N_16147);
and U16414 (N_16414,N_16162,N_16052);
nand U16415 (N_16415,N_15817,N_15933);
xnor U16416 (N_16416,N_16197,N_15886);
xnor U16417 (N_16417,N_15775,N_15734);
nor U16418 (N_16418,N_15667,N_16170);
xor U16419 (N_16419,N_16010,N_15628);
nand U16420 (N_16420,N_16041,N_15813);
and U16421 (N_16421,N_15855,N_16224);
or U16422 (N_16422,N_16120,N_15983);
nor U16423 (N_16423,N_15830,N_15970);
or U16424 (N_16424,N_15746,N_16006);
xor U16425 (N_16425,N_16103,N_15721);
nor U16426 (N_16426,N_15844,N_16115);
xnor U16427 (N_16427,N_15904,N_16229);
nor U16428 (N_16428,N_16126,N_15901);
nand U16429 (N_16429,N_15695,N_15791);
nand U16430 (N_16430,N_16174,N_15748);
nand U16431 (N_16431,N_16076,N_16203);
xnor U16432 (N_16432,N_16196,N_16239);
xor U16433 (N_16433,N_16108,N_16183);
nand U16434 (N_16434,N_15722,N_15682);
nand U16435 (N_16435,N_16035,N_16007);
nand U16436 (N_16436,N_15860,N_15994);
nand U16437 (N_16437,N_16175,N_15776);
nand U16438 (N_16438,N_15675,N_15826);
and U16439 (N_16439,N_16008,N_16047);
nand U16440 (N_16440,N_15926,N_16193);
or U16441 (N_16441,N_15783,N_15796);
or U16442 (N_16442,N_15997,N_16025);
nand U16443 (N_16443,N_15637,N_16037);
nor U16444 (N_16444,N_15960,N_15837);
nand U16445 (N_16445,N_15954,N_16016);
or U16446 (N_16446,N_15822,N_15804);
and U16447 (N_16447,N_16083,N_15677);
or U16448 (N_16448,N_16038,N_15898);
xnor U16449 (N_16449,N_16000,N_16009);
nand U16450 (N_16450,N_16228,N_15937);
and U16451 (N_16451,N_16058,N_16201);
xor U16452 (N_16452,N_15948,N_15631);
nor U16453 (N_16453,N_15731,N_15973);
and U16454 (N_16454,N_15657,N_15833);
or U16455 (N_16455,N_15757,N_16091);
xnor U16456 (N_16456,N_16132,N_15838);
nor U16457 (N_16457,N_16068,N_15832);
nor U16458 (N_16458,N_15897,N_15691);
nor U16459 (N_16459,N_15836,N_15726);
or U16460 (N_16460,N_15929,N_16199);
xor U16461 (N_16461,N_15742,N_15809);
and U16462 (N_16462,N_16018,N_15661);
xnor U16463 (N_16463,N_16097,N_16223);
xnor U16464 (N_16464,N_16001,N_15906);
or U16465 (N_16465,N_16173,N_15881);
xor U16466 (N_16466,N_16121,N_15827);
nor U16467 (N_16467,N_16221,N_15769);
and U16468 (N_16468,N_15940,N_16156);
nor U16469 (N_16469,N_16059,N_15799);
xnor U16470 (N_16470,N_16192,N_16118);
or U16471 (N_16471,N_16113,N_16082);
nor U16472 (N_16472,N_16164,N_15758);
or U16473 (N_16473,N_16048,N_16028);
nor U16474 (N_16474,N_16114,N_15788);
xor U16475 (N_16475,N_16135,N_15982);
or U16476 (N_16476,N_15888,N_16116);
or U16477 (N_16477,N_15702,N_15992);
xnor U16478 (N_16478,N_15991,N_15956);
nor U16479 (N_16479,N_16158,N_15672);
or U16480 (N_16480,N_16017,N_15767);
or U16481 (N_16481,N_15670,N_15980);
or U16482 (N_16482,N_15632,N_15656);
or U16483 (N_16483,N_16182,N_16216);
and U16484 (N_16484,N_15941,N_15959);
or U16485 (N_16485,N_16098,N_15990);
nand U16486 (N_16486,N_16130,N_15849);
nand U16487 (N_16487,N_15697,N_16178);
nand U16488 (N_16488,N_15957,N_16092);
or U16489 (N_16489,N_15710,N_16206);
xor U16490 (N_16490,N_15671,N_15669);
nor U16491 (N_16491,N_16095,N_15728);
nand U16492 (N_16492,N_15666,N_15663);
xnor U16493 (N_16493,N_15658,N_15872);
and U16494 (N_16494,N_16131,N_15698);
nor U16495 (N_16495,N_15753,N_16245);
nand U16496 (N_16496,N_16014,N_16220);
or U16497 (N_16497,N_15936,N_15841);
or U16498 (N_16498,N_15845,N_15877);
and U16499 (N_16499,N_16043,N_15730);
or U16500 (N_16500,N_15981,N_15863);
or U16501 (N_16501,N_16042,N_16154);
nor U16502 (N_16502,N_15919,N_15950);
and U16503 (N_16503,N_15634,N_16034);
nand U16504 (N_16504,N_16005,N_16168);
and U16505 (N_16505,N_15944,N_15751);
nand U16506 (N_16506,N_15707,N_15892);
xor U16507 (N_16507,N_16078,N_15934);
nand U16508 (N_16508,N_15650,N_15951);
nor U16509 (N_16509,N_16218,N_15735);
or U16510 (N_16510,N_15921,N_15922);
nor U16511 (N_16511,N_16087,N_15625);
and U16512 (N_16512,N_15869,N_15766);
nand U16513 (N_16513,N_15843,N_15999);
nor U16514 (N_16514,N_16089,N_16127);
or U16515 (N_16515,N_16050,N_15744);
nor U16516 (N_16516,N_15764,N_15808);
and U16517 (N_16517,N_16074,N_15740);
and U16518 (N_16518,N_16106,N_16026);
nor U16519 (N_16519,N_15737,N_16143);
nor U16520 (N_16520,N_15903,N_15971);
or U16521 (N_16521,N_15820,N_15763);
nand U16522 (N_16522,N_15928,N_15846);
xnor U16523 (N_16523,N_15984,N_16030);
nor U16524 (N_16524,N_16212,N_16119);
nor U16525 (N_16525,N_15756,N_15866);
and U16526 (N_16526,N_15770,N_15905);
or U16527 (N_16527,N_16191,N_16045);
and U16528 (N_16528,N_16171,N_15795);
and U16529 (N_16529,N_15680,N_15867);
and U16530 (N_16530,N_15645,N_16093);
or U16531 (N_16531,N_16063,N_15975);
or U16532 (N_16532,N_15736,N_15873);
and U16533 (N_16533,N_16159,N_16169);
or U16534 (N_16534,N_15800,N_15760);
or U16535 (N_16535,N_15900,N_15871);
xnor U16536 (N_16536,N_16177,N_16023);
or U16537 (N_16537,N_16110,N_15839);
nor U16538 (N_16538,N_15823,N_15890);
or U16539 (N_16539,N_16205,N_16105);
nor U16540 (N_16540,N_15816,N_16027);
or U16541 (N_16541,N_16140,N_15891);
and U16542 (N_16542,N_16149,N_15927);
nor U16543 (N_16543,N_15723,N_15699);
or U16544 (N_16544,N_16029,N_16150);
xor U16545 (N_16545,N_16099,N_16066);
and U16546 (N_16546,N_16064,N_15995);
nand U16547 (N_16547,N_15889,N_15662);
and U16548 (N_16548,N_15771,N_15966);
xor U16549 (N_16549,N_15989,N_16090);
xor U16550 (N_16550,N_15895,N_15792);
nor U16551 (N_16551,N_16040,N_16031);
and U16552 (N_16552,N_15681,N_16020);
xor U16553 (N_16553,N_15805,N_16233);
nand U16554 (N_16554,N_15825,N_15745);
nor U16555 (N_16555,N_15814,N_15811);
nand U16556 (N_16556,N_16185,N_15908);
nand U16557 (N_16557,N_15646,N_16248);
nor U16558 (N_16558,N_16069,N_16208);
nand U16559 (N_16559,N_16053,N_15850);
and U16560 (N_16560,N_15862,N_16194);
nand U16561 (N_16561,N_15909,N_16198);
or U16562 (N_16562,N_16084,N_16148);
nand U16563 (N_16563,N_15914,N_15630);
xor U16564 (N_16564,N_15808,N_15777);
xnor U16565 (N_16565,N_16201,N_15731);
nand U16566 (N_16566,N_15661,N_15837);
nand U16567 (N_16567,N_15654,N_16059);
xor U16568 (N_16568,N_16099,N_15853);
xnor U16569 (N_16569,N_15935,N_16181);
nor U16570 (N_16570,N_15819,N_15689);
and U16571 (N_16571,N_16009,N_16092);
xnor U16572 (N_16572,N_15712,N_15855);
nand U16573 (N_16573,N_15899,N_16042);
or U16574 (N_16574,N_16039,N_16155);
xnor U16575 (N_16575,N_16033,N_15824);
nor U16576 (N_16576,N_15773,N_16059);
xnor U16577 (N_16577,N_16186,N_15797);
xor U16578 (N_16578,N_16209,N_16035);
nor U16579 (N_16579,N_16125,N_16080);
or U16580 (N_16580,N_16015,N_16033);
nor U16581 (N_16581,N_15706,N_15748);
xnor U16582 (N_16582,N_16156,N_15910);
or U16583 (N_16583,N_15799,N_15705);
nor U16584 (N_16584,N_15950,N_15836);
xnor U16585 (N_16585,N_15966,N_15838);
xor U16586 (N_16586,N_16238,N_15877);
xnor U16587 (N_16587,N_16187,N_15864);
and U16588 (N_16588,N_15936,N_15918);
nand U16589 (N_16589,N_16118,N_15961);
nand U16590 (N_16590,N_16206,N_15838);
nand U16591 (N_16591,N_16147,N_15960);
nand U16592 (N_16592,N_15962,N_16242);
nor U16593 (N_16593,N_15684,N_16104);
xor U16594 (N_16594,N_15660,N_16054);
nand U16595 (N_16595,N_15646,N_15877);
and U16596 (N_16596,N_16214,N_16083);
xnor U16597 (N_16597,N_15901,N_15643);
xor U16598 (N_16598,N_15700,N_15933);
nor U16599 (N_16599,N_15749,N_15881);
nand U16600 (N_16600,N_15753,N_15720);
nand U16601 (N_16601,N_16224,N_15941);
xor U16602 (N_16602,N_15798,N_15748);
or U16603 (N_16603,N_15671,N_16024);
or U16604 (N_16604,N_15677,N_15765);
or U16605 (N_16605,N_16088,N_15876);
nor U16606 (N_16606,N_15726,N_15725);
nor U16607 (N_16607,N_16216,N_15822);
or U16608 (N_16608,N_16060,N_15885);
nand U16609 (N_16609,N_16023,N_16123);
nor U16610 (N_16610,N_16245,N_15685);
or U16611 (N_16611,N_16149,N_16211);
xor U16612 (N_16612,N_16081,N_16144);
nand U16613 (N_16613,N_15707,N_15974);
or U16614 (N_16614,N_15880,N_16057);
xor U16615 (N_16615,N_16240,N_16222);
or U16616 (N_16616,N_15754,N_16089);
nand U16617 (N_16617,N_16173,N_16147);
and U16618 (N_16618,N_16136,N_15940);
nor U16619 (N_16619,N_15954,N_16082);
xor U16620 (N_16620,N_15658,N_15849);
nor U16621 (N_16621,N_16080,N_15823);
xnor U16622 (N_16622,N_15762,N_16110);
nor U16623 (N_16623,N_16042,N_15873);
nand U16624 (N_16624,N_15769,N_16119);
nor U16625 (N_16625,N_16203,N_15718);
or U16626 (N_16626,N_16181,N_16191);
xnor U16627 (N_16627,N_16018,N_15996);
or U16628 (N_16628,N_15797,N_15640);
nor U16629 (N_16629,N_15977,N_15664);
or U16630 (N_16630,N_15714,N_15923);
or U16631 (N_16631,N_16099,N_15789);
and U16632 (N_16632,N_16082,N_15815);
and U16633 (N_16633,N_15861,N_15682);
nor U16634 (N_16634,N_16212,N_16248);
nor U16635 (N_16635,N_16133,N_15839);
nand U16636 (N_16636,N_15986,N_15746);
nor U16637 (N_16637,N_16083,N_15762);
xor U16638 (N_16638,N_15646,N_16183);
nor U16639 (N_16639,N_15733,N_15809);
and U16640 (N_16640,N_15917,N_15807);
and U16641 (N_16641,N_16061,N_15792);
nand U16642 (N_16642,N_15638,N_15745);
xnor U16643 (N_16643,N_15910,N_16128);
nor U16644 (N_16644,N_16216,N_15821);
or U16645 (N_16645,N_15863,N_15717);
and U16646 (N_16646,N_15923,N_15715);
nor U16647 (N_16647,N_15694,N_16202);
or U16648 (N_16648,N_16179,N_16077);
or U16649 (N_16649,N_15991,N_15884);
xnor U16650 (N_16650,N_16245,N_15955);
xnor U16651 (N_16651,N_15812,N_15686);
nor U16652 (N_16652,N_15756,N_16024);
xnor U16653 (N_16653,N_16067,N_16127);
nand U16654 (N_16654,N_16104,N_15745);
nor U16655 (N_16655,N_16127,N_15856);
nand U16656 (N_16656,N_15766,N_15676);
nand U16657 (N_16657,N_15779,N_15685);
xor U16658 (N_16658,N_15888,N_16231);
xnor U16659 (N_16659,N_16011,N_16187);
nand U16660 (N_16660,N_15654,N_16170);
nor U16661 (N_16661,N_15898,N_15681);
nor U16662 (N_16662,N_15828,N_15626);
or U16663 (N_16663,N_15631,N_15763);
or U16664 (N_16664,N_15960,N_15885);
or U16665 (N_16665,N_15796,N_16044);
nand U16666 (N_16666,N_16020,N_15776);
and U16667 (N_16667,N_16125,N_15735);
and U16668 (N_16668,N_16008,N_16116);
nand U16669 (N_16669,N_16243,N_15912);
or U16670 (N_16670,N_15903,N_16237);
xor U16671 (N_16671,N_15777,N_15725);
nand U16672 (N_16672,N_15751,N_16032);
or U16673 (N_16673,N_15636,N_16075);
xor U16674 (N_16674,N_15882,N_16198);
nand U16675 (N_16675,N_15892,N_16168);
xor U16676 (N_16676,N_16101,N_15948);
nand U16677 (N_16677,N_16030,N_15972);
nand U16678 (N_16678,N_15871,N_16203);
xnor U16679 (N_16679,N_16055,N_15898);
or U16680 (N_16680,N_15641,N_15666);
xnor U16681 (N_16681,N_15995,N_16186);
xor U16682 (N_16682,N_15678,N_16103);
nor U16683 (N_16683,N_15800,N_16209);
and U16684 (N_16684,N_15694,N_15932);
xnor U16685 (N_16685,N_15664,N_15856);
xnor U16686 (N_16686,N_16111,N_16213);
nor U16687 (N_16687,N_15967,N_15969);
and U16688 (N_16688,N_15858,N_16221);
and U16689 (N_16689,N_16032,N_15790);
xnor U16690 (N_16690,N_15658,N_15955);
xnor U16691 (N_16691,N_15930,N_15968);
and U16692 (N_16692,N_15706,N_16128);
nand U16693 (N_16693,N_15744,N_16047);
nand U16694 (N_16694,N_15941,N_15771);
or U16695 (N_16695,N_16006,N_16132);
nor U16696 (N_16696,N_15671,N_15745);
nand U16697 (N_16697,N_16134,N_15729);
or U16698 (N_16698,N_15937,N_15816);
xor U16699 (N_16699,N_15830,N_15769);
and U16700 (N_16700,N_16136,N_15892);
nor U16701 (N_16701,N_15732,N_16231);
xnor U16702 (N_16702,N_16033,N_15772);
xnor U16703 (N_16703,N_15919,N_15815);
or U16704 (N_16704,N_15758,N_16126);
or U16705 (N_16705,N_15843,N_15870);
nand U16706 (N_16706,N_16152,N_16019);
xnor U16707 (N_16707,N_16196,N_15801);
xor U16708 (N_16708,N_15825,N_16141);
nor U16709 (N_16709,N_16099,N_15857);
and U16710 (N_16710,N_15897,N_15639);
and U16711 (N_16711,N_15906,N_15705);
and U16712 (N_16712,N_16234,N_16050);
and U16713 (N_16713,N_16160,N_15877);
and U16714 (N_16714,N_16179,N_16034);
xnor U16715 (N_16715,N_15955,N_15793);
or U16716 (N_16716,N_15704,N_15905);
or U16717 (N_16717,N_15721,N_15832);
xor U16718 (N_16718,N_15795,N_15652);
nor U16719 (N_16719,N_16022,N_15970);
and U16720 (N_16720,N_15992,N_15989);
nor U16721 (N_16721,N_15880,N_15865);
xor U16722 (N_16722,N_15977,N_15965);
nor U16723 (N_16723,N_15743,N_15625);
or U16724 (N_16724,N_16203,N_15719);
and U16725 (N_16725,N_16170,N_15725);
nor U16726 (N_16726,N_16042,N_15933);
nor U16727 (N_16727,N_15636,N_16175);
nor U16728 (N_16728,N_16162,N_15671);
xor U16729 (N_16729,N_15975,N_15822);
or U16730 (N_16730,N_15981,N_15781);
and U16731 (N_16731,N_16027,N_15789);
or U16732 (N_16732,N_15852,N_15983);
and U16733 (N_16733,N_15863,N_15656);
xor U16734 (N_16734,N_15984,N_15801);
or U16735 (N_16735,N_15788,N_15900);
and U16736 (N_16736,N_16235,N_16218);
and U16737 (N_16737,N_16159,N_15720);
xnor U16738 (N_16738,N_15633,N_15812);
or U16739 (N_16739,N_15929,N_16204);
or U16740 (N_16740,N_15920,N_15820);
nor U16741 (N_16741,N_15823,N_16120);
xnor U16742 (N_16742,N_15725,N_15728);
or U16743 (N_16743,N_16217,N_15776);
nand U16744 (N_16744,N_16088,N_15777);
and U16745 (N_16745,N_15772,N_15994);
nand U16746 (N_16746,N_15897,N_16059);
nand U16747 (N_16747,N_15951,N_15953);
xor U16748 (N_16748,N_15997,N_15629);
or U16749 (N_16749,N_16220,N_16023);
nand U16750 (N_16750,N_16115,N_16150);
xnor U16751 (N_16751,N_16210,N_16072);
nand U16752 (N_16752,N_15876,N_15869);
nor U16753 (N_16753,N_15983,N_16213);
nor U16754 (N_16754,N_15779,N_16211);
and U16755 (N_16755,N_16203,N_15924);
or U16756 (N_16756,N_16099,N_15625);
and U16757 (N_16757,N_16085,N_15784);
nand U16758 (N_16758,N_15696,N_15810);
nand U16759 (N_16759,N_16095,N_15808);
and U16760 (N_16760,N_15808,N_16102);
nor U16761 (N_16761,N_16005,N_16180);
and U16762 (N_16762,N_15652,N_15769);
and U16763 (N_16763,N_15993,N_16188);
xnor U16764 (N_16764,N_16072,N_16218);
and U16765 (N_16765,N_15706,N_16228);
nor U16766 (N_16766,N_15655,N_16199);
xor U16767 (N_16767,N_15891,N_16049);
nand U16768 (N_16768,N_15674,N_16225);
or U16769 (N_16769,N_15860,N_15976);
nor U16770 (N_16770,N_16062,N_16192);
nand U16771 (N_16771,N_16018,N_15697);
xnor U16772 (N_16772,N_16027,N_15815);
nand U16773 (N_16773,N_15748,N_15862);
xor U16774 (N_16774,N_15655,N_15970);
or U16775 (N_16775,N_15809,N_16214);
nor U16776 (N_16776,N_16221,N_16020);
xor U16777 (N_16777,N_15894,N_16008);
and U16778 (N_16778,N_16010,N_15651);
or U16779 (N_16779,N_16043,N_15754);
or U16780 (N_16780,N_16055,N_15857);
and U16781 (N_16781,N_15658,N_15910);
and U16782 (N_16782,N_15882,N_16162);
and U16783 (N_16783,N_15790,N_15997);
and U16784 (N_16784,N_15994,N_16054);
or U16785 (N_16785,N_16064,N_16106);
xor U16786 (N_16786,N_15973,N_16136);
nand U16787 (N_16787,N_15906,N_15996);
xnor U16788 (N_16788,N_15791,N_16245);
nor U16789 (N_16789,N_15891,N_16231);
nor U16790 (N_16790,N_15706,N_15907);
nand U16791 (N_16791,N_16229,N_15867);
or U16792 (N_16792,N_15934,N_15689);
nor U16793 (N_16793,N_16238,N_15794);
nor U16794 (N_16794,N_15853,N_16086);
xor U16795 (N_16795,N_16070,N_15720);
nand U16796 (N_16796,N_15847,N_16197);
or U16797 (N_16797,N_15654,N_15777);
nand U16798 (N_16798,N_15995,N_16005);
and U16799 (N_16799,N_15796,N_15844);
and U16800 (N_16800,N_16035,N_15958);
nor U16801 (N_16801,N_16082,N_15735);
nand U16802 (N_16802,N_16033,N_15677);
nand U16803 (N_16803,N_15823,N_15694);
xor U16804 (N_16804,N_15816,N_15685);
nor U16805 (N_16805,N_16093,N_15643);
or U16806 (N_16806,N_15637,N_15920);
nand U16807 (N_16807,N_16020,N_16085);
nor U16808 (N_16808,N_16057,N_16160);
xnor U16809 (N_16809,N_15888,N_15781);
xnor U16810 (N_16810,N_16237,N_15684);
xnor U16811 (N_16811,N_15892,N_15834);
nor U16812 (N_16812,N_15946,N_15839);
xnor U16813 (N_16813,N_15823,N_16071);
xor U16814 (N_16814,N_16001,N_16061);
nor U16815 (N_16815,N_16101,N_15695);
nand U16816 (N_16816,N_15768,N_15900);
nand U16817 (N_16817,N_16139,N_15942);
nor U16818 (N_16818,N_16179,N_15778);
xor U16819 (N_16819,N_15755,N_15932);
and U16820 (N_16820,N_15889,N_15689);
or U16821 (N_16821,N_16065,N_16196);
and U16822 (N_16822,N_15717,N_15804);
and U16823 (N_16823,N_16025,N_16081);
xnor U16824 (N_16824,N_15630,N_15852);
nand U16825 (N_16825,N_15809,N_15972);
xnor U16826 (N_16826,N_15836,N_16076);
and U16827 (N_16827,N_15844,N_15657);
or U16828 (N_16828,N_15978,N_15649);
nor U16829 (N_16829,N_15698,N_15695);
or U16830 (N_16830,N_15984,N_15944);
or U16831 (N_16831,N_15629,N_16221);
nand U16832 (N_16832,N_16195,N_15662);
or U16833 (N_16833,N_15885,N_15972);
nor U16834 (N_16834,N_16080,N_15833);
nand U16835 (N_16835,N_16011,N_15814);
or U16836 (N_16836,N_15939,N_15773);
or U16837 (N_16837,N_16204,N_15886);
nand U16838 (N_16838,N_16111,N_16230);
xnor U16839 (N_16839,N_15691,N_15880);
or U16840 (N_16840,N_15640,N_16229);
and U16841 (N_16841,N_15872,N_16206);
nand U16842 (N_16842,N_15952,N_15943);
nor U16843 (N_16843,N_15845,N_15829);
xnor U16844 (N_16844,N_15800,N_15727);
nor U16845 (N_16845,N_16184,N_16061);
and U16846 (N_16846,N_15923,N_16026);
and U16847 (N_16847,N_15897,N_16187);
nand U16848 (N_16848,N_15793,N_15646);
or U16849 (N_16849,N_16188,N_15900);
xor U16850 (N_16850,N_15834,N_16108);
or U16851 (N_16851,N_16002,N_16247);
nor U16852 (N_16852,N_16046,N_16177);
nand U16853 (N_16853,N_15679,N_16088);
nor U16854 (N_16854,N_16000,N_15842);
or U16855 (N_16855,N_16034,N_16124);
nand U16856 (N_16856,N_15872,N_15675);
nand U16857 (N_16857,N_16070,N_15994);
nand U16858 (N_16858,N_15948,N_15679);
nand U16859 (N_16859,N_16190,N_16119);
or U16860 (N_16860,N_15937,N_15703);
nand U16861 (N_16861,N_16165,N_15936);
or U16862 (N_16862,N_15729,N_16146);
or U16863 (N_16863,N_15959,N_16199);
xor U16864 (N_16864,N_15720,N_16051);
nor U16865 (N_16865,N_15792,N_15795);
and U16866 (N_16866,N_15926,N_15755);
xnor U16867 (N_16867,N_16209,N_15842);
and U16868 (N_16868,N_15920,N_15709);
and U16869 (N_16869,N_15854,N_15970);
or U16870 (N_16870,N_16014,N_16050);
nand U16871 (N_16871,N_15646,N_15801);
xnor U16872 (N_16872,N_15916,N_16213);
or U16873 (N_16873,N_16077,N_15741);
and U16874 (N_16874,N_15894,N_15943);
xor U16875 (N_16875,N_16737,N_16493);
nand U16876 (N_16876,N_16814,N_16730);
xnor U16877 (N_16877,N_16425,N_16822);
or U16878 (N_16878,N_16422,N_16476);
nor U16879 (N_16879,N_16804,N_16679);
xor U16880 (N_16880,N_16395,N_16328);
nor U16881 (N_16881,N_16472,N_16464);
or U16882 (N_16882,N_16580,N_16776);
xor U16883 (N_16883,N_16640,N_16429);
or U16884 (N_16884,N_16346,N_16707);
nor U16885 (N_16885,N_16303,N_16269);
nor U16886 (N_16886,N_16528,N_16529);
xnor U16887 (N_16887,N_16443,N_16811);
nor U16888 (N_16888,N_16389,N_16274);
nor U16889 (N_16889,N_16576,N_16742);
nand U16890 (N_16890,N_16584,N_16265);
nand U16891 (N_16891,N_16502,N_16579);
nand U16892 (N_16892,N_16668,N_16763);
or U16893 (N_16893,N_16681,N_16499);
nor U16894 (N_16894,N_16733,N_16673);
or U16895 (N_16895,N_16504,N_16526);
or U16896 (N_16896,N_16294,N_16571);
nand U16897 (N_16897,N_16678,N_16827);
or U16898 (N_16898,N_16390,N_16541);
xnor U16899 (N_16899,N_16857,N_16451);
nand U16900 (N_16900,N_16849,N_16563);
nand U16901 (N_16901,N_16364,N_16470);
nor U16902 (N_16902,N_16825,N_16802);
and U16903 (N_16903,N_16765,N_16672);
nand U16904 (N_16904,N_16700,N_16310);
or U16905 (N_16905,N_16292,N_16725);
and U16906 (N_16906,N_16358,N_16869);
nand U16907 (N_16907,N_16257,N_16585);
and U16908 (N_16908,N_16551,N_16850);
nand U16909 (N_16909,N_16354,N_16340);
or U16910 (N_16910,N_16839,N_16626);
and U16911 (N_16911,N_16759,N_16782);
nor U16912 (N_16912,N_16637,N_16515);
xnor U16913 (N_16913,N_16342,N_16512);
or U16914 (N_16914,N_16773,N_16721);
nand U16915 (N_16915,N_16578,N_16345);
or U16916 (N_16916,N_16293,N_16307);
xnor U16917 (N_16917,N_16468,N_16666);
or U16918 (N_16918,N_16692,N_16736);
or U16919 (N_16919,N_16517,N_16750);
nor U16920 (N_16920,N_16557,N_16483);
nand U16921 (N_16921,N_16271,N_16683);
and U16922 (N_16922,N_16829,N_16255);
nand U16923 (N_16923,N_16462,N_16300);
or U16924 (N_16924,N_16491,N_16795);
xor U16925 (N_16925,N_16769,N_16705);
and U16926 (N_16926,N_16812,N_16560);
or U16927 (N_16927,N_16383,N_16756);
nor U16928 (N_16928,N_16416,N_16531);
and U16929 (N_16929,N_16800,N_16538);
and U16930 (N_16930,N_16284,N_16537);
nand U16931 (N_16931,N_16507,N_16665);
and U16932 (N_16932,N_16868,N_16315);
and U16933 (N_16933,N_16574,N_16497);
or U16934 (N_16934,N_16290,N_16494);
or U16935 (N_16935,N_16412,N_16847);
and U16936 (N_16936,N_16682,N_16696);
or U16937 (N_16937,N_16394,N_16319);
or U16938 (N_16938,N_16349,N_16510);
and U16939 (N_16939,N_16282,N_16837);
nand U16940 (N_16940,N_16691,N_16758);
xnor U16941 (N_16941,N_16323,N_16550);
nor U16942 (N_16942,N_16455,N_16488);
nand U16943 (N_16943,N_16598,N_16757);
nand U16944 (N_16944,N_16820,N_16302);
xnor U16945 (N_16945,N_16411,N_16748);
or U16946 (N_16946,N_16465,N_16806);
and U16947 (N_16947,N_16830,N_16701);
and U16948 (N_16948,N_16370,N_16699);
or U16949 (N_16949,N_16309,N_16546);
or U16950 (N_16950,N_16562,N_16365);
or U16951 (N_16951,N_16657,N_16709);
nor U16952 (N_16952,N_16771,N_16596);
or U16953 (N_16953,N_16329,N_16287);
nor U16954 (N_16954,N_16407,N_16556);
and U16955 (N_16955,N_16259,N_16306);
nand U16956 (N_16956,N_16481,N_16577);
and U16957 (N_16957,N_16836,N_16446);
and U16958 (N_16958,N_16608,N_16856);
nand U16959 (N_16959,N_16522,N_16703);
nor U16960 (N_16960,N_16855,N_16559);
xor U16961 (N_16961,N_16713,N_16660);
xor U16962 (N_16962,N_16723,N_16607);
and U16963 (N_16963,N_16648,N_16780);
nor U16964 (N_16964,N_16376,N_16508);
xnor U16965 (N_16965,N_16469,N_16454);
nand U16966 (N_16966,N_16788,N_16357);
nor U16967 (N_16967,N_16663,N_16409);
xnor U16968 (N_16968,N_16266,N_16420);
or U16969 (N_16969,N_16430,N_16459);
or U16970 (N_16970,N_16369,N_16728);
xnor U16971 (N_16971,N_16783,N_16513);
xor U16972 (N_16972,N_16487,N_16819);
nor U16973 (N_16973,N_16646,N_16263);
nor U16974 (N_16974,N_16642,N_16661);
and U16975 (N_16975,N_16729,N_16521);
or U16976 (N_16976,N_16397,N_16654);
or U16977 (N_16977,N_16359,N_16414);
xor U16978 (N_16978,N_16356,N_16784);
and U16979 (N_16979,N_16866,N_16588);
or U16980 (N_16980,N_16438,N_16623);
nand U16981 (N_16981,N_16644,N_16848);
and U16982 (N_16982,N_16523,N_16870);
nor U16983 (N_16983,N_16832,N_16851);
or U16984 (N_16984,N_16272,N_16859);
or U16985 (N_16985,N_16872,N_16698);
nand U16986 (N_16986,N_16382,N_16308);
xor U16987 (N_16987,N_16778,N_16317);
or U16988 (N_16988,N_16344,N_16643);
xnor U16989 (N_16989,N_16413,N_16432);
xor U16990 (N_16990,N_16313,N_16500);
nand U16991 (N_16991,N_16400,N_16594);
xnor U16992 (N_16992,N_16418,N_16867);
xnor U16993 (N_16993,N_16461,N_16600);
xnor U16994 (N_16994,N_16658,N_16480);
nor U16995 (N_16995,N_16296,N_16599);
nand U16996 (N_16996,N_16575,N_16860);
or U16997 (N_16997,N_16656,N_16690);
nand U16998 (N_16998,N_16402,N_16677);
nor U16999 (N_16999,N_16466,N_16388);
or U17000 (N_17000,N_16817,N_16536);
xor U17001 (N_17001,N_16570,N_16670);
nand U17002 (N_17002,N_16652,N_16372);
nand U17003 (N_17003,N_16410,N_16612);
xnor U17004 (N_17004,N_16366,N_16337);
or U17005 (N_17005,N_16798,N_16331);
and U17006 (N_17006,N_16447,N_16601);
nor U17007 (N_17007,N_16613,N_16761);
nor U17008 (N_17008,N_16264,N_16277);
xnor U17009 (N_17009,N_16726,N_16740);
nor U17010 (N_17010,N_16650,N_16821);
nor U17011 (N_17011,N_16715,N_16281);
xnor U17012 (N_17012,N_16327,N_16621);
and U17013 (N_17013,N_16831,N_16635);
xor U17014 (N_17014,N_16602,N_16473);
or U17015 (N_17015,N_16714,N_16338);
or U17016 (N_17016,N_16744,N_16341);
nand U17017 (N_17017,N_16605,N_16445);
or U17018 (N_17018,N_16863,N_16801);
nor U17019 (N_17019,N_16318,N_16506);
nor U17020 (N_17020,N_16297,N_16826);
or U17021 (N_17021,N_16845,N_16371);
nand U17022 (N_17022,N_16322,N_16535);
and U17023 (N_17023,N_16336,N_16270);
xnor U17024 (N_17024,N_16375,N_16693);
or U17025 (N_17025,N_16450,N_16633);
or U17026 (N_17026,N_16316,N_16791);
and U17027 (N_17027,N_16841,N_16620);
nor U17028 (N_17028,N_16655,N_16355);
nor U17029 (N_17029,N_16734,N_16424);
or U17030 (N_17030,N_16545,N_16645);
nor U17031 (N_17031,N_16628,N_16311);
or U17032 (N_17032,N_16632,N_16647);
xor U17033 (N_17033,N_16518,N_16779);
or U17034 (N_17034,N_16485,N_16426);
nand U17035 (N_17035,N_16511,N_16764);
xnor U17036 (N_17036,N_16732,N_16343);
nor U17037 (N_17037,N_16428,N_16254);
xnor U17038 (N_17038,N_16564,N_16482);
nor U17039 (N_17039,N_16840,N_16842);
xor U17040 (N_17040,N_16838,N_16735);
nor U17041 (N_17041,N_16865,N_16630);
or U17042 (N_17042,N_16688,N_16398);
xnor U17043 (N_17043,N_16492,N_16267);
nand U17044 (N_17044,N_16680,N_16694);
or U17045 (N_17045,N_16717,N_16258);
and U17046 (N_17046,N_16671,N_16861);
nand U17047 (N_17047,N_16285,N_16864);
nor U17048 (N_17048,N_16770,N_16361);
and U17049 (N_17049,N_16572,N_16467);
nor U17050 (N_17050,N_16835,N_16458);
or U17051 (N_17051,N_16475,N_16796);
nand U17052 (N_17052,N_16794,N_16609);
nor U17053 (N_17053,N_16495,N_16435);
xor U17054 (N_17054,N_16568,N_16706);
nand U17055 (N_17055,N_16716,N_16874);
and U17056 (N_17056,N_16719,N_16675);
xor U17057 (N_17057,N_16423,N_16766);
and U17058 (N_17058,N_16738,N_16543);
nor U17059 (N_17059,N_16415,N_16380);
nand U17060 (N_17060,N_16253,N_16363);
or U17061 (N_17061,N_16404,N_16421);
or U17062 (N_17062,N_16772,N_16697);
xor U17063 (N_17063,N_16662,N_16743);
and U17064 (N_17064,N_16790,N_16519);
xor U17065 (N_17065,N_16751,N_16843);
nor U17066 (N_17066,N_16573,N_16616);
nor U17067 (N_17067,N_16614,N_16619);
and U17068 (N_17068,N_16664,N_16419);
nor U17069 (N_17069,N_16540,N_16604);
xnor U17070 (N_17070,N_16289,N_16286);
nor U17071 (N_17071,N_16745,N_16676);
nor U17072 (N_17072,N_16813,N_16325);
nor U17073 (N_17073,N_16542,N_16288);
and U17074 (N_17074,N_16718,N_16687);
and U17075 (N_17075,N_16797,N_16332);
nor U17076 (N_17076,N_16651,N_16440);
nand U17077 (N_17077,N_16314,N_16312);
nand U17078 (N_17078,N_16828,N_16787);
nand U17079 (N_17079,N_16275,N_16752);
nor U17080 (N_17080,N_16622,N_16674);
and U17081 (N_17081,N_16582,N_16471);
and U17082 (N_17082,N_16815,N_16378);
and U17083 (N_17083,N_16393,N_16304);
nand U17084 (N_17084,N_16280,N_16548);
xnor U17085 (N_17085,N_16478,N_16854);
nor U17086 (N_17086,N_16767,N_16639);
nand U17087 (N_17087,N_16659,N_16603);
nand U17088 (N_17088,N_16809,N_16268);
xor U17089 (N_17089,N_16256,N_16509);
or U17090 (N_17090,N_16610,N_16374);
nand U17091 (N_17091,N_16449,N_16786);
nand U17092 (N_17092,N_16641,N_16534);
or U17093 (N_17093,N_16305,N_16514);
nor U17094 (N_17094,N_16689,N_16373);
xor U17095 (N_17095,N_16739,N_16260);
nor U17096 (N_17096,N_16516,N_16777);
nand U17097 (N_17097,N_16808,N_16334);
nand U17098 (N_17098,N_16871,N_16524);
nand U17099 (N_17099,N_16362,N_16544);
nor U17100 (N_17100,N_16252,N_16460);
nor U17101 (N_17101,N_16749,N_16846);
xnor U17102 (N_17102,N_16406,N_16486);
nand U17103 (N_17103,N_16417,N_16781);
nand U17104 (N_17104,N_16427,N_16439);
nand U17105 (N_17105,N_16554,N_16368);
nor U17106 (N_17106,N_16532,N_16477);
xor U17107 (N_17107,N_16589,N_16834);
nand U17108 (N_17108,N_16629,N_16333);
nor U17109 (N_17109,N_16792,N_16261);
nand U17110 (N_17110,N_16347,N_16724);
nor U17111 (N_17111,N_16527,N_16754);
and U17112 (N_17112,N_16753,N_16324);
or U17113 (N_17113,N_16384,N_16503);
xor U17114 (N_17114,N_16789,N_16597);
or U17115 (N_17115,N_16401,N_16624);
nand U17116 (N_17116,N_16442,N_16377);
or U17117 (N_17117,N_16591,N_16561);
or U17118 (N_17118,N_16379,N_16391);
and U17119 (N_17119,N_16403,N_16539);
nand U17120 (N_17120,N_16436,N_16649);
nand U17121 (N_17121,N_16712,N_16853);
xnor U17122 (N_17122,N_16452,N_16685);
nand U17123 (N_17123,N_16823,N_16279);
nand U17124 (N_17124,N_16708,N_16533);
xor U17125 (N_17125,N_16722,N_16810);
or U17126 (N_17126,N_16775,N_16731);
and U17127 (N_17127,N_16484,N_16755);
nand U17128 (N_17128,N_16456,N_16262);
or U17129 (N_17129,N_16530,N_16760);
nor U17130 (N_17130,N_16392,N_16321);
and U17131 (N_17131,N_16553,N_16453);
and U17132 (N_17132,N_16295,N_16552);
or U17133 (N_17133,N_16489,N_16405);
nor U17134 (N_17134,N_16833,N_16567);
nor U17135 (N_17135,N_16824,N_16555);
and U17136 (N_17136,N_16704,N_16581);
nor U17137 (N_17137,N_16348,N_16520);
and U17138 (N_17138,N_16593,N_16352);
nor U17139 (N_17139,N_16768,N_16501);
nand U17140 (N_17140,N_16448,N_16862);
nor U17141 (N_17141,N_16844,N_16618);
or U17142 (N_17142,N_16463,N_16278);
nor U17143 (N_17143,N_16565,N_16431);
or U17144 (N_17144,N_16805,N_16852);
nand U17145 (N_17145,N_16762,N_16399);
and U17146 (N_17146,N_16434,N_16276);
or U17147 (N_17147,N_16339,N_16615);
or U17148 (N_17148,N_16818,N_16433);
nor U17149 (N_17149,N_16686,N_16525);
nor U17150 (N_17150,N_16505,N_16496);
nand U17151 (N_17151,N_16360,N_16479);
and U17152 (N_17152,N_16606,N_16350);
and U17153 (N_17153,N_16695,N_16335);
and U17154 (N_17154,N_16387,N_16558);
nand U17155 (N_17155,N_16586,N_16627);
or U17156 (N_17156,N_16741,N_16547);
nor U17157 (N_17157,N_16638,N_16273);
and U17158 (N_17158,N_16711,N_16569);
xor U17159 (N_17159,N_16298,N_16595);
xor U17160 (N_17160,N_16611,N_16634);
nand U17161 (N_17161,N_16386,N_16250);
or U17162 (N_17162,N_16720,N_16631);
nor U17163 (N_17163,N_16549,N_16653);
nand U17164 (N_17164,N_16587,N_16441);
and U17165 (N_17165,N_16299,N_16408);
nor U17166 (N_17166,N_16437,N_16873);
and U17167 (N_17167,N_16474,N_16283);
and U17168 (N_17168,N_16803,N_16381);
xor U17169 (N_17169,N_16590,N_16774);
xor U17170 (N_17170,N_16793,N_16746);
xor U17171 (N_17171,N_16353,N_16684);
nor U17172 (N_17172,N_16251,N_16444);
nand U17173 (N_17173,N_16807,N_16367);
or U17174 (N_17174,N_16799,N_16301);
nor U17175 (N_17175,N_16667,N_16727);
nand U17176 (N_17176,N_16625,N_16291);
or U17177 (N_17177,N_16583,N_16858);
nand U17178 (N_17178,N_16702,N_16669);
nand U17179 (N_17179,N_16330,N_16396);
xor U17180 (N_17180,N_16636,N_16490);
and U17181 (N_17181,N_16816,N_16617);
and U17182 (N_17182,N_16351,N_16710);
and U17183 (N_17183,N_16747,N_16457);
xnor U17184 (N_17184,N_16592,N_16566);
xor U17185 (N_17185,N_16498,N_16785);
or U17186 (N_17186,N_16320,N_16326);
nor U17187 (N_17187,N_16385,N_16755);
xnor U17188 (N_17188,N_16379,N_16314);
nand U17189 (N_17189,N_16773,N_16744);
xor U17190 (N_17190,N_16699,N_16842);
and U17191 (N_17191,N_16497,N_16308);
and U17192 (N_17192,N_16831,N_16400);
or U17193 (N_17193,N_16517,N_16808);
or U17194 (N_17194,N_16823,N_16491);
and U17195 (N_17195,N_16740,N_16790);
nor U17196 (N_17196,N_16296,N_16749);
and U17197 (N_17197,N_16380,N_16381);
xnor U17198 (N_17198,N_16823,N_16446);
nor U17199 (N_17199,N_16708,N_16454);
or U17200 (N_17200,N_16264,N_16859);
and U17201 (N_17201,N_16469,N_16821);
or U17202 (N_17202,N_16773,N_16726);
nor U17203 (N_17203,N_16573,N_16423);
or U17204 (N_17204,N_16617,N_16772);
nand U17205 (N_17205,N_16709,N_16382);
nor U17206 (N_17206,N_16589,N_16733);
and U17207 (N_17207,N_16451,N_16637);
nand U17208 (N_17208,N_16794,N_16473);
or U17209 (N_17209,N_16467,N_16673);
or U17210 (N_17210,N_16544,N_16682);
nand U17211 (N_17211,N_16592,N_16697);
nor U17212 (N_17212,N_16700,N_16450);
and U17213 (N_17213,N_16279,N_16818);
and U17214 (N_17214,N_16796,N_16536);
nor U17215 (N_17215,N_16506,N_16366);
nor U17216 (N_17216,N_16546,N_16791);
nand U17217 (N_17217,N_16436,N_16555);
and U17218 (N_17218,N_16257,N_16747);
nand U17219 (N_17219,N_16421,N_16265);
xor U17220 (N_17220,N_16584,N_16822);
or U17221 (N_17221,N_16440,N_16291);
or U17222 (N_17222,N_16325,N_16308);
or U17223 (N_17223,N_16691,N_16841);
xnor U17224 (N_17224,N_16430,N_16381);
and U17225 (N_17225,N_16590,N_16537);
or U17226 (N_17226,N_16706,N_16672);
nor U17227 (N_17227,N_16361,N_16601);
or U17228 (N_17228,N_16293,N_16607);
xnor U17229 (N_17229,N_16271,N_16867);
and U17230 (N_17230,N_16723,N_16510);
nor U17231 (N_17231,N_16307,N_16546);
nand U17232 (N_17232,N_16369,N_16721);
xnor U17233 (N_17233,N_16368,N_16557);
nor U17234 (N_17234,N_16545,N_16534);
nand U17235 (N_17235,N_16832,N_16315);
xnor U17236 (N_17236,N_16426,N_16725);
xnor U17237 (N_17237,N_16400,N_16852);
nor U17238 (N_17238,N_16567,N_16407);
nor U17239 (N_17239,N_16815,N_16744);
or U17240 (N_17240,N_16307,N_16487);
nand U17241 (N_17241,N_16602,N_16343);
xor U17242 (N_17242,N_16366,N_16363);
nor U17243 (N_17243,N_16834,N_16411);
and U17244 (N_17244,N_16862,N_16574);
or U17245 (N_17245,N_16496,N_16589);
nand U17246 (N_17246,N_16420,N_16654);
nand U17247 (N_17247,N_16512,N_16693);
and U17248 (N_17248,N_16303,N_16618);
or U17249 (N_17249,N_16587,N_16554);
nand U17250 (N_17250,N_16658,N_16783);
xnor U17251 (N_17251,N_16464,N_16785);
or U17252 (N_17252,N_16362,N_16497);
nor U17253 (N_17253,N_16790,N_16509);
nor U17254 (N_17254,N_16682,N_16495);
xor U17255 (N_17255,N_16563,N_16776);
and U17256 (N_17256,N_16497,N_16619);
nand U17257 (N_17257,N_16824,N_16357);
nand U17258 (N_17258,N_16667,N_16277);
and U17259 (N_17259,N_16561,N_16312);
nand U17260 (N_17260,N_16810,N_16747);
or U17261 (N_17261,N_16616,N_16597);
xor U17262 (N_17262,N_16545,N_16313);
nand U17263 (N_17263,N_16398,N_16706);
xor U17264 (N_17264,N_16564,N_16871);
and U17265 (N_17265,N_16427,N_16616);
nor U17266 (N_17266,N_16704,N_16462);
and U17267 (N_17267,N_16268,N_16664);
nand U17268 (N_17268,N_16351,N_16598);
xor U17269 (N_17269,N_16753,N_16430);
nand U17270 (N_17270,N_16690,N_16868);
nand U17271 (N_17271,N_16378,N_16586);
and U17272 (N_17272,N_16646,N_16357);
xor U17273 (N_17273,N_16318,N_16251);
xnor U17274 (N_17274,N_16841,N_16333);
or U17275 (N_17275,N_16762,N_16805);
nor U17276 (N_17276,N_16599,N_16595);
xnor U17277 (N_17277,N_16515,N_16737);
nand U17278 (N_17278,N_16801,N_16465);
nor U17279 (N_17279,N_16540,N_16605);
nand U17280 (N_17280,N_16857,N_16747);
nand U17281 (N_17281,N_16411,N_16573);
or U17282 (N_17282,N_16825,N_16565);
or U17283 (N_17283,N_16771,N_16857);
nand U17284 (N_17284,N_16646,N_16288);
or U17285 (N_17285,N_16453,N_16333);
or U17286 (N_17286,N_16385,N_16669);
xnor U17287 (N_17287,N_16639,N_16376);
and U17288 (N_17288,N_16629,N_16421);
xor U17289 (N_17289,N_16324,N_16733);
or U17290 (N_17290,N_16416,N_16667);
and U17291 (N_17291,N_16679,N_16723);
and U17292 (N_17292,N_16447,N_16384);
or U17293 (N_17293,N_16430,N_16274);
and U17294 (N_17294,N_16540,N_16503);
nor U17295 (N_17295,N_16589,N_16640);
or U17296 (N_17296,N_16570,N_16445);
and U17297 (N_17297,N_16497,N_16487);
xor U17298 (N_17298,N_16797,N_16345);
and U17299 (N_17299,N_16779,N_16748);
and U17300 (N_17300,N_16740,N_16486);
nand U17301 (N_17301,N_16739,N_16255);
xnor U17302 (N_17302,N_16559,N_16637);
xor U17303 (N_17303,N_16839,N_16645);
and U17304 (N_17304,N_16300,N_16785);
xor U17305 (N_17305,N_16381,N_16774);
or U17306 (N_17306,N_16264,N_16428);
and U17307 (N_17307,N_16831,N_16839);
xor U17308 (N_17308,N_16728,N_16692);
nor U17309 (N_17309,N_16402,N_16511);
and U17310 (N_17310,N_16644,N_16410);
or U17311 (N_17311,N_16836,N_16867);
xnor U17312 (N_17312,N_16478,N_16561);
or U17313 (N_17313,N_16577,N_16633);
or U17314 (N_17314,N_16850,N_16265);
and U17315 (N_17315,N_16817,N_16379);
nor U17316 (N_17316,N_16500,N_16559);
or U17317 (N_17317,N_16364,N_16712);
nor U17318 (N_17318,N_16326,N_16817);
or U17319 (N_17319,N_16503,N_16814);
or U17320 (N_17320,N_16655,N_16450);
nand U17321 (N_17321,N_16422,N_16469);
or U17322 (N_17322,N_16536,N_16259);
and U17323 (N_17323,N_16515,N_16779);
xnor U17324 (N_17324,N_16576,N_16706);
xor U17325 (N_17325,N_16659,N_16469);
xnor U17326 (N_17326,N_16864,N_16368);
xor U17327 (N_17327,N_16801,N_16530);
or U17328 (N_17328,N_16523,N_16287);
nor U17329 (N_17329,N_16787,N_16584);
nor U17330 (N_17330,N_16509,N_16530);
nor U17331 (N_17331,N_16736,N_16783);
and U17332 (N_17332,N_16459,N_16766);
nor U17333 (N_17333,N_16328,N_16804);
and U17334 (N_17334,N_16734,N_16570);
and U17335 (N_17335,N_16826,N_16557);
nand U17336 (N_17336,N_16456,N_16559);
or U17337 (N_17337,N_16591,N_16377);
and U17338 (N_17338,N_16367,N_16612);
or U17339 (N_17339,N_16852,N_16662);
nor U17340 (N_17340,N_16456,N_16653);
xor U17341 (N_17341,N_16527,N_16263);
nand U17342 (N_17342,N_16588,N_16257);
or U17343 (N_17343,N_16476,N_16658);
and U17344 (N_17344,N_16851,N_16420);
and U17345 (N_17345,N_16834,N_16782);
xnor U17346 (N_17346,N_16533,N_16781);
nand U17347 (N_17347,N_16733,N_16404);
and U17348 (N_17348,N_16332,N_16386);
nor U17349 (N_17349,N_16844,N_16866);
nand U17350 (N_17350,N_16656,N_16649);
xnor U17351 (N_17351,N_16423,N_16542);
or U17352 (N_17352,N_16702,N_16641);
or U17353 (N_17353,N_16256,N_16663);
nand U17354 (N_17354,N_16772,N_16310);
and U17355 (N_17355,N_16640,N_16330);
or U17356 (N_17356,N_16383,N_16347);
nand U17357 (N_17357,N_16795,N_16428);
xor U17358 (N_17358,N_16726,N_16706);
or U17359 (N_17359,N_16863,N_16398);
or U17360 (N_17360,N_16431,N_16587);
nand U17361 (N_17361,N_16566,N_16451);
xor U17362 (N_17362,N_16285,N_16724);
and U17363 (N_17363,N_16745,N_16809);
and U17364 (N_17364,N_16327,N_16407);
or U17365 (N_17365,N_16626,N_16545);
nor U17366 (N_17366,N_16380,N_16607);
nand U17367 (N_17367,N_16266,N_16458);
xnor U17368 (N_17368,N_16394,N_16792);
and U17369 (N_17369,N_16856,N_16314);
xor U17370 (N_17370,N_16811,N_16682);
or U17371 (N_17371,N_16493,N_16568);
nand U17372 (N_17372,N_16764,N_16474);
and U17373 (N_17373,N_16594,N_16498);
and U17374 (N_17374,N_16696,N_16431);
nand U17375 (N_17375,N_16661,N_16409);
and U17376 (N_17376,N_16607,N_16268);
xor U17377 (N_17377,N_16628,N_16321);
nor U17378 (N_17378,N_16393,N_16485);
and U17379 (N_17379,N_16801,N_16719);
or U17380 (N_17380,N_16472,N_16432);
or U17381 (N_17381,N_16773,N_16811);
nor U17382 (N_17382,N_16260,N_16769);
or U17383 (N_17383,N_16315,N_16709);
nand U17384 (N_17384,N_16362,N_16712);
nor U17385 (N_17385,N_16800,N_16722);
nand U17386 (N_17386,N_16262,N_16459);
xor U17387 (N_17387,N_16713,N_16824);
xor U17388 (N_17388,N_16310,N_16695);
nor U17389 (N_17389,N_16653,N_16406);
nand U17390 (N_17390,N_16706,N_16377);
nor U17391 (N_17391,N_16616,N_16361);
or U17392 (N_17392,N_16286,N_16707);
xnor U17393 (N_17393,N_16864,N_16586);
xor U17394 (N_17394,N_16780,N_16607);
and U17395 (N_17395,N_16866,N_16736);
xor U17396 (N_17396,N_16671,N_16661);
nand U17397 (N_17397,N_16279,N_16303);
and U17398 (N_17398,N_16261,N_16372);
nand U17399 (N_17399,N_16668,N_16460);
or U17400 (N_17400,N_16372,N_16358);
or U17401 (N_17401,N_16712,N_16448);
xor U17402 (N_17402,N_16338,N_16443);
or U17403 (N_17403,N_16708,N_16824);
or U17404 (N_17404,N_16741,N_16521);
nor U17405 (N_17405,N_16513,N_16631);
nand U17406 (N_17406,N_16641,N_16650);
nor U17407 (N_17407,N_16682,N_16638);
nor U17408 (N_17408,N_16376,N_16360);
nor U17409 (N_17409,N_16436,N_16671);
or U17410 (N_17410,N_16837,N_16665);
nand U17411 (N_17411,N_16301,N_16410);
xor U17412 (N_17412,N_16637,N_16688);
or U17413 (N_17413,N_16382,N_16632);
and U17414 (N_17414,N_16431,N_16739);
nor U17415 (N_17415,N_16645,N_16779);
and U17416 (N_17416,N_16836,N_16796);
and U17417 (N_17417,N_16803,N_16425);
nor U17418 (N_17418,N_16728,N_16808);
xnor U17419 (N_17419,N_16392,N_16327);
nor U17420 (N_17420,N_16469,N_16740);
nand U17421 (N_17421,N_16605,N_16695);
and U17422 (N_17422,N_16727,N_16339);
xor U17423 (N_17423,N_16543,N_16707);
or U17424 (N_17424,N_16728,N_16442);
nand U17425 (N_17425,N_16813,N_16283);
nand U17426 (N_17426,N_16652,N_16426);
nand U17427 (N_17427,N_16641,N_16664);
nor U17428 (N_17428,N_16476,N_16288);
nand U17429 (N_17429,N_16400,N_16497);
and U17430 (N_17430,N_16754,N_16337);
and U17431 (N_17431,N_16273,N_16556);
nand U17432 (N_17432,N_16439,N_16677);
or U17433 (N_17433,N_16743,N_16523);
and U17434 (N_17434,N_16733,N_16375);
xor U17435 (N_17435,N_16462,N_16627);
nand U17436 (N_17436,N_16327,N_16705);
nor U17437 (N_17437,N_16870,N_16276);
and U17438 (N_17438,N_16514,N_16679);
or U17439 (N_17439,N_16457,N_16450);
nor U17440 (N_17440,N_16806,N_16549);
or U17441 (N_17441,N_16490,N_16549);
or U17442 (N_17442,N_16734,N_16257);
nor U17443 (N_17443,N_16287,N_16863);
nor U17444 (N_17444,N_16288,N_16375);
and U17445 (N_17445,N_16625,N_16556);
and U17446 (N_17446,N_16518,N_16613);
xor U17447 (N_17447,N_16556,N_16575);
nand U17448 (N_17448,N_16490,N_16415);
or U17449 (N_17449,N_16543,N_16784);
and U17450 (N_17450,N_16861,N_16563);
nor U17451 (N_17451,N_16297,N_16475);
xor U17452 (N_17452,N_16376,N_16594);
and U17453 (N_17453,N_16444,N_16288);
xor U17454 (N_17454,N_16448,N_16689);
nor U17455 (N_17455,N_16605,N_16684);
nor U17456 (N_17456,N_16413,N_16359);
and U17457 (N_17457,N_16761,N_16691);
nand U17458 (N_17458,N_16616,N_16413);
or U17459 (N_17459,N_16852,N_16447);
nand U17460 (N_17460,N_16586,N_16486);
nor U17461 (N_17461,N_16696,N_16508);
nor U17462 (N_17462,N_16613,N_16331);
nor U17463 (N_17463,N_16629,N_16708);
nor U17464 (N_17464,N_16806,N_16667);
or U17465 (N_17465,N_16323,N_16677);
nand U17466 (N_17466,N_16773,N_16638);
and U17467 (N_17467,N_16511,N_16520);
xnor U17468 (N_17468,N_16843,N_16688);
xnor U17469 (N_17469,N_16466,N_16432);
nand U17470 (N_17470,N_16347,N_16734);
xor U17471 (N_17471,N_16870,N_16261);
or U17472 (N_17472,N_16413,N_16523);
and U17473 (N_17473,N_16741,N_16811);
nand U17474 (N_17474,N_16600,N_16503);
xor U17475 (N_17475,N_16493,N_16627);
and U17476 (N_17476,N_16361,N_16794);
nor U17477 (N_17477,N_16428,N_16788);
nor U17478 (N_17478,N_16412,N_16627);
and U17479 (N_17479,N_16303,N_16287);
nor U17480 (N_17480,N_16364,N_16416);
nor U17481 (N_17481,N_16680,N_16604);
and U17482 (N_17482,N_16490,N_16576);
nand U17483 (N_17483,N_16811,N_16406);
xor U17484 (N_17484,N_16315,N_16769);
or U17485 (N_17485,N_16850,N_16530);
and U17486 (N_17486,N_16626,N_16558);
xnor U17487 (N_17487,N_16387,N_16580);
or U17488 (N_17488,N_16694,N_16402);
nor U17489 (N_17489,N_16529,N_16452);
xor U17490 (N_17490,N_16529,N_16739);
nand U17491 (N_17491,N_16614,N_16454);
nor U17492 (N_17492,N_16346,N_16820);
nor U17493 (N_17493,N_16578,N_16264);
xnor U17494 (N_17494,N_16664,N_16759);
or U17495 (N_17495,N_16537,N_16768);
nor U17496 (N_17496,N_16736,N_16773);
and U17497 (N_17497,N_16827,N_16330);
nor U17498 (N_17498,N_16546,N_16658);
and U17499 (N_17499,N_16449,N_16318);
nand U17500 (N_17500,N_17329,N_17430);
and U17501 (N_17501,N_17062,N_16946);
xor U17502 (N_17502,N_17120,N_16995);
or U17503 (N_17503,N_17354,N_17210);
and U17504 (N_17504,N_16997,N_17350);
nor U17505 (N_17505,N_17428,N_17466);
and U17506 (N_17506,N_16983,N_17098);
and U17507 (N_17507,N_17280,N_17105);
and U17508 (N_17508,N_17290,N_17419);
xor U17509 (N_17509,N_17009,N_17154);
and U17510 (N_17510,N_17401,N_17447);
nor U17511 (N_17511,N_17153,N_17285);
nor U17512 (N_17512,N_17383,N_16987);
or U17513 (N_17513,N_16936,N_17181);
or U17514 (N_17514,N_17315,N_17099);
xnor U17515 (N_17515,N_16977,N_17405);
nand U17516 (N_17516,N_17398,N_17452);
or U17517 (N_17517,N_17194,N_17433);
and U17518 (N_17518,N_17249,N_17030);
nor U17519 (N_17519,N_17361,N_17253);
or U17520 (N_17520,N_16999,N_17384);
and U17521 (N_17521,N_17027,N_17381);
xor U17522 (N_17522,N_16990,N_17054);
xnor U17523 (N_17523,N_17060,N_17128);
or U17524 (N_17524,N_17295,N_17113);
nand U17525 (N_17525,N_17330,N_16961);
nor U17526 (N_17526,N_17310,N_16988);
nor U17527 (N_17527,N_17243,N_17038);
and U17528 (N_17528,N_17326,N_17208);
and U17529 (N_17529,N_17161,N_17051);
nand U17530 (N_17530,N_17132,N_17474);
and U17531 (N_17531,N_16996,N_16918);
nor U17532 (N_17532,N_17166,N_17495);
or U17533 (N_17533,N_17008,N_17072);
or U17534 (N_17534,N_17061,N_17052);
nand U17535 (N_17535,N_16901,N_16939);
nor U17536 (N_17536,N_17411,N_17050);
xnor U17537 (N_17537,N_16962,N_17019);
nor U17538 (N_17538,N_17198,N_17087);
or U17539 (N_17539,N_16891,N_17313);
and U17540 (N_17540,N_17215,N_16966);
and U17541 (N_17541,N_17133,N_17497);
nor U17542 (N_17542,N_17164,N_17115);
or U17543 (N_17543,N_17229,N_17341);
nand U17544 (N_17544,N_17311,N_17325);
or U17545 (N_17545,N_17085,N_16951);
xor U17546 (N_17546,N_17231,N_17424);
or U17547 (N_17547,N_17021,N_16913);
nor U17548 (N_17548,N_17273,N_16947);
nor U17549 (N_17549,N_17162,N_17138);
xor U17550 (N_17550,N_17455,N_16973);
xor U17551 (N_17551,N_17141,N_16949);
or U17552 (N_17552,N_16896,N_17260);
nor U17553 (N_17553,N_17366,N_17192);
nor U17554 (N_17554,N_17404,N_17074);
nor U17555 (N_17555,N_17055,N_16910);
and U17556 (N_17556,N_17331,N_16985);
nand U17557 (N_17557,N_17291,N_17429);
nand U17558 (N_17558,N_17396,N_17139);
and U17559 (N_17559,N_17413,N_17368);
and U17560 (N_17560,N_17477,N_17137);
xor U17561 (N_17561,N_17416,N_17304);
xor U17562 (N_17562,N_16964,N_17190);
nor U17563 (N_17563,N_17233,N_16920);
nor U17564 (N_17564,N_17016,N_17111);
and U17565 (N_17565,N_17343,N_17459);
and U17566 (N_17566,N_17183,N_17207);
xor U17567 (N_17567,N_16978,N_17252);
or U17568 (N_17568,N_17044,N_17205);
nand U17569 (N_17569,N_17298,N_17148);
nand U17570 (N_17570,N_17490,N_16878);
nor U17571 (N_17571,N_17212,N_17004);
xor U17572 (N_17572,N_17439,N_17178);
nand U17573 (N_17573,N_17235,N_16928);
or U17574 (N_17574,N_17118,N_17450);
and U17575 (N_17575,N_17492,N_17349);
and U17576 (N_17576,N_17493,N_17213);
nor U17577 (N_17577,N_17143,N_16994);
or U17578 (N_17578,N_17374,N_17244);
or U17579 (N_17579,N_16909,N_17180);
nand U17580 (N_17580,N_17024,N_17306);
or U17581 (N_17581,N_17068,N_16963);
nor U17582 (N_17582,N_16885,N_17499);
and U17583 (N_17583,N_17032,N_16927);
and U17584 (N_17584,N_16991,N_16895);
nand U17585 (N_17585,N_16965,N_17234);
xor U17586 (N_17586,N_17156,N_16915);
nor U17587 (N_17587,N_17059,N_17241);
or U17588 (N_17588,N_17250,N_17432);
or U17589 (N_17589,N_17408,N_17042);
or U17590 (N_17590,N_17079,N_17461);
and U17591 (N_17591,N_16886,N_17367);
and U17592 (N_17592,N_16917,N_17245);
nor U17593 (N_17593,N_17028,N_17070);
nand U17594 (N_17594,N_17491,N_16960);
xnor U17595 (N_17595,N_17026,N_16898);
nor U17596 (N_17596,N_16968,N_17391);
xnor U17597 (N_17597,N_17223,N_17332);
or U17598 (N_17598,N_17093,N_17457);
and U17599 (N_17599,N_16981,N_17443);
or U17600 (N_17600,N_17365,N_17409);
and U17601 (N_17601,N_17160,N_17063);
and U17602 (N_17602,N_17182,N_17057);
nor U17603 (N_17603,N_16922,N_17053);
nor U17604 (N_17604,N_17399,N_17193);
or U17605 (N_17605,N_17380,N_17216);
nor U17606 (N_17606,N_17155,N_17000);
nor U17607 (N_17607,N_17171,N_16926);
nand U17608 (N_17608,N_17127,N_16902);
and U17609 (N_17609,N_17270,N_17043);
nand U17610 (N_17610,N_17344,N_17251);
nor U17611 (N_17611,N_16941,N_17096);
or U17612 (N_17612,N_17114,N_17097);
nand U17613 (N_17613,N_17257,N_16986);
nand U17614 (N_17614,N_17297,N_17091);
and U17615 (N_17615,N_17206,N_17395);
nor U17616 (N_17616,N_17420,N_17084);
and U17617 (N_17617,N_17121,N_17112);
or U17618 (N_17618,N_16993,N_17486);
or U17619 (N_17619,N_17471,N_16907);
xor U17620 (N_17620,N_17488,N_17119);
or U17621 (N_17621,N_17364,N_17134);
and U17622 (N_17622,N_16942,N_17440);
nand U17623 (N_17623,N_17056,N_16933);
or U17624 (N_17624,N_17266,N_16921);
xor U17625 (N_17625,N_17415,N_17240);
and U17626 (N_17626,N_17149,N_17264);
nand U17627 (N_17627,N_17382,N_17279);
and U17628 (N_17628,N_17302,N_17372);
and U17629 (N_17629,N_16998,N_16894);
xnor U17630 (N_17630,N_17351,N_17412);
and U17631 (N_17631,N_17135,N_17454);
and U17632 (N_17632,N_17140,N_17323);
or U17633 (N_17633,N_17246,N_16897);
and U17634 (N_17634,N_16903,N_17029);
xnor U17635 (N_17635,N_17169,N_17468);
nand U17636 (N_17636,N_17108,N_17189);
nand U17637 (N_17637,N_17371,N_17464);
and U17638 (N_17638,N_16950,N_17126);
xnor U17639 (N_17639,N_17336,N_16953);
or U17640 (N_17640,N_17438,N_17358);
nand U17641 (N_17641,N_17202,N_17214);
or U17642 (N_17642,N_17001,N_17066);
and U17643 (N_17643,N_17048,N_17259);
nor U17644 (N_17644,N_17089,N_17011);
and U17645 (N_17645,N_16883,N_17427);
xnor U17646 (N_17646,N_17006,N_17345);
xnor U17647 (N_17647,N_17479,N_17248);
nand U17648 (N_17648,N_17073,N_17204);
xor U17649 (N_17649,N_17142,N_17263);
xor U17650 (N_17650,N_17159,N_16930);
nand U17651 (N_17651,N_17301,N_16948);
nor U17652 (N_17652,N_17230,N_17335);
or U17653 (N_17653,N_16935,N_17258);
and U17654 (N_17654,N_17226,N_17356);
xnor U17655 (N_17655,N_17237,N_17375);
and U17656 (N_17656,N_17065,N_17017);
or U17657 (N_17657,N_16982,N_17224);
nor U17658 (N_17658,N_16893,N_17437);
or U17659 (N_17659,N_17386,N_17035);
nor U17660 (N_17660,N_17308,N_16980);
and U17661 (N_17661,N_17232,N_17076);
or U17662 (N_17662,N_17448,N_17463);
nor U17663 (N_17663,N_17123,N_17077);
nand U17664 (N_17664,N_16944,N_17136);
or U17665 (N_17665,N_16945,N_17034);
nand U17666 (N_17666,N_17129,N_17125);
and U17667 (N_17667,N_17092,N_17388);
nand U17668 (N_17668,N_17163,N_17378);
nor U17669 (N_17669,N_17015,N_16971);
nand U17670 (N_17670,N_17067,N_17431);
or U17671 (N_17671,N_17151,N_16975);
xnor U17672 (N_17672,N_17261,N_16887);
and U17673 (N_17673,N_17238,N_17324);
nand U17674 (N_17674,N_17348,N_17445);
nand U17675 (N_17675,N_17045,N_17353);
nor U17676 (N_17676,N_17394,N_17100);
or U17677 (N_17677,N_17275,N_16970);
and U17678 (N_17678,N_17172,N_17106);
nor U17679 (N_17679,N_17018,N_17094);
nand U17680 (N_17680,N_17292,N_17037);
nand U17681 (N_17681,N_17470,N_17462);
xnor U17682 (N_17682,N_17426,N_17397);
nand U17683 (N_17683,N_17318,N_17347);
and U17684 (N_17684,N_17482,N_17489);
nor U17685 (N_17685,N_16929,N_17316);
xnor U17686 (N_17686,N_17338,N_17392);
or U17687 (N_17687,N_16958,N_16955);
xor U17688 (N_17688,N_17451,N_17086);
and U17689 (N_17689,N_17219,N_17170);
nand U17690 (N_17690,N_16931,N_17305);
nor U17691 (N_17691,N_17370,N_16923);
or U17692 (N_17692,N_16905,N_17255);
xor U17693 (N_17693,N_17047,N_17480);
or U17694 (N_17694,N_16984,N_16969);
nand U17695 (N_17695,N_17406,N_17188);
and U17696 (N_17696,N_17071,N_17269);
or U17697 (N_17697,N_17373,N_17124);
nand U17698 (N_17698,N_16943,N_17435);
and U17699 (N_17699,N_17236,N_17217);
nor U17700 (N_17700,N_17058,N_16900);
and U17701 (N_17701,N_16919,N_17458);
and U17702 (N_17702,N_17483,N_17012);
or U17703 (N_17703,N_17369,N_16875);
or U17704 (N_17704,N_17078,N_17165);
and U17705 (N_17705,N_16937,N_17359);
and U17706 (N_17706,N_17307,N_17337);
nand U17707 (N_17707,N_17107,N_17173);
or U17708 (N_17708,N_17002,N_17110);
xor U17709 (N_17709,N_17444,N_17101);
and U17710 (N_17710,N_17147,N_17104);
nand U17711 (N_17711,N_17039,N_17352);
nand U17712 (N_17712,N_16892,N_16932);
and U17713 (N_17713,N_17225,N_17080);
and U17714 (N_17714,N_17247,N_17402);
nand U17715 (N_17715,N_16911,N_17303);
nor U17716 (N_17716,N_17276,N_17081);
xor U17717 (N_17717,N_16976,N_17033);
or U17718 (N_17718,N_16952,N_16974);
nand U17719 (N_17719,N_17103,N_17300);
or U17720 (N_17720,N_16957,N_17288);
xnor U17721 (N_17721,N_17465,N_17453);
xnor U17722 (N_17722,N_17176,N_17342);
xor U17723 (N_17723,N_16992,N_17442);
nand U17724 (N_17724,N_17377,N_17167);
nand U17725 (N_17725,N_17496,N_17265);
and U17726 (N_17726,N_17007,N_16972);
or U17727 (N_17727,N_17175,N_17179);
or U17728 (N_17728,N_17157,N_17242);
nor U17729 (N_17729,N_17456,N_17469);
and U17730 (N_17730,N_17075,N_16882);
nand U17731 (N_17731,N_17201,N_17283);
or U17732 (N_17732,N_17403,N_17421);
xnor U17733 (N_17733,N_17168,N_16899);
and U17734 (N_17734,N_17362,N_17389);
xnor U17735 (N_17735,N_17145,N_17195);
nand U17736 (N_17736,N_17436,N_17363);
xor U17737 (N_17737,N_17387,N_17284);
or U17738 (N_17738,N_17239,N_17003);
and U17739 (N_17739,N_17289,N_17320);
nor U17740 (N_17740,N_17268,N_17196);
nand U17741 (N_17741,N_17340,N_17487);
nor U17742 (N_17742,N_17475,N_16888);
nand U17743 (N_17743,N_17434,N_17197);
xor U17744 (N_17744,N_17186,N_17174);
nand U17745 (N_17745,N_17339,N_17473);
or U17746 (N_17746,N_17481,N_16924);
and U17747 (N_17747,N_17199,N_16914);
nor U17748 (N_17748,N_17187,N_17267);
or U17749 (N_17749,N_17425,N_17262);
or U17750 (N_17750,N_17256,N_16889);
or U17751 (N_17751,N_17334,N_17322);
nor U17752 (N_17752,N_16890,N_17327);
or U17753 (N_17753,N_17446,N_16880);
or U17754 (N_17754,N_17150,N_17376);
and U17755 (N_17755,N_17346,N_17109);
xor U17756 (N_17756,N_17158,N_16906);
and U17757 (N_17757,N_17146,N_17271);
and U17758 (N_17758,N_17130,N_17319);
and U17759 (N_17759,N_16876,N_17294);
nand U17760 (N_17760,N_17069,N_17200);
nand U17761 (N_17761,N_17272,N_17041);
nor U17762 (N_17762,N_17254,N_17441);
and U17763 (N_17763,N_16956,N_17116);
or U17764 (N_17764,N_17220,N_17218);
xnor U17765 (N_17765,N_17277,N_16940);
nor U17766 (N_17766,N_17418,N_17184);
nand U17767 (N_17767,N_16916,N_17005);
or U17768 (N_17768,N_17131,N_17122);
nor U17769 (N_17769,N_16954,N_17144);
nor U17770 (N_17770,N_17379,N_17314);
xnor U17771 (N_17771,N_17023,N_17417);
nand U17772 (N_17772,N_16879,N_16925);
nor U17773 (N_17773,N_17296,N_17274);
nor U17774 (N_17774,N_17309,N_16881);
or U17775 (N_17775,N_17191,N_17117);
and U17776 (N_17776,N_17476,N_17203);
nor U17777 (N_17777,N_17020,N_17278);
or U17778 (N_17778,N_17393,N_17049);
and U17779 (N_17779,N_17478,N_17357);
nand U17780 (N_17780,N_17422,N_17013);
xor U17781 (N_17781,N_17385,N_17328);
and U17782 (N_17782,N_17498,N_17222);
xor U17783 (N_17783,N_17390,N_17209);
and U17784 (N_17784,N_17449,N_17494);
xor U17785 (N_17785,N_17227,N_17321);
and U17786 (N_17786,N_17281,N_17014);
and U17787 (N_17787,N_17090,N_17102);
nor U17788 (N_17788,N_16912,N_17025);
or U17789 (N_17789,N_17360,N_17317);
nand U17790 (N_17790,N_17484,N_16908);
nor U17791 (N_17791,N_17282,N_17083);
or U17792 (N_17792,N_17221,N_17082);
nor U17793 (N_17793,N_17355,N_16934);
or U17794 (N_17794,N_16967,N_17031);
nor U17795 (N_17795,N_16884,N_17036);
xnor U17796 (N_17796,N_17010,N_17333);
nor U17797 (N_17797,N_17022,N_17046);
and U17798 (N_17798,N_17040,N_17287);
or U17799 (N_17799,N_17177,N_17472);
nand U17800 (N_17800,N_17095,N_17460);
nor U17801 (N_17801,N_16959,N_16904);
nor U17802 (N_17802,N_16877,N_17407);
nor U17803 (N_17803,N_17400,N_16979);
or U17804 (N_17804,N_17312,N_16938);
or U17805 (N_17805,N_17423,N_16989);
nand U17806 (N_17806,N_17410,N_17152);
nor U17807 (N_17807,N_17299,N_17414);
and U17808 (N_17808,N_17064,N_17211);
nor U17809 (N_17809,N_17088,N_17185);
and U17810 (N_17810,N_17293,N_17485);
nand U17811 (N_17811,N_17467,N_17286);
and U17812 (N_17812,N_17228,N_17248);
nand U17813 (N_17813,N_17197,N_17361);
or U17814 (N_17814,N_17267,N_16999);
and U17815 (N_17815,N_17269,N_17458);
and U17816 (N_17816,N_17398,N_16950);
xor U17817 (N_17817,N_17471,N_17413);
or U17818 (N_17818,N_17254,N_17171);
nor U17819 (N_17819,N_16899,N_17479);
nand U17820 (N_17820,N_17307,N_17181);
nor U17821 (N_17821,N_17210,N_16985);
xnor U17822 (N_17822,N_16877,N_17077);
xnor U17823 (N_17823,N_17279,N_17019);
nand U17824 (N_17824,N_17294,N_17495);
xor U17825 (N_17825,N_17187,N_17236);
or U17826 (N_17826,N_16997,N_17481);
nand U17827 (N_17827,N_17166,N_17228);
and U17828 (N_17828,N_17382,N_17176);
xor U17829 (N_17829,N_16969,N_17003);
nand U17830 (N_17830,N_17046,N_17157);
and U17831 (N_17831,N_17415,N_17148);
or U17832 (N_17832,N_16894,N_17282);
nand U17833 (N_17833,N_16968,N_17479);
nand U17834 (N_17834,N_17149,N_17157);
and U17835 (N_17835,N_17070,N_17015);
or U17836 (N_17836,N_17184,N_16915);
and U17837 (N_17837,N_17101,N_17035);
or U17838 (N_17838,N_17246,N_17028);
nor U17839 (N_17839,N_17366,N_16939);
and U17840 (N_17840,N_16923,N_17115);
or U17841 (N_17841,N_16914,N_16919);
nor U17842 (N_17842,N_17408,N_16976);
nor U17843 (N_17843,N_17226,N_17390);
nand U17844 (N_17844,N_17051,N_17469);
nor U17845 (N_17845,N_17452,N_17034);
and U17846 (N_17846,N_17197,N_17415);
or U17847 (N_17847,N_17139,N_17398);
nand U17848 (N_17848,N_17365,N_17464);
or U17849 (N_17849,N_16909,N_17028);
or U17850 (N_17850,N_16993,N_17110);
nand U17851 (N_17851,N_17165,N_16934);
and U17852 (N_17852,N_16904,N_17111);
or U17853 (N_17853,N_16927,N_17441);
nor U17854 (N_17854,N_17136,N_17049);
or U17855 (N_17855,N_16965,N_16975);
xor U17856 (N_17856,N_17048,N_17415);
xor U17857 (N_17857,N_17470,N_17254);
or U17858 (N_17858,N_17440,N_17491);
and U17859 (N_17859,N_17338,N_16936);
or U17860 (N_17860,N_17498,N_17143);
and U17861 (N_17861,N_17460,N_16876);
xnor U17862 (N_17862,N_16892,N_17181);
or U17863 (N_17863,N_17115,N_16998);
nor U17864 (N_17864,N_17219,N_17360);
xor U17865 (N_17865,N_17062,N_17449);
and U17866 (N_17866,N_17268,N_16985);
nor U17867 (N_17867,N_16953,N_17285);
nor U17868 (N_17868,N_17138,N_17475);
nand U17869 (N_17869,N_16927,N_17112);
nor U17870 (N_17870,N_17325,N_17380);
or U17871 (N_17871,N_17447,N_16965);
xor U17872 (N_17872,N_17312,N_17150);
and U17873 (N_17873,N_17418,N_16914);
or U17874 (N_17874,N_17462,N_16955);
or U17875 (N_17875,N_16922,N_17102);
xnor U17876 (N_17876,N_17367,N_16929);
nor U17877 (N_17877,N_17070,N_17002);
and U17878 (N_17878,N_17443,N_17468);
nor U17879 (N_17879,N_17335,N_17159);
nand U17880 (N_17880,N_17021,N_16908);
xnor U17881 (N_17881,N_17286,N_17051);
and U17882 (N_17882,N_17245,N_17182);
or U17883 (N_17883,N_16979,N_17215);
nand U17884 (N_17884,N_17263,N_16935);
or U17885 (N_17885,N_17118,N_17369);
or U17886 (N_17886,N_17449,N_17044);
and U17887 (N_17887,N_17004,N_17277);
nand U17888 (N_17888,N_17130,N_17460);
nand U17889 (N_17889,N_17040,N_17247);
xor U17890 (N_17890,N_17121,N_17288);
and U17891 (N_17891,N_17377,N_17072);
and U17892 (N_17892,N_17217,N_17487);
or U17893 (N_17893,N_17223,N_17098);
nor U17894 (N_17894,N_17215,N_17206);
nor U17895 (N_17895,N_17158,N_17075);
and U17896 (N_17896,N_17390,N_16996);
and U17897 (N_17897,N_17002,N_16924);
nor U17898 (N_17898,N_17234,N_17308);
xor U17899 (N_17899,N_17301,N_17448);
xor U17900 (N_17900,N_17112,N_17068);
and U17901 (N_17901,N_17099,N_16984);
or U17902 (N_17902,N_17118,N_17373);
nor U17903 (N_17903,N_17191,N_17174);
nor U17904 (N_17904,N_16886,N_17037);
and U17905 (N_17905,N_16931,N_17417);
nor U17906 (N_17906,N_17032,N_17083);
xnor U17907 (N_17907,N_17122,N_17042);
and U17908 (N_17908,N_16944,N_16908);
nand U17909 (N_17909,N_17135,N_17097);
or U17910 (N_17910,N_17244,N_17096);
and U17911 (N_17911,N_16930,N_16924);
xor U17912 (N_17912,N_17022,N_16996);
nand U17913 (N_17913,N_17265,N_17445);
and U17914 (N_17914,N_16893,N_17067);
nand U17915 (N_17915,N_17099,N_17103);
nand U17916 (N_17916,N_17496,N_16982);
or U17917 (N_17917,N_17000,N_17172);
or U17918 (N_17918,N_17235,N_17259);
xor U17919 (N_17919,N_17012,N_17248);
nand U17920 (N_17920,N_17097,N_17492);
and U17921 (N_17921,N_17162,N_17196);
xnor U17922 (N_17922,N_16914,N_17133);
or U17923 (N_17923,N_17232,N_17455);
xor U17924 (N_17924,N_17098,N_17072);
nand U17925 (N_17925,N_17213,N_17052);
nand U17926 (N_17926,N_17079,N_17470);
nand U17927 (N_17927,N_17333,N_16927);
nor U17928 (N_17928,N_17215,N_17395);
or U17929 (N_17929,N_17121,N_17065);
nor U17930 (N_17930,N_16984,N_17197);
xor U17931 (N_17931,N_16897,N_17457);
or U17932 (N_17932,N_16969,N_17129);
nand U17933 (N_17933,N_17356,N_17051);
or U17934 (N_17934,N_17031,N_17057);
or U17935 (N_17935,N_17003,N_16963);
and U17936 (N_17936,N_17021,N_17314);
or U17937 (N_17937,N_16877,N_17425);
and U17938 (N_17938,N_17021,N_17178);
and U17939 (N_17939,N_17318,N_17009);
nor U17940 (N_17940,N_17347,N_17300);
nand U17941 (N_17941,N_17021,N_17295);
and U17942 (N_17942,N_17007,N_16882);
xor U17943 (N_17943,N_16929,N_17485);
nor U17944 (N_17944,N_17374,N_17345);
nand U17945 (N_17945,N_16881,N_16957);
xnor U17946 (N_17946,N_17110,N_17432);
or U17947 (N_17947,N_17339,N_17286);
and U17948 (N_17948,N_16998,N_17179);
nor U17949 (N_17949,N_17272,N_17309);
xor U17950 (N_17950,N_17075,N_17055);
nand U17951 (N_17951,N_17293,N_16923);
nor U17952 (N_17952,N_17129,N_17040);
and U17953 (N_17953,N_16887,N_17462);
xor U17954 (N_17954,N_17198,N_17463);
nor U17955 (N_17955,N_17485,N_17192);
nand U17956 (N_17956,N_16909,N_17476);
nor U17957 (N_17957,N_17168,N_17359);
nor U17958 (N_17958,N_17352,N_17446);
nand U17959 (N_17959,N_16893,N_17011);
and U17960 (N_17960,N_16945,N_16974);
xor U17961 (N_17961,N_17382,N_17302);
xor U17962 (N_17962,N_17471,N_16891);
xnor U17963 (N_17963,N_17252,N_17128);
xor U17964 (N_17964,N_17342,N_17028);
nand U17965 (N_17965,N_17190,N_17084);
and U17966 (N_17966,N_17393,N_17004);
or U17967 (N_17967,N_17004,N_17318);
and U17968 (N_17968,N_17420,N_16936);
nand U17969 (N_17969,N_17319,N_17041);
nand U17970 (N_17970,N_16894,N_17115);
or U17971 (N_17971,N_17361,N_17230);
or U17972 (N_17972,N_17190,N_17110);
nor U17973 (N_17973,N_17263,N_16934);
nand U17974 (N_17974,N_17273,N_17354);
xor U17975 (N_17975,N_17444,N_16939);
nand U17976 (N_17976,N_17107,N_17499);
or U17977 (N_17977,N_17370,N_16979);
or U17978 (N_17978,N_17140,N_17303);
nor U17979 (N_17979,N_17202,N_17301);
xor U17980 (N_17980,N_16928,N_17138);
nor U17981 (N_17981,N_16975,N_17181);
xor U17982 (N_17982,N_16892,N_17492);
nor U17983 (N_17983,N_17442,N_17017);
and U17984 (N_17984,N_17482,N_17331);
or U17985 (N_17985,N_16929,N_17416);
or U17986 (N_17986,N_17452,N_17092);
or U17987 (N_17987,N_17147,N_17058);
or U17988 (N_17988,N_17202,N_17423);
and U17989 (N_17989,N_16921,N_17334);
xor U17990 (N_17990,N_17392,N_17006);
nand U17991 (N_17991,N_17135,N_16947);
xnor U17992 (N_17992,N_17044,N_17057);
nand U17993 (N_17993,N_17024,N_16990);
nor U17994 (N_17994,N_17108,N_17364);
nor U17995 (N_17995,N_17409,N_17435);
and U17996 (N_17996,N_16971,N_17439);
or U17997 (N_17997,N_17402,N_17477);
and U17998 (N_17998,N_17129,N_17215);
and U17999 (N_17999,N_16975,N_17012);
or U18000 (N_18000,N_16932,N_17018);
nand U18001 (N_18001,N_17020,N_17333);
nor U18002 (N_18002,N_17121,N_16905);
and U18003 (N_18003,N_17072,N_16966);
nand U18004 (N_18004,N_16951,N_17260);
and U18005 (N_18005,N_17193,N_17026);
xor U18006 (N_18006,N_17115,N_17407);
nor U18007 (N_18007,N_17175,N_17440);
and U18008 (N_18008,N_17282,N_16980);
nor U18009 (N_18009,N_17122,N_17154);
or U18010 (N_18010,N_17375,N_17155);
nor U18011 (N_18011,N_16913,N_16998);
xor U18012 (N_18012,N_16976,N_17342);
nor U18013 (N_18013,N_16940,N_17160);
nor U18014 (N_18014,N_16962,N_16987);
or U18015 (N_18015,N_17278,N_17251);
xnor U18016 (N_18016,N_17332,N_16922);
xnor U18017 (N_18017,N_17162,N_17298);
nand U18018 (N_18018,N_17089,N_17095);
or U18019 (N_18019,N_16972,N_16890);
and U18020 (N_18020,N_17328,N_17227);
nor U18021 (N_18021,N_17376,N_16923);
or U18022 (N_18022,N_17280,N_17224);
nand U18023 (N_18023,N_17347,N_17327);
nand U18024 (N_18024,N_17279,N_17479);
or U18025 (N_18025,N_16912,N_17064);
xnor U18026 (N_18026,N_17058,N_16939);
or U18027 (N_18027,N_17062,N_17103);
or U18028 (N_18028,N_17498,N_16921);
xor U18029 (N_18029,N_17402,N_16968);
nand U18030 (N_18030,N_16889,N_17061);
and U18031 (N_18031,N_17322,N_17364);
nand U18032 (N_18032,N_16977,N_17424);
xor U18033 (N_18033,N_16935,N_17060);
xnor U18034 (N_18034,N_16943,N_17499);
and U18035 (N_18035,N_17058,N_17421);
nand U18036 (N_18036,N_16887,N_17328);
nor U18037 (N_18037,N_17303,N_17353);
nor U18038 (N_18038,N_17484,N_17393);
or U18039 (N_18039,N_17203,N_17038);
xnor U18040 (N_18040,N_17352,N_16976);
or U18041 (N_18041,N_17453,N_17183);
and U18042 (N_18042,N_17431,N_17459);
nand U18043 (N_18043,N_17397,N_16924);
and U18044 (N_18044,N_16990,N_17262);
xor U18045 (N_18045,N_17236,N_17437);
or U18046 (N_18046,N_17162,N_17153);
and U18047 (N_18047,N_17054,N_17033);
nor U18048 (N_18048,N_17392,N_17461);
and U18049 (N_18049,N_17402,N_17030);
nand U18050 (N_18050,N_17061,N_17156);
nand U18051 (N_18051,N_17261,N_17307);
and U18052 (N_18052,N_17439,N_16889);
nor U18053 (N_18053,N_17244,N_17116);
nand U18054 (N_18054,N_17075,N_17125);
and U18055 (N_18055,N_17080,N_17476);
xnor U18056 (N_18056,N_17051,N_17100);
xnor U18057 (N_18057,N_17433,N_17400);
xor U18058 (N_18058,N_17477,N_17105);
or U18059 (N_18059,N_17104,N_17372);
nand U18060 (N_18060,N_16929,N_17147);
or U18061 (N_18061,N_16932,N_17162);
xnor U18062 (N_18062,N_17335,N_17029);
and U18063 (N_18063,N_17497,N_17059);
xnor U18064 (N_18064,N_16941,N_16980);
nand U18065 (N_18065,N_17193,N_17413);
or U18066 (N_18066,N_16976,N_17108);
nor U18067 (N_18067,N_17057,N_17118);
nor U18068 (N_18068,N_16891,N_17208);
xnor U18069 (N_18069,N_17165,N_17241);
nand U18070 (N_18070,N_17038,N_17233);
nor U18071 (N_18071,N_17224,N_17440);
or U18072 (N_18072,N_16959,N_17097);
or U18073 (N_18073,N_16929,N_17360);
or U18074 (N_18074,N_17242,N_17307);
xnor U18075 (N_18075,N_17187,N_16889);
and U18076 (N_18076,N_16961,N_16988);
or U18077 (N_18077,N_17350,N_17408);
nor U18078 (N_18078,N_16919,N_17372);
xnor U18079 (N_18079,N_16912,N_17497);
and U18080 (N_18080,N_17161,N_17159);
nor U18081 (N_18081,N_17169,N_17098);
xor U18082 (N_18082,N_17304,N_17330);
nand U18083 (N_18083,N_17416,N_17200);
and U18084 (N_18084,N_16967,N_17362);
or U18085 (N_18085,N_17058,N_17300);
or U18086 (N_18086,N_16901,N_17268);
or U18087 (N_18087,N_17465,N_17323);
or U18088 (N_18088,N_17124,N_17115);
or U18089 (N_18089,N_17365,N_17027);
nor U18090 (N_18090,N_16917,N_17165);
and U18091 (N_18091,N_17483,N_17078);
or U18092 (N_18092,N_17449,N_17418);
nand U18093 (N_18093,N_17319,N_17434);
and U18094 (N_18094,N_17331,N_16876);
xnor U18095 (N_18095,N_17298,N_17391);
or U18096 (N_18096,N_17311,N_17313);
nand U18097 (N_18097,N_17263,N_17231);
xor U18098 (N_18098,N_17073,N_16895);
xnor U18099 (N_18099,N_17342,N_17395);
xor U18100 (N_18100,N_17287,N_16948);
or U18101 (N_18101,N_17158,N_17166);
nor U18102 (N_18102,N_16916,N_17025);
and U18103 (N_18103,N_17217,N_17132);
nor U18104 (N_18104,N_17107,N_17237);
nand U18105 (N_18105,N_17429,N_17165);
xnor U18106 (N_18106,N_17143,N_17433);
nand U18107 (N_18107,N_16961,N_17083);
nand U18108 (N_18108,N_17210,N_17353);
or U18109 (N_18109,N_17415,N_16993);
or U18110 (N_18110,N_17202,N_17456);
or U18111 (N_18111,N_16979,N_17428);
or U18112 (N_18112,N_17363,N_17365);
xnor U18113 (N_18113,N_16905,N_16946);
nor U18114 (N_18114,N_16922,N_17274);
nand U18115 (N_18115,N_16980,N_17459);
and U18116 (N_18116,N_17401,N_17353);
nand U18117 (N_18117,N_17079,N_17209);
and U18118 (N_18118,N_17457,N_16890);
and U18119 (N_18119,N_17076,N_17160);
nor U18120 (N_18120,N_17286,N_16934);
or U18121 (N_18121,N_16945,N_17281);
xnor U18122 (N_18122,N_17316,N_17075);
and U18123 (N_18123,N_17405,N_17274);
or U18124 (N_18124,N_16972,N_17014);
nor U18125 (N_18125,N_17756,N_17745);
nand U18126 (N_18126,N_17914,N_17862);
or U18127 (N_18127,N_18081,N_18123);
or U18128 (N_18128,N_17636,N_17705);
xnor U18129 (N_18129,N_17655,N_17529);
nand U18130 (N_18130,N_17912,N_17552);
xor U18131 (N_18131,N_17839,N_18060);
or U18132 (N_18132,N_18083,N_18061);
and U18133 (N_18133,N_17743,N_17808);
xnor U18134 (N_18134,N_17754,N_17604);
nor U18135 (N_18135,N_17879,N_17648);
nor U18136 (N_18136,N_17586,N_17973);
or U18137 (N_18137,N_17541,N_17974);
and U18138 (N_18138,N_17926,N_17704);
nor U18139 (N_18139,N_17840,N_17778);
and U18140 (N_18140,N_18009,N_17728);
nand U18141 (N_18141,N_17519,N_17640);
nor U18142 (N_18142,N_17751,N_17844);
or U18143 (N_18143,N_17890,N_17511);
xor U18144 (N_18144,N_17799,N_17601);
and U18145 (N_18145,N_17989,N_18018);
nor U18146 (N_18146,N_17520,N_17795);
nand U18147 (N_18147,N_17528,N_18029);
nor U18148 (N_18148,N_17698,N_17797);
or U18149 (N_18149,N_17607,N_17677);
nor U18150 (N_18150,N_17544,N_17638);
or U18151 (N_18151,N_17847,N_17939);
nand U18152 (N_18152,N_17582,N_17709);
nand U18153 (N_18153,N_17576,N_17644);
or U18154 (N_18154,N_17632,N_17894);
nand U18155 (N_18155,N_18047,N_17932);
and U18156 (N_18156,N_17920,N_17899);
nor U18157 (N_18157,N_17590,N_17700);
nor U18158 (N_18158,N_17739,N_17666);
xnor U18159 (N_18159,N_18032,N_17738);
xor U18160 (N_18160,N_18003,N_18120);
and U18161 (N_18161,N_18107,N_18118);
and U18162 (N_18162,N_17887,N_17831);
and U18163 (N_18163,N_17958,N_17506);
nand U18164 (N_18164,N_17896,N_17803);
nand U18165 (N_18165,N_17810,N_17575);
and U18166 (N_18166,N_17913,N_17993);
nor U18167 (N_18167,N_17750,N_17950);
nand U18168 (N_18168,N_18058,N_18034);
nor U18169 (N_18169,N_17781,N_17804);
and U18170 (N_18170,N_17849,N_17904);
xnor U18171 (N_18171,N_17692,N_18014);
nor U18172 (N_18172,N_17843,N_17864);
nand U18173 (N_18173,N_17583,N_18078);
or U18174 (N_18174,N_18030,N_18010);
nand U18175 (N_18175,N_18068,N_17717);
nand U18176 (N_18176,N_17612,N_17516);
nor U18177 (N_18177,N_17559,N_17554);
xnor U18178 (N_18178,N_17714,N_17652);
xor U18179 (N_18179,N_17665,N_17654);
nand U18180 (N_18180,N_17757,N_17600);
xnor U18181 (N_18181,N_17727,N_17905);
nor U18182 (N_18182,N_17962,N_17955);
xnor U18183 (N_18183,N_18089,N_18093);
nand U18184 (N_18184,N_17703,N_17518);
and U18185 (N_18185,N_17574,N_17760);
nor U18186 (N_18186,N_17673,N_18063);
xor U18187 (N_18187,N_17551,N_17748);
xnor U18188 (N_18188,N_17690,N_17774);
nor U18189 (N_18189,N_17538,N_17884);
or U18190 (N_18190,N_17512,N_17531);
and U18191 (N_18191,N_17813,N_17992);
or U18192 (N_18192,N_17943,N_18006);
or U18193 (N_18193,N_17959,N_17622);
nor U18194 (N_18194,N_18045,N_17610);
or U18195 (N_18195,N_17647,N_17602);
nor U18196 (N_18196,N_17819,N_18049);
and U18197 (N_18197,N_17807,N_17557);
xor U18198 (N_18198,N_17581,N_17987);
or U18199 (N_18199,N_17597,N_17791);
nand U18200 (N_18200,N_17599,N_17759);
xor U18201 (N_18201,N_18076,N_18062);
or U18202 (N_18202,N_17558,N_18114);
nand U18203 (N_18203,N_17822,N_17620);
xor U18204 (N_18204,N_17867,N_17977);
xor U18205 (N_18205,N_17567,N_17618);
or U18206 (N_18206,N_17817,N_17545);
or U18207 (N_18207,N_17971,N_17829);
nor U18208 (N_18208,N_17776,N_17928);
nor U18209 (N_18209,N_17539,N_18096);
nand U18210 (N_18210,N_17861,N_17758);
and U18211 (N_18211,N_17566,N_18109);
nand U18212 (N_18212,N_17659,N_17821);
nand U18213 (N_18213,N_17838,N_17645);
and U18214 (N_18214,N_17577,N_17708);
xor U18215 (N_18215,N_17967,N_17854);
or U18216 (N_18216,N_17850,N_17951);
nand U18217 (N_18217,N_17685,N_17777);
and U18218 (N_18218,N_17701,N_17882);
xor U18219 (N_18219,N_17903,N_17689);
and U18220 (N_18220,N_17956,N_17938);
or U18221 (N_18221,N_17683,N_17584);
and U18222 (N_18222,N_17981,N_17830);
xor U18223 (N_18223,N_17684,N_17623);
nand U18224 (N_18224,N_17515,N_17883);
or U18225 (N_18225,N_18036,N_17783);
xor U18226 (N_18226,N_18119,N_17790);
and U18227 (N_18227,N_17753,N_18027);
nand U18228 (N_18228,N_18012,N_17934);
nand U18229 (N_18229,N_17814,N_18023);
xnor U18230 (N_18230,N_17787,N_17982);
and U18231 (N_18231,N_17898,N_17869);
or U18232 (N_18232,N_18033,N_17980);
and U18233 (N_18233,N_17579,N_17832);
and U18234 (N_18234,N_17729,N_18056);
and U18235 (N_18235,N_17860,N_17536);
xnor U18236 (N_18236,N_18090,N_17936);
and U18237 (N_18237,N_17929,N_17572);
and U18238 (N_18238,N_17979,N_17766);
xnor U18239 (N_18239,N_17872,N_18042);
nor U18240 (N_18240,N_17578,N_18065);
and U18241 (N_18241,N_18038,N_18087);
nand U18242 (N_18242,N_17837,N_18002);
and U18243 (N_18243,N_18016,N_18048);
or U18244 (N_18244,N_18072,N_17818);
xor U18245 (N_18245,N_17911,N_17816);
xnor U18246 (N_18246,N_17919,N_18015);
or U18247 (N_18247,N_17960,N_17761);
or U18248 (N_18248,N_17719,N_17857);
nand U18249 (N_18249,N_17556,N_17945);
nor U18250 (N_18250,N_17990,N_17796);
nand U18251 (N_18251,N_17637,N_17606);
and U18252 (N_18252,N_17889,N_17957);
xor U18253 (N_18253,N_17909,N_17994);
nand U18254 (N_18254,N_17963,N_17851);
and U18255 (N_18255,N_17532,N_17866);
xnor U18256 (N_18256,N_17853,N_17771);
and U18257 (N_18257,N_18094,N_17710);
or U18258 (N_18258,N_17877,N_17835);
nand U18259 (N_18259,N_17931,N_17731);
xor U18260 (N_18260,N_17616,N_17734);
nor U18261 (N_18261,N_17678,N_18088);
xnor U18262 (N_18262,N_17718,N_17617);
nand U18263 (N_18263,N_17667,N_17681);
xor U18264 (N_18264,N_17635,N_17824);
xor U18265 (N_18265,N_17846,N_17985);
and U18266 (N_18266,N_17646,N_17741);
and U18267 (N_18267,N_17711,N_17933);
nand U18268 (N_18268,N_17779,N_17863);
nor U18269 (N_18269,N_17841,N_17630);
nor U18270 (N_18270,N_17629,N_17649);
nor U18271 (N_18271,N_17561,N_17921);
nor U18272 (N_18272,N_17619,N_17769);
and U18273 (N_18273,N_17798,N_18071);
nand U18274 (N_18274,N_17540,N_17664);
nor U18275 (N_18275,N_17868,N_17508);
xnor U18276 (N_18276,N_17671,N_17686);
xor U18277 (N_18277,N_17725,N_18121);
nand U18278 (N_18278,N_17712,N_18099);
and U18279 (N_18279,N_17972,N_17679);
or U18280 (N_18280,N_17716,N_17715);
and U18281 (N_18281,N_17513,N_17916);
nor U18282 (N_18282,N_18082,N_17687);
xor U18283 (N_18283,N_17876,N_17706);
nor U18284 (N_18284,N_17676,N_17997);
nand U18285 (N_18285,N_17792,N_17949);
nor U18286 (N_18286,N_18086,N_17517);
and U18287 (N_18287,N_17902,N_17588);
and U18288 (N_18288,N_17806,N_18084);
and U18289 (N_18289,N_17788,N_17553);
xor U18290 (N_18290,N_18050,N_17733);
xor U18291 (N_18291,N_17625,N_17952);
nand U18292 (N_18292,N_17895,N_17651);
nand U18293 (N_18293,N_17875,N_17827);
xor U18294 (N_18294,N_17873,N_18085);
and U18295 (N_18295,N_17770,N_17737);
nor U18296 (N_18296,N_17713,N_18101);
and U18297 (N_18297,N_17611,N_17550);
and U18298 (N_18298,N_17772,N_17746);
and U18299 (N_18299,N_17674,N_18080);
nand U18300 (N_18300,N_18046,N_17762);
nand U18301 (N_18301,N_17848,N_17744);
and U18302 (N_18302,N_17961,N_17947);
or U18303 (N_18303,N_17500,N_17888);
or U18304 (N_18304,N_17680,N_17591);
or U18305 (N_18305,N_18075,N_17815);
nand U18306 (N_18306,N_17927,N_17688);
and U18307 (N_18307,N_18020,N_18000);
or U18308 (N_18308,N_17596,N_18055);
and U18309 (N_18309,N_18067,N_17918);
nor U18310 (N_18310,N_17735,N_17812);
xor U18311 (N_18311,N_17537,N_18017);
nor U18312 (N_18312,N_17624,N_17663);
nor U18313 (N_18313,N_17609,N_18026);
nor U18314 (N_18314,N_18103,N_17749);
nor U18315 (N_18315,N_17670,N_17970);
or U18316 (N_18316,N_17907,N_18105);
and U18317 (N_18317,N_17811,N_18111);
or U18318 (N_18318,N_17723,N_18064);
nor U18319 (N_18319,N_18113,N_17794);
xnor U18320 (N_18320,N_17641,N_18059);
nand U18321 (N_18321,N_17852,N_17585);
nor U18322 (N_18322,N_17983,N_18035);
xor U18323 (N_18323,N_17521,N_17917);
nand U18324 (N_18324,N_18043,N_17732);
nor U18325 (N_18325,N_17966,N_18095);
nand U18326 (N_18326,N_17747,N_18021);
nor U18327 (N_18327,N_17800,N_17998);
and U18328 (N_18328,N_17507,N_17908);
xnor U18329 (N_18329,N_17660,N_17805);
and U18330 (N_18330,N_17859,N_17563);
nand U18331 (N_18331,N_17721,N_17595);
xor U18332 (N_18332,N_17662,N_17548);
nor U18333 (N_18333,N_18057,N_17661);
and U18334 (N_18334,N_17740,N_17634);
xor U18335 (N_18335,N_17580,N_17555);
or U18336 (N_18336,N_17504,N_18013);
or U18337 (N_18337,N_17874,N_17569);
and U18338 (N_18338,N_17886,N_17656);
and U18339 (N_18339,N_18079,N_17773);
nand U18340 (N_18340,N_17722,N_18102);
and U18341 (N_18341,N_17871,N_17720);
or U18342 (N_18342,N_17786,N_17940);
nor U18343 (N_18343,N_18053,N_18037);
nor U18344 (N_18344,N_17568,N_17834);
nor U18345 (N_18345,N_17964,N_18040);
and U18346 (N_18346,N_17525,N_17878);
nand U18347 (N_18347,N_17802,N_17924);
nor U18348 (N_18348,N_17828,N_18041);
and U18349 (N_18349,N_18069,N_17650);
xnor U18350 (N_18350,N_17763,N_18110);
xnor U18351 (N_18351,N_17941,N_17954);
nor U18352 (N_18352,N_17605,N_18091);
and U18353 (N_18353,N_17530,N_18077);
and U18354 (N_18354,N_17855,N_17668);
xor U18355 (N_18355,N_17639,N_17880);
nor U18356 (N_18356,N_18024,N_17675);
nand U18357 (N_18357,N_17643,N_18001);
nand U18358 (N_18358,N_17615,N_17526);
and U18359 (N_18359,N_17845,N_17823);
nand U18360 (N_18360,N_17589,N_17897);
nor U18361 (N_18361,N_17833,N_17592);
or U18362 (N_18362,N_17767,N_17653);
nand U18363 (N_18363,N_17535,N_17631);
or U18364 (N_18364,N_18011,N_17503);
nand U18365 (N_18365,N_17642,N_17825);
and U18366 (N_18366,N_17527,N_17672);
or U18367 (N_18367,N_18073,N_17657);
nor U18368 (N_18368,N_17820,N_17842);
and U18369 (N_18369,N_17682,N_17944);
and U18370 (N_18370,N_18005,N_17502);
and U18371 (N_18371,N_17598,N_17885);
xor U18372 (N_18372,N_17699,N_17893);
and U18373 (N_18373,N_17780,N_17906);
or U18374 (N_18374,N_17693,N_17509);
and U18375 (N_18375,N_17564,N_17627);
or U18376 (N_18376,N_17547,N_18066);
or U18377 (N_18377,N_17946,N_17533);
nor U18378 (N_18378,N_17881,N_17991);
nor U18379 (N_18379,N_18108,N_17995);
nand U18380 (N_18380,N_18054,N_17614);
xnor U18381 (N_18381,N_17626,N_17726);
xnor U18382 (N_18382,N_18004,N_17522);
nor U18383 (N_18383,N_17984,N_17562);
xor U18384 (N_18384,N_17570,N_17910);
xnor U18385 (N_18385,N_17510,N_17594);
xnor U18386 (N_18386,N_17542,N_17935);
and U18387 (N_18387,N_17789,N_18112);
or U18388 (N_18388,N_17793,N_17768);
and U18389 (N_18389,N_17836,N_17633);
or U18390 (N_18390,N_17923,N_17999);
nand U18391 (N_18391,N_18031,N_17901);
nand U18392 (N_18392,N_17801,N_17892);
xor U18393 (N_18393,N_17696,N_17965);
nor U18394 (N_18394,N_17826,N_17942);
nor U18395 (N_18395,N_18117,N_17724);
and U18396 (N_18396,N_17784,N_17986);
or U18397 (N_18397,N_17930,N_17976);
or U18398 (N_18398,N_17782,N_17628);
xor U18399 (N_18399,N_17856,N_18008);
nand U18400 (N_18400,N_17514,N_17523);
nor U18401 (N_18401,N_17765,N_18052);
and U18402 (N_18402,N_17702,N_18106);
xnor U18403 (N_18403,N_17603,N_17891);
nor U18404 (N_18404,N_17501,N_18019);
nor U18405 (N_18405,N_17613,N_18122);
nand U18406 (N_18406,N_17764,N_18097);
or U18407 (N_18407,N_17858,N_18039);
and U18408 (N_18408,N_17736,N_17621);
nor U18409 (N_18409,N_18074,N_17571);
xor U18410 (N_18410,N_18124,N_17695);
nor U18411 (N_18411,N_18104,N_17658);
xnor U18412 (N_18412,N_17925,N_18022);
nand U18413 (N_18413,N_18116,N_17900);
and U18414 (N_18414,N_17752,N_17543);
nand U18415 (N_18415,N_17505,N_17953);
and U18416 (N_18416,N_17524,N_17691);
or U18417 (N_18417,N_17755,N_17565);
or U18418 (N_18418,N_17573,N_18100);
and U18419 (N_18419,N_17988,N_18051);
nand U18420 (N_18420,N_17669,N_17865);
nand U18421 (N_18421,N_18098,N_17915);
or U18422 (N_18422,N_17697,N_18070);
nand U18423 (N_18423,N_17978,N_17587);
xor U18424 (N_18424,N_17969,N_17968);
nor U18425 (N_18425,N_17922,N_17870);
nor U18426 (N_18426,N_18115,N_17742);
nand U18427 (N_18427,N_17730,N_17775);
or U18428 (N_18428,N_17549,N_17534);
nand U18429 (N_18429,N_18007,N_17937);
nor U18430 (N_18430,N_17809,N_17996);
nand U18431 (N_18431,N_18028,N_17593);
or U18432 (N_18432,N_17560,N_17785);
nand U18433 (N_18433,N_17694,N_18044);
and U18434 (N_18434,N_17975,N_17608);
or U18435 (N_18435,N_18092,N_17546);
nand U18436 (N_18436,N_17707,N_17948);
or U18437 (N_18437,N_18025,N_17925);
xnor U18438 (N_18438,N_17578,N_17996);
nor U18439 (N_18439,N_17726,N_17898);
and U18440 (N_18440,N_17930,N_17969);
or U18441 (N_18441,N_18087,N_17709);
and U18442 (N_18442,N_17836,N_17646);
xor U18443 (N_18443,N_17658,N_17696);
nor U18444 (N_18444,N_17649,N_17664);
nand U18445 (N_18445,N_17704,N_17712);
or U18446 (N_18446,N_17546,N_17650);
nor U18447 (N_18447,N_17785,N_17746);
or U18448 (N_18448,N_17538,N_17641);
and U18449 (N_18449,N_17753,N_17509);
and U18450 (N_18450,N_17833,N_17863);
nor U18451 (N_18451,N_17719,N_17699);
or U18452 (N_18452,N_17820,N_18007);
nor U18453 (N_18453,N_17943,N_17514);
and U18454 (N_18454,N_18020,N_17868);
and U18455 (N_18455,N_18024,N_17541);
nor U18456 (N_18456,N_17668,N_18032);
xnor U18457 (N_18457,N_17713,N_17883);
nor U18458 (N_18458,N_17596,N_18089);
xnor U18459 (N_18459,N_17613,N_17548);
or U18460 (N_18460,N_17984,N_18008);
xnor U18461 (N_18461,N_17977,N_17754);
nor U18462 (N_18462,N_17879,N_18112);
and U18463 (N_18463,N_17561,N_17904);
nor U18464 (N_18464,N_17594,N_17952);
nor U18465 (N_18465,N_17616,N_17684);
or U18466 (N_18466,N_17837,N_17505);
or U18467 (N_18467,N_18015,N_17726);
nor U18468 (N_18468,N_17806,N_17567);
nand U18469 (N_18469,N_18067,N_17670);
or U18470 (N_18470,N_17831,N_17661);
and U18471 (N_18471,N_18065,N_17942);
nand U18472 (N_18472,N_17915,N_17634);
and U18473 (N_18473,N_17872,N_17899);
nor U18474 (N_18474,N_17555,N_17673);
or U18475 (N_18475,N_17865,N_17503);
or U18476 (N_18476,N_18041,N_17652);
or U18477 (N_18477,N_17712,N_17542);
nand U18478 (N_18478,N_17937,N_18110);
xor U18479 (N_18479,N_17803,N_17654);
nor U18480 (N_18480,N_17591,N_17922);
and U18481 (N_18481,N_18010,N_17878);
nor U18482 (N_18482,N_17670,N_17882);
nand U18483 (N_18483,N_18027,N_17635);
and U18484 (N_18484,N_17715,N_17826);
nand U18485 (N_18485,N_17717,N_17649);
or U18486 (N_18486,N_17652,N_17990);
or U18487 (N_18487,N_18058,N_17637);
nor U18488 (N_18488,N_17646,N_17640);
and U18489 (N_18489,N_17912,N_17822);
or U18490 (N_18490,N_17625,N_17805);
and U18491 (N_18491,N_17733,N_18016);
nand U18492 (N_18492,N_18058,N_18057);
nor U18493 (N_18493,N_17568,N_17683);
and U18494 (N_18494,N_17590,N_17514);
and U18495 (N_18495,N_18053,N_17781);
and U18496 (N_18496,N_17718,N_17867);
xor U18497 (N_18497,N_18103,N_17817);
and U18498 (N_18498,N_17866,N_17533);
or U18499 (N_18499,N_17536,N_17800);
or U18500 (N_18500,N_18082,N_17836);
or U18501 (N_18501,N_17758,N_17955);
xor U18502 (N_18502,N_17615,N_17850);
and U18503 (N_18503,N_17570,N_17919);
nand U18504 (N_18504,N_17985,N_17527);
nor U18505 (N_18505,N_17588,N_17699);
xor U18506 (N_18506,N_17635,N_17948);
nor U18507 (N_18507,N_17757,N_17878);
nand U18508 (N_18508,N_17606,N_17779);
nor U18509 (N_18509,N_17752,N_17611);
nand U18510 (N_18510,N_17813,N_17725);
or U18511 (N_18511,N_17593,N_17686);
and U18512 (N_18512,N_17871,N_17803);
xnor U18513 (N_18513,N_17903,N_18031);
or U18514 (N_18514,N_17650,N_17592);
or U18515 (N_18515,N_17929,N_17623);
and U18516 (N_18516,N_17556,N_18053);
and U18517 (N_18517,N_17976,N_17623);
nand U18518 (N_18518,N_17668,N_18075);
or U18519 (N_18519,N_18072,N_17681);
nand U18520 (N_18520,N_18048,N_17855);
and U18521 (N_18521,N_17590,N_17746);
or U18522 (N_18522,N_17559,N_17635);
xor U18523 (N_18523,N_18050,N_17570);
nand U18524 (N_18524,N_18028,N_17905);
or U18525 (N_18525,N_17633,N_17638);
nand U18526 (N_18526,N_17921,N_17989);
or U18527 (N_18527,N_17730,N_17811);
nand U18528 (N_18528,N_17604,N_17913);
xnor U18529 (N_18529,N_17880,N_18051);
or U18530 (N_18530,N_17525,N_18033);
and U18531 (N_18531,N_17674,N_17899);
nor U18532 (N_18532,N_17966,N_17703);
and U18533 (N_18533,N_17895,N_17778);
nand U18534 (N_18534,N_17794,N_18005);
xor U18535 (N_18535,N_17642,N_17962);
and U18536 (N_18536,N_17663,N_18049);
nand U18537 (N_18537,N_17837,N_17582);
nand U18538 (N_18538,N_17944,N_17568);
nand U18539 (N_18539,N_17750,N_17699);
or U18540 (N_18540,N_17943,N_17620);
xor U18541 (N_18541,N_17556,N_17686);
xor U18542 (N_18542,N_17761,N_18035);
and U18543 (N_18543,N_17710,N_17616);
or U18544 (N_18544,N_17598,N_18078);
nand U18545 (N_18545,N_17627,N_17977);
or U18546 (N_18546,N_17603,N_17626);
or U18547 (N_18547,N_17911,N_17841);
nand U18548 (N_18548,N_17791,N_17647);
xnor U18549 (N_18549,N_17877,N_17852);
or U18550 (N_18550,N_17931,N_17629);
and U18551 (N_18551,N_17880,N_18119);
xor U18552 (N_18552,N_17743,N_18038);
xor U18553 (N_18553,N_18009,N_17812);
nor U18554 (N_18554,N_17795,N_18076);
nor U18555 (N_18555,N_18085,N_18094);
and U18556 (N_18556,N_17808,N_17920);
nand U18557 (N_18557,N_17663,N_17606);
nor U18558 (N_18558,N_17532,N_17985);
nand U18559 (N_18559,N_18041,N_17598);
nor U18560 (N_18560,N_17650,N_18121);
and U18561 (N_18561,N_18047,N_17718);
nor U18562 (N_18562,N_17682,N_17796);
or U18563 (N_18563,N_17822,N_17873);
nor U18564 (N_18564,N_17806,N_17519);
or U18565 (N_18565,N_17505,N_17754);
nand U18566 (N_18566,N_17978,N_17977);
xnor U18567 (N_18567,N_17850,N_17582);
nor U18568 (N_18568,N_17742,N_17699);
and U18569 (N_18569,N_18001,N_17749);
xor U18570 (N_18570,N_17905,N_18091);
and U18571 (N_18571,N_17610,N_17934);
nand U18572 (N_18572,N_17868,N_17750);
and U18573 (N_18573,N_17852,N_18021);
and U18574 (N_18574,N_17951,N_17555);
xnor U18575 (N_18575,N_17883,N_17685);
nor U18576 (N_18576,N_18060,N_18004);
and U18577 (N_18577,N_17999,N_18074);
xnor U18578 (N_18578,N_17912,N_17505);
or U18579 (N_18579,N_17845,N_17738);
or U18580 (N_18580,N_17997,N_17746);
and U18581 (N_18581,N_17941,N_17781);
nand U18582 (N_18582,N_17810,N_17667);
or U18583 (N_18583,N_18024,N_18036);
xor U18584 (N_18584,N_18111,N_17801);
or U18585 (N_18585,N_17742,N_18050);
nor U18586 (N_18586,N_17576,N_18019);
or U18587 (N_18587,N_17958,N_17523);
or U18588 (N_18588,N_17552,N_17669);
nor U18589 (N_18589,N_17770,N_17994);
or U18590 (N_18590,N_17937,N_17788);
nand U18591 (N_18591,N_17984,N_18041);
or U18592 (N_18592,N_17656,N_17565);
nand U18593 (N_18593,N_17601,N_17655);
xnor U18594 (N_18594,N_17523,N_17899);
xnor U18595 (N_18595,N_17880,N_17528);
nand U18596 (N_18596,N_17579,N_17958);
or U18597 (N_18597,N_18025,N_17926);
nor U18598 (N_18598,N_17953,N_18085);
nor U18599 (N_18599,N_17812,N_18108);
nor U18600 (N_18600,N_18040,N_18116);
and U18601 (N_18601,N_17811,N_18045);
nand U18602 (N_18602,N_17917,N_18061);
nor U18603 (N_18603,N_18031,N_17826);
xnor U18604 (N_18604,N_17708,N_18054);
or U18605 (N_18605,N_18015,N_17997);
xnor U18606 (N_18606,N_17883,N_17943);
xor U18607 (N_18607,N_17589,N_18045);
xor U18608 (N_18608,N_17870,N_18079);
or U18609 (N_18609,N_17849,N_17884);
nor U18610 (N_18610,N_17545,N_17699);
and U18611 (N_18611,N_18077,N_17588);
or U18612 (N_18612,N_17777,N_17714);
nor U18613 (N_18613,N_17908,N_17689);
or U18614 (N_18614,N_17505,N_17984);
xor U18615 (N_18615,N_17734,N_17590);
and U18616 (N_18616,N_17593,N_17708);
and U18617 (N_18617,N_18095,N_17588);
nor U18618 (N_18618,N_17825,N_17703);
or U18619 (N_18619,N_17910,N_17676);
xor U18620 (N_18620,N_17632,N_17513);
nor U18621 (N_18621,N_17971,N_17755);
nand U18622 (N_18622,N_18123,N_17825);
nand U18623 (N_18623,N_17727,N_17920);
or U18624 (N_18624,N_17584,N_17925);
nor U18625 (N_18625,N_18063,N_17911);
xnor U18626 (N_18626,N_17945,N_17530);
and U18627 (N_18627,N_17592,N_18080);
or U18628 (N_18628,N_18027,N_17709);
nand U18629 (N_18629,N_17700,N_17942);
and U18630 (N_18630,N_17867,N_17687);
and U18631 (N_18631,N_17657,N_17662);
nor U18632 (N_18632,N_17734,N_17918);
nor U18633 (N_18633,N_17962,N_17659);
or U18634 (N_18634,N_18093,N_17746);
nand U18635 (N_18635,N_17939,N_17933);
and U18636 (N_18636,N_17704,N_17632);
or U18637 (N_18637,N_17752,N_17620);
nand U18638 (N_18638,N_18081,N_18087);
or U18639 (N_18639,N_17577,N_17641);
xnor U18640 (N_18640,N_17921,N_17588);
nor U18641 (N_18641,N_18004,N_17631);
or U18642 (N_18642,N_17649,N_17727);
and U18643 (N_18643,N_18019,N_17963);
or U18644 (N_18644,N_18075,N_17743);
or U18645 (N_18645,N_17964,N_17708);
xnor U18646 (N_18646,N_17539,N_17702);
and U18647 (N_18647,N_18121,N_17704);
or U18648 (N_18648,N_17846,N_17925);
and U18649 (N_18649,N_17604,N_18028);
and U18650 (N_18650,N_17975,N_17737);
nor U18651 (N_18651,N_17954,N_18026);
and U18652 (N_18652,N_17520,N_17655);
nand U18653 (N_18653,N_17651,N_17641);
nand U18654 (N_18654,N_17861,N_17931);
nand U18655 (N_18655,N_17609,N_17819);
nand U18656 (N_18656,N_17741,N_17594);
xor U18657 (N_18657,N_17904,N_17567);
nor U18658 (N_18658,N_18087,N_17572);
and U18659 (N_18659,N_17682,N_17591);
and U18660 (N_18660,N_18064,N_18089);
xor U18661 (N_18661,N_17993,N_17878);
nand U18662 (N_18662,N_17887,N_17536);
or U18663 (N_18663,N_17917,N_18018);
and U18664 (N_18664,N_17679,N_18076);
nor U18665 (N_18665,N_17899,N_17730);
nor U18666 (N_18666,N_17878,N_17913);
nor U18667 (N_18667,N_18010,N_17900);
and U18668 (N_18668,N_17662,N_17775);
nand U18669 (N_18669,N_17792,N_17601);
nor U18670 (N_18670,N_17506,N_17940);
and U18671 (N_18671,N_17665,N_17612);
or U18672 (N_18672,N_17841,N_17529);
xor U18673 (N_18673,N_18017,N_17843);
nand U18674 (N_18674,N_18105,N_17804);
xor U18675 (N_18675,N_17762,N_17564);
xnor U18676 (N_18676,N_18032,N_18075);
xor U18677 (N_18677,N_17630,N_17576);
nand U18678 (N_18678,N_17579,N_17518);
xnor U18679 (N_18679,N_18108,N_17582);
xor U18680 (N_18680,N_17832,N_18032);
and U18681 (N_18681,N_18000,N_17687);
nand U18682 (N_18682,N_17943,N_18085);
nand U18683 (N_18683,N_17811,N_17967);
and U18684 (N_18684,N_17641,N_18033);
nand U18685 (N_18685,N_17515,N_17892);
or U18686 (N_18686,N_17622,N_18025);
and U18687 (N_18687,N_17915,N_17622);
nand U18688 (N_18688,N_17798,N_17548);
nand U18689 (N_18689,N_17887,N_17981);
or U18690 (N_18690,N_17794,N_17755);
nand U18691 (N_18691,N_17645,N_17594);
xor U18692 (N_18692,N_17848,N_17601);
and U18693 (N_18693,N_18087,N_17734);
xor U18694 (N_18694,N_18072,N_18012);
xor U18695 (N_18695,N_18027,N_18102);
and U18696 (N_18696,N_17908,N_17672);
nand U18697 (N_18697,N_17989,N_17869);
nor U18698 (N_18698,N_17522,N_17996);
and U18699 (N_18699,N_17555,N_18008);
and U18700 (N_18700,N_17607,N_17649);
nor U18701 (N_18701,N_17714,N_17669);
or U18702 (N_18702,N_18101,N_17570);
xnor U18703 (N_18703,N_17631,N_17565);
nor U18704 (N_18704,N_17763,N_17560);
nor U18705 (N_18705,N_18043,N_17594);
nor U18706 (N_18706,N_17913,N_18026);
nor U18707 (N_18707,N_18036,N_17525);
or U18708 (N_18708,N_17613,N_17969);
and U18709 (N_18709,N_17946,N_17564);
xnor U18710 (N_18710,N_17539,N_17804);
nor U18711 (N_18711,N_17771,N_17677);
nand U18712 (N_18712,N_17662,N_17643);
or U18713 (N_18713,N_17738,N_17778);
or U18714 (N_18714,N_18029,N_17930);
or U18715 (N_18715,N_17935,N_17835);
nor U18716 (N_18716,N_17884,N_17897);
nand U18717 (N_18717,N_18082,N_17960);
and U18718 (N_18718,N_17961,N_17716);
nor U18719 (N_18719,N_17923,N_18012);
nor U18720 (N_18720,N_17934,N_17870);
and U18721 (N_18721,N_17508,N_18026);
or U18722 (N_18722,N_17821,N_18022);
nand U18723 (N_18723,N_17984,N_17786);
nor U18724 (N_18724,N_18124,N_17891);
and U18725 (N_18725,N_17945,N_17585);
and U18726 (N_18726,N_17926,N_17757);
xor U18727 (N_18727,N_17876,N_18067);
or U18728 (N_18728,N_17588,N_17946);
and U18729 (N_18729,N_18122,N_17845);
xor U18730 (N_18730,N_17845,N_17724);
and U18731 (N_18731,N_17892,N_17566);
nand U18732 (N_18732,N_17546,N_17961);
xnor U18733 (N_18733,N_17665,N_17734);
nand U18734 (N_18734,N_17888,N_17699);
nor U18735 (N_18735,N_17702,N_17853);
nand U18736 (N_18736,N_17581,N_17776);
or U18737 (N_18737,N_18077,N_17996);
nor U18738 (N_18738,N_17837,N_17965);
xor U18739 (N_18739,N_17910,N_17986);
nand U18740 (N_18740,N_17827,N_17519);
and U18741 (N_18741,N_17891,N_18118);
nand U18742 (N_18742,N_17615,N_17726);
and U18743 (N_18743,N_17906,N_17502);
and U18744 (N_18744,N_17725,N_17690);
xor U18745 (N_18745,N_17944,N_17971);
and U18746 (N_18746,N_17958,N_18059);
nor U18747 (N_18747,N_18041,N_17902);
xnor U18748 (N_18748,N_17801,N_17639);
nand U18749 (N_18749,N_18020,N_17851);
nand U18750 (N_18750,N_18399,N_18186);
or U18751 (N_18751,N_18244,N_18324);
and U18752 (N_18752,N_18700,N_18320);
xor U18753 (N_18753,N_18631,N_18139);
and U18754 (N_18754,N_18705,N_18422);
and U18755 (N_18755,N_18668,N_18734);
nand U18756 (N_18756,N_18493,N_18731);
and U18757 (N_18757,N_18430,N_18174);
or U18758 (N_18758,N_18628,N_18382);
nand U18759 (N_18759,N_18485,N_18612);
xnor U18760 (N_18760,N_18397,N_18685);
nand U18761 (N_18761,N_18605,N_18189);
nor U18762 (N_18762,N_18423,N_18130);
or U18763 (N_18763,N_18603,N_18249);
xor U18764 (N_18764,N_18720,N_18175);
nor U18765 (N_18765,N_18405,N_18489);
nor U18766 (N_18766,N_18352,N_18235);
or U18767 (N_18767,N_18208,N_18245);
nand U18768 (N_18768,N_18665,N_18209);
and U18769 (N_18769,N_18125,N_18184);
nor U18770 (N_18770,N_18657,N_18435);
nor U18771 (N_18771,N_18254,N_18514);
xnor U18772 (N_18772,N_18210,N_18718);
or U18773 (N_18773,N_18313,N_18323);
nor U18774 (N_18774,N_18142,N_18398);
xnor U18775 (N_18775,N_18539,N_18149);
nor U18776 (N_18776,N_18617,N_18201);
and U18777 (N_18777,N_18523,N_18265);
nand U18778 (N_18778,N_18616,N_18376);
or U18779 (N_18779,N_18503,N_18241);
xnor U18780 (N_18780,N_18452,N_18296);
or U18781 (N_18781,N_18721,N_18146);
nor U18782 (N_18782,N_18145,N_18273);
and U18783 (N_18783,N_18333,N_18574);
nand U18784 (N_18784,N_18411,N_18308);
nor U18785 (N_18785,N_18153,N_18219);
and U18786 (N_18786,N_18613,N_18699);
and U18787 (N_18787,N_18159,N_18297);
nor U18788 (N_18788,N_18476,N_18334);
or U18789 (N_18789,N_18369,N_18483);
xor U18790 (N_18790,N_18715,N_18164);
xor U18791 (N_18791,N_18500,N_18739);
xor U18792 (N_18792,N_18545,N_18428);
or U18793 (N_18793,N_18622,N_18177);
or U18794 (N_18794,N_18306,N_18325);
and U18795 (N_18795,N_18623,N_18740);
or U18796 (N_18796,N_18591,N_18566);
nand U18797 (N_18797,N_18392,N_18698);
and U18798 (N_18798,N_18330,N_18446);
nor U18799 (N_18799,N_18374,N_18196);
nor U18800 (N_18800,N_18311,N_18237);
and U18801 (N_18801,N_18161,N_18275);
and U18802 (N_18802,N_18318,N_18451);
nand U18803 (N_18803,N_18144,N_18732);
or U18804 (N_18804,N_18637,N_18517);
or U18805 (N_18805,N_18513,N_18327);
nor U18806 (N_18806,N_18129,N_18687);
nand U18807 (N_18807,N_18194,N_18638);
nor U18808 (N_18808,N_18415,N_18172);
nor U18809 (N_18809,N_18480,N_18585);
nor U18810 (N_18810,N_18437,N_18512);
nand U18811 (N_18811,N_18378,N_18364);
nand U18812 (N_18812,N_18542,N_18266);
and U18813 (N_18813,N_18494,N_18738);
xnor U18814 (N_18814,N_18213,N_18419);
nor U18815 (N_18815,N_18239,N_18733);
or U18816 (N_18816,N_18525,N_18182);
nor U18817 (N_18817,N_18580,N_18280);
or U18818 (N_18818,N_18586,N_18233);
and U18819 (N_18819,N_18564,N_18462);
nand U18820 (N_18820,N_18328,N_18302);
and U18821 (N_18821,N_18481,N_18474);
nand U18822 (N_18822,N_18171,N_18472);
nand U18823 (N_18823,N_18455,N_18625);
or U18824 (N_18824,N_18238,N_18644);
and U18825 (N_18825,N_18300,N_18589);
or U18826 (N_18826,N_18424,N_18304);
nor U18827 (N_18827,N_18659,N_18127);
nand U18828 (N_18828,N_18348,N_18597);
nand U18829 (N_18829,N_18363,N_18741);
and U18830 (N_18830,N_18457,N_18742);
or U18831 (N_18831,N_18290,N_18258);
nand U18832 (N_18832,N_18601,N_18147);
or U18833 (N_18833,N_18632,N_18389);
nor U18834 (N_18834,N_18203,N_18530);
xnor U18835 (N_18835,N_18349,N_18450);
xor U18836 (N_18836,N_18285,N_18669);
nor U18837 (N_18837,N_18608,N_18402);
nor U18838 (N_18838,N_18384,N_18640);
nor U18839 (N_18839,N_18747,N_18132);
xnor U18840 (N_18840,N_18646,N_18690);
nand U18841 (N_18841,N_18188,N_18575);
and U18842 (N_18842,N_18307,N_18614);
nand U18843 (N_18843,N_18261,N_18710);
nand U18844 (N_18844,N_18256,N_18284);
nand U18845 (N_18845,N_18192,N_18507);
or U18846 (N_18846,N_18353,N_18588);
xor U18847 (N_18847,N_18448,N_18596);
or U18848 (N_18848,N_18367,N_18473);
nand U18849 (N_18849,N_18169,N_18453);
and U18850 (N_18850,N_18620,N_18178);
nor U18851 (N_18851,N_18426,N_18711);
or U18852 (N_18852,N_18358,N_18317);
and U18853 (N_18853,N_18412,N_18624);
or U18854 (N_18854,N_18381,N_18135);
and U18855 (N_18855,N_18548,N_18357);
nand U18856 (N_18856,N_18314,N_18294);
and U18857 (N_18857,N_18240,N_18534);
nand U18858 (N_18858,N_18630,N_18354);
xor U18859 (N_18859,N_18425,N_18730);
nor U18860 (N_18860,N_18185,N_18745);
and U18861 (N_18861,N_18243,N_18224);
nand U18862 (N_18862,N_18658,N_18642);
or U18863 (N_18863,N_18331,N_18247);
or U18864 (N_18864,N_18277,N_18554);
or U18865 (N_18865,N_18373,N_18414);
nor U18866 (N_18866,N_18743,N_18216);
nand U18867 (N_18867,N_18326,N_18447);
xor U18868 (N_18868,N_18694,N_18166);
or U18869 (N_18869,N_18270,N_18684);
and U18870 (N_18870,N_18579,N_18592);
nand U18871 (N_18871,N_18410,N_18491);
nand U18872 (N_18872,N_18394,N_18681);
and U18873 (N_18873,N_18140,N_18420);
nor U18874 (N_18874,N_18242,N_18533);
nand U18875 (N_18875,N_18482,N_18496);
nand U18876 (N_18876,N_18499,N_18683);
or U18877 (N_18877,N_18281,N_18246);
nor U18878 (N_18878,N_18636,N_18571);
xor U18879 (N_18879,N_18553,N_18214);
and U18880 (N_18880,N_18652,N_18168);
and U18881 (N_18881,N_18527,N_18726);
and U18882 (N_18882,N_18322,N_18519);
nand U18883 (N_18883,N_18439,N_18343);
or U18884 (N_18884,N_18627,N_18529);
or U18885 (N_18885,N_18160,N_18618);
nor U18886 (N_18886,N_18193,N_18639);
or U18887 (N_18887,N_18305,N_18163);
xor U18888 (N_18888,N_18634,N_18152);
xnor U18889 (N_18889,N_18274,N_18647);
nand U18890 (N_18890,N_18744,N_18408);
or U18891 (N_18891,N_18283,N_18427);
or U18892 (N_18892,N_18502,N_18377);
nand U18893 (N_18893,N_18299,N_18362);
nor U18894 (N_18894,N_18716,N_18371);
nor U18895 (N_18895,N_18128,N_18561);
nand U18896 (N_18896,N_18212,N_18136);
and U18897 (N_18897,N_18475,N_18292);
or U18898 (N_18898,N_18309,N_18717);
or U18899 (N_18899,N_18547,N_18355);
xnor U18900 (N_18900,N_18736,N_18471);
and U18901 (N_18901,N_18436,N_18440);
nand U18902 (N_18902,N_18599,N_18590);
xnor U18903 (N_18903,N_18498,N_18255);
nor U18904 (N_18904,N_18445,N_18339);
nor U18905 (N_18905,N_18651,N_18342);
nand U18906 (N_18906,N_18151,N_18312);
and U18907 (N_18907,N_18133,N_18449);
nor U18908 (N_18908,N_18198,N_18505);
and U18909 (N_18909,N_18315,N_18225);
xor U18910 (N_18910,N_18158,N_18336);
and U18911 (N_18911,N_18218,N_18458);
or U18912 (N_18912,N_18269,N_18704);
nand U18913 (N_18913,N_18137,N_18391);
and U18914 (N_18914,N_18727,N_18217);
and U18915 (N_18915,N_18584,N_18538);
nor U18916 (N_18916,N_18433,N_18663);
nor U18917 (N_18917,N_18434,N_18583);
nor U18918 (N_18918,N_18234,N_18543);
nor U18919 (N_18919,N_18165,N_18679);
and U18920 (N_18920,N_18131,N_18735);
xor U18921 (N_18921,N_18386,N_18197);
xor U18922 (N_18922,N_18232,N_18372);
xor U18923 (N_18923,N_18662,N_18673);
xnor U18924 (N_18924,N_18350,N_18515);
xnor U18925 (N_18925,N_18401,N_18709);
nor U18926 (N_18926,N_18466,N_18697);
and U18927 (N_18927,N_18677,N_18220);
nor U18928 (N_18928,N_18746,N_18495);
xor U18929 (N_18929,N_18286,N_18725);
and U18930 (N_18930,N_18595,N_18737);
nand U18931 (N_18931,N_18464,N_18582);
xnor U18932 (N_18932,N_18712,N_18470);
nor U18933 (N_18933,N_18332,N_18497);
nor U18934 (N_18934,N_18602,N_18385);
nand U18935 (N_18935,N_18520,N_18691);
nor U18936 (N_18936,N_18594,N_18484);
and U18937 (N_18937,N_18526,N_18532);
or U18938 (N_18938,N_18406,N_18228);
or U18939 (N_18939,N_18337,N_18393);
xnor U18940 (N_18940,N_18199,N_18600);
or U18941 (N_18941,N_18703,N_18508);
or U18942 (N_18942,N_18252,N_18154);
xnor U18943 (N_18943,N_18356,N_18674);
xnor U18944 (N_18944,N_18649,N_18442);
nor U18945 (N_18945,N_18516,N_18215);
nor U18946 (N_18946,N_18250,N_18276);
and U18947 (N_18947,N_18572,N_18728);
and U18948 (N_18948,N_18609,N_18682);
nor U18949 (N_18949,N_18672,N_18461);
nor U18950 (N_18950,N_18549,N_18492);
nand U18951 (N_18951,N_18635,N_18263);
xnor U18952 (N_18952,N_18223,N_18230);
xor U18953 (N_18953,N_18541,N_18301);
nor U18954 (N_18954,N_18438,N_18559);
nor U18955 (N_18955,N_18345,N_18141);
nand U18956 (N_18956,N_18407,N_18176);
nand U18957 (N_18957,N_18417,N_18179);
xnor U18958 (N_18958,N_18504,N_18573);
or U18959 (N_18959,N_18714,N_18706);
nand U18960 (N_18960,N_18678,N_18722);
and U18961 (N_18961,N_18211,N_18578);
xnor U18962 (N_18962,N_18469,N_18404);
and U18963 (N_18963,N_18289,N_18156);
or U18964 (N_18964,N_18552,N_18205);
or U18965 (N_18965,N_18170,N_18604);
nor U18966 (N_18966,N_18335,N_18581);
xor U18967 (N_18967,N_18167,N_18524);
nand U18968 (N_18968,N_18465,N_18248);
xnor U18969 (N_18969,N_18531,N_18670);
nor U18970 (N_18970,N_18390,N_18431);
and U18971 (N_18971,N_18567,N_18251);
nand U18972 (N_18972,N_18221,N_18303);
xor U18973 (N_18973,N_18558,N_18259);
xor U18974 (N_18974,N_18676,N_18329);
xor U18975 (N_18975,N_18551,N_18138);
nand U18976 (N_18976,N_18346,N_18187);
nand U18977 (N_18977,N_18207,N_18191);
nor U18978 (N_18978,N_18593,N_18680);
nand U18979 (N_18979,N_18380,N_18368);
or U18980 (N_18980,N_18360,N_18459);
or U18981 (N_18981,N_18229,N_18282);
nor U18982 (N_18982,N_18660,N_18231);
nand U18983 (N_18983,N_18695,N_18319);
or U18984 (N_18984,N_18563,N_18157);
nor U18985 (N_18985,N_18370,N_18359);
and U18986 (N_18986,N_18366,N_18291);
and U18987 (N_18987,N_18645,N_18713);
or U18988 (N_18988,N_18454,N_18162);
xnor U18989 (N_18989,N_18190,N_18236);
nand U18990 (N_18990,N_18226,N_18126);
nor U18991 (N_18991,N_18615,N_18701);
nor U18992 (N_18992,N_18432,N_18650);
nor U18993 (N_18993,N_18383,N_18268);
xnor U18994 (N_18994,N_18488,N_18460);
xor U18995 (N_18995,N_18260,N_18688);
or U18996 (N_18996,N_18155,N_18467);
or U18997 (N_18997,N_18293,N_18375);
nand U18998 (N_18998,N_18724,N_18267);
nand U18999 (N_18999,N_18478,N_18379);
or U19000 (N_19000,N_18347,N_18555);
xnor U19001 (N_19001,N_18344,N_18202);
nor U19002 (N_19002,N_18418,N_18490);
nor U19003 (N_19003,N_18568,N_18748);
or U19004 (N_19004,N_18653,N_18257);
or U19005 (N_19005,N_18463,N_18506);
xor U19006 (N_19006,N_18173,N_18253);
nand U19007 (N_19007,N_18598,N_18629);
or U19008 (N_19008,N_18708,N_18723);
xor U19009 (N_19009,N_18501,N_18456);
or U19010 (N_19010,N_18468,N_18689);
or U19011 (N_19011,N_18528,N_18643);
or U19012 (N_19012,N_18656,N_18621);
nor U19013 (N_19013,N_18556,N_18562);
nand U19014 (N_19014,N_18641,N_18606);
nand U19015 (N_19015,N_18321,N_18413);
or U19016 (N_19016,N_18416,N_18654);
xor U19017 (N_19017,N_18633,N_18619);
or U19018 (N_19018,N_18403,N_18222);
and U19019 (N_19019,N_18429,N_18666);
or U19020 (N_19020,N_18509,N_18535);
nand U19021 (N_19021,N_18693,N_18546);
and U19022 (N_19022,N_18648,N_18664);
xnor U19023 (N_19023,N_18387,N_18536);
xnor U19024 (N_19024,N_18341,N_18227);
xor U19025 (N_19025,N_18486,N_18479);
or U19026 (N_19026,N_18444,N_18729);
and U19027 (N_19027,N_18361,N_18298);
or U19028 (N_19028,N_18570,N_18204);
or U19029 (N_19029,N_18287,N_18271);
nand U19030 (N_19030,N_18544,N_18421);
xor U19031 (N_19031,N_18521,N_18278);
nand U19032 (N_19032,N_18487,N_18587);
xnor U19033 (N_19033,N_18611,N_18560);
nand U19034 (N_19034,N_18134,N_18206);
or U19035 (N_19035,N_18719,N_18692);
or U19036 (N_19036,N_18667,N_18477);
xnor U19037 (N_19037,N_18576,N_18409);
nor U19038 (N_19038,N_18395,N_18400);
nor U19039 (N_19039,N_18550,N_18511);
xor U19040 (N_19040,N_18181,N_18510);
nor U19041 (N_19041,N_18143,N_18518);
or U19042 (N_19042,N_18522,N_18195);
and U19043 (N_19043,N_18661,N_18262);
or U19044 (N_19044,N_18675,N_18200);
xor U19045 (N_19045,N_18365,N_18607);
or U19046 (N_19046,N_18288,N_18626);
xnor U19047 (N_19047,N_18180,N_18150);
nor U19048 (N_19048,N_18655,N_18396);
nand U19049 (N_19049,N_18696,N_18686);
or U19050 (N_19050,N_18540,N_18610);
nor U19051 (N_19051,N_18148,N_18272);
nor U19052 (N_19052,N_18279,N_18537);
nand U19053 (N_19053,N_18295,N_18707);
nand U19054 (N_19054,N_18351,N_18565);
nor U19055 (N_19055,N_18338,N_18310);
nor U19056 (N_19056,N_18441,N_18316);
and U19057 (N_19057,N_18340,N_18388);
and U19058 (N_19058,N_18671,N_18264);
or U19059 (N_19059,N_18557,N_18569);
or U19060 (N_19060,N_18577,N_18183);
xnor U19061 (N_19061,N_18702,N_18443);
xnor U19062 (N_19062,N_18749,N_18660);
or U19063 (N_19063,N_18326,N_18555);
and U19064 (N_19064,N_18733,N_18253);
nor U19065 (N_19065,N_18537,N_18357);
nand U19066 (N_19066,N_18493,N_18332);
and U19067 (N_19067,N_18215,N_18448);
nand U19068 (N_19068,N_18208,N_18495);
xor U19069 (N_19069,N_18580,N_18451);
nand U19070 (N_19070,N_18348,N_18267);
nand U19071 (N_19071,N_18582,N_18366);
xnor U19072 (N_19072,N_18131,N_18471);
and U19073 (N_19073,N_18477,N_18211);
nand U19074 (N_19074,N_18500,N_18610);
nor U19075 (N_19075,N_18583,N_18552);
xnor U19076 (N_19076,N_18728,N_18677);
and U19077 (N_19077,N_18249,N_18422);
nand U19078 (N_19078,N_18480,N_18555);
nor U19079 (N_19079,N_18671,N_18288);
or U19080 (N_19080,N_18737,N_18312);
and U19081 (N_19081,N_18177,N_18208);
nor U19082 (N_19082,N_18635,N_18395);
and U19083 (N_19083,N_18486,N_18574);
or U19084 (N_19084,N_18474,N_18593);
nand U19085 (N_19085,N_18443,N_18496);
nand U19086 (N_19086,N_18451,N_18527);
xor U19087 (N_19087,N_18488,N_18256);
or U19088 (N_19088,N_18481,N_18555);
or U19089 (N_19089,N_18371,N_18564);
or U19090 (N_19090,N_18562,N_18524);
or U19091 (N_19091,N_18622,N_18396);
nor U19092 (N_19092,N_18599,N_18270);
or U19093 (N_19093,N_18171,N_18624);
xnor U19094 (N_19094,N_18428,N_18341);
and U19095 (N_19095,N_18597,N_18437);
and U19096 (N_19096,N_18265,N_18594);
nor U19097 (N_19097,N_18733,N_18594);
nand U19098 (N_19098,N_18595,N_18363);
nor U19099 (N_19099,N_18376,N_18478);
or U19100 (N_19100,N_18537,N_18624);
and U19101 (N_19101,N_18523,N_18354);
nand U19102 (N_19102,N_18644,N_18546);
or U19103 (N_19103,N_18552,N_18255);
nand U19104 (N_19104,N_18724,N_18563);
xor U19105 (N_19105,N_18543,N_18353);
or U19106 (N_19106,N_18438,N_18341);
and U19107 (N_19107,N_18225,N_18749);
xor U19108 (N_19108,N_18246,N_18333);
nand U19109 (N_19109,N_18546,N_18376);
or U19110 (N_19110,N_18537,N_18633);
or U19111 (N_19111,N_18362,N_18422);
or U19112 (N_19112,N_18474,N_18696);
or U19113 (N_19113,N_18541,N_18516);
and U19114 (N_19114,N_18151,N_18138);
xnor U19115 (N_19115,N_18144,N_18701);
or U19116 (N_19116,N_18428,N_18321);
nor U19117 (N_19117,N_18524,N_18252);
or U19118 (N_19118,N_18232,N_18436);
or U19119 (N_19119,N_18646,N_18602);
xor U19120 (N_19120,N_18595,N_18171);
nor U19121 (N_19121,N_18251,N_18166);
and U19122 (N_19122,N_18551,N_18262);
nand U19123 (N_19123,N_18530,N_18369);
nor U19124 (N_19124,N_18361,N_18367);
xnor U19125 (N_19125,N_18354,N_18357);
or U19126 (N_19126,N_18581,N_18742);
nand U19127 (N_19127,N_18576,N_18222);
nand U19128 (N_19128,N_18674,N_18384);
nand U19129 (N_19129,N_18323,N_18596);
nand U19130 (N_19130,N_18625,N_18277);
or U19131 (N_19131,N_18605,N_18207);
xnor U19132 (N_19132,N_18255,N_18436);
nor U19133 (N_19133,N_18362,N_18455);
nand U19134 (N_19134,N_18283,N_18154);
nor U19135 (N_19135,N_18132,N_18314);
nor U19136 (N_19136,N_18184,N_18620);
nor U19137 (N_19137,N_18380,N_18524);
nand U19138 (N_19138,N_18663,N_18214);
nor U19139 (N_19139,N_18737,N_18169);
xnor U19140 (N_19140,N_18417,N_18667);
xor U19141 (N_19141,N_18666,N_18369);
nor U19142 (N_19142,N_18190,N_18349);
or U19143 (N_19143,N_18152,N_18603);
nand U19144 (N_19144,N_18459,N_18711);
nand U19145 (N_19145,N_18462,N_18540);
or U19146 (N_19146,N_18271,N_18285);
nand U19147 (N_19147,N_18520,N_18300);
nor U19148 (N_19148,N_18724,N_18411);
nor U19149 (N_19149,N_18675,N_18399);
nor U19150 (N_19150,N_18263,N_18719);
nor U19151 (N_19151,N_18230,N_18596);
and U19152 (N_19152,N_18368,N_18291);
nor U19153 (N_19153,N_18168,N_18238);
or U19154 (N_19154,N_18564,N_18454);
xnor U19155 (N_19155,N_18567,N_18459);
or U19156 (N_19156,N_18295,N_18294);
and U19157 (N_19157,N_18305,N_18574);
xor U19158 (N_19158,N_18602,N_18307);
and U19159 (N_19159,N_18647,N_18440);
nor U19160 (N_19160,N_18336,N_18508);
or U19161 (N_19161,N_18290,N_18512);
xnor U19162 (N_19162,N_18251,N_18619);
and U19163 (N_19163,N_18293,N_18514);
nor U19164 (N_19164,N_18462,N_18180);
nand U19165 (N_19165,N_18336,N_18277);
and U19166 (N_19166,N_18574,N_18618);
nor U19167 (N_19167,N_18397,N_18261);
and U19168 (N_19168,N_18601,N_18196);
xnor U19169 (N_19169,N_18257,N_18742);
or U19170 (N_19170,N_18176,N_18431);
or U19171 (N_19171,N_18291,N_18654);
xor U19172 (N_19172,N_18211,N_18618);
or U19173 (N_19173,N_18280,N_18171);
and U19174 (N_19174,N_18179,N_18214);
nor U19175 (N_19175,N_18600,N_18362);
xnor U19176 (N_19176,N_18358,N_18395);
nor U19177 (N_19177,N_18717,N_18579);
or U19178 (N_19178,N_18349,N_18571);
xor U19179 (N_19179,N_18181,N_18679);
or U19180 (N_19180,N_18279,N_18356);
xnor U19181 (N_19181,N_18699,N_18722);
and U19182 (N_19182,N_18295,N_18610);
and U19183 (N_19183,N_18651,N_18703);
or U19184 (N_19184,N_18528,N_18149);
nor U19185 (N_19185,N_18242,N_18229);
and U19186 (N_19186,N_18696,N_18495);
nor U19187 (N_19187,N_18456,N_18653);
nor U19188 (N_19188,N_18186,N_18134);
or U19189 (N_19189,N_18716,N_18622);
xnor U19190 (N_19190,N_18559,N_18160);
xor U19191 (N_19191,N_18699,N_18731);
and U19192 (N_19192,N_18321,N_18640);
nand U19193 (N_19193,N_18266,N_18241);
nor U19194 (N_19194,N_18562,N_18618);
nor U19195 (N_19195,N_18725,N_18126);
xnor U19196 (N_19196,N_18281,N_18593);
nand U19197 (N_19197,N_18677,N_18419);
nand U19198 (N_19198,N_18187,N_18333);
nand U19199 (N_19199,N_18590,N_18699);
nor U19200 (N_19200,N_18376,N_18351);
nor U19201 (N_19201,N_18521,N_18264);
and U19202 (N_19202,N_18500,N_18657);
nand U19203 (N_19203,N_18256,N_18739);
and U19204 (N_19204,N_18542,N_18432);
or U19205 (N_19205,N_18707,N_18588);
xnor U19206 (N_19206,N_18602,N_18464);
nand U19207 (N_19207,N_18478,N_18517);
and U19208 (N_19208,N_18455,N_18488);
or U19209 (N_19209,N_18226,N_18426);
nor U19210 (N_19210,N_18476,N_18729);
nand U19211 (N_19211,N_18289,N_18432);
and U19212 (N_19212,N_18535,N_18662);
xor U19213 (N_19213,N_18681,N_18176);
or U19214 (N_19214,N_18699,N_18324);
or U19215 (N_19215,N_18283,N_18245);
nor U19216 (N_19216,N_18241,N_18636);
xor U19217 (N_19217,N_18413,N_18175);
and U19218 (N_19218,N_18294,N_18292);
nor U19219 (N_19219,N_18617,N_18196);
nand U19220 (N_19220,N_18193,N_18661);
nor U19221 (N_19221,N_18433,N_18475);
xnor U19222 (N_19222,N_18276,N_18584);
or U19223 (N_19223,N_18722,N_18719);
and U19224 (N_19224,N_18386,N_18682);
nand U19225 (N_19225,N_18187,N_18386);
nor U19226 (N_19226,N_18587,N_18669);
or U19227 (N_19227,N_18310,N_18382);
nor U19228 (N_19228,N_18355,N_18594);
and U19229 (N_19229,N_18622,N_18282);
or U19230 (N_19230,N_18423,N_18635);
xor U19231 (N_19231,N_18478,N_18185);
or U19232 (N_19232,N_18692,N_18625);
or U19233 (N_19233,N_18411,N_18288);
or U19234 (N_19234,N_18249,N_18720);
and U19235 (N_19235,N_18274,N_18719);
and U19236 (N_19236,N_18689,N_18225);
nor U19237 (N_19237,N_18449,N_18204);
xor U19238 (N_19238,N_18189,N_18297);
or U19239 (N_19239,N_18303,N_18240);
and U19240 (N_19240,N_18449,N_18476);
or U19241 (N_19241,N_18166,N_18428);
xnor U19242 (N_19242,N_18445,N_18333);
xor U19243 (N_19243,N_18359,N_18656);
or U19244 (N_19244,N_18487,N_18315);
xnor U19245 (N_19245,N_18291,N_18441);
xnor U19246 (N_19246,N_18261,N_18601);
and U19247 (N_19247,N_18184,N_18494);
and U19248 (N_19248,N_18613,N_18411);
nor U19249 (N_19249,N_18573,N_18292);
xor U19250 (N_19250,N_18358,N_18146);
nand U19251 (N_19251,N_18405,N_18199);
nor U19252 (N_19252,N_18176,N_18365);
or U19253 (N_19253,N_18183,N_18429);
nor U19254 (N_19254,N_18549,N_18565);
nor U19255 (N_19255,N_18457,N_18348);
or U19256 (N_19256,N_18304,N_18741);
and U19257 (N_19257,N_18673,N_18352);
nor U19258 (N_19258,N_18687,N_18653);
nor U19259 (N_19259,N_18150,N_18547);
nor U19260 (N_19260,N_18465,N_18367);
nor U19261 (N_19261,N_18420,N_18489);
nand U19262 (N_19262,N_18363,N_18738);
nand U19263 (N_19263,N_18307,N_18341);
nor U19264 (N_19264,N_18570,N_18461);
nor U19265 (N_19265,N_18738,N_18283);
nand U19266 (N_19266,N_18617,N_18475);
or U19267 (N_19267,N_18462,N_18333);
nor U19268 (N_19268,N_18282,N_18249);
or U19269 (N_19269,N_18187,N_18127);
xnor U19270 (N_19270,N_18493,N_18336);
or U19271 (N_19271,N_18586,N_18349);
xnor U19272 (N_19272,N_18673,N_18427);
nor U19273 (N_19273,N_18572,N_18318);
or U19274 (N_19274,N_18355,N_18283);
or U19275 (N_19275,N_18687,N_18334);
or U19276 (N_19276,N_18557,N_18610);
and U19277 (N_19277,N_18346,N_18569);
or U19278 (N_19278,N_18347,N_18418);
or U19279 (N_19279,N_18585,N_18289);
or U19280 (N_19280,N_18507,N_18573);
xnor U19281 (N_19281,N_18543,N_18513);
nor U19282 (N_19282,N_18202,N_18515);
nand U19283 (N_19283,N_18545,N_18425);
nand U19284 (N_19284,N_18352,N_18528);
nand U19285 (N_19285,N_18478,N_18234);
nor U19286 (N_19286,N_18664,N_18608);
xnor U19287 (N_19287,N_18316,N_18331);
and U19288 (N_19288,N_18146,N_18629);
or U19289 (N_19289,N_18636,N_18471);
and U19290 (N_19290,N_18471,N_18385);
xnor U19291 (N_19291,N_18561,N_18702);
nand U19292 (N_19292,N_18366,N_18680);
xnor U19293 (N_19293,N_18341,N_18126);
or U19294 (N_19294,N_18340,N_18491);
and U19295 (N_19295,N_18453,N_18735);
or U19296 (N_19296,N_18705,N_18529);
and U19297 (N_19297,N_18485,N_18358);
nor U19298 (N_19298,N_18685,N_18460);
nand U19299 (N_19299,N_18202,N_18474);
nand U19300 (N_19300,N_18638,N_18527);
xnor U19301 (N_19301,N_18540,N_18154);
nand U19302 (N_19302,N_18173,N_18337);
xnor U19303 (N_19303,N_18630,N_18181);
and U19304 (N_19304,N_18329,N_18303);
nand U19305 (N_19305,N_18154,N_18233);
nand U19306 (N_19306,N_18407,N_18291);
and U19307 (N_19307,N_18669,N_18447);
or U19308 (N_19308,N_18213,N_18608);
and U19309 (N_19309,N_18199,N_18134);
or U19310 (N_19310,N_18230,N_18733);
xnor U19311 (N_19311,N_18482,N_18722);
or U19312 (N_19312,N_18187,N_18240);
or U19313 (N_19313,N_18257,N_18150);
and U19314 (N_19314,N_18288,N_18577);
xor U19315 (N_19315,N_18285,N_18745);
and U19316 (N_19316,N_18749,N_18578);
xor U19317 (N_19317,N_18148,N_18444);
nand U19318 (N_19318,N_18298,N_18715);
nor U19319 (N_19319,N_18569,N_18375);
xor U19320 (N_19320,N_18642,N_18714);
nor U19321 (N_19321,N_18149,N_18723);
nand U19322 (N_19322,N_18319,N_18231);
xnor U19323 (N_19323,N_18363,N_18502);
nor U19324 (N_19324,N_18398,N_18228);
nand U19325 (N_19325,N_18142,N_18411);
xnor U19326 (N_19326,N_18629,N_18371);
nand U19327 (N_19327,N_18443,N_18745);
or U19328 (N_19328,N_18505,N_18578);
xnor U19329 (N_19329,N_18683,N_18246);
or U19330 (N_19330,N_18529,N_18272);
and U19331 (N_19331,N_18478,N_18552);
nand U19332 (N_19332,N_18736,N_18710);
nor U19333 (N_19333,N_18141,N_18463);
nand U19334 (N_19334,N_18163,N_18563);
nand U19335 (N_19335,N_18581,N_18384);
or U19336 (N_19336,N_18724,N_18389);
xor U19337 (N_19337,N_18650,N_18444);
nand U19338 (N_19338,N_18411,N_18341);
nand U19339 (N_19339,N_18310,N_18146);
and U19340 (N_19340,N_18221,N_18196);
nor U19341 (N_19341,N_18292,N_18610);
nor U19342 (N_19342,N_18263,N_18176);
nor U19343 (N_19343,N_18626,N_18454);
or U19344 (N_19344,N_18639,N_18540);
nand U19345 (N_19345,N_18743,N_18288);
nor U19346 (N_19346,N_18328,N_18372);
and U19347 (N_19347,N_18135,N_18338);
nand U19348 (N_19348,N_18562,N_18209);
nor U19349 (N_19349,N_18722,N_18647);
and U19350 (N_19350,N_18532,N_18632);
and U19351 (N_19351,N_18596,N_18357);
xnor U19352 (N_19352,N_18173,N_18175);
xor U19353 (N_19353,N_18281,N_18272);
and U19354 (N_19354,N_18467,N_18663);
or U19355 (N_19355,N_18403,N_18589);
nand U19356 (N_19356,N_18516,N_18387);
nand U19357 (N_19357,N_18540,N_18680);
or U19358 (N_19358,N_18345,N_18501);
xnor U19359 (N_19359,N_18242,N_18279);
or U19360 (N_19360,N_18594,N_18683);
nand U19361 (N_19361,N_18190,N_18166);
xor U19362 (N_19362,N_18595,N_18576);
and U19363 (N_19363,N_18299,N_18385);
and U19364 (N_19364,N_18265,N_18744);
nand U19365 (N_19365,N_18635,N_18499);
and U19366 (N_19366,N_18701,N_18162);
and U19367 (N_19367,N_18285,N_18267);
xnor U19368 (N_19368,N_18640,N_18393);
nor U19369 (N_19369,N_18366,N_18209);
nor U19370 (N_19370,N_18453,N_18476);
or U19371 (N_19371,N_18537,N_18559);
and U19372 (N_19372,N_18526,N_18300);
or U19373 (N_19373,N_18546,N_18170);
xnor U19374 (N_19374,N_18389,N_18291);
nand U19375 (N_19375,N_19278,N_18970);
nand U19376 (N_19376,N_19114,N_18884);
or U19377 (N_19377,N_18929,N_19356);
xor U19378 (N_19378,N_19218,N_18973);
nor U19379 (N_19379,N_18943,N_18924);
nand U19380 (N_19380,N_18855,N_19062);
and U19381 (N_19381,N_18859,N_19214);
and U19382 (N_19382,N_18996,N_19051);
or U19383 (N_19383,N_19290,N_19272);
and U19384 (N_19384,N_18875,N_19192);
xor U19385 (N_19385,N_19220,N_19074);
xnor U19386 (N_19386,N_18988,N_19287);
or U19387 (N_19387,N_18945,N_19171);
nand U19388 (N_19388,N_19132,N_19135);
nor U19389 (N_19389,N_18926,N_19265);
or U19390 (N_19390,N_19305,N_19107);
xor U19391 (N_19391,N_19008,N_18785);
xnor U19392 (N_19392,N_18967,N_19322);
nand U19393 (N_19393,N_19295,N_18830);
xnor U19394 (N_19394,N_18920,N_19369);
nand U19395 (N_19395,N_19228,N_18824);
xnor U19396 (N_19396,N_18754,N_19089);
or U19397 (N_19397,N_18962,N_19041);
nor U19398 (N_19398,N_19108,N_19053);
nand U19399 (N_19399,N_18896,N_18792);
nand U19400 (N_19400,N_18872,N_19082);
nor U19401 (N_19401,N_18815,N_19020);
and U19402 (N_19402,N_19345,N_19194);
and U19403 (N_19403,N_19170,N_19306);
and U19404 (N_19404,N_19307,N_18771);
nand U19405 (N_19405,N_18981,N_19365);
nand U19406 (N_19406,N_18763,N_18964);
and U19407 (N_19407,N_19124,N_18874);
nand U19408 (N_19408,N_18909,N_19248);
nor U19409 (N_19409,N_19260,N_18858);
or U19410 (N_19410,N_19340,N_18787);
and U19411 (N_19411,N_18805,N_19167);
and U19412 (N_19412,N_18833,N_19316);
nand U19413 (N_19413,N_19002,N_19269);
nand U19414 (N_19414,N_18794,N_19252);
nor U19415 (N_19415,N_19088,N_18903);
nand U19416 (N_19416,N_19054,N_18880);
nor U19417 (N_19417,N_18827,N_19156);
nor U19418 (N_19418,N_18977,N_18760);
xnor U19419 (N_19419,N_19077,N_18863);
nor U19420 (N_19420,N_19099,N_19208);
xnor U19421 (N_19421,N_19258,N_18915);
nor U19422 (N_19422,N_19025,N_19188);
nand U19423 (N_19423,N_19043,N_18819);
xor U19424 (N_19424,N_19288,N_19106);
xnor U19425 (N_19425,N_19183,N_18839);
nand U19426 (N_19426,N_18759,N_18906);
xnor U19427 (N_19427,N_18832,N_19354);
nand U19428 (N_19428,N_18914,N_19215);
nor U19429 (N_19429,N_19009,N_19297);
or U19430 (N_19430,N_19312,N_19111);
xnor U19431 (N_19431,N_19225,N_18940);
nor U19432 (N_19432,N_19174,N_18756);
nor U19433 (N_19433,N_18841,N_19056);
nand U19434 (N_19434,N_19035,N_19261);
and U19435 (N_19435,N_19187,N_19096);
and U19436 (N_19436,N_19285,N_18922);
and U19437 (N_19437,N_19245,N_18993);
nor U19438 (N_19438,N_18971,N_19205);
nand U19439 (N_19439,N_18803,N_19332);
xor U19440 (N_19440,N_18991,N_18867);
xor U19441 (N_19441,N_19113,N_19121);
xor U19442 (N_19442,N_19159,N_19022);
and U19443 (N_19443,N_18857,N_19267);
or U19444 (N_19444,N_19204,N_18976);
and U19445 (N_19445,N_18910,N_19224);
xnor U19446 (N_19446,N_18823,N_19296);
nor U19447 (N_19447,N_18776,N_18947);
and U19448 (N_19448,N_18844,N_18817);
nand U19449 (N_19449,N_19370,N_19199);
nand U19450 (N_19450,N_19076,N_19353);
or U19451 (N_19451,N_18790,N_19223);
nand U19452 (N_19452,N_19263,N_19133);
and U19453 (N_19453,N_19085,N_19317);
nand U19454 (N_19454,N_19029,N_18797);
or U19455 (N_19455,N_19289,N_19055);
xnor U19456 (N_19456,N_18835,N_18985);
or U19457 (N_19457,N_18886,N_18974);
nor U19458 (N_19458,N_19037,N_19311);
xnor U19459 (N_19459,N_19068,N_19105);
xnor U19460 (N_19460,N_19014,N_19044);
or U19461 (N_19461,N_19367,N_19255);
nor U19462 (N_19462,N_18795,N_19018);
or U19463 (N_19463,N_19348,N_18767);
nor U19464 (N_19464,N_18818,N_19264);
or U19465 (N_19465,N_19058,N_19362);
and U19466 (N_19466,N_18758,N_18798);
nand U19467 (N_19467,N_19244,N_18762);
nand U19468 (N_19468,N_19091,N_19197);
xnor U19469 (N_19469,N_18912,N_18822);
and U19470 (N_19470,N_19090,N_18949);
nor U19471 (N_19471,N_18921,N_19161);
and U19472 (N_19472,N_18897,N_19160);
nand U19473 (N_19473,N_19072,N_18898);
nor U19474 (N_19474,N_18948,N_19122);
and U19475 (N_19475,N_19097,N_19326);
or U19476 (N_19476,N_19176,N_19047);
nand U19477 (N_19477,N_19003,N_19284);
xor U19478 (N_19478,N_18881,N_19095);
nand U19479 (N_19479,N_18957,N_19011);
xor U19480 (N_19480,N_18895,N_19268);
xor U19481 (N_19481,N_19092,N_18804);
and U19482 (N_19482,N_19064,N_19331);
nand U19483 (N_19483,N_18999,N_18994);
nand U19484 (N_19484,N_18821,N_18975);
xnor U19485 (N_19485,N_19172,N_18944);
xnor U19486 (N_19486,N_19222,N_18904);
and U19487 (N_19487,N_19158,N_19241);
nand U19488 (N_19488,N_19327,N_19190);
nor U19489 (N_19489,N_18869,N_19315);
nor U19490 (N_19490,N_19127,N_19182);
and U19491 (N_19491,N_19350,N_18887);
or U19492 (N_19492,N_19237,N_19007);
or U19493 (N_19493,N_19173,N_19254);
and U19494 (N_19494,N_19004,N_18969);
xnor U19495 (N_19495,N_19137,N_19328);
and U19496 (N_19496,N_19081,N_19017);
xnor U19497 (N_19497,N_18955,N_18780);
nand U19498 (N_19498,N_18845,N_19103);
nor U19499 (N_19499,N_19116,N_19325);
and U19500 (N_19500,N_18876,N_19136);
nand U19501 (N_19501,N_18885,N_18960);
xnor U19502 (N_19502,N_19262,N_18764);
and U19503 (N_19503,N_19334,N_18978);
nor U19504 (N_19504,N_18772,N_19293);
or U19505 (N_19505,N_18865,N_18984);
nand U19506 (N_19506,N_18963,N_18765);
nand U19507 (N_19507,N_18983,N_18807);
nor U19508 (N_19508,N_19084,N_19238);
and U19509 (N_19509,N_19200,N_19217);
nor U19510 (N_19510,N_19213,N_18861);
or U19511 (N_19511,N_18786,N_19071);
nor U19512 (N_19512,N_19080,N_19109);
xnor U19513 (N_19513,N_18900,N_18927);
xnor U19514 (N_19514,N_19175,N_19128);
and U19515 (N_19515,N_19368,N_19164);
or U19516 (N_19516,N_19335,N_19276);
or U19517 (N_19517,N_19216,N_18777);
xor U19518 (N_19518,N_18843,N_19229);
and U19519 (N_19519,N_18752,N_18916);
and U19520 (N_19520,N_19141,N_19036);
nor U19521 (N_19521,N_19015,N_19112);
nand U19522 (N_19522,N_18814,N_19052);
and U19523 (N_19523,N_19010,N_19363);
and U19524 (N_19524,N_19023,N_18837);
nor U19525 (N_19525,N_19125,N_19360);
xor U19526 (N_19526,N_19211,N_18751);
or U19527 (N_19527,N_19243,N_19361);
or U19528 (N_19528,N_18800,N_19079);
nand U19529 (N_19529,N_19166,N_18851);
nand U19530 (N_19530,N_18862,N_19155);
or U19531 (N_19531,N_19016,N_18965);
nand U19532 (N_19532,N_19130,N_19343);
xor U19533 (N_19533,N_18781,N_19337);
xor U19534 (N_19534,N_19249,N_19157);
and U19535 (N_19535,N_19239,N_18968);
nor U19536 (N_19536,N_18778,N_18826);
nor U19537 (N_19537,N_19061,N_18879);
and U19538 (N_19538,N_19299,N_18773);
nor U19539 (N_19539,N_18882,N_19012);
nor U19540 (N_19540,N_19318,N_18933);
xnor U19541 (N_19541,N_19291,N_18799);
xnor U19542 (N_19542,N_19232,N_19338);
xnor U19543 (N_19543,N_19021,N_18810);
nand U19544 (N_19544,N_19031,N_18766);
or U19545 (N_19545,N_19026,N_18919);
xor U19546 (N_19546,N_18989,N_19153);
nand U19547 (N_19547,N_18873,N_19069);
and U19548 (N_19548,N_18825,N_19013);
nand U19549 (N_19549,N_19303,N_19046);
xnor U19550 (N_19550,N_19301,N_19186);
and U19551 (N_19551,N_19351,N_19027);
xor U19552 (N_19552,N_18834,N_18959);
and U19553 (N_19553,N_19134,N_19000);
nand U19554 (N_19554,N_19319,N_18925);
xor U19555 (N_19555,N_19251,N_18936);
xnor U19556 (N_19556,N_19352,N_18911);
nor U19557 (N_19557,N_19034,N_19206);
nor U19558 (N_19558,N_18990,N_18793);
nand U19559 (N_19559,N_18811,N_19179);
nor U19560 (N_19560,N_18901,N_19330);
xnor U19561 (N_19561,N_18998,N_18812);
xnor U19562 (N_19562,N_19165,N_19118);
nand U19563 (N_19563,N_19101,N_19282);
nor U19564 (N_19564,N_18779,N_18980);
xor U19565 (N_19565,N_19304,N_19250);
nor U19566 (N_19566,N_19094,N_19341);
nand U19567 (N_19567,N_19185,N_19049);
nand U19568 (N_19568,N_19372,N_19087);
and U19569 (N_19569,N_19048,N_18934);
nand U19570 (N_19570,N_18997,N_18950);
and U19571 (N_19571,N_19280,N_18956);
xnor U19572 (N_19572,N_18995,N_18789);
nand U19573 (N_19573,N_19032,N_19227);
and U19574 (N_19574,N_18768,N_19024);
nor U19575 (N_19575,N_19298,N_18761);
xnor U19576 (N_19576,N_19057,N_18979);
nor U19577 (N_19577,N_19279,N_19309);
xnor U19578 (N_19578,N_19207,N_19181);
nand U19579 (N_19579,N_19039,N_18961);
xor U19580 (N_19580,N_19203,N_19073);
nand U19581 (N_19581,N_18918,N_19120);
nor U19582 (N_19582,N_18937,N_18774);
and U19583 (N_19583,N_19163,N_19075);
and U19584 (N_19584,N_19067,N_18958);
and U19585 (N_19585,N_18923,N_19152);
or U19586 (N_19586,N_19346,N_18842);
xnor U19587 (N_19587,N_18870,N_19143);
nand U19588 (N_19588,N_19275,N_19257);
nand U19589 (N_19589,N_18890,N_19006);
nand U19590 (N_19590,N_18899,N_19247);
or U19591 (N_19591,N_18770,N_18853);
nand U19592 (N_19592,N_18808,N_18954);
and U19593 (N_19593,N_19151,N_19235);
xor U19594 (N_19594,N_19310,N_19313);
and U19595 (N_19595,N_19050,N_19321);
or U19596 (N_19596,N_19119,N_18828);
nor U19597 (N_19597,N_18953,N_18788);
xor U19598 (N_19598,N_19139,N_19274);
xnor U19599 (N_19599,N_18883,N_19283);
and U19600 (N_19600,N_18860,N_19131);
and U19601 (N_19601,N_18782,N_19202);
and U19602 (N_19602,N_18769,N_19195);
nand U19603 (N_19603,N_19040,N_18848);
or U19604 (N_19604,N_18917,N_19019);
xor U19605 (N_19605,N_19102,N_19256);
nand U19606 (N_19606,N_19140,N_18753);
nor U19607 (N_19607,N_19129,N_18840);
nand U19608 (N_19608,N_19300,N_18829);
and U19609 (N_19609,N_18966,N_19115);
nand U19610 (N_19610,N_18932,N_18907);
and U19611 (N_19611,N_18849,N_19246);
or U19612 (N_19612,N_19148,N_19138);
nand U19613 (N_19613,N_18783,N_19083);
nor U19614 (N_19614,N_19098,N_19221);
or U19615 (N_19615,N_18941,N_19142);
xor U19616 (N_19616,N_19271,N_18942);
xor U19617 (N_19617,N_19357,N_19201);
nand U19618 (N_19618,N_19323,N_19294);
nor U19619 (N_19619,N_19374,N_19308);
or U19620 (N_19620,N_18856,N_18935);
and U19621 (N_19621,N_18852,N_19028);
nor U19622 (N_19622,N_19324,N_19344);
nor U19623 (N_19623,N_18972,N_18755);
nor U19624 (N_19624,N_19038,N_19233);
nand U19625 (N_19625,N_19066,N_19302);
nor U19626 (N_19626,N_18864,N_18987);
nor U19627 (N_19627,N_19371,N_19292);
or U19628 (N_19628,N_18928,N_19231);
xor U19629 (N_19629,N_19196,N_19336);
xnor U19630 (N_19630,N_19033,N_18784);
nor U19631 (N_19631,N_19286,N_18775);
nor U19632 (N_19632,N_18847,N_19329);
xnor U19633 (N_19633,N_18952,N_18992);
nor U19634 (N_19634,N_18913,N_19104);
nand U19635 (N_19635,N_19147,N_18877);
nor U19636 (N_19636,N_19001,N_18854);
and U19637 (N_19637,N_19193,N_19355);
nor U19638 (N_19638,N_19314,N_18893);
xnor U19639 (N_19639,N_19242,N_19065);
or U19640 (N_19640,N_19191,N_19059);
xor U19641 (N_19641,N_18938,N_18878);
or U19642 (N_19642,N_19266,N_18946);
xor U19643 (N_19643,N_19184,N_19212);
nand U19644 (N_19644,N_19117,N_19273);
xnor U19645 (N_19645,N_18820,N_19045);
xor U19646 (N_19646,N_18894,N_19126);
nor U19647 (N_19647,N_19042,N_19270);
nor U19648 (N_19648,N_18796,N_19146);
and U19649 (N_19649,N_19178,N_19198);
or U19650 (N_19650,N_19240,N_19277);
or U19651 (N_19651,N_19253,N_18801);
or U19652 (N_19652,N_18982,N_18816);
nor U19653 (N_19653,N_18888,N_19373);
nand U19654 (N_19654,N_19086,N_18930);
nor U19655 (N_19655,N_19219,N_19230);
nor U19656 (N_19656,N_19359,N_19030);
and U19657 (N_19657,N_18939,N_19060);
and U19658 (N_19658,N_18850,N_18838);
or U19659 (N_19659,N_18750,N_19123);
nand U19660 (N_19660,N_18846,N_19168);
nor U19661 (N_19661,N_19364,N_19149);
and U19662 (N_19662,N_19005,N_18931);
and U19663 (N_19663,N_19320,N_19144);
nand U19664 (N_19664,N_19339,N_18892);
nor U19665 (N_19665,N_19078,N_18802);
and U19666 (N_19666,N_18836,N_19234);
or U19667 (N_19667,N_19189,N_19366);
nand U19668 (N_19668,N_19347,N_18868);
xnor U19669 (N_19669,N_19210,N_18866);
or U19670 (N_19670,N_19063,N_18813);
nor U19671 (N_19671,N_18831,N_19110);
xnor U19672 (N_19672,N_18809,N_19180);
nor U19673 (N_19673,N_18871,N_19358);
nand U19674 (N_19674,N_19333,N_19281);
or U19675 (N_19675,N_19093,N_18905);
and U19676 (N_19676,N_18908,N_19177);
nor U19677 (N_19677,N_18806,N_19236);
or U19678 (N_19678,N_18891,N_19150);
nor U19679 (N_19679,N_19226,N_19145);
nor U19680 (N_19680,N_19169,N_18902);
or U19681 (N_19681,N_19100,N_19070);
xor U19682 (N_19682,N_19154,N_19209);
nand U19683 (N_19683,N_18757,N_18986);
and U19684 (N_19684,N_19342,N_19349);
xnor U19685 (N_19685,N_19259,N_18889);
nand U19686 (N_19686,N_18951,N_18791);
xnor U19687 (N_19687,N_19162,N_18806);
nor U19688 (N_19688,N_19069,N_19227);
nor U19689 (N_19689,N_18936,N_18754);
or U19690 (N_19690,N_19359,N_18892);
xnor U19691 (N_19691,N_19054,N_18976);
xor U19692 (N_19692,N_18799,N_19120);
nand U19693 (N_19693,N_19030,N_19334);
nor U19694 (N_19694,N_18754,N_19139);
nor U19695 (N_19695,N_19332,N_19142);
nor U19696 (N_19696,N_18828,N_19146);
xor U19697 (N_19697,N_19047,N_19149);
and U19698 (N_19698,N_19108,N_19004);
nand U19699 (N_19699,N_19030,N_19323);
nor U19700 (N_19700,N_19018,N_18772);
or U19701 (N_19701,N_18781,N_19262);
xnor U19702 (N_19702,N_19286,N_19147);
and U19703 (N_19703,N_19072,N_19057);
and U19704 (N_19704,N_18970,N_19102);
nand U19705 (N_19705,N_19073,N_18887);
and U19706 (N_19706,N_18889,N_19221);
or U19707 (N_19707,N_18957,N_19093);
and U19708 (N_19708,N_18939,N_19350);
nand U19709 (N_19709,N_18806,N_19071);
nand U19710 (N_19710,N_19211,N_19069);
nand U19711 (N_19711,N_19277,N_19095);
nor U19712 (N_19712,N_18874,N_18802);
or U19713 (N_19713,N_18830,N_19149);
or U19714 (N_19714,N_19279,N_19193);
or U19715 (N_19715,N_18939,N_19334);
or U19716 (N_19716,N_19340,N_18956);
nand U19717 (N_19717,N_19133,N_19246);
nor U19718 (N_19718,N_19042,N_18983);
and U19719 (N_19719,N_19199,N_18894);
or U19720 (N_19720,N_19021,N_19257);
xnor U19721 (N_19721,N_19310,N_18996);
and U19722 (N_19722,N_19116,N_18910);
or U19723 (N_19723,N_19176,N_19230);
nand U19724 (N_19724,N_19366,N_19239);
or U19725 (N_19725,N_19068,N_18933);
xnor U19726 (N_19726,N_18811,N_18879);
or U19727 (N_19727,N_18997,N_18878);
nand U19728 (N_19728,N_18868,N_18829);
xnor U19729 (N_19729,N_18923,N_18973);
xor U19730 (N_19730,N_18858,N_19347);
or U19731 (N_19731,N_18987,N_19066);
and U19732 (N_19732,N_19211,N_19173);
and U19733 (N_19733,N_18988,N_18823);
nand U19734 (N_19734,N_19168,N_18764);
or U19735 (N_19735,N_19071,N_19061);
or U19736 (N_19736,N_19174,N_19054);
nand U19737 (N_19737,N_19123,N_18876);
nand U19738 (N_19738,N_18791,N_18981);
and U19739 (N_19739,N_18848,N_18787);
nor U19740 (N_19740,N_18934,N_19050);
nor U19741 (N_19741,N_18926,N_18786);
or U19742 (N_19742,N_19131,N_18893);
or U19743 (N_19743,N_19319,N_18932);
or U19744 (N_19744,N_19034,N_19327);
nor U19745 (N_19745,N_18800,N_19363);
and U19746 (N_19746,N_19292,N_18888);
nor U19747 (N_19747,N_19195,N_19340);
xor U19748 (N_19748,N_18896,N_19305);
or U19749 (N_19749,N_19311,N_19166);
nor U19750 (N_19750,N_19343,N_19066);
xnor U19751 (N_19751,N_19065,N_18934);
xor U19752 (N_19752,N_19313,N_18805);
xor U19753 (N_19753,N_18925,N_19169);
nand U19754 (N_19754,N_18944,N_18995);
nor U19755 (N_19755,N_19023,N_19124);
xor U19756 (N_19756,N_19023,N_18960);
nand U19757 (N_19757,N_19271,N_18988);
and U19758 (N_19758,N_18809,N_19220);
nor U19759 (N_19759,N_18944,N_18813);
nand U19760 (N_19760,N_19154,N_19242);
or U19761 (N_19761,N_19034,N_19277);
or U19762 (N_19762,N_18798,N_18913);
nand U19763 (N_19763,N_18836,N_18956);
or U19764 (N_19764,N_18865,N_18795);
nand U19765 (N_19765,N_19006,N_19362);
xor U19766 (N_19766,N_19047,N_18886);
and U19767 (N_19767,N_19217,N_18880);
nand U19768 (N_19768,N_19188,N_19058);
nand U19769 (N_19769,N_18968,N_19170);
xor U19770 (N_19770,N_18948,N_19363);
nand U19771 (N_19771,N_19153,N_18983);
or U19772 (N_19772,N_19103,N_18944);
and U19773 (N_19773,N_19295,N_19344);
nand U19774 (N_19774,N_19266,N_19115);
or U19775 (N_19775,N_19279,N_19159);
xor U19776 (N_19776,N_18872,N_19321);
nor U19777 (N_19777,N_19242,N_19223);
nor U19778 (N_19778,N_19067,N_19253);
nand U19779 (N_19779,N_19256,N_18882);
nor U19780 (N_19780,N_19248,N_19372);
nand U19781 (N_19781,N_18781,N_19180);
and U19782 (N_19782,N_19342,N_19218);
nand U19783 (N_19783,N_19080,N_19061);
or U19784 (N_19784,N_18858,N_18835);
and U19785 (N_19785,N_19096,N_19344);
or U19786 (N_19786,N_19296,N_18984);
or U19787 (N_19787,N_18926,N_18989);
xor U19788 (N_19788,N_18971,N_19135);
xnor U19789 (N_19789,N_19157,N_18959);
xnor U19790 (N_19790,N_18906,N_19124);
or U19791 (N_19791,N_19371,N_18942);
xnor U19792 (N_19792,N_19142,N_19233);
nor U19793 (N_19793,N_19236,N_18851);
or U19794 (N_19794,N_19267,N_19179);
nand U19795 (N_19795,N_18938,N_18797);
nor U19796 (N_19796,N_18812,N_18928);
nand U19797 (N_19797,N_18864,N_19355);
xnor U19798 (N_19798,N_19271,N_18879);
nand U19799 (N_19799,N_18785,N_19284);
nor U19800 (N_19800,N_18847,N_19341);
xnor U19801 (N_19801,N_19016,N_19191);
or U19802 (N_19802,N_18767,N_18870);
xor U19803 (N_19803,N_19240,N_19304);
nand U19804 (N_19804,N_19240,N_18782);
nand U19805 (N_19805,N_18945,N_18832);
xnor U19806 (N_19806,N_18837,N_19198);
nand U19807 (N_19807,N_19364,N_19089);
xnor U19808 (N_19808,N_19294,N_19287);
nor U19809 (N_19809,N_19161,N_18766);
xnor U19810 (N_19810,N_18755,N_18871);
or U19811 (N_19811,N_19123,N_19057);
and U19812 (N_19812,N_19229,N_19012);
xnor U19813 (N_19813,N_19339,N_18766);
nand U19814 (N_19814,N_18888,N_18862);
nor U19815 (N_19815,N_19349,N_19107);
or U19816 (N_19816,N_19350,N_19211);
nand U19817 (N_19817,N_19055,N_19069);
nor U19818 (N_19818,N_19264,N_18819);
and U19819 (N_19819,N_19369,N_19275);
nor U19820 (N_19820,N_19043,N_18871);
nand U19821 (N_19821,N_19164,N_18846);
or U19822 (N_19822,N_19194,N_18775);
nor U19823 (N_19823,N_19089,N_18904);
or U19824 (N_19824,N_19160,N_18937);
and U19825 (N_19825,N_19315,N_19052);
xnor U19826 (N_19826,N_18827,N_19323);
nor U19827 (N_19827,N_18824,N_18974);
or U19828 (N_19828,N_19257,N_19042);
xor U19829 (N_19829,N_19147,N_18859);
xnor U19830 (N_19830,N_19299,N_18900);
xnor U19831 (N_19831,N_19208,N_19333);
xnor U19832 (N_19832,N_19214,N_19265);
or U19833 (N_19833,N_19044,N_19332);
or U19834 (N_19834,N_18963,N_19359);
nor U19835 (N_19835,N_19351,N_19104);
or U19836 (N_19836,N_18869,N_19227);
nand U19837 (N_19837,N_18819,N_19073);
and U19838 (N_19838,N_18803,N_19304);
nor U19839 (N_19839,N_18834,N_19003);
nand U19840 (N_19840,N_19219,N_18865);
or U19841 (N_19841,N_19344,N_19168);
xor U19842 (N_19842,N_18866,N_19038);
nand U19843 (N_19843,N_19162,N_18940);
nand U19844 (N_19844,N_18788,N_19177);
nor U19845 (N_19845,N_19093,N_18839);
and U19846 (N_19846,N_18780,N_18953);
nor U19847 (N_19847,N_19275,N_19278);
or U19848 (N_19848,N_19312,N_18830);
or U19849 (N_19849,N_18907,N_18753);
nand U19850 (N_19850,N_18997,N_18770);
nor U19851 (N_19851,N_18940,N_18773);
or U19852 (N_19852,N_18848,N_18754);
xnor U19853 (N_19853,N_19210,N_19247);
or U19854 (N_19854,N_19001,N_18983);
and U19855 (N_19855,N_18807,N_19293);
nand U19856 (N_19856,N_19269,N_19221);
nand U19857 (N_19857,N_19106,N_18813);
nand U19858 (N_19858,N_18935,N_18962);
xor U19859 (N_19859,N_19115,N_19027);
or U19860 (N_19860,N_19034,N_18794);
xor U19861 (N_19861,N_19142,N_19158);
xnor U19862 (N_19862,N_19088,N_18915);
or U19863 (N_19863,N_18797,N_19150);
nand U19864 (N_19864,N_18998,N_18828);
nand U19865 (N_19865,N_18944,N_19047);
or U19866 (N_19866,N_19039,N_18920);
nand U19867 (N_19867,N_18824,N_19358);
and U19868 (N_19868,N_19094,N_18841);
or U19869 (N_19869,N_19319,N_19280);
and U19870 (N_19870,N_18763,N_18787);
and U19871 (N_19871,N_19368,N_19167);
and U19872 (N_19872,N_19299,N_19091);
nor U19873 (N_19873,N_19248,N_18761);
or U19874 (N_19874,N_18868,N_19203);
or U19875 (N_19875,N_18759,N_19304);
or U19876 (N_19876,N_18923,N_18976);
xnor U19877 (N_19877,N_19105,N_19278);
and U19878 (N_19878,N_19359,N_18775);
and U19879 (N_19879,N_19228,N_19125);
or U19880 (N_19880,N_19269,N_18967);
nand U19881 (N_19881,N_18839,N_19269);
or U19882 (N_19882,N_19215,N_19148);
or U19883 (N_19883,N_19260,N_19000);
xor U19884 (N_19884,N_19174,N_19330);
and U19885 (N_19885,N_19090,N_19003);
nand U19886 (N_19886,N_19174,N_19006);
xnor U19887 (N_19887,N_18968,N_18897);
and U19888 (N_19888,N_19172,N_19317);
xor U19889 (N_19889,N_19039,N_18975);
nor U19890 (N_19890,N_19088,N_19148);
and U19891 (N_19891,N_19096,N_18793);
nand U19892 (N_19892,N_18792,N_18987);
xor U19893 (N_19893,N_18809,N_19176);
nand U19894 (N_19894,N_18768,N_19187);
or U19895 (N_19895,N_19259,N_18964);
nor U19896 (N_19896,N_19368,N_19019);
nand U19897 (N_19897,N_19262,N_19290);
nor U19898 (N_19898,N_19224,N_18813);
and U19899 (N_19899,N_18762,N_19233);
nor U19900 (N_19900,N_18829,N_19218);
nand U19901 (N_19901,N_19122,N_19248);
or U19902 (N_19902,N_19217,N_19082);
and U19903 (N_19903,N_19262,N_18867);
or U19904 (N_19904,N_19359,N_18870);
xnor U19905 (N_19905,N_18966,N_19273);
or U19906 (N_19906,N_19254,N_18854);
xor U19907 (N_19907,N_18966,N_19098);
and U19908 (N_19908,N_18956,N_18947);
and U19909 (N_19909,N_19195,N_18916);
and U19910 (N_19910,N_19098,N_19299);
nand U19911 (N_19911,N_18896,N_19135);
nor U19912 (N_19912,N_18925,N_19034);
nor U19913 (N_19913,N_18770,N_19185);
or U19914 (N_19914,N_19360,N_19140);
and U19915 (N_19915,N_19308,N_18761);
or U19916 (N_19916,N_19349,N_19362);
and U19917 (N_19917,N_19277,N_18895);
nor U19918 (N_19918,N_18913,N_19263);
nand U19919 (N_19919,N_18803,N_19066);
nor U19920 (N_19920,N_18812,N_19146);
and U19921 (N_19921,N_18770,N_19371);
and U19922 (N_19922,N_18882,N_19303);
xnor U19923 (N_19923,N_18992,N_19143);
and U19924 (N_19924,N_19285,N_19151);
xnor U19925 (N_19925,N_18831,N_19287);
xor U19926 (N_19926,N_18803,N_18935);
and U19927 (N_19927,N_19077,N_19090);
or U19928 (N_19928,N_18969,N_19279);
and U19929 (N_19929,N_19099,N_19220);
and U19930 (N_19930,N_18912,N_19249);
or U19931 (N_19931,N_19339,N_19238);
and U19932 (N_19932,N_19024,N_19033);
and U19933 (N_19933,N_18756,N_19049);
nor U19934 (N_19934,N_18958,N_19306);
nor U19935 (N_19935,N_19156,N_19045);
or U19936 (N_19936,N_18934,N_19245);
nand U19937 (N_19937,N_19129,N_18974);
nand U19938 (N_19938,N_18822,N_19014);
nor U19939 (N_19939,N_19067,N_19296);
and U19940 (N_19940,N_18962,N_18982);
or U19941 (N_19941,N_19074,N_19134);
xor U19942 (N_19942,N_19082,N_18808);
or U19943 (N_19943,N_19216,N_18887);
nor U19944 (N_19944,N_18784,N_18859);
nand U19945 (N_19945,N_19333,N_19071);
and U19946 (N_19946,N_18892,N_19116);
and U19947 (N_19947,N_19350,N_19015);
nor U19948 (N_19948,N_19032,N_19155);
nor U19949 (N_19949,N_19098,N_18986);
or U19950 (N_19950,N_19248,N_19365);
xor U19951 (N_19951,N_19102,N_18803);
nor U19952 (N_19952,N_19050,N_18878);
nand U19953 (N_19953,N_19033,N_19265);
nand U19954 (N_19954,N_18903,N_18920);
and U19955 (N_19955,N_18903,N_18753);
xor U19956 (N_19956,N_19371,N_19014);
nand U19957 (N_19957,N_19155,N_18955);
nand U19958 (N_19958,N_19000,N_19081);
nor U19959 (N_19959,N_19052,N_18837);
nor U19960 (N_19960,N_19033,N_19209);
and U19961 (N_19961,N_18785,N_18784);
nand U19962 (N_19962,N_19008,N_19134);
nor U19963 (N_19963,N_19059,N_19264);
nand U19964 (N_19964,N_19151,N_19033);
and U19965 (N_19965,N_19031,N_18750);
or U19966 (N_19966,N_18846,N_19374);
or U19967 (N_19967,N_19003,N_18956);
xnor U19968 (N_19968,N_18911,N_18865);
xnor U19969 (N_19969,N_19268,N_19129);
nand U19970 (N_19970,N_18863,N_19338);
xor U19971 (N_19971,N_19004,N_19130);
nand U19972 (N_19972,N_18892,N_18987);
nand U19973 (N_19973,N_18875,N_18783);
nand U19974 (N_19974,N_18960,N_18990);
and U19975 (N_19975,N_19043,N_18934);
nand U19976 (N_19976,N_18852,N_18833);
xor U19977 (N_19977,N_18963,N_19057);
and U19978 (N_19978,N_19040,N_19032);
nor U19979 (N_19979,N_18931,N_18957);
nor U19980 (N_19980,N_19149,N_19175);
nor U19981 (N_19981,N_19214,N_19070);
xnor U19982 (N_19982,N_19326,N_19170);
and U19983 (N_19983,N_18981,N_18952);
or U19984 (N_19984,N_19196,N_19328);
xnor U19985 (N_19985,N_19244,N_19173);
or U19986 (N_19986,N_18893,N_19230);
nand U19987 (N_19987,N_19251,N_19050);
nor U19988 (N_19988,N_19076,N_18886);
and U19989 (N_19989,N_18849,N_18971);
nor U19990 (N_19990,N_18789,N_18775);
nand U19991 (N_19991,N_19133,N_19349);
nand U19992 (N_19992,N_19302,N_19081);
xor U19993 (N_19993,N_19114,N_18912);
xor U19994 (N_19994,N_18806,N_19134);
xnor U19995 (N_19995,N_19004,N_19313);
xnor U19996 (N_19996,N_19293,N_19166);
and U19997 (N_19997,N_19236,N_18889);
and U19998 (N_19998,N_18803,N_18862);
and U19999 (N_19999,N_18946,N_19062);
or U20000 (N_20000,N_19808,N_19858);
nand U20001 (N_20001,N_19943,N_19555);
nor U20002 (N_20002,N_19459,N_19481);
and U20003 (N_20003,N_19627,N_19628);
nor U20004 (N_20004,N_19738,N_19997);
nand U20005 (N_20005,N_19438,N_19647);
nor U20006 (N_20006,N_19847,N_19565);
and U20007 (N_20007,N_19967,N_19614);
nand U20008 (N_20008,N_19879,N_19390);
or U20009 (N_20009,N_19630,N_19440);
nor U20010 (N_20010,N_19785,N_19993);
and U20011 (N_20011,N_19391,N_19940);
xnor U20012 (N_20012,N_19831,N_19846);
nand U20013 (N_20013,N_19712,N_19533);
nor U20014 (N_20014,N_19706,N_19723);
nand U20015 (N_20015,N_19609,N_19758);
or U20016 (N_20016,N_19931,N_19950);
xor U20017 (N_20017,N_19749,N_19849);
nand U20018 (N_20018,N_19934,N_19543);
nor U20019 (N_20019,N_19770,N_19494);
or U20020 (N_20020,N_19376,N_19691);
xor U20021 (N_20021,N_19973,N_19988);
xor U20022 (N_20022,N_19528,N_19745);
or U20023 (N_20023,N_19439,N_19479);
nor U20024 (N_20024,N_19495,N_19673);
and U20025 (N_20025,N_19883,N_19915);
or U20026 (N_20026,N_19492,N_19780);
nor U20027 (N_20027,N_19919,N_19425);
and U20028 (N_20028,N_19935,N_19748);
or U20029 (N_20029,N_19821,N_19660);
or U20030 (N_20030,N_19818,N_19897);
nor U20031 (N_20031,N_19421,N_19728);
nor U20032 (N_20032,N_19717,N_19526);
nor U20033 (N_20033,N_19431,N_19804);
and U20034 (N_20034,N_19407,N_19841);
nor U20035 (N_20035,N_19870,N_19653);
nor U20036 (N_20036,N_19907,N_19602);
or U20037 (N_20037,N_19828,N_19774);
nor U20038 (N_20038,N_19856,N_19799);
and U20039 (N_20039,N_19592,N_19531);
nor U20040 (N_20040,N_19900,N_19589);
nor U20041 (N_20041,N_19619,N_19827);
nand U20042 (N_20042,N_19772,N_19595);
and U20043 (N_20043,N_19633,N_19835);
xnor U20044 (N_20044,N_19722,N_19581);
nor U20045 (N_20045,N_19864,N_19582);
nor U20046 (N_20046,N_19980,N_19670);
nor U20047 (N_20047,N_19701,N_19966);
or U20048 (N_20048,N_19777,N_19979);
nor U20049 (N_20049,N_19876,N_19845);
nor U20050 (N_20050,N_19601,N_19715);
nor U20051 (N_20051,N_19585,N_19648);
nand U20052 (N_20052,N_19392,N_19987);
and U20053 (N_20053,N_19505,N_19552);
and U20054 (N_20054,N_19939,N_19877);
or U20055 (N_20055,N_19755,N_19735);
nand U20056 (N_20056,N_19468,N_19450);
nand U20057 (N_20057,N_19751,N_19557);
xor U20058 (N_20058,N_19575,N_19588);
xor U20059 (N_20059,N_19913,N_19613);
and U20060 (N_20060,N_19923,N_19382);
and U20061 (N_20061,N_19594,N_19961);
nor U20062 (N_20062,N_19607,N_19960);
nand U20063 (N_20063,N_19556,N_19747);
xor U20064 (N_20064,N_19662,N_19805);
and U20065 (N_20065,N_19677,N_19655);
xor U20066 (N_20066,N_19882,N_19576);
nor U20067 (N_20067,N_19823,N_19529);
and U20068 (N_20068,N_19457,N_19649);
xor U20069 (N_20069,N_19536,N_19472);
nand U20070 (N_20070,N_19410,N_19416);
nand U20071 (N_20071,N_19986,N_19800);
nor U20072 (N_20072,N_19832,N_19636);
and U20073 (N_20073,N_19704,N_19461);
xor U20074 (N_20074,N_19600,N_19697);
nor U20075 (N_20075,N_19473,N_19626);
nand U20076 (N_20076,N_19801,N_19675);
nor U20077 (N_20077,N_19642,N_19475);
nor U20078 (N_20078,N_19519,N_19843);
xor U20079 (N_20079,N_19646,N_19788);
or U20080 (N_20080,N_19941,N_19978);
or U20081 (N_20081,N_19857,N_19426);
or U20082 (N_20082,N_19571,N_19658);
nand U20083 (N_20083,N_19509,N_19781);
nor U20084 (N_20084,N_19507,N_19558);
xor U20085 (N_20085,N_19891,N_19419);
xor U20086 (N_20086,N_19949,N_19656);
and U20087 (N_20087,N_19682,N_19631);
nand U20088 (N_20088,N_19895,N_19460);
or U20089 (N_20089,N_19463,N_19469);
nor U20090 (N_20090,N_19810,N_19448);
nand U20091 (N_20091,N_19963,N_19638);
xnor U20092 (N_20092,N_19922,N_19844);
and U20093 (N_20093,N_19692,N_19523);
nand U20094 (N_20094,N_19707,N_19579);
and U20095 (N_20095,N_19502,N_19834);
or U20096 (N_20096,N_19784,N_19766);
nand U20097 (N_20097,N_19713,N_19868);
xnor U20098 (N_20098,N_19930,N_19905);
nor U20099 (N_20099,N_19423,N_19942);
nor U20100 (N_20100,N_19737,N_19500);
xor U20101 (N_20101,N_19694,N_19616);
and U20102 (N_20102,N_19976,N_19449);
nand U20103 (N_20103,N_19503,N_19819);
and U20104 (N_20104,N_19708,N_19861);
nor U20105 (N_20105,N_19397,N_19926);
nand U20106 (N_20106,N_19802,N_19947);
nand U20107 (N_20107,N_19637,N_19957);
nor U20108 (N_20108,N_19786,N_19726);
nand U20109 (N_20109,N_19990,N_19865);
nor U20110 (N_20110,N_19487,N_19887);
nor U20111 (N_20111,N_19992,N_19603);
xor U20112 (N_20112,N_19659,N_19667);
nand U20113 (N_20113,N_19550,N_19453);
nor U20114 (N_20114,N_19880,N_19984);
and U20115 (N_20115,N_19508,N_19488);
xnor U20116 (N_20116,N_19791,N_19484);
xnor U20117 (N_20117,N_19635,N_19608);
nand U20118 (N_20118,N_19776,N_19620);
or U20119 (N_20119,N_19501,N_19486);
and U20120 (N_20120,N_19377,N_19605);
and U20121 (N_20121,N_19386,N_19918);
xnor U20122 (N_20122,N_19560,N_19518);
or U20123 (N_20123,N_19890,N_19688);
xor U20124 (N_20124,N_19937,N_19643);
nor U20125 (N_20125,N_19753,N_19437);
nor U20126 (N_20126,N_19447,N_19898);
nand U20127 (N_20127,N_19510,N_19577);
nor U20128 (N_20128,N_19482,N_19666);
xnor U20129 (N_20129,N_19686,N_19914);
nand U20130 (N_20130,N_19393,N_19962);
nor U20131 (N_20131,N_19970,N_19545);
or U20132 (N_20132,N_19379,N_19756);
xor U20133 (N_20133,N_19395,N_19885);
or U20134 (N_20134,N_19862,N_19665);
xnor U20135 (N_20135,N_19794,N_19549);
xor U20136 (N_20136,N_19398,N_19956);
xor U20137 (N_20137,N_19792,N_19491);
nor U20138 (N_20138,N_19597,N_19743);
or U20139 (N_20139,N_19902,N_19744);
xnor U20140 (N_20140,N_19764,N_19807);
nand U20141 (N_20141,N_19720,N_19977);
nor U20142 (N_20142,N_19452,N_19454);
or U20143 (N_20143,N_19586,N_19933);
nand U20144 (N_20144,N_19681,N_19520);
and U20145 (N_20145,N_19981,N_19816);
and U20146 (N_20146,N_19496,N_19467);
nor U20147 (N_20147,N_19892,N_19672);
nor U20148 (N_20148,N_19664,N_19991);
nor U20149 (N_20149,N_19850,N_19955);
and U20150 (N_20150,N_19563,N_19583);
nor U20151 (N_20151,N_19652,N_19532);
nor U20152 (N_20152,N_19465,N_19783);
xor U20153 (N_20153,N_19559,N_19553);
or U20154 (N_20154,N_19401,N_19871);
nand U20155 (N_20155,N_19964,N_19860);
xor U20156 (N_20156,N_19702,N_19402);
nor U20157 (N_20157,N_19497,N_19951);
or U20158 (N_20158,N_19428,N_19873);
xor U20159 (N_20159,N_19842,N_19797);
nor U20160 (N_20160,N_19859,N_19750);
nor U20161 (N_20161,N_19610,N_19483);
nor U20162 (N_20162,N_19663,N_19411);
or U20163 (N_20163,N_19669,N_19718);
or U20164 (N_20164,N_19727,N_19615);
xor U20165 (N_20165,N_19969,N_19760);
or U20166 (N_20166,N_19538,N_19551);
nand U20167 (N_20167,N_19640,N_19629);
or U20168 (N_20168,N_19757,N_19462);
xor U20169 (N_20169,N_19932,N_19710);
or U20170 (N_20170,N_19954,N_19464);
xor U20171 (N_20171,N_19734,N_19668);
or U20172 (N_20172,N_19739,N_19546);
xor U20173 (N_20173,N_19434,N_19485);
nor U20174 (N_20174,N_19671,N_19412);
xor U20175 (N_20175,N_19938,N_19769);
xor U20176 (N_20176,N_19474,N_19886);
nand U20177 (N_20177,N_19789,N_19378);
and U20178 (N_20178,N_19917,N_19674);
or U20179 (N_20179,N_19654,N_19644);
xnor U20180 (N_20180,N_19541,N_19684);
xnor U20181 (N_20181,N_19683,N_19623);
nor U20182 (N_20182,N_19417,N_19752);
nand U20183 (N_20183,N_19403,N_19953);
nand U20184 (N_20184,N_19912,N_19685);
nand U20185 (N_20185,N_19763,N_19539);
xnor U20186 (N_20186,N_19471,N_19948);
nand U20187 (N_20187,N_19921,N_19436);
nand U20188 (N_20188,N_19590,N_19490);
nand U20189 (N_20189,N_19830,N_19394);
xnor U20190 (N_20190,N_19995,N_19548);
and U20191 (N_20191,N_19840,N_19420);
xnor U20192 (N_20192,N_19498,N_19478);
nand U20193 (N_20193,N_19598,N_19773);
nor U20194 (N_20194,N_19888,N_19554);
nor U20195 (N_20195,N_19853,N_19515);
or U20196 (N_20196,N_19927,N_19470);
nand U20197 (N_20197,N_19893,N_19855);
nand U20198 (N_20198,N_19444,N_19989);
and U20199 (N_20199,N_19689,N_19716);
nand U20200 (N_20200,N_19432,N_19829);
nor U20201 (N_20201,N_19809,N_19771);
xnor U20202 (N_20202,N_19920,N_19599);
nand U20203 (N_20203,N_19971,N_19721);
xnor U20204 (N_20204,N_19387,N_19514);
or U20205 (N_20205,N_19906,N_19404);
nand U20206 (N_20206,N_19511,N_19945);
or U20207 (N_20207,N_19936,N_19889);
nor U20208 (N_20208,N_19443,N_19430);
xor U20209 (N_20209,N_19825,N_19901);
and U20210 (N_20210,N_19779,N_19729);
xor U20211 (N_20211,N_19813,N_19812);
and U20212 (N_20212,N_19612,N_19826);
nor U20213 (N_20213,N_19380,N_19916);
nor U20214 (N_20214,N_19740,N_19896);
nand U20215 (N_20215,N_19946,N_19820);
xor U20216 (N_20216,N_19639,N_19578);
xnor U20217 (N_20217,N_19854,N_19869);
nand U20218 (N_20218,N_19544,N_19974);
nand U20219 (N_20219,N_19574,N_19504);
and U20220 (N_20220,N_19566,N_19924);
and U20221 (N_20221,N_19903,N_19837);
or U20222 (N_20222,N_19695,N_19928);
nand U20223 (N_20223,N_19513,N_19451);
and U20224 (N_20224,N_19848,N_19904);
or U20225 (N_20225,N_19894,N_19522);
and U20226 (N_20226,N_19568,N_19782);
and U20227 (N_20227,N_19817,N_19982);
or U20228 (N_20228,N_19687,N_19445);
nand U20229 (N_20229,N_19641,N_19591);
or U20230 (N_20230,N_19433,N_19573);
and U20231 (N_20231,N_19908,N_19765);
and U20232 (N_20232,N_19838,N_19867);
nand U20233 (N_20233,N_19994,N_19476);
nor U20234 (N_20234,N_19778,N_19796);
or U20235 (N_20235,N_19998,N_19851);
nand U20236 (N_20236,N_19881,N_19540);
nor U20237 (N_20237,N_19506,N_19696);
xnor U20238 (N_20238,N_19719,N_19661);
nand U20239 (N_20239,N_19516,N_19746);
nand U20240 (N_20240,N_19709,N_19442);
and U20241 (N_20241,N_19385,N_19406);
or U20242 (N_20242,N_19679,N_19676);
nand U20243 (N_20243,N_19572,N_19547);
xnor U20244 (N_20244,N_19878,N_19732);
nor U20245 (N_20245,N_19775,N_19972);
or U20246 (N_20246,N_19527,N_19383);
or U20247 (N_20247,N_19884,N_19564);
and U20248 (N_20248,N_19703,N_19985);
nand U20249 (N_20249,N_19409,N_19711);
or U20250 (N_20250,N_19632,N_19759);
and U20251 (N_20251,N_19621,N_19534);
nor U20252 (N_20252,N_19606,N_19767);
or U20253 (N_20253,N_19725,N_19657);
nand U20254 (N_20254,N_19787,N_19811);
xnor U20255 (N_20255,N_19618,N_19815);
and U20256 (N_20256,N_19418,N_19730);
and U20257 (N_20257,N_19733,N_19803);
xor U20258 (N_20258,N_19731,N_19567);
nand U20259 (N_20259,N_19795,N_19645);
or U20260 (N_20260,N_19793,N_19700);
nor U20261 (N_20261,N_19814,N_19381);
nand U20262 (N_20262,N_19839,N_19836);
or U20263 (N_20263,N_19584,N_19678);
nor U20264 (N_20264,N_19824,N_19952);
xor U20265 (N_20265,N_19480,N_19996);
xor U20266 (N_20266,N_19524,N_19875);
or U20267 (N_20267,N_19790,N_19910);
xor U20268 (N_20268,N_19622,N_19863);
nor U20269 (N_20269,N_19441,N_19761);
and U20270 (N_20270,N_19604,N_19415);
and U20271 (N_20271,N_19999,N_19396);
nand U20272 (N_20272,N_19699,N_19611);
xnor U20273 (N_20273,N_19429,N_19408);
or U20274 (N_20274,N_19625,N_19562);
nand U20275 (N_20275,N_19422,N_19530);
and U20276 (N_20276,N_19570,N_19899);
or U20277 (N_20277,N_19736,N_19489);
xnor U20278 (N_20278,N_19714,N_19959);
or U20279 (N_20279,N_19968,N_19680);
nor U20280 (N_20280,N_19535,N_19872);
or U20281 (N_20281,N_19651,N_19435);
and U20282 (N_20282,N_19911,N_19384);
and U20283 (N_20283,N_19624,N_19617);
xor U20284 (N_20284,N_19768,N_19975);
nor U20285 (N_20285,N_19388,N_19852);
nor U20286 (N_20286,N_19798,N_19521);
nand U20287 (N_20287,N_19833,N_19958);
and U20288 (N_20288,N_19693,N_19400);
xnor U20289 (N_20289,N_19874,N_19596);
or U20290 (N_20290,N_19822,N_19944);
or U20291 (N_20291,N_19705,N_19965);
nand U20292 (N_20292,N_19650,N_19909);
nor U20293 (N_20293,N_19587,N_19446);
and U20294 (N_20294,N_19414,N_19537);
nand U20295 (N_20295,N_19542,N_19424);
and U20296 (N_20296,N_19690,N_19925);
nand U20297 (N_20297,N_19466,N_19561);
nand U20298 (N_20298,N_19762,N_19698);
nand U20299 (N_20299,N_19866,N_19569);
nand U20300 (N_20300,N_19724,N_19499);
nand U20301 (N_20301,N_19754,N_19806);
nand U20302 (N_20302,N_19455,N_19413);
and U20303 (N_20303,N_19389,N_19512);
xnor U20304 (N_20304,N_19456,N_19580);
nand U20305 (N_20305,N_19427,N_19375);
and U20306 (N_20306,N_19634,N_19525);
or U20307 (N_20307,N_19405,N_19929);
xor U20308 (N_20308,N_19477,N_19458);
xor U20309 (N_20309,N_19983,N_19493);
nor U20310 (N_20310,N_19742,N_19399);
nand U20311 (N_20311,N_19517,N_19741);
xor U20312 (N_20312,N_19593,N_19832);
xnor U20313 (N_20313,N_19740,N_19879);
or U20314 (N_20314,N_19635,N_19380);
xor U20315 (N_20315,N_19672,N_19511);
and U20316 (N_20316,N_19375,N_19686);
xor U20317 (N_20317,N_19447,N_19417);
and U20318 (N_20318,N_19872,N_19694);
or U20319 (N_20319,N_19969,N_19819);
nand U20320 (N_20320,N_19774,N_19728);
nand U20321 (N_20321,N_19698,N_19381);
nor U20322 (N_20322,N_19887,N_19410);
and U20323 (N_20323,N_19445,N_19462);
xnor U20324 (N_20324,N_19487,N_19475);
or U20325 (N_20325,N_19689,N_19795);
or U20326 (N_20326,N_19879,N_19827);
nand U20327 (N_20327,N_19575,N_19957);
and U20328 (N_20328,N_19943,N_19444);
xor U20329 (N_20329,N_19912,N_19428);
nor U20330 (N_20330,N_19939,N_19968);
xor U20331 (N_20331,N_19669,N_19904);
nor U20332 (N_20332,N_19719,N_19947);
and U20333 (N_20333,N_19441,N_19828);
nand U20334 (N_20334,N_19670,N_19659);
or U20335 (N_20335,N_19932,N_19654);
or U20336 (N_20336,N_19585,N_19709);
xor U20337 (N_20337,N_19962,N_19887);
or U20338 (N_20338,N_19376,N_19628);
nand U20339 (N_20339,N_19615,N_19399);
nor U20340 (N_20340,N_19536,N_19975);
and U20341 (N_20341,N_19415,N_19414);
nor U20342 (N_20342,N_19809,N_19846);
or U20343 (N_20343,N_19618,N_19392);
nor U20344 (N_20344,N_19560,N_19627);
nand U20345 (N_20345,N_19434,N_19451);
and U20346 (N_20346,N_19419,N_19492);
nor U20347 (N_20347,N_19621,N_19631);
xnor U20348 (N_20348,N_19476,N_19713);
nor U20349 (N_20349,N_19806,N_19879);
xor U20350 (N_20350,N_19642,N_19437);
and U20351 (N_20351,N_19927,N_19702);
and U20352 (N_20352,N_19474,N_19391);
nand U20353 (N_20353,N_19928,N_19686);
and U20354 (N_20354,N_19511,N_19731);
nor U20355 (N_20355,N_19796,N_19435);
xnor U20356 (N_20356,N_19895,N_19510);
and U20357 (N_20357,N_19628,N_19818);
or U20358 (N_20358,N_19468,N_19626);
xor U20359 (N_20359,N_19391,N_19680);
nand U20360 (N_20360,N_19500,N_19930);
xor U20361 (N_20361,N_19440,N_19441);
nor U20362 (N_20362,N_19424,N_19776);
or U20363 (N_20363,N_19672,N_19408);
nor U20364 (N_20364,N_19668,N_19777);
and U20365 (N_20365,N_19738,N_19580);
and U20366 (N_20366,N_19677,N_19845);
xnor U20367 (N_20367,N_19696,N_19430);
xnor U20368 (N_20368,N_19517,N_19719);
nor U20369 (N_20369,N_19795,N_19454);
xnor U20370 (N_20370,N_19825,N_19582);
xnor U20371 (N_20371,N_19938,N_19863);
or U20372 (N_20372,N_19861,N_19852);
xor U20373 (N_20373,N_19736,N_19854);
and U20374 (N_20374,N_19783,N_19821);
and U20375 (N_20375,N_19683,N_19875);
xor U20376 (N_20376,N_19855,N_19877);
and U20377 (N_20377,N_19418,N_19428);
nor U20378 (N_20378,N_19956,N_19893);
and U20379 (N_20379,N_19427,N_19558);
nor U20380 (N_20380,N_19911,N_19412);
nor U20381 (N_20381,N_19647,N_19421);
and U20382 (N_20382,N_19773,N_19805);
or U20383 (N_20383,N_19938,N_19765);
or U20384 (N_20384,N_19820,N_19738);
nand U20385 (N_20385,N_19589,N_19752);
nor U20386 (N_20386,N_19399,N_19536);
nor U20387 (N_20387,N_19412,N_19521);
and U20388 (N_20388,N_19497,N_19811);
xor U20389 (N_20389,N_19820,N_19742);
and U20390 (N_20390,N_19873,N_19477);
nand U20391 (N_20391,N_19801,N_19912);
nor U20392 (N_20392,N_19919,N_19543);
or U20393 (N_20393,N_19637,N_19848);
xnor U20394 (N_20394,N_19941,N_19708);
or U20395 (N_20395,N_19883,N_19476);
nor U20396 (N_20396,N_19538,N_19553);
or U20397 (N_20397,N_19635,N_19840);
nand U20398 (N_20398,N_19997,N_19521);
or U20399 (N_20399,N_19953,N_19721);
or U20400 (N_20400,N_19554,N_19575);
nand U20401 (N_20401,N_19549,N_19386);
nor U20402 (N_20402,N_19390,N_19860);
xnor U20403 (N_20403,N_19674,N_19840);
or U20404 (N_20404,N_19795,N_19890);
or U20405 (N_20405,N_19851,N_19523);
or U20406 (N_20406,N_19628,N_19970);
and U20407 (N_20407,N_19851,N_19864);
xor U20408 (N_20408,N_19941,N_19710);
or U20409 (N_20409,N_19568,N_19726);
or U20410 (N_20410,N_19920,N_19723);
xor U20411 (N_20411,N_19465,N_19839);
nor U20412 (N_20412,N_19443,N_19389);
nor U20413 (N_20413,N_19407,N_19895);
nor U20414 (N_20414,N_19692,N_19708);
or U20415 (N_20415,N_19397,N_19527);
nor U20416 (N_20416,N_19597,N_19475);
nand U20417 (N_20417,N_19683,N_19796);
nand U20418 (N_20418,N_19717,N_19701);
nand U20419 (N_20419,N_19988,N_19548);
or U20420 (N_20420,N_19508,N_19867);
xnor U20421 (N_20421,N_19700,N_19716);
nand U20422 (N_20422,N_19880,N_19788);
nand U20423 (N_20423,N_19504,N_19745);
nand U20424 (N_20424,N_19428,N_19588);
and U20425 (N_20425,N_19396,N_19411);
nand U20426 (N_20426,N_19757,N_19811);
nand U20427 (N_20427,N_19629,N_19891);
xnor U20428 (N_20428,N_19617,N_19968);
and U20429 (N_20429,N_19587,N_19634);
nor U20430 (N_20430,N_19705,N_19949);
xor U20431 (N_20431,N_19871,N_19438);
nand U20432 (N_20432,N_19842,N_19935);
xnor U20433 (N_20433,N_19579,N_19534);
nor U20434 (N_20434,N_19418,N_19765);
and U20435 (N_20435,N_19631,N_19426);
xnor U20436 (N_20436,N_19974,N_19429);
xnor U20437 (N_20437,N_19713,N_19508);
nor U20438 (N_20438,N_19840,N_19439);
and U20439 (N_20439,N_19642,N_19683);
or U20440 (N_20440,N_19614,N_19686);
nand U20441 (N_20441,N_19707,N_19664);
nor U20442 (N_20442,N_19620,N_19773);
and U20443 (N_20443,N_19534,N_19968);
nand U20444 (N_20444,N_19874,N_19492);
or U20445 (N_20445,N_19593,N_19932);
xnor U20446 (N_20446,N_19552,N_19711);
and U20447 (N_20447,N_19875,N_19422);
or U20448 (N_20448,N_19734,N_19885);
nor U20449 (N_20449,N_19994,N_19888);
nor U20450 (N_20450,N_19599,N_19857);
and U20451 (N_20451,N_19386,N_19380);
nand U20452 (N_20452,N_19653,N_19737);
and U20453 (N_20453,N_19877,N_19985);
nand U20454 (N_20454,N_19854,N_19794);
nand U20455 (N_20455,N_19921,N_19839);
or U20456 (N_20456,N_19860,N_19556);
nor U20457 (N_20457,N_19807,N_19854);
xnor U20458 (N_20458,N_19721,N_19585);
nor U20459 (N_20459,N_19438,N_19508);
and U20460 (N_20460,N_19997,N_19592);
xor U20461 (N_20461,N_19654,N_19715);
or U20462 (N_20462,N_19812,N_19376);
nand U20463 (N_20463,N_19742,N_19463);
xnor U20464 (N_20464,N_19823,N_19868);
xnor U20465 (N_20465,N_19560,N_19437);
and U20466 (N_20466,N_19859,N_19554);
or U20467 (N_20467,N_19378,N_19609);
xor U20468 (N_20468,N_19740,N_19835);
and U20469 (N_20469,N_19533,N_19500);
and U20470 (N_20470,N_19732,N_19907);
nand U20471 (N_20471,N_19988,N_19816);
xnor U20472 (N_20472,N_19922,N_19644);
and U20473 (N_20473,N_19552,N_19838);
or U20474 (N_20474,N_19817,N_19652);
nand U20475 (N_20475,N_19948,N_19536);
or U20476 (N_20476,N_19551,N_19595);
nor U20477 (N_20477,N_19552,N_19779);
nand U20478 (N_20478,N_19829,N_19972);
or U20479 (N_20479,N_19444,N_19880);
or U20480 (N_20480,N_19703,N_19523);
nand U20481 (N_20481,N_19870,N_19907);
xor U20482 (N_20482,N_19740,N_19814);
xor U20483 (N_20483,N_19873,N_19905);
and U20484 (N_20484,N_19726,N_19989);
xnor U20485 (N_20485,N_19743,N_19727);
and U20486 (N_20486,N_19869,N_19552);
nand U20487 (N_20487,N_19754,N_19454);
nand U20488 (N_20488,N_19745,N_19505);
xor U20489 (N_20489,N_19923,N_19727);
nor U20490 (N_20490,N_19528,N_19665);
nand U20491 (N_20491,N_19450,N_19998);
xor U20492 (N_20492,N_19558,N_19627);
and U20493 (N_20493,N_19723,N_19984);
and U20494 (N_20494,N_19928,N_19619);
xor U20495 (N_20495,N_19748,N_19508);
and U20496 (N_20496,N_19992,N_19897);
nor U20497 (N_20497,N_19836,N_19592);
nor U20498 (N_20498,N_19421,N_19868);
or U20499 (N_20499,N_19383,N_19596);
or U20500 (N_20500,N_19929,N_19386);
nand U20501 (N_20501,N_19428,N_19666);
nor U20502 (N_20502,N_19833,N_19653);
nor U20503 (N_20503,N_19530,N_19390);
or U20504 (N_20504,N_19404,N_19494);
and U20505 (N_20505,N_19579,N_19486);
and U20506 (N_20506,N_19602,N_19879);
nand U20507 (N_20507,N_19784,N_19929);
and U20508 (N_20508,N_19745,N_19640);
xor U20509 (N_20509,N_19854,N_19899);
and U20510 (N_20510,N_19671,N_19878);
or U20511 (N_20511,N_19633,N_19794);
or U20512 (N_20512,N_19986,N_19617);
or U20513 (N_20513,N_19916,N_19731);
and U20514 (N_20514,N_19928,N_19578);
and U20515 (N_20515,N_19406,N_19524);
or U20516 (N_20516,N_19527,N_19791);
or U20517 (N_20517,N_19750,N_19950);
or U20518 (N_20518,N_19535,N_19851);
nand U20519 (N_20519,N_19892,N_19661);
and U20520 (N_20520,N_19709,N_19833);
xnor U20521 (N_20521,N_19444,N_19877);
nand U20522 (N_20522,N_19450,N_19829);
nand U20523 (N_20523,N_19401,N_19916);
nor U20524 (N_20524,N_19452,N_19815);
or U20525 (N_20525,N_19798,N_19385);
nor U20526 (N_20526,N_19592,N_19767);
xor U20527 (N_20527,N_19444,N_19468);
and U20528 (N_20528,N_19983,N_19485);
or U20529 (N_20529,N_19607,N_19479);
nor U20530 (N_20530,N_19840,N_19488);
and U20531 (N_20531,N_19902,N_19816);
or U20532 (N_20532,N_19437,N_19469);
and U20533 (N_20533,N_19646,N_19821);
nand U20534 (N_20534,N_19764,N_19644);
or U20535 (N_20535,N_19504,N_19805);
xnor U20536 (N_20536,N_19532,N_19634);
or U20537 (N_20537,N_19447,N_19922);
and U20538 (N_20538,N_19965,N_19885);
or U20539 (N_20539,N_19390,N_19792);
nand U20540 (N_20540,N_19427,N_19635);
or U20541 (N_20541,N_19651,N_19974);
nand U20542 (N_20542,N_19791,N_19879);
nand U20543 (N_20543,N_19788,N_19935);
xnor U20544 (N_20544,N_19712,N_19643);
xnor U20545 (N_20545,N_19818,N_19704);
or U20546 (N_20546,N_19484,N_19676);
and U20547 (N_20547,N_19894,N_19519);
xnor U20548 (N_20548,N_19983,N_19686);
and U20549 (N_20549,N_19746,N_19934);
nand U20550 (N_20550,N_19711,N_19392);
nand U20551 (N_20551,N_19467,N_19587);
and U20552 (N_20552,N_19531,N_19832);
nand U20553 (N_20553,N_19709,N_19835);
and U20554 (N_20554,N_19646,N_19512);
or U20555 (N_20555,N_19688,N_19790);
xor U20556 (N_20556,N_19625,N_19957);
xor U20557 (N_20557,N_19975,N_19749);
xnor U20558 (N_20558,N_19702,N_19968);
nand U20559 (N_20559,N_19742,N_19995);
or U20560 (N_20560,N_19924,N_19636);
nor U20561 (N_20561,N_19547,N_19624);
or U20562 (N_20562,N_19481,N_19663);
xor U20563 (N_20563,N_19906,N_19558);
xnor U20564 (N_20564,N_19691,N_19426);
nor U20565 (N_20565,N_19556,N_19413);
and U20566 (N_20566,N_19604,N_19786);
xnor U20567 (N_20567,N_19611,N_19445);
nand U20568 (N_20568,N_19943,N_19685);
nand U20569 (N_20569,N_19670,N_19956);
nor U20570 (N_20570,N_19448,N_19551);
and U20571 (N_20571,N_19808,N_19414);
and U20572 (N_20572,N_19977,N_19709);
xor U20573 (N_20573,N_19725,N_19843);
or U20574 (N_20574,N_19982,N_19422);
or U20575 (N_20575,N_19880,N_19811);
nand U20576 (N_20576,N_19902,N_19381);
or U20577 (N_20577,N_19862,N_19498);
xnor U20578 (N_20578,N_19890,N_19968);
nor U20579 (N_20579,N_19977,N_19799);
xnor U20580 (N_20580,N_19732,N_19955);
xnor U20581 (N_20581,N_19986,N_19746);
xor U20582 (N_20582,N_19901,N_19630);
or U20583 (N_20583,N_19942,N_19687);
xnor U20584 (N_20584,N_19448,N_19614);
nor U20585 (N_20585,N_19979,N_19516);
xor U20586 (N_20586,N_19771,N_19877);
or U20587 (N_20587,N_19584,N_19377);
nand U20588 (N_20588,N_19470,N_19970);
or U20589 (N_20589,N_19905,N_19817);
nand U20590 (N_20590,N_19414,N_19791);
xnor U20591 (N_20591,N_19751,N_19916);
xnor U20592 (N_20592,N_19651,N_19768);
nor U20593 (N_20593,N_19971,N_19589);
xnor U20594 (N_20594,N_19690,N_19446);
nor U20595 (N_20595,N_19896,N_19773);
and U20596 (N_20596,N_19825,N_19974);
and U20597 (N_20597,N_19725,N_19691);
nor U20598 (N_20598,N_19577,N_19517);
xor U20599 (N_20599,N_19467,N_19547);
or U20600 (N_20600,N_19849,N_19594);
or U20601 (N_20601,N_19942,N_19526);
nand U20602 (N_20602,N_19787,N_19562);
xnor U20603 (N_20603,N_19537,N_19731);
xor U20604 (N_20604,N_19508,N_19828);
or U20605 (N_20605,N_19753,N_19813);
nand U20606 (N_20606,N_19865,N_19708);
nand U20607 (N_20607,N_19562,N_19972);
nor U20608 (N_20608,N_19715,N_19477);
or U20609 (N_20609,N_19743,N_19752);
nor U20610 (N_20610,N_19777,N_19914);
or U20611 (N_20611,N_19678,N_19518);
nand U20612 (N_20612,N_19520,N_19742);
and U20613 (N_20613,N_19643,N_19919);
or U20614 (N_20614,N_19403,N_19419);
and U20615 (N_20615,N_19831,N_19813);
xor U20616 (N_20616,N_19765,N_19823);
xnor U20617 (N_20617,N_19864,N_19592);
nand U20618 (N_20618,N_19843,N_19447);
and U20619 (N_20619,N_19406,N_19469);
nand U20620 (N_20620,N_19725,N_19998);
nor U20621 (N_20621,N_19734,N_19933);
and U20622 (N_20622,N_19497,N_19656);
and U20623 (N_20623,N_19970,N_19607);
and U20624 (N_20624,N_19773,N_19820);
nand U20625 (N_20625,N_20605,N_20273);
or U20626 (N_20626,N_20322,N_20381);
nor U20627 (N_20627,N_20043,N_20317);
xor U20628 (N_20628,N_20556,N_20230);
nand U20629 (N_20629,N_20595,N_20136);
xnor U20630 (N_20630,N_20284,N_20597);
and U20631 (N_20631,N_20165,N_20151);
and U20632 (N_20632,N_20326,N_20430);
and U20633 (N_20633,N_20333,N_20563);
xnor U20634 (N_20634,N_20603,N_20443);
nand U20635 (N_20635,N_20371,N_20542);
xnor U20636 (N_20636,N_20211,N_20616);
or U20637 (N_20637,N_20120,N_20567);
nor U20638 (N_20638,N_20503,N_20184);
or U20639 (N_20639,N_20152,N_20299);
nand U20640 (N_20640,N_20548,N_20046);
xnor U20641 (N_20641,N_20144,N_20604);
nand U20642 (N_20642,N_20358,N_20301);
nand U20643 (N_20643,N_20335,N_20412);
xor U20644 (N_20644,N_20400,N_20467);
and U20645 (N_20645,N_20027,N_20159);
xnor U20646 (N_20646,N_20235,N_20303);
nand U20647 (N_20647,N_20613,N_20300);
and U20648 (N_20648,N_20294,N_20247);
and U20649 (N_20649,N_20407,N_20615);
and U20650 (N_20650,N_20296,N_20608);
or U20651 (N_20651,N_20111,N_20137);
nand U20652 (N_20652,N_20025,N_20426);
nand U20653 (N_20653,N_20492,N_20131);
nor U20654 (N_20654,N_20589,N_20479);
and U20655 (N_20655,N_20188,N_20341);
xor U20656 (N_20656,N_20254,N_20245);
and U20657 (N_20657,N_20419,N_20310);
xnor U20658 (N_20658,N_20531,N_20553);
or U20659 (N_20659,N_20013,N_20576);
or U20660 (N_20660,N_20231,N_20432);
xor U20661 (N_20661,N_20440,N_20242);
or U20662 (N_20662,N_20620,N_20126);
and U20663 (N_20663,N_20028,N_20601);
and U20664 (N_20664,N_20219,N_20554);
nor U20665 (N_20665,N_20007,N_20033);
nand U20666 (N_20666,N_20324,N_20173);
nand U20667 (N_20667,N_20463,N_20591);
xnor U20668 (N_20668,N_20030,N_20402);
and U20669 (N_20669,N_20186,N_20337);
xnor U20670 (N_20670,N_20011,N_20330);
nor U20671 (N_20671,N_20427,N_20020);
nand U20672 (N_20672,N_20372,N_20157);
xor U20673 (N_20673,N_20285,N_20134);
nor U20674 (N_20674,N_20583,N_20228);
xnor U20675 (N_20675,N_20225,N_20023);
and U20676 (N_20676,N_20451,N_20405);
nor U20677 (N_20677,N_20218,N_20229);
nand U20678 (N_20678,N_20562,N_20175);
nand U20679 (N_20679,N_20431,N_20507);
or U20680 (N_20680,N_20267,N_20316);
xnor U20681 (N_20681,N_20297,N_20077);
or U20682 (N_20682,N_20318,N_20329);
nand U20683 (N_20683,N_20001,N_20521);
or U20684 (N_20684,N_20308,N_20256);
or U20685 (N_20685,N_20206,N_20176);
nand U20686 (N_20686,N_20534,N_20529);
or U20687 (N_20687,N_20018,N_20055);
or U20688 (N_20688,N_20403,N_20573);
or U20689 (N_20689,N_20350,N_20449);
or U20690 (N_20690,N_20113,N_20362);
or U20691 (N_20691,N_20085,N_20196);
and U20692 (N_20692,N_20496,N_20532);
or U20693 (N_20693,N_20410,N_20281);
nor U20694 (N_20694,N_20227,N_20074);
and U20695 (N_20695,N_20088,N_20476);
nand U20696 (N_20696,N_20581,N_20278);
and U20697 (N_20697,N_20580,N_20309);
nand U20698 (N_20698,N_20209,N_20455);
nor U20699 (N_20699,N_20109,N_20079);
xor U20700 (N_20700,N_20050,N_20198);
or U20701 (N_20701,N_20374,N_20295);
nand U20702 (N_20702,N_20552,N_20068);
nor U20703 (N_20703,N_20090,N_20586);
and U20704 (N_20704,N_20272,N_20514);
nand U20705 (N_20705,N_20446,N_20429);
nand U20706 (N_20706,N_20289,N_20205);
xnor U20707 (N_20707,N_20389,N_20453);
and U20708 (N_20708,N_20384,N_20445);
or U20709 (N_20709,N_20009,N_20448);
nand U20710 (N_20710,N_20064,N_20210);
xor U20711 (N_20711,N_20288,N_20142);
xor U20712 (N_20712,N_20150,N_20207);
or U20713 (N_20713,N_20197,N_20490);
and U20714 (N_20714,N_20241,N_20060);
or U20715 (N_20715,N_20199,N_20240);
xnor U20716 (N_20716,N_20472,N_20355);
or U20717 (N_20717,N_20481,N_20038);
xor U20718 (N_20718,N_20270,N_20559);
or U20719 (N_20719,N_20332,N_20338);
nor U20720 (N_20720,N_20202,N_20590);
xnor U20721 (N_20721,N_20408,N_20065);
nor U20722 (N_20722,N_20238,N_20364);
or U20723 (N_20723,N_20571,N_20100);
and U20724 (N_20724,N_20162,N_20261);
and U20725 (N_20725,N_20491,N_20139);
nor U20726 (N_20726,N_20266,N_20054);
and U20727 (N_20727,N_20457,N_20473);
and U20728 (N_20728,N_20411,N_20342);
nor U20729 (N_20729,N_20171,N_20462);
xor U20730 (N_20730,N_20089,N_20086);
or U20731 (N_20731,N_20524,N_20480);
nor U20732 (N_20732,N_20359,N_20452);
and U20733 (N_20733,N_20437,N_20494);
xor U20734 (N_20734,N_20406,N_20127);
and U20735 (N_20735,N_20118,N_20277);
nor U20736 (N_20736,N_20083,N_20026);
and U20737 (N_20737,N_20203,N_20349);
or U20738 (N_20738,N_20078,N_20062);
or U20739 (N_20739,N_20216,N_20268);
nand U20740 (N_20740,N_20459,N_20502);
and U20741 (N_20741,N_20593,N_20170);
nor U20742 (N_20742,N_20376,N_20510);
nand U20743 (N_20743,N_20233,N_20153);
nand U20744 (N_20744,N_20505,N_20387);
xor U20745 (N_20745,N_20485,N_20380);
and U20746 (N_20746,N_20409,N_20461);
xor U20747 (N_20747,N_20114,N_20577);
or U20748 (N_20748,N_20515,N_20558);
nand U20749 (N_20749,N_20262,N_20071);
nand U20750 (N_20750,N_20061,N_20423);
nand U20751 (N_20751,N_20167,N_20444);
nand U20752 (N_20752,N_20325,N_20339);
nor U20753 (N_20753,N_20464,N_20069);
nor U20754 (N_20754,N_20477,N_20222);
xnor U20755 (N_20755,N_20178,N_20257);
nor U20756 (N_20756,N_20253,N_20331);
xnor U20757 (N_20757,N_20200,N_20124);
xnor U20758 (N_20758,N_20236,N_20279);
and U20759 (N_20759,N_20094,N_20450);
xor U20760 (N_20760,N_20536,N_20592);
nor U20761 (N_20761,N_20187,N_20441);
xnor U20762 (N_20762,N_20158,N_20223);
nor U20763 (N_20763,N_20504,N_20495);
or U20764 (N_20764,N_20140,N_20067);
nor U20765 (N_20765,N_20422,N_20511);
xnor U20766 (N_20766,N_20195,N_20311);
and U20767 (N_20767,N_20383,N_20382);
or U20768 (N_20768,N_20081,N_20470);
and U20769 (N_20769,N_20221,N_20006);
nor U20770 (N_20770,N_20123,N_20133);
xor U20771 (N_20771,N_20180,N_20312);
or U20772 (N_20772,N_20397,N_20469);
and U20773 (N_20773,N_20447,N_20465);
and U20774 (N_20774,N_20214,N_20049);
nor U20775 (N_20775,N_20244,N_20174);
nand U20776 (N_20776,N_20039,N_20621);
nor U20777 (N_20777,N_20500,N_20304);
nor U20778 (N_20778,N_20599,N_20122);
nor U20779 (N_20779,N_20129,N_20293);
xnor U20780 (N_20780,N_20141,N_20594);
or U20781 (N_20781,N_20442,N_20414);
or U20782 (N_20782,N_20066,N_20619);
nor U20783 (N_20783,N_20258,N_20572);
xnor U20784 (N_20784,N_20008,N_20164);
nor U20785 (N_20785,N_20399,N_20569);
or U20786 (N_20786,N_20475,N_20428);
xnor U20787 (N_20787,N_20080,N_20566);
nand U20788 (N_20788,N_20119,N_20624);
and U20789 (N_20789,N_20377,N_20353);
xor U20790 (N_20790,N_20224,N_20533);
nor U20791 (N_20791,N_20024,N_20356);
nand U20792 (N_20792,N_20550,N_20468);
xnor U20793 (N_20793,N_20386,N_20501);
nand U20794 (N_20794,N_20488,N_20348);
or U20795 (N_20795,N_20498,N_20345);
xnor U20796 (N_20796,N_20147,N_20314);
and U20797 (N_20797,N_20249,N_20103);
or U20798 (N_20798,N_20075,N_20041);
nand U20799 (N_20799,N_20280,N_20252);
and U20800 (N_20800,N_20555,N_20105);
or U20801 (N_20801,N_20226,N_20582);
nor U20802 (N_20802,N_20395,N_20035);
nor U20803 (N_20803,N_20194,N_20436);
nand U20804 (N_20804,N_20037,N_20019);
nor U20805 (N_20805,N_20336,N_20042);
or U20806 (N_20806,N_20574,N_20396);
xor U20807 (N_20807,N_20513,N_20421);
xnor U20808 (N_20808,N_20177,N_20357);
and U20809 (N_20809,N_20528,N_20286);
and U20810 (N_20810,N_20391,N_20320);
nor U20811 (N_20811,N_20466,N_20096);
and U20812 (N_20812,N_20438,N_20092);
and U20813 (N_20813,N_20319,N_20204);
nor U20814 (N_20814,N_20185,N_20526);
and U20815 (N_20815,N_20212,N_20146);
and U20816 (N_20816,N_20598,N_20036);
nor U20817 (N_20817,N_20541,N_20328);
xor U20818 (N_20818,N_20539,N_20366);
and U20819 (N_20819,N_20456,N_20535);
xnor U20820 (N_20820,N_20302,N_20561);
or U20821 (N_20821,N_20298,N_20259);
xor U20822 (N_20822,N_20220,N_20327);
and U20823 (N_20823,N_20022,N_20243);
and U20824 (N_20824,N_20138,N_20029);
nand U20825 (N_20825,N_20208,N_20557);
or U20826 (N_20826,N_20568,N_20365);
xor U20827 (N_20827,N_20392,N_20570);
or U20828 (N_20828,N_20232,N_20527);
nor U20829 (N_20829,N_20191,N_20073);
and U20830 (N_20830,N_20263,N_20082);
or U20831 (N_20831,N_20367,N_20506);
nor U20832 (N_20832,N_20084,N_20596);
and U20833 (N_20833,N_20003,N_20032);
and U20834 (N_20834,N_20095,N_20606);
xnor U20835 (N_20835,N_20537,N_20201);
nor U20836 (N_20836,N_20179,N_20315);
and U20837 (N_20837,N_20617,N_20148);
nand U20838 (N_20838,N_20340,N_20017);
and U20839 (N_20839,N_20239,N_20250);
xor U20840 (N_20840,N_20493,N_20121);
and U20841 (N_20841,N_20360,N_20434);
or U20842 (N_20842,N_20474,N_20471);
xor U20843 (N_20843,N_20487,N_20149);
nand U20844 (N_20844,N_20394,N_20098);
and U20845 (N_20845,N_20363,N_20093);
nor U20846 (N_20846,N_20269,N_20588);
nand U20847 (N_20847,N_20587,N_20519);
or U20848 (N_20848,N_20047,N_20565);
nand U20849 (N_20849,N_20313,N_20016);
and U20850 (N_20850,N_20489,N_20482);
xnor U20851 (N_20851,N_20217,N_20040);
nand U20852 (N_20852,N_20305,N_20540);
and U20853 (N_20853,N_20622,N_20215);
and U20854 (N_20854,N_20101,N_20497);
nor U20855 (N_20855,N_20546,N_20059);
xnor U20856 (N_20856,N_20015,N_20156);
and U20857 (N_20857,N_20182,N_20373);
nor U20858 (N_20858,N_20145,N_20610);
or U20859 (N_20859,N_20237,N_20058);
and U20860 (N_20860,N_20416,N_20183);
nor U20861 (N_20861,N_20192,N_20125);
or U20862 (N_20862,N_20307,N_20002);
nor U20863 (N_20863,N_20160,N_20344);
or U20864 (N_20864,N_20021,N_20255);
or U20865 (N_20865,N_20271,N_20602);
nand U20866 (N_20866,N_20614,N_20623);
or U20867 (N_20867,N_20169,N_20283);
and U20868 (N_20868,N_20045,N_20545);
and U20869 (N_20869,N_20117,N_20306);
and U20870 (N_20870,N_20135,N_20520);
nand U20871 (N_20871,N_20274,N_20424);
xnor U20872 (N_20872,N_20034,N_20385);
or U20873 (N_20873,N_20347,N_20251);
or U20874 (N_20874,N_20612,N_20560);
or U20875 (N_20875,N_20234,N_20106);
or U20876 (N_20876,N_20110,N_20609);
nand U20877 (N_20877,N_20478,N_20053);
nand U20878 (N_20878,N_20418,N_20010);
and U20879 (N_20879,N_20543,N_20091);
or U20880 (N_20880,N_20014,N_20275);
nand U20881 (N_20881,N_20172,N_20549);
nand U20882 (N_20882,N_20458,N_20056);
nor U20883 (N_20883,N_20530,N_20070);
nand U20884 (N_20884,N_20213,N_20130);
xor U20885 (N_20885,N_20525,N_20343);
and U20886 (N_20886,N_20404,N_20107);
xor U20887 (N_20887,N_20097,N_20163);
xor U20888 (N_20888,N_20181,N_20460);
or U20889 (N_20889,N_20099,N_20516);
nor U20890 (N_20890,N_20352,N_20547);
or U20891 (N_20891,N_20102,N_20484);
xnor U20892 (N_20892,N_20260,N_20522);
and U20893 (N_20893,N_20415,N_20076);
nor U20894 (N_20894,N_20551,N_20005);
nor U20895 (N_20895,N_20143,N_20112);
nand U20896 (N_20896,N_20057,N_20004);
nor U20897 (N_20897,N_20413,N_20265);
or U20898 (N_20898,N_20439,N_20499);
or U20899 (N_20899,N_20323,N_20585);
and U20900 (N_20900,N_20321,N_20607);
and U20901 (N_20901,N_20104,N_20346);
xnor U20902 (N_20902,N_20388,N_20051);
xor U20903 (N_20903,N_20509,N_20115);
xnor U20904 (N_20904,N_20287,N_20128);
or U20905 (N_20905,N_20370,N_20190);
xnor U20906 (N_20906,N_20564,N_20048);
or U20907 (N_20907,N_20401,N_20155);
nor U20908 (N_20908,N_20378,N_20282);
nand U20909 (N_20909,N_20417,N_20486);
or U20910 (N_20910,N_20246,N_20575);
nor U20911 (N_20911,N_20063,N_20512);
nand U20912 (N_20912,N_20523,N_20368);
nand U20913 (N_20913,N_20264,N_20618);
or U20914 (N_20914,N_20454,N_20334);
nor U20915 (N_20915,N_20390,N_20248);
nand U20916 (N_20916,N_20012,N_20579);
xnor U20917 (N_20917,N_20544,N_20369);
nand U20918 (N_20918,N_20398,N_20168);
xnor U20919 (N_20919,N_20578,N_20351);
nand U20920 (N_20920,N_20600,N_20154);
xor U20921 (N_20921,N_20518,N_20087);
or U20922 (N_20922,N_20193,N_20276);
nor U20923 (N_20923,N_20291,N_20483);
or U20924 (N_20924,N_20031,N_20354);
and U20925 (N_20925,N_20072,N_20166);
and U20926 (N_20926,N_20116,N_20161);
xor U20927 (N_20927,N_20433,N_20189);
and U20928 (N_20928,N_20052,N_20508);
or U20929 (N_20929,N_20290,N_20538);
xor U20930 (N_20930,N_20000,N_20584);
and U20931 (N_20931,N_20361,N_20132);
or U20932 (N_20932,N_20375,N_20435);
nand U20933 (N_20933,N_20292,N_20108);
xnor U20934 (N_20934,N_20393,N_20379);
or U20935 (N_20935,N_20517,N_20611);
nor U20936 (N_20936,N_20425,N_20420);
nand U20937 (N_20937,N_20044,N_20386);
or U20938 (N_20938,N_20228,N_20092);
or U20939 (N_20939,N_20535,N_20373);
or U20940 (N_20940,N_20385,N_20102);
nor U20941 (N_20941,N_20160,N_20156);
xnor U20942 (N_20942,N_20367,N_20031);
xnor U20943 (N_20943,N_20370,N_20525);
nand U20944 (N_20944,N_20422,N_20258);
or U20945 (N_20945,N_20143,N_20188);
or U20946 (N_20946,N_20016,N_20354);
nand U20947 (N_20947,N_20552,N_20261);
xor U20948 (N_20948,N_20280,N_20411);
or U20949 (N_20949,N_20074,N_20172);
nor U20950 (N_20950,N_20125,N_20213);
xnor U20951 (N_20951,N_20594,N_20542);
or U20952 (N_20952,N_20045,N_20396);
and U20953 (N_20953,N_20044,N_20470);
xor U20954 (N_20954,N_20098,N_20113);
nor U20955 (N_20955,N_20141,N_20244);
xor U20956 (N_20956,N_20575,N_20509);
nor U20957 (N_20957,N_20257,N_20436);
or U20958 (N_20958,N_20502,N_20015);
xor U20959 (N_20959,N_20160,N_20312);
nor U20960 (N_20960,N_20235,N_20149);
and U20961 (N_20961,N_20572,N_20381);
xor U20962 (N_20962,N_20023,N_20531);
or U20963 (N_20963,N_20174,N_20055);
xnor U20964 (N_20964,N_20479,N_20323);
or U20965 (N_20965,N_20574,N_20264);
nor U20966 (N_20966,N_20302,N_20375);
xor U20967 (N_20967,N_20190,N_20199);
nor U20968 (N_20968,N_20078,N_20298);
nand U20969 (N_20969,N_20615,N_20032);
xnor U20970 (N_20970,N_20431,N_20274);
xnor U20971 (N_20971,N_20456,N_20116);
or U20972 (N_20972,N_20198,N_20375);
or U20973 (N_20973,N_20150,N_20033);
nand U20974 (N_20974,N_20198,N_20097);
nand U20975 (N_20975,N_20186,N_20531);
and U20976 (N_20976,N_20365,N_20351);
nand U20977 (N_20977,N_20452,N_20252);
and U20978 (N_20978,N_20511,N_20514);
and U20979 (N_20979,N_20009,N_20058);
or U20980 (N_20980,N_20586,N_20325);
and U20981 (N_20981,N_20134,N_20535);
and U20982 (N_20982,N_20003,N_20533);
and U20983 (N_20983,N_20425,N_20203);
and U20984 (N_20984,N_20002,N_20415);
nand U20985 (N_20985,N_20556,N_20219);
xnor U20986 (N_20986,N_20223,N_20377);
nor U20987 (N_20987,N_20363,N_20095);
nand U20988 (N_20988,N_20211,N_20265);
nor U20989 (N_20989,N_20328,N_20276);
or U20990 (N_20990,N_20455,N_20129);
or U20991 (N_20991,N_20182,N_20158);
nand U20992 (N_20992,N_20255,N_20393);
xnor U20993 (N_20993,N_20458,N_20424);
or U20994 (N_20994,N_20550,N_20578);
nor U20995 (N_20995,N_20496,N_20082);
and U20996 (N_20996,N_20290,N_20389);
and U20997 (N_20997,N_20550,N_20330);
and U20998 (N_20998,N_20087,N_20434);
and U20999 (N_20999,N_20409,N_20298);
nor U21000 (N_21000,N_20016,N_20364);
or U21001 (N_21001,N_20025,N_20431);
and U21002 (N_21002,N_20037,N_20337);
and U21003 (N_21003,N_20565,N_20407);
nand U21004 (N_21004,N_20159,N_20026);
and U21005 (N_21005,N_20497,N_20202);
and U21006 (N_21006,N_20448,N_20218);
and U21007 (N_21007,N_20303,N_20270);
and U21008 (N_21008,N_20387,N_20225);
xor U21009 (N_21009,N_20548,N_20614);
nand U21010 (N_21010,N_20355,N_20136);
or U21011 (N_21011,N_20551,N_20084);
and U21012 (N_21012,N_20008,N_20457);
xnor U21013 (N_21013,N_20566,N_20260);
and U21014 (N_21014,N_20335,N_20529);
xnor U21015 (N_21015,N_20275,N_20461);
nand U21016 (N_21016,N_20036,N_20138);
and U21017 (N_21017,N_20312,N_20428);
or U21018 (N_21018,N_20012,N_20462);
xor U21019 (N_21019,N_20332,N_20311);
nand U21020 (N_21020,N_20357,N_20611);
and U21021 (N_21021,N_20324,N_20488);
and U21022 (N_21022,N_20031,N_20593);
xnor U21023 (N_21023,N_20036,N_20002);
and U21024 (N_21024,N_20613,N_20023);
or U21025 (N_21025,N_20330,N_20099);
xnor U21026 (N_21026,N_20270,N_20213);
nor U21027 (N_21027,N_20048,N_20599);
and U21028 (N_21028,N_20066,N_20589);
xor U21029 (N_21029,N_20362,N_20329);
xnor U21030 (N_21030,N_20017,N_20388);
and U21031 (N_21031,N_20171,N_20115);
nand U21032 (N_21032,N_20436,N_20540);
nor U21033 (N_21033,N_20056,N_20307);
and U21034 (N_21034,N_20556,N_20118);
or U21035 (N_21035,N_20170,N_20351);
and U21036 (N_21036,N_20191,N_20037);
nor U21037 (N_21037,N_20549,N_20416);
xor U21038 (N_21038,N_20374,N_20335);
xnor U21039 (N_21039,N_20443,N_20323);
and U21040 (N_21040,N_20050,N_20511);
nand U21041 (N_21041,N_20160,N_20269);
and U21042 (N_21042,N_20365,N_20489);
xnor U21043 (N_21043,N_20420,N_20439);
nand U21044 (N_21044,N_20620,N_20130);
xor U21045 (N_21045,N_20504,N_20083);
nand U21046 (N_21046,N_20049,N_20272);
and U21047 (N_21047,N_20262,N_20000);
and U21048 (N_21048,N_20555,N_20587);
nand U21049 (N_21049,N_20196,N_20121);
or U21050 (N_21050,N_20025,N_20347);
xnor U21051 (N_21051,N_20287,N_20404);
nor U21052 (N_21052,N_20452,N_20516);
nand U21053 (N_21053,N_20179,N_20251);
or U21054 (N_21054,N_20440,N_20337);
or U21055 (N_21055,N_20594,N_20089);
or U21056 (N_21056,N_20200,N_20345);
nand U21057 (N_21057,N_20186,N_20134);
and U21058 (N_21058,N_20015,N_20049);
xnor U21059 (N_21059,N_20162,N_20015);
or U21060 (N_21060,N_20006,N_20594);
xor U21061 (N_21061,N_20356,N_20329);
nand U21062 (N_21062,N_20316,N_20000);
or U21063 (N_21063,N_20605,N_20193);
nand U21064 (N_21064,N_20228,N_20456);
nor U21065 (N_21065,N_20251,N_20442);
nor U21066 (N_21066,N_20046,N_20417);
nor U21067 (N_21067,N_20471,N_20189);
nor U21068 (N_21068,N_20151,N_20364);
and U21069 (N_21069,N_20276,N_20103);
or U21070 (N_21070,N_20066,N_20582);
and U21071 (N_21071,N_20203,N_20008);
xor U21072 (N_21072,N_20473,N_20439);
nand U21073 (N_21073,N_20195,N_20529);
xnor U21074 (N_21074,N_20531,N_20165);
xnor U21075 (N_21075,N_20283,N_20476);
nand U21076 (N_21076,N_20196,N_20289);
xnor U21077 (N_21077,N_20118,N_20081);
nand U21078 (N_21078,N_20250,N_20535);
nor U21079 (N_21079,N_20571,N_20545);
nand U21080 (N_21080,N_20440,N_20158);
nor U21081 (N_21081,N_20216,N_20073);
xor U21082 (N_21082,N_20614,N_20500);
or U21083 (N_21083,N_20516,N_20496);
nand U21084 (N_21084,N_20406,N_20289);
nor U21085 (N_21085,N_20172,N_20623);
and U21086 (N_21086,N_20168,N_20359);
nand U21087 (N_21087,N_20376,N_20356);
or U21088 (N_21088,N_20428,N_20370);
xor U21089 (N_21089,N_20250,N_20068);
and U21090 (N_21090,N_20548,N_20295);
xor U21091 (N_21091,N_20233,N_20498);
nand U21092 (N_21092,N_20153,N_20307);
xnor U21093 (N_21093,N_20298,N_20290);
nand U21094 (N_21094,N_20315,N_20408);
and U21095 (N_21095,N_20592,N_20463);
and U21096 (N_21096,N_20121,N_20104);
nand U21097 (N_21097,N_20395,N_20412);
nor U21098 (N_21098,N_20315,N_20519);
xor U21099 (N_21099,N_20059,N_20291);
and U21100 (N_21100,N_20559,N_20206);
and U21101 (N_21101,N_20284,N_20585);
or U21102 (N_21102,N_20062,N_20175);
xnor U21103 (N_21103,N_20552,N_20604);
xor U21104 (N_21104,N_20477,N_20473);
and U21105 (N_21105,N_20571,N_20601);
xor U21106 (N_21106,N_20494,N_20429);
nor U21107 (N_21107,N_20498,N_20347);
nor U21108 (N_21108,N_20437,N_20252);
and U21109 (N_21109,N_20624,N_20558);
or U21110 (N_21110,N_20422,N_20467);
nor U21111 (N_21111,N_20493,N_20613);
nor U21112 (N_21112,N_20080,N_20212);
nand U21113 (N_21113,N_20232,N_20536);
xnor U21114 (N_21114,N_20122,N_20002);
or U21115 (N_21115,N_20613,N_20246);
nor U21116 (N_21116,N_20279,N_20546);
xor U21117 (N_21117,N_20215,N_20369);
or U21118 (N_21118,N_20339,N_20257);
nor U21119 (N_21119,N_20071,N_20529);
nor U21120 (N_21120,N_20066,N_20378);
nand U21121 (N_21121,N_20481,N_20555);
and U21122 (N_21122,N_20571,N_20466);
nor U21123 (N_21123,N_20396,N_20458);
xnor U21124 (N_21124,N_20575,N_20338);
nor U21125 (N_21125,N_20041,N_20296);
nand U21126 (N_21126,N_20469,N_20527);
xnor U21127 (N_21127,N_20527,N_20479);
nor U21128 (N_21128,N_20406,N_20475);
and U21129 (N_21129,N_20575,N_20352);
xor U21130 (N_21130,N_20585,N_20282);
xnor U21131 (N_21131,N_20423,N_20208);
xor U21132 (N_21132,N_20089,N_20255);
and U21133 (N_21133,N_20299,N_20069);
xnor U21134 (N_21134,N_20055,N_20540);
nand U21135 (N_21135,N_20109,N_20038);
and U21136 (N_21136,N_20578,N_20144);
or U21137 (N_21137,N_20300,N_20255);
or U21138 (N_21138,N_20323,N_20091);
xnor U21139 (N_21139,N_20582,N_20420);
nor U21140 (N_21140,N_20164,N_20078);
nor U21141 (N_21141,N_20584,N_20161);
xor U21142 (N_21142,N_20502,N_20117);
or U21143 (N_21143,N_20535,N_20122);
nor U21144 (N_21144,N_20270,N_20006);
nand U21145 (N_21145,N_20533,N_20036);
nor U21146 (N_21146,N_20143,N_20545);
and U21147 (N_21147,N_20141,N_20618);
and U21148 (N_21148,N_20201,N_20507);
xor U21149 (N_21149,N_20103,N_20389);
nor U21150 (N_21150,N_20114,N_20208);
or U21151 (N_21151,N_20583,N_20096);
and U21152 (N_21152,N_20406,N_20257);
and U21153 (N_21153,N_20162,N_20242);
nand U21154 (N_21154,N_20608,N_20430);
or U21155 (N_21155,N_20388,N_20381);
and U21156 (N_21156,N_20461,N_20555);
nor U21157 (N_21157,N_20263,N_20496);
nor U21158 (N_21158,N_20136,N_20224);
xnor U21159 (N_21159,N_20482,N_20126);
nor U21160 (N_21160,N_20237,N_20206);
nand U21161 (N_21161,N_20482,N_20500);
xor U21162 (N_21162,N_20591,N_20464);
xor U21163 (N_21163,N_20358,N_20609);
and U21164 (N_21164,N_20427,N_20189);
or U21165 (N_21165,N_20624,N_20259);
and U21166 (N_21166,N_20348,N_20495);
nor U21167 (N_21167,N_20415,N_20305);
and U21168 (N_21168,N_20139,N_20455);
or U21169 (N_21169,N_20020,N_20360);
and U21170 (N_21170,N_20456,N_20488);
and U21171 (N_21171,N_20198,N_20341);
xnor U21172 (N_21172,N_20161,N_20162);
xor U21173 (N_21173,N_20054,N_20062);
xor U21174 (N_21174,N_20269,N_20242);
nand U21175 (N_21175,N_20304,N_20355);
and U21176 (N_21176,N_20519,N_20091);
xor U21177 (N_21177,N_20409,N_20144);
nor U21178 (N_21178,N_20531,N_20592);
and U21179 (N_21179,N_20240,N_20481);
and U21180 (N_21180,N_20175,N_20050);
xnor U21181 (N_21181,N_20254,N_20004);
or U21182 (N_21182,N_20277,N_20216);
and U21183 (N_21183,N_20287,N_20234);
xnor U21184 (N_21184,N_20166,N_20075);
xnor U21185 (N_21185,N_20391,N_20319);
and U21186 (N_21186,N_20518,N_20091);
nor U21187 (N_21187,N_20046,N_20073);
and U21188 (N_21188,N_20553,N_20079);
and U21189 (N_21189,N_20111,N_20231);
nor U21190 (N_21190,N_20619,N_20048);
nor U21191 (N_21191,N_20113,N_20101);
nor U21192 (N_21192,N_20110,N_20460);
xor U21193 (N_21193,N_20165,N_20262);
or U21194 (N_21194,N_20136,N_20377);
nor U21195 (N_21195,N_20046,N_20542);
nand U21196 (N_21196,N_20370,N_20582);
xnor U21197 (N_21197,N_20051,N_20042);
or U21198 (N_21198,N_20516,N_20507);
nand U21199 (N_21199,N_20263,N_20602);
and U21200 (N_21200,N_20419,N_20022);
xnor U21201 (N_21201,N_20172,N_20237);
nor U21202 (N_21202,N_20396,N_20602);
xnor U21203 (N_21203,N_20616,N_20090);
or U21204 (N_21204,N_20283,N_20009);
nand U21205 (N_21205,N_20228,N_20291);
nor U21206 (N_21206,N_20012,N_20219);
and U21207 (N_21207,N_20316,N_20455);
or U21208 (N_21208,N_20212,N_20549);
or U21209 (N_21209,N_20344,N_20483);
and U21210 (N_21210,N_20184,N_20573);
nand U21211 (N_21211,N_20098,N_20018);
nor U21212 (N_21212,N_20214,N_20486);
and U21213 (N_21213,N_20234,N_20077);
and U21214 (N_21214,N_20183,N_20469);
and U21215 (N_21215,N_20457,N_20421);
xnor U21216 (N_21216,N_20381,N_20161);
xnor U21217 (N_21217,N_20478,N_20335);
nor U21218 (N_21218,N_20189,N_20512);
nor U21219 (N_21219,N_20205,N_20039);
nand U21220 (N_21220,N_20060,N_20191);
or U21221 (N_21221,N_20618,N_20006);
xor U21222 (N_21222,N_20140,N_20548);
and U21223 (N_21223,N_20484,N_20379);
nand U21224 (N_21224,N_20426,N_20330);
nor U21225 (N_21225,N_20305,N_20077);
and U21226 (N_21226,N_20293,N_20166);
and U21227 (N_21227,N_20219,N_20326);
nor U21228 (N_21228,N_20387,N_20176);
xor U21229 (N_21229,N_20046,N_20209);
xnor U21230 (N_21230,N_20572,N_20101);
xnor U21231 (N_21231,N_20555,N_20319);
or U21232 (N_21232,N_20193,N_20333);
and U21233 (N_21233,N_20468,N_20139);
or U21234 (N_21234,N_20360,N_20194);
or U21235 (N_21235,N_20116,N_20138);
nor U21236 (N_21236,N_20337,N_20587);
nor U21237 (N_21237,N_20513,N_20470);
nand U21238 (N_21238,N_20009,N_20446);
nor U21239 (N_21239,N_20354,N_20042);
nor U21240 (N_21240,N_20585,N_20445);
nor U21241 (N_21241,N_20100,N_20246);
xor U21242 (N_21242,N_20330,N_20322);
or U21243 (N_21243,N_20617,N_20116);
nand U21244 (N_21244,N_20283,N_20459);
nand U21245 (N_21245,N_20585,N_20174);
and U21246 (N_21246,N_20020,N_20027);
or U21247 (N_21247,N_20251,N_20268);
or U21248 (N_21248,N_20431,N_20446);
or U21249 (N_21249,N_20291,N_20555);
and U21250 (N_21250,N_20969,N_20930);
nor U21251 (N_21251,N_21015,N_20861);
and U21252 (N_21252,N_20862,N_20640);
and U21253 (N_21253,N_20763,N_20849);
nand U21254 (N_21254,N_20769,N_21069);
and U21255 (N_21255,N_20725,N_20895);
nand U21256 (N_21256,N_21071,N_20952);
or U21257 (N_21257,N_20652,N_20950);
nor U21258 (N_21258,N_21023,N_20958);
nand U21259 (N_21259,N_20778,N_20834);
nand U21260 (N_21260,N_21065,N_21246);
nor U21261 (N_21261,N_20721,N_20870);
nand U21262 (N_21262,N_20893,N_20888);
nand U21263 (N_21263,N_20634,N_20845);
or U21264 (N_21264,N_20799,N_20875);
and U21265 (N_21265,N_20859,N_21085);
nor U21266 (N_21266,N_21201,N_21185);
or U21267 (N_21267,N_20768,N_21152);
nor U21268 (N_21268,N_20703,N_21012);
or U21269 (N_21269,N_21043,N_20673);
or U21270 (N_21270,N_20663,N_20696);
nor U21271 (N_21271,N_20788,N_20814);
or U21272 (N_21272,N_20737,N_20986);
nand U21273 (N_21273,N_20934,N_20997);
xnor U21274 (N_21274,N_20776,N_20835);
or U21275 (N_21275,N_20828,N_20842);
nor U21276 (N_21276,N_21086,N_21045);
nor U21277 (N_21277,N_20743,N_21180);
or U21278 (N_21278,N_21159,N_20771);
and U21279 (N_21279,N_20912,N_20773);
xnor U21280 (N_21280,N_20797,N_20823);
nand U21281 (N_21281,N_20729,N_21026);
and U21282 (N_21282,N_20745,N_21112);
xor U21283 (N_21283,N_20671,N_20841);
nand U21284 (N_21284,N_21111,N_21144);
xor U21285 (N_21285,N_20960,N_21224);
and U21286 (N_21286,N_20880,N_20804);
xnor U21287 (N_21287,N_20962,N_21237);
and U21288 (N_21288,N_20942,N_21156);
nor U21289 (N_21289,N_20949,N_20976);
and U21290 (N_21290,N_20672,N_20818);
or U21291 (N_21291,N_21054,N_21155);
xor U21292 (N_21292,N_21082,N_21179);
xor U21293 (N_21293,N_20863,N_20808);
or U21294 (N_21294,N_20753,N_20687);
nor U21295 (N_21295,N_20712,N_20813);
nor U21296 (N_21296,N_20898,N_20767);
xor U21297 (N_21297,N_21076,N_21247);
nand U21298 (N_21298,N_20682,N_20750);
xnor U21299 (N_21299,N_21027,N_21164);
or U21300 (N_21300,N_20754,N_20765);
xor U21301 (N_21301,N_21133,N_20921);
and U21302 (N_21302,N_21038,N_21230);
xor U21303 (N_21303,N_21091,N_20832);
nor U21304 (N_21304,N_20747,N_21098);
nor U21305 (N_21305,N_20783,N_20955);
nand U21306 (N_21306,N_20943,N_21048);
or U21307 (N_21307,N_20787,N_21183);
xor U21308 (N_21308,N_20642,N_20654);
nand U21309 (N_21309,N_21209,N_21193);
nor U21310 (N_21310,N_20770,N_21101);
and U21311 (N_21311,N_20900,N_20953);
or U21312 (N_21312,N_21046,N_20857);
nor U21313 (N_21313,N_21149,N_21196);
and U21314 (N_21314,N_20637,N_21050);
and U21315 (N_21315,N_20793,N_21108);
xor U21316 (N_21316,N_21234,N_21088);
and U21317 (N_21317,N_21216,N_21142);
or U21318 (N_21318,N_20669,N_21009);
nor U21319 (N_21319,N_20851,N_20951);
or U21320 (N_21320,N_21102,N_21089);
nor U21321 (N_21321,N_20829,N_20739);
or U21322 (N_21322,N_20760,N_20990);
or U21323 (N_21323,N_20651,N_20931);
xnor U21324 (N_21324,N_20833,N_21211);
or U21325 (N_21325,N_20744,N_21081);
nor U21326 (N_21326,N_20968,N_21030);
nor U21327 (N_21327,N_21148,N_20852);
xnor U21328 (N_21328,N_20944,N_20805);
xnor U21329 (N_21329,N_20741,N_21213);
nand U21330 (N_21330,N_20819,N_21079);
xor U21331 (N_21331,N_21161,N_20831);
nor U21332 (N_21332,N_20702,N_21137);
nand U21333 (N_21333,N_20865,N_21113);
or U21334 (N_21334,N_20887,N_21225);
nor U21335 (N_21335,N_21123,N_20988);
and U21336 (N_21336,N_20885,N_20850);
or U21337 (N_21337,N_20918,N_21244);
nor U21338 (N_21338,N_20653,N_21181);
xor U21339 (N_21339,N_20731,N_21227);
nor U21340 (N_21340,N_21068,N_20670);
or U21341 (N_21341,N_20647,N_21096);
xor U21342 (N_21342,N_20630,N_20704);
nand U21343 (N_21343,N_21075,N_20762);
nand U21344 (N_21344,N_21221,N_20994);
or U21345 (N_21345,N_21125,N_20728);
or U21346 (N_21346,N_21067,N_21190);
nand U21347 (N_21347,N_20959,N_20809);
xor U21348 (N_21348,N_21202,N_21151);
and U21349 (N_21349,N_20926,N_20662);
nor U21350 (N_21350,N_21062,N_20719);
nor U21351 (N_21351,N_20646,N_21210);
nor U21352 (N_21352,N_20800,N_21220);
or U21353 (N_21353,N_20920,N_21172);
or U21354 (N_21354,N_21019,N_21037);
and U21355 (N_21355,N_20681,N_21191);
nand U21356 (N_21356,N_20947,N_20645);
or U21357 (N_21357,N_20825,N_20735);
and U21358 (N_21358,N_20711,N_21212);
and U21359 (N_21359,N_20869,N_21243);
nor U21360 (N_21360,N_21154,N_21014);
or U21361 (N_21361,N_20989,N_20956);
or U21362 (N_21362,N_20977,N_21090);
nor U21363 (N_21363,N_20941,N_21057);
or U21364 (N_21364,N_21248,N_21165);
nand U21365 (N_21365,N_21061,N_20935);
and U21366 (N_21366,N_20734,N_20802);
and U21367 (N_21367,N_20854,N_21004);
xor U21368 (N_21368,N_21130,N_21241);
nand U21369 (N_21369,N_20700,N_21029);
or U21370 (N_21370,N_20812,N_20840);
and U21371 (N_21371,N_21025,N_21117);
nand U21372 (N_21372,N_21097,N_20998);
nand U21373 (N_21373,N_21005,N_20718);
nand U21374 (N_21374,N_21049,N_20925);
xor U21375 (N_21375,N_20665,N_21031);
and U21376 (N_21376,N_21087,N_21240);
and U21377 (N_21377,N_20755,N_20838);
xnor U21378 (N_21378,N_20985,N_21233);
or U21379 (N_21379,N_20633,N_21115);
nor U21380 (N_21380,N_20923,N_20780);
and U21381 (N_21381,N_20713,N_20911);
and U21382 (N_21382,N_21053,N_21018);
and U21383 (N_21383,N_20676,N_20806);
or U21384 (N_21384,N_20684,N_21007);
and U21385 (N_21385,N_21132,N_20904);
xnor U21386 (N_21386,N_20786,N_20933);
xnor U21387 (N_21387,N_20656,N_21214);
nor U21388 (N_21388,N_21093,N_20648);
xnor U21389 (N_21389,N_21083,N_21208);
nor U21390 (N_21390,N_21074,N_21094);
and U21391 (N_21391,N_20903,N_20844);
or U21392 (N_21392,N_20973,N_21186);
nor U21393 (N_21393,N_21135,N_20693);
nor U21394 (N_21394,N_20641,N_20858);
nor U21395 (N_21395,N_20650,N_20864);
xnor U21396 (N_21396,N_21134,N_20679);
or U21397 (N_21397,N_20932,N_21040);
or U21398 (N_21398,N_20625,N_21139);
nand U21399 (N_21399,N_20946,N_20699);
and U21400 (N_21400,N_21016,N_20860);
nor U21401 (N_21401,N_20816,N_21182);
nor U21402 (N_21402,N_20777,N_21175);
and U21403 (N_21403,N_21226,N_20638);
or U21404 (N_21404,N_20709,N_20736);
or U21405 (N_21405,N_21109,N_20766);
xnor U21406 (N_21406,N_21041,N_20678);
nand U21407 (N_21407,N_21222,N_20824);
xnor U21408 (N_21408,N_21022,N_20627);
nand U21409 (N_21409,N_20782,N_20867);
and U21410 (N_21410,N_20698,N_21239);
nand U21411 (N_21411,N_21021,N_20707);
nor U21412 (N_21412,N_20881,N_20720);
and U21413 (N_21413,N_20983,N_20724);
and U21414 (N_21414,N_20631,N_20938);
and U21415 (N_21415,N_20848,N_20928);
nand U21416 (N_21416,N_20655,N_20677);
and U21417 (N_21417,N_20905,N_21160);
xnor U21418 (N_21418,N_20810,N_21052);
nor U21419 (N_21419,N_20674,N_20733);
nor U21420 (N_21420,N_20846,N_20980);
xor U21421 (N_21421,N_20792,N_21072);
and U21422 (N_21422,N_20948,N_20661);
nand U21423 (N_21423,N_21070,N_20784);
xor U21424 (N_21424,N_21080,N_20815);
nand U21425 (N_21425,N_20970,N_20629);
nand U21426 (N_21426,N_20751,N_21105);
nand U21427 (N_21427,N_20664,N_20891);
and U21428 (N_21428,N_20884,N_20966);
or U21429 (N_21429,N_20781,N_21127);
or U21430 (N_21430,N_20710,N_20701);
xor U21431 (N_21431,N_20758,N_20847);
nand U21432 (N_21432,N_20752,N_21114);
nor U21433 (N_21433,N_21146,N_20822);
xor U21434 (N_21434,N_20993,N_20639);
or U21435 (N_21435,N_20685,N_20984);
xnor U21436 (N_21436,N_20872,N_21170);
or U21437 (N_21437,N_21189,N_20902);
nor U21438 (N_21438,N_21228,N_21157);
or U21439 (N_21439,N_20957,N_20961);
nand U21440 (N_21440,N_20853,N_21205);
nor U21441 (N_21441,N_20791,N_20686);
nor U21442 (N_21442,N_20726,N_20981);
xor U21443 (N_21443,N_20979,N_21118);
nor U21444 (N_21444,N_20971,N_20632);
or U21445 (N_21445,N_20873,N_21235);
or U21446 (N_21446,N_20992,N_21198);
or U21447 (N_21447,N_21063,N_20856);
nand U21448 (N_21448,N_20757,N_20742);
xor U21449 (N_21449,N_21238,N_20830);
nor U21450 (N_21450,N_20715,N_20628);
nand U21451 (N_21451,N_21000,N_21188);
or U21452 (N_21452,N_21099,N_20772);
xnor U21453 (N_21453,N_20803,N_21059);
nand U21454 (N_21454,N_20866,N_20764);
nand U21455 (N_21455,N_20798,N_21171);
nor U21456 (N_21456,N_20929,N_20964);
nand U21457 (N_21457,N_20644,N_20913);
xor U21458 (N_21458,N_21206,N_21249);
nor U21459 (N_21459,N_20680,N_21197);
nor U21460 (N_21460,N_20692,N_21028);
xnor U21461 (N_21461,N_20871,N_21055);
xor U21462 (N_21462,N_20790,N_21162);
and U21463 (N_21463,N_21141,N_20683);
or U21464 (N_21464,N_21060,N_20982);
xnor U21465 (N_21465,N_20821,N_20668);
xnor U21466 (N_21466,N_21124,N_20658);
xor U21467 (N_21467,N_20826,N_20667);
and U21468 (N_21468,N_20716,N_20978);
and U21469 (N_21469,N_20868,N_20759);
or U21470 (N_21470,N_20789,N_20635);
nand U21471 (N_21471,N_21158,N_20740);
xnor U21472 (N_21472,N_21104,N_20974);
and U21473 (N_21473,N_21042,N_20748);
nand U21474 (N_21474,N_21095,N_20940);
nor U21475 (N_21475,N_21058,N_21008);
nor U21476 (N_21476,N_20839,N_21034);
xnor U21477 (N_21477,N_21013,N_20714);
and U21478 (N_21478,N_20690,N_21173);
nor U21479 (N_21479,N_20909,N_20890);
nor U21480 (N_21480,N_21039,N_20897);
or U21481 (N_21481,N_21195,N_20924);
nor U21482 (N_21482,N_20939,N_21017);
and U21483 (N_21483,N_20836,N_21092);
and U21484 (N_21484,N_20794,N_21232);
nor U21485 (N_21485,N_20820,N_20732);
nor U21486 (N_21486,N_20811,N_20675);
nor U21487 (N_21487,N_21231,N_21207);
and U21488 (N_21488,N_20876,N_20706);
and U21489 (N_21489,N_21242,N_21035);
nand U21490 (N_21490,N_21126,N_20907);
or U21491 (N_21491,N_21166,N_21200);
xnor U21492 (N_21492,N_20738,N_20817);
nand U21493 (N_21493,N_20795,N_21184);
and U21494 (N_21494,N_21236,N_21215);
or U21495 (N_21495,N_21103,N_21120);
nand U21496 (N_21496,N_21194,N_21078);
and U21497 (N_21497,N_20965,N_21084);
or U21498 (N_21498,N_20837,N_20899);
and U21499 (N_21499,N_20991,N_20660);
and U21500 (N_21500,N_20691,N_21056);
or U21501 (N_21501,N_20746,N_21174);
and U21502 (N_21502,N_21245,N_20827);
and U21503 (N_21503,N_20967,N_21167);
nor U21504 (N_21504,N_20882,N_20919);
xnor U21505 (N_21505,N_20657,N_21204);
and U21506 (N_21506,N_21131,N_21153);
nor U21507 (N_21507,N_21119,N_21011);
or U21508 (N_21508,N_20915,N_20659);
and U21509 (N_21509,N_20927,N_21006);
nand U21510 (N_21510,N_20730,N_20883);
or U21511 (N_21511,N_21033,N_20801);
and U21512 (N_21512,N_20779,N_21143);
or U21513 (N_21513,N_20908,N_20723);
xnor U21514 (N_21514,N_20626,N_21192);
nand U21515 (N_21515,N_21001,N_21073);
xnor U21516 (N_21516,N_21150,N_20775);
nand U21517 (N_21517,N_20666,N_20922);
xor U21518 (N_21518,N_20689,N_21116);
xor U21519 (N_21519,N_20649,N_20878);
nand U21520 (N_21520,N_21163,N_21147);
nand U21521 (N_21521,N_21064,N_20785);
nor U21522 (N_21522,N_21036,N_20999);
or U21523 (N_21523,N_21051,N_20855);
xnor U21524 (N_21524,N_21122,N_21145);
or U21525 (N_21525,N_21003,N_21066);
xor U21526 (N_21526,N_20761,N_21203);
xor U21527 (N_21527,N_20874,N_21176);
and U21528 (N_21528,N_20936,N_20892);
or U21529 (N_21529,N_20756,N_20916);
nor U21530 (N_21530,N_20717,N_20917);
xor U21531 (N_21531,N_21002,N_20894);
or U21532 (N_21532,N_20727,N_21217);
or U21533 (N_21533,N_20695,N_21187);
or U21534 (N_21534,N_20945,N_21178);
xor U21535 (N_21535,N_20996,N_21199);
or U21536 (N_21536,N_20636,N_21106);
nor U21537 (N_21537,N_21024,N_21121);
xnor U21538 (N_21538,N_20697,N_21168);
or U21539 (N_21539,N_20910,N_21128);
and U21540 (N_21540,N_20643,N_20722);
and U21541 (N_21541,N_20889,N_21110);
and U21542 (N_21542,N_20972,N_20774);
or U21543 (N_21543,N_21169,N_21218);
or U21544 (N_21544,N_20705,N_20879);
or U21545 (N_21545,N_20877,N_20749);
nand U21546 (N_21546,N_20843,N_21100);
or U21547 (N_21547,N_21229,N_20688);
or U21548 (N_21548,N_20906,N_21138);
nand U21549 (N_21549,N_20708,N_21077);
or U21550 (N_21550,N_20975,N_20937);
xor U21551 (N_21551,N_21129,N_20896);
nor U21552 (N_21552,N_20963,N_20807);
nand U21553 (N_21553,N_21136,N_20995);
nor U21554 (N_21554,N_20914,N_20796);
nand U21555 (N_21555,N_20694,N_20987);
or U21556 (N_21556,N_21032,N_20901);
xnor U21557 (N_21557,N_21020,N_21140);
nand U21558 (N_21558,N_20954,N_21107);
and U21559 (N_21559,N_21010,N_21219);
nand U21560 (N_21560,N_20886,N_21223);
nor U21561 (N_21561,N_21177,N_21047);
nor U21562 (N_21562,N_21044,N_21128);
nand U21563 (N_21563,N_21213,N_21058);
and U21564 (N_21564,N_21232,N_20916);
or U21565 (N_21565,N_21213,N_21228);
or U21566 (N_21566,N_20785,N_20761);
nand U21567 (N_21567,N_20953,N_20859);
or U21568 (N_21568,N_20974,N_20923);
nor U21569 (N_21569,N_21137,N_20715);
nor U21570 (N_21570,N_21213,N_20685);
nor U21571 (N_21571,N_21229,N_21025);
nand U21572 (N_21572,N_21123,N_20751);
and U21573 (N_21573,N_20791,N_21245);
nand U21574 (N_21574,N_20673,N_20679);
nor U21575 (N_21575,N_21240,N_20899);
xnor U21576 (N_21576,N_21157,N_20817);
and U21577 (N_21577,N_20925,N_20672);
nand U21578 (N_21578,N_20920,N_20935);
or U21579 (N_21579,N_21233,N_20854);
xnor U21580 (N_21580,N_20998,N_21057);
and U21581 (N_21581,N_20625,N_21090);
and U21582 (N_21582,N_20680,N_20934);
nor U21583 (N_21583,N_20774,N_21182);
or U21584 (N_21584,N_20643,N_21221);
and U21585 (N_21585,N_20791,N_20793);
nand U21586 (N_21586,N_20798,N_21005);
nor U21587 (N_21587,N_21106,N_20901);
nand U21588 (N_21588,N_20779,N_21009);
nand U21589 (N_21589,N_20863,N_20956);
xnor U21590 (N_21590,N_21110,N_20864);
nand U21591 (N_21591,N_20753,N_20691);
or U21592 (N_21592,N_20899,N_20773);
or U21593 (N_21593,N_20924,N_21237);
nor U21594 (N_21594,N_20798,N_21156);
nor U21595 (N_21595,N_20854,N_20880);
or U21596 (N_21596,N_21034,N_20796);
xor U21597 (N_21597,N_21214,N_20687);
xor U21598 (N_21598,N_21025,N_20745);
or U21599 (N_21599,N_21068,N_21207);
and U21600 (N_21600,N_20955,N_20954);
and U21601 (N_21601,N_20968,N_21199);
nand U21602 (N_21602,N_20893,N_20686);
and U21603 (N_21603,N_20991,N_21027);
or U21604 (N_21604,N_20887,N_20780);
and U21605 (N_21605,N_20849,N_20854);
nand U21606 (N_21606,N_20699,N_20983);
nand U21607 (N_21607,N_21215,N_20788);
nand U21608 (N_21608,N_21116,N_20903);
and U21609 (N_21609,N_20739,N_20686);
xnor U21610 (N_21610,N_21218,N_21133);
nand U21611 (N_21611,N_21064,N_20994);
and U21612 (N_21612,N_21018,N_20691);
nand U21613 (N_21613,N_20967,N_20697);
xor U21614 (N_21614,N_21010,N_20991);
xnor U21615 (N_21615,N_21170,N_21046);
xor U21616 (N_21616,N_20630,N_21177);
and U21617 (N_21617,N_20798,N_21185);
and U21618 (N_21618,N_20640,N_20733);
and U21619 (N_21619,N_20926,N_20795);
and U21620 (N_21620,N_20636,N_20886);
xnor U21621 (N_21621,N_20748,N_21133);
or U21622 (N_21622,N_21211,N_20733);
nor U21623 (N_21623,N_21119,N_21198);
xnor U21624 (N_21624,N_21239,N_21152);
xor U21625 (N_21625,N_20816,N_20654);
xor U21626 (N_21626,N_20896,N_21195);
nor U21627 (N_21627,N_20940,N_20911);
nand U21628 (N_21628,N_20943,N_20986);
or U21629 (N_21629,N_21013,N_20901);
nand U21630 (N_21630,N_20948,N_20961);
nor U21631 (N_21631,N_20919,N_20659);
nand U21632 (N_21632,N_20951,N_20982);
or U21633 (N_21633,N_20819,N_20749);
nor U21634 (N_21634,N_20815,N_21009);
nand U21635 (N_21635,N_20910,N_20814);
nand U21636 (N_21636,N_20829,N_20822);
nand U21637 (N_21637,N_21237,N_20659);
nand U21638 (N_21638,N_21098,N_20646);
xor U21639 (N_21639,N_21058,N_20679);
and U21640 (N_21640,N_20789,N_20843);
nand U21641 (N_21641,N_21198,N_20839);
or U21642 (N_21642,N_21102,N_21088);
nand U21643 (N_21643,N_21095,N_20785);
nor U21644 (N_21644,N_21040,N_20920);
nand U21645 (N_21645,N_21082,N_20900);
xnor U21646 (N_21646,N_20693,N_21031);
xor U21647 (N_21647,N_20673,N_21202);
nand U21648 (N_21648,N_21143,N_21190);
and U21649 (N_21649,N_20738,N_20802);
or U21650 (N_21650,N_20933,N_20931);
or U21651 (N_21651,N_20983,N_20804);
nand U21652 (N_21652,N_21180,N_20764);
or U21653 (N_21653,N_21098,N_21143);
nor U21654 (N_21654,N_21062,N_21140);
and U21655 (N_21655,N_20702,N_20644);
or U21656 (N_21656,N_21124,N_20771);
nor U21657 (N_21657,N_20959,N_20924);
and U21658 (N_21658,N_20812,N_20942);
or U21659 (N_21659,N_21016,N_21199);
nor U21660 (N_21660,N_21113,N_20876);
nor U21661 (N_21661,N_21043,N_20871);
and U21662 (N_21662,N_21162,N_20931);
nor U21663 (N_21663,N_20878,N_20806);
xnor U21664 (N_21664,N_20626,N_20999);
xnor U21665 (N_21665,N_20858,N_20763);
nor U21666 (N_21666,N_20841,N_21131);
nand U21667 (N_21667,N_20882,N_20941);
nand U21668 (N_21668,N_20914,N_21131);
nor U21669 (N_21669,N_21114,N_20835);
and U21670 (N_21670,N_20693,N_21214);
nand U21671 (N_21671,N_21175,N_20646);
nor U21672 (N_21672,N_20854,N_21201);
nor U21673 (N_21673,N_21160,N_21028);
xor U21674 (N_21674,N_20683,N_20672);
xor U21675 (N_21675,N_21116,N_21118);
nand U21676 (N_21676,N_21221,N_20678);
nor U21677 (N_21677,N_20850,N_21167);
or U21678 (N_21678,N_21175,N_20742);
nor U21679 (N_21679,N_20785,N_20801);
xor U21680 (N_21680,N_20661,N_21222);
xor U21681 (N_21681,N_20845,N_20939);
xor U21682 (N_21682,N_20702,N_21198);
and U21683 (N_21683,N_20955,N_20671);
xnor U21684 (N_21684,N_21183,N_21116);
nand U21685 (N_21685,N_21072,N_21061);
and U21686 (N_21686,N_21239,N_21071);
nand U21687 (N_21687,N_20677,N_20799);
nand U21688 (N_21688,N_21067,N_21225);
or U21689 (N_21689,N_21014,N_20815);
xnor U21690 (N_21690,N_21068,N_20727);
xnor U21691 (N_21691,N_20874,N_21006);
or U21692 (N_21692,N_21174,N_21093);
nor U21693 (N_21693,N_20960,N_20823);
nor U21694 (N_21694,N_21078,N_20872);
nand U21695 (N_21695,N_20800,N_21130);
and U21696 (N_21696,N_20912,N_20789);
xor U21697 (N_21697,N_20634,N_21179);
nand U21698 (N_21698,N_21188,N_21247);
or U21699 (N_21699,N_20867,N_20706);
or U21700 (N_21700,N_20862,N_20900);
xor U21701 (N_21701,N_21030,N_21106);
xnor U21702 (N_21702,N_21213,N_20693);
or U21703 (N_21703,N_20676,N_20690);
xnor U21704 (N_21704,N_20986,N_20714);
or U21705 (N_21705,N_20867,N_20784);
and U21706 (N_21706,N_21025,N_21036);
nor U21707 (N_21707,N_20860,N_20882);
xor U21708 (N_21708,N_21045,N_21196);
or U21709 (N_21709,N_20651,N_21224);
xnor U21710 (N_21710,N_21055,N_21221);
nand U21711 (N_21711,N_20704,N_20717);
xor U21712 (N_21712,N_20822,N_20890);
nand U21713 (N_21713,N_20972,N_21219);
or U21714 (N_21714,N_21100,N_21080);
and U21715 (N_21715,N_20909,N_21230);
or U21716 (N_21716,N_20933,N_21030);
nor U21717 (N_21717,N_20724,N_20843);
nand U21718 (N_21718,N_21220,N_21243);
or U21719 (N_21719,N_20976,N_21233);
xnor U21720 (N_21720,N_20989,N_21125);
xnor U21721 (N_21721,N_21140,N_20787);
xor U21722 (N_21722,N_21126,N_20771);
nor U21723 (N_21723,N_21165,N_20735);
or U21724 (N_21724,N_20638,N_20961);
nor U21725 (N_21725,N_20944,N_20748);
or U21726 (N_21726,N_21237,N_21139);
nor U21727 (N_21727,N_20758,N_20806);
nor U21728 (N_21728,N_21151,N_20809);
nand U21729 (N_21729,N_20904,N_20770);
nor U21730 (N_21730,N_20917,N_21200);
and U21731 (N_21731,N_20812,N_21123);
nor U21732 (N_21732,N_20657,N_21115);
or U21733 (N_21733,N_21055,N_20680);
or U21734 (N_21734,N_21231,N_20730);
nand U21735 (N_21735,N_20717,N_21044);
and U21736 (N_21736,N_21023,N_20975);
nor U21737 (N_21737,N_20855,N_21249);
nor U21738 (N_21738,N_20894,N_20648);
nand U21739 (N_21739,N_20634,N_21013);
and U21740 (N_21740,N_20766,N_20828);
nand U21741 (N_21741,N_21068,N_21146);
or U21742 (N_21742,N_20915,N_21214);
xor U21743 (N_21743,N_21024,N_21111);
or U21744 (N_21744,N_21237,N_21147);
and U21745 (N_21745,N_20684,N_20835);
xnor U21746 (N_21746,N_20880,N_20968);
or U21747 (N_21747,N_20793,N_20710);
and U21748 (N_21748,N_20734,N_20943);
nand U21749 (N_21749,N_21184,N_21116);
nand U21750 (N_21750,N_20641,N_21141);
nand U21751 (N_21751,N_21012,N_20807);
nor U21752 (N_21752,N_21208,N_20788);
and U21753 (N_21753,N_20774,N_20684);
and U21754 (N_21754,N_21132,N_21081);
nor U21755 (N_21755,N_20771,N_21016);
and U21756 (N_21756,N_20970,N_20744);
nor U21757 (N_21757,N_20826,N_20684);
or U21758 (N_21758,N_20829,N_20903);
and U21759 (N_21759,N_21242,N_21066);
or U21760 (N_21760,N_20694,N_21219);
nand U21761 (N_21761,N_21003,N_21116);
or U21762 (N_21762,N_20966,N_20669);
xnor U21763 (N_21763,N_21176,N_20658);
xor U21764 (N_21764,N_20690,N_21023);
nor U21765 (N_21765,N_20958,N_20792);
or U21766 (N_21766,N_20971,N_20625);
nor U21767 (N_21767,N_20688,N_20789);
nand U21768 (N_21768,N_21065,N_20689);
xor U21769 (N_21769,N_20888,N_21175);
nor U21770 (N_21770,N_20889,N_21233);
xnor U21771 (N_21771,N_21105,N_21171);
nor U21772 (N_21772,N_20676,N_20774);
xnor U21773 (N_21773,N_20704,N_20957);
nor U21774 (N_21774,N_21086,N_21176);
and U21775 (N_21775,N_20727,N_20923);
nand U21776 (N_21776,N_21129,N_20848);
or U21777 (N_21777,N_20655,N_21156);
nor U21778 (N_21778,N_20981,N_20649);
and U21779 (N_21779,N_20948,N_21127);
or U21780 (N_21780,N_20838,N_21079);
or U21781 (N_21781,N_21024,N_20709);
xnor U21782 (N_21782,N_20892,N_21028);
nor U21783 (N_21783,N_20932,N_21018);
nor U21784 (N_21784,N_21125,N_20707);
xnor U21785 (N_21785,N_21117,N_20786);
nand U21786 (N_21786,N_21238,N_20743);
nor U21787 (N_21787,N_21032,N_21128);
xor U21788 (N_21788,N_20872,N_20968);
or U21789 (N_21789,N_21051,N_20656);
and U21790 (N_21790,N_21044,N_20948);
xnor U21791 (N_21791,N_20848,N_20735);
nor U21792 (N_21792,N_21033,N_21042);
nand U21793 (N_21793,N_20831,N_21221);
and U21794 (N_21794,N_20733,N_20965);
nor U21795 (N_21795,N_20704,N_20810);
nor U21796 (N_21796,N_20823,N_20827);
nand U21797 (N_21797,N_21031,N_21246);
or U21798 (N_21798,N_21101,N_21107);
xor U21799 (N_21799,N_20898,N_21192);
nor U21800 (N_21800,N_20960,N_21120);
nor U21801 (N_21801,N_21116,N_21181);
nand U21802 (N_21802,N_20941,N_21060);
xnor U21803 (N_21803,N_20669,N_20703);
nand U21804 (N_21804,N_20794,N_20896);
nand U21805 (N_21805,N_21210,N_20980);
and U21806 (N_21806,N_21013,N_21079);
xor U21807 (N_21807,N_21235,N_20650);
xor U21808 (N_21808,N_20996,N_20789);
or U21809 (N_21809,N_20873,N_20714);
nor U21810 (N_21810,N_20845,N_20635);
nor U21811 (N_21811,N_20850,N_20972);
and U21812 (N_21812,N_21001,N_20862);
nor U21813 (N_21813,N_20855,N_21031);
and U21814 (N_21814,N_21048,N_20954);
xor U21815 (N_21815,N_20874,N_21057);
nor U21816 (N_21816,N_20917,N_20934);
and U21817 (N_21817,N_20932,N_20805);
nor U21818 (N_21818,N_21089,N_20774);
and U21819 (N_21819,N_21007,N_20743);
or U21820 (N_21820,N_20685,N_21159);
and U21821 (N_21821,N_21139,N_20800);
nor U21822 (N_21822,N_21083,N_21167);
nand U21823 (N_21823,N_21226,N_20636);
or U21824 (N_21824,N_20801,N_20869);
and U21825 (N_21825,N_21169,N_20966);
nand U21826 (N_21826,N_21217,N_20832);
and U21827 (N_21827,N_21136,N_21171);
nor U21828 (N_21828,N_20841,N_21068);
or U21829 (N_21829,N_20729,N_20712);
or U21830 (N_21830,N_20819,N_20872);
nand U21831 (N_21831,N_21121,N_20641);
xnor U21832 (N_21832,N_20857,N_20661);
and U21833 (N_21833,N_20644,N_20780);
and U21834 (N_21834,N_20965,N_21185);
nor U21835 (N_21835,N_20821,N_21015);
and U21836 (N_21836,N_20970,N_20812);
xor U21837 (N_21837,N_21098,N_20850);
and U21838 (N_21838,N_21060,N_20782);
nor U21839 (N_21839,N_21169,N_20705);
or U21840 (N_21840,N_20965,N_21246);
xor U21841 (N_21841,N_20825,N_20766);
or U21842 (N_21842,N_20833,N_20785);
or U21843 (N_21843,N_20678,N_20776);
and U21844 (N_21844,N_21233,N_20763);
xnor U21845 (N_21845,N_21190,N_20627);
xnor U21846 (N_21846,N_20713,N_20725);
xor U21847 (N_21847,N_20675,N_21115);
nand U21848 (N_21848,N_21011,N_21097);
nor U21849 (N_21849,N_21028,N_20927);
and U21850 (N_21850,N_20938,N_21210);
xor U21851 (N_21851,N_20998,N_20713);
and U21852 (N_21852,N_20847,N_20857);
and U21853 (N_21853,N_21107,N_20999);
or U21854 (N_21854,N_20738,N_20778);
nor U21855 (N_21855,N_20919,N_21229);
nor U21856 (N_21856,N_20675,N_20931);
or U21857 (N_21857,N_20686,N_20926);
nand U21858 (N_21858,N_20626,N_21080);
nor U21859 (N_21859,N_21136,N_21011);
or U21860 (N_21860,N_20667,N_20922);
nor U21861 (N_21861,N_21018,N_21093);
or U21862 (N_21862,N_20639,N_21031);
and U21863 (N_21863,N_20806,N_20650);
nand U21864 (N_21864,N_20961,N_21222);
xnor U21865 (N_21865,N_20906,N_21066);
nand U21866 (N_21866,N_21157,N_21213);
nand U21867 (N_21867,N_20796,N_20658);
xor U21868 (N_21868,N_21052,N_20917);
nand U21869 (N_21869,N_21015,N_20866);
and U21870 (N_21870,N_21045,N_20859);
nor U21871 (N_21871,N_21092,N_21223);
or U21872 (N_21872,N_21085,N_20703);
and U21873 (N_21873,N_21236,N_20908);
and U21874 (N_21874,N_21083,N_21039);
nor U21875 (N_21875,N_21467,N_21324);
and U21876 (N_21876,N_21498,N_21624);
xnor U21877 (N_21877,N_21349,N_21452);
xnor U21878 (N_21878,N_21725,N_21537);
or U21879 (N_21879,N_21346,N_21716);
and U21880 (N_21880,N_21345,N_21434);
xor U21881 (N_21881,N_21618,N_21389);
nand U21882 (N_21882,N_21741,N_21719);
xor U21883 (N_21883,N_21531,N_21302);
or U21884 (N_21884,N_21567,N_21577);
and U21885 (N_21885,N_21608,N_21401);
xnor U21886 (N_21886,N_21762,N_21444);
or U21887 (N_21887,N_21621,N_21536);
and U21888 (N_21888,N_21406,N_21559);
nor U21889 (N_21889,N_21449,N_21427);
and U21890 (N_21890,N_21832,N_21315);
and U21891 (N_21891,N_21822,N_21689);
nand U21892 (N_21892,N_21425,N_21326);
xnor U21893 (N_21893,N_21544,N_21554);
or U21894 (N_21894,N_21610,N_21705);
nor U21895 (N_21895,N_21416,N_21343);
nand U21896 (N_21896,N_21506,N_21623);
nand U21897 (N_21897,N_21671,N_21767);
xor U21898 (N_21898,N_21474,N_21672);
xor U21899 (N_21899,N_21321,N_21590);
xor U21900 (N_21900,N_21863,N_21338);
xnor U21901 (N_21901,N_21335,N_21553);
and U21902 (N_21902,N_21825,N_21469);
xnor U21903 (N_21903,N_21639,N_21276);
xor U21904 (N_21904,N_21541,N_21446);
nor U21905 (N_21905,N_21582,N_21297);
and U21906 (N_21906,N_21835,N_21684);
nor U21907 (N_21907,N_21394,N_21695);
nand U21908 (N_21908,N_21795,N_21319);
nor U21909 (N_21909,N_21735,N_21815);
xor U21910 (N_21910,N_21723,N_21512);
nand U21911 (N_21911,N_21337,N_21391);
nor U21912 (N_21912,N_21518,N_21779);
or U21913 (N_21913,N_21367,N_21558);
and U21914 (N_21914,N_21404,N_21816);
nor U21915 (N_21915,N_21399,N_21385);
xnor U21916 (N_21916,N_21682,N_21379);
xor U21917 (N_21917,N_21584,N_21633);
nor U21918 (N_21918,N_21329,N_21647);
and U21919 (N_21919,N_21722,N_21766);
nor U21920 (N_21920,N_21826,N_21311);
and U21921 (N_21921,N_21727,N_21448);
or U21922 (N_21922,N_21871,N_21793);
and U21923 (N_21923,N_21428,N_21614);
xnor U21924 (N_21924,N_21694,N_21412);
xnor U21925 (N_21925,N_21461,N_21630);
or U21926 (N_21926,N_21411,N_21360);
nand U21927 (N_21927,N_21515,N_21362);
nor U21928 (N_21928,N_21540,N_21830);
and U21929 (N_21929,N_21644,N_21460);
and U21930 (N_21930,N_21844,N_21805);
nand U21931 (N_21931,N_21602,N_21706);
or U21932 (N_21932,N_21642,N_21625);
and U21933 (N_21933,N_21847,N_21365);
or U21934 (N_21934,N_21468,N_21369);
nor U21935 (N_21935,N_21291,N_21521);
or U21936 (N_21936,N_21552,N_21317);
nor U21937 (N_21937,N_21670,N_21342);
xnor U21938 (N_21938,N_21638,N_21481);
nand U21939 (N_21939,N_21504,N_21569);
xnor U21940 (N_21940,N_21445,N_21688);
and U21941 (N_21941,N_21358,N_21818);
and U21942 (N_21942,N_21803,N_21737);
nor U21943 (N_21943,N_21351,N_21388);
xnor U21944 (N_21944,N_21294,N_21692);
xor U21945 (N_21945,N_21415,N_21619);
nand U21946 (N_21946,N_21405,N_21457);
or U21947 (N_21947,N_21796,N_21508);
nor U21948 (N_21948,N_21597,N_21479);
nand U21949 (N_21949,N_21437,N_21780);
nand U21950 (N_21950,N_21857,N_21866);
xnor U21951 (N_21951,N_21462,N_21836);
and U21952 (N_21952,N_21856,N_21659);
nand U21953 (N_21953,N_21340,N_21864);
and U21954 (N_21954,N_21591,N_21418);
nand U21955 (N_21955,N_21661,N_21528);
nand U21956 (N_21956,N_21598,N_21852);
and U21957 (N_21957,N_21426,N_21331);
or U21958 (N_21958,N_21606,N_21484);
or U21959 (N_21959,N_21547,N_21256);
or U21960 (N_21960,N_21842,N_21786);
nor U21961 (N_21961,N_21287,N_21356);
nand U21962 (N_21962,N_21505,N_21740);
and U21963 (N_21963,N_21398,N_21765);
nor U21964 (N_21964,N_21328,N_21586);
nor U21965 (N_21965,N_21579,N_21396);
nand U21966 (N_21966,N_21667,N_21292);
nand U21967 (N_21967,N_21703,N_21407);
nor U21968 (N_21968,N_21529,N_21333);
or U21969 (N_21969,N_21441,N_21378);
or U21970 (N_21970,N_21746,N_21278);
nor U21971 (N_21971,N_21353,N_21650);
nand U21972 (N_21972,N_21702,N_21861);
xnor U21973 (N_21973,N_21691,N_21601);
or U21974 (N_21974,N_21698,N_21447);
or U21975 (N_21975,N_21806,N_21564);
nor U21976 (N_21976,N_21493,N_21592);
and U21977 (N_21977,N_21542,N_21649);
nor U21978 (N_21978,N_21566,N_21611);
nand U21979 (N_21979,N_21872,N_21262);
and U21980 (N_21980,N_21733,N_21768);
nor U21981 (N_21981,N_21734,N_21574);
and U21982 (N_21982,N_21675,N_21257);
and U21983 (N_21983,N_21402,N_21383);
nor U21984 (N_21984,N_21289,N_21681);
nor U21985 (N_21985,N_21583,N_21458);
or U21986 (N_21986,N_21259,N_21299);
xor U21987 (N_21987,N_21466,N_21422);
nand U21988 (N_21988,N_21539,N_21252);
nor U21989 (N_21989,N_21419,N_21264);
xor U21990 (N_21990,N_21332,N_21673);
nand U21991 (N_21991,N_21386,N_21485);
nand U21992 (N_21992,N_21433,N_21867);
xor U21993 (N_21993,N_21748,N_21785);
nand U21994 (N_21994,N_21470,N_21439);
or U21995 (N_21995,N_21686,N_21543);
and U21996 (N_21996,N_21492,N_21862);
xnor U21997 (N_21997,N_21400,N_21507);
nand U21998 (N_21998,N_21849,N_21525);
and U21999 (N_21999,N_21534,N_21770);
nand U22000 (N_22000,N_21640,N_21593);
or U22001 (N_22001,N_21387,N_21381);
nand U22002 (N_22002,N_21293,N_21473);
nor U22003 (N_22003,N_21565,N_21423);
xnor U22004 (N_22004,N_21480,N_21858);
and U22005 (N_22005,N_21420,N_21373);
nand U22006 (N_22006,N_21730,N_21296);
xor U22007 (N_22007,N_21634,N_21424);
xnor U22008 (N_22008,N_21489,N_21873);
nor U22009 (N_22009,N_21773,N_21812);
or U22010 (N_22010,N_21341,N_21840);
or U22011 (N_22011,N_21496,N_21472);
nand U22012 (N_22012,N_21350,N_21410);
nand U22013 (N_22013,N_21581,N_21511);
nand U22014 (N_22014,N_21305,N_21318);
nor U22015 (N_22015,N_21599,N_21578);
nor U22016 (N_22016,N_21440,N_21545);
and U22017 (N_22017,N_21306,N_21550);
xor U22018 (N_22018,N_21755,N_21509);
xor U22019 (N_22019,N_21513,N_21589);
nand U22020 (N_22020,N_21334,N_21769);
nand U22021 (N_22021,N_21707,N_21514);
nand U22022 (N_22022,N_21546,N_21393);
xnor U22023 (N_22023,N_21314,N_21652);
nand U22024 (N_22024,N_21573,N_21376);
and U22025 (N_22025,N_21798,N_21637);
or U22026 (N_22026,N_21745,N_21371);
nand U22027 (N_22027,N_21710,N_21323);
and U22028 (N_22028,N_21366,N_21656);
nor U22029 (N_22029,N_21585,N_21283);
nand U22030 (N_22030,N_21853,N_21561);
and U22031 (N_22031,N_21253,N_21772);
nand U22032 (N_22032,N_21450,N_21501);
xnor U22033 (N_22033,N_21459,N_21678);
nand U22034 (N_22034,N_21685,N_21322);
nand U22035 (N_22035,N_21403,N_21813);
xnor U22036 (N_22036,N_21680,N_21551);
xnor U22037 (N_22037,N_21330,N_21266);
nor U22038 (N_22038,N_21641,N_21497);
or U22039 (N_22039,N_21265,N_21657);
xnor U22040 (N_22040,N_21414,N_21303);
and U22041 (N_22041,N_21743,N_21848);
and U22042 (N_22042,N_21568,N_21571);
nand U22043 (N_22043,N_21756,N_21603);
nor U22044 (N_22044,N_21281,N_21635);
xor U22045 (N_22045,N_21488,N_21288);
or U22046 (N_22046,N_21258,N_21778);
or U22047 (N_22047,N_21774,N_21463);
and U22048 (N_22048,N_21575,N_21273);
nand U22049 (N_22049,N_21254,N_21776);
nor U22050 (N_22050,N_21761,N_21609);
and U22051 (N_22051,N_21382,N_21438);
nand U22052 (N_22052,N_21286,N_21503);
xnor U22053 (N_22053,N_21653,N_21738);
nand U22054 (N_22054,N_21777,N_21482);
nand U22055 (N_22055,N_21417,N_21261);
and U22056 (N_22056,N_21364,N_21313);
xnor U22057 (N_22057,N_21846,N_21658);
nor U22058 (N_22058,N_21519,N_21749);
or U22059 (N_22059,N_21804,N_21841);
or U22060 (N_22060,N_21347,N_21595);
and U22061 (N_22061,N_21782,N_21838);
and U22062 (N_22062,N_21845,N_21801);
or U22063 (N_22063,N_21701,N_21352);
nor U22064 (N_22064,N_21298,N_21712);
xor U22065 (N_22065,N_21660,N_21431);
or U22066 (N_22066,N_21833,N_21819);
xor U22067 (N_22067,N_21478,N_21556);
xnor U22068 (N_22068,N_21664,N_21742);
nand U22069 (N_22069,N_21628,N_21392);
nand U22070 (N_22070,N_21309,N_21285);
or U22071 (N_22071,N_21275,N_21729);
nor U22072 (N_22072,N_21700,N_21357);
or U22073 (N_22073,N_21697,N_21821);
and U22074 (N_22074,N_21409,N_21348);
and U22075 (N_22075,N_21272,N_21533);
xnor U22076 (N_22076,N_21791,N_21295);
nor U22077 (N_22077,N_21487,N_21336);
nor U22078 (N_22078,N_21607,N_21636);
nand U22079 (N_22079,N_21374,N_21308);
or U22080 (N_22080,N_21802,N_21683);
and U22081 (N_22081,N_21491,N_21435);
nor U22082 (N_22082,N_21271,N_21455);
or U22083 (N_22083,N_21363,N_21523);
nor U22084 (N_22084,N_21714,N_21549);
xor U22085 (N_22085,N_21851,N_21829);
xnor U22086 (N_22086,N_21429,N_21526);
nor U22087 (N_22087,N_21736,N_21250);
nor U22088 (N_22088,N_21588,N_21532);
xnor U22089 (N_22089,N_21612,N_21465);
xnor U22090 (N_22090,N_21715,N_21375);
nor U22091 (N_22091,N_21708,N_21760);
xor U22092 (N_22092,N_21654,N_21728);
nand U22093 (N_22093,N_21316,N_21724);
nand U22094 (N_22094,N_21693,N_21837);
and U22095 (N_22095,N_21269,N_21797);
nor U22096 (N_22096,N_21300,N_21339);
nand U22097 (N_22097,N_21739,N_21442);
xnor U22098 (N_22098,N_21810,N_21709);
nor U22099 (N_22099,N_21807,N_21731);
nor U22100 (N_22100,N_21408,N_21270);
xnor U22101 (N_22101,N_21477,N_21604);
xor U22102 (N_22102,N_21390,N_21843);
nand U22103 (N_22103,N_21620,N_21794);
nand U22104 (N_22104,N_21535,N_21372);
xor U22105 (N_22105,N_21563,N_21320);
xnor U22106 (N_22106,N_21666,N_21790);
nand U22107 (N_22107,N_21430,N_21282);
nor U22108 (N_22108,N_21645,N_21655);
nor U22109 (N_22109,N_21600,N_21814);
and U22110 (N_22110,N_21277,N_21676);
xnor U22111 (N_22111,N_21744,N_21354);
xor U22112 (N_22112,N_21255,N_21869);
nor U22113 (N_22113,N_21527,N_21855);
xor U22114 (N_22114,N_21763,N_21750);
or U22115 (N_22115,N_21717,N_21486);
and U22116 (N_22116,N_21524,N_21704);
and U22117 (N_22117,N_21451,N_21668);
or U22118 (N_22118,N_21594,N_21260);
nor U22119 (N_22119,N_21456,N_21799);
nand U22120 (N_22120,N_21510,N_21368);
and U22121 (N_22121,N_21792,N_21310);
xnor U22122 (N_22122,N_21570,N_21674);
or U22123 (N_22123,N_21752,N_21530);
nor U22124 (N_22124,N_21267,N_21711);
nand U22125 (N_22125,N_21483,N_21732);
and U22126 (N_22126,N_21718,N_21643);
and U22127 (N_22127,N_21520,N_21679);
and U22128 (N_22128,N_21870,N_21677);
nand U22129 (N_22129,N_21280,N_21538);
or U22130 (N_22130,N_21500,N_21831);
nand U22131 (N_22131,N_21263,N_21312);
or U22132 (N_22132,N_21860,N_21629);
xnor U22133 (N_22133,N_21865,N_21759);
and U22134 (N_22134,N_21370,N_21436);
nor U22135 (N_22135,N_21476,N_21787);
or U22136 (N_22136,N_21557,N_21301);
nand U22137 (N_22137,N_21834,N_21576);
or U22138 (N_22138,N_21783,N_21788);
xnor U22139 (N_22139,N_21384,N_21651);
and U22140 (N_22140,N_21817,N_21720);
xor U22141 (N_22141,N_21344,N_21397);
nor U22142 (N_22142,N_21646,N_21758);
nor U22143 (N_22143,N_21454,N_21380);
nor U22144 (N_22144,N_21850,N_21771);
nand U22145 (N_22145,N_21764,N_21517);
and U22146 (N_22146,N_21307,N_21475);
nor U22147 (N_22147,N_21268,N_21626);
nor U22148 (N_22148,N_21361,N_21432);
nor U22149 (N_22149,N_21548,N_21753);
and U22150 (N_22150,N_21687,N_21631);
and U22151 (N_22151,N_21471,N_21824);
xnor U22152 (N_22152,N_21809,N_21662);
and U22153 (N_22153,N_21757,N_21751);
nand U22154 (N_22154,N_21304,N_21453);
xor U22155 (N_22155,N_21874,N_21632);
nand U22156 (N_22156,N_21274,N_21359);
nand U22157 (N_22157,N_21443,N_21868);
nor U22158 (N_22158,N_21696,N_21775);
or U22159 (N_22159,N_21839,N_21490);
xnor U22160 (N_22160,N_21516,N_21781);
nor U22161 (N_22161,N_21859,N_21377);
nand U22162 (N_22162,N_21648,N_21605);
or U22163 (N_22163,N_21325,N_21522);
or U22164 (N_22164,N_21560,N_21699);
nor U22165 (N_22165,N_21502,N_21413);
or U22166 (N_22166,N_21828,N_21395);
nand U22167 (N_22167,N_21627,N_21617);
or U22168 (N_22168,N_21721,N_21284);
nor U22169 (N_22169,N_21495,N_21499);
and U22170 (N_22170,N_21290,N_21596);
nor U22171 (N_22171,N_21820,N_21421);
xor U22172 (N_22172,N_21279,N_21800);
xnor U22173 (N_22173,N_21616,N_21789);
nor U22174 (N_22174,N_21754,N_21663);
nor U22175 (N_22175,N_21811,N_21823);
xnor U22176 (N_22176,N_21587,N_21355);
nor U22177 (N_22177,N_21665,N_21726);
nand U22178 (N_22178,N_21572,N_21713);
and U22179 (N_22179,N_21690,N_21669);
and U22180 (N_22180,N_21464,N_21555);
xor U22181 (N_22181,N_21327,N_21580);
nand U22182 (N_22182,N_21615,N_21251);
nor U22183 (N_22183,N_21622,N_21808);
or U22184 (N_22184,N_21827,N_21854);
nor U22185 (N_22185,N_21747,N_21562);
xor U22186 (N_22186,N_21784,N_21494);
and U22187 (N_22187,N_21613,N_21514);
nor U22188 (N_22188,N_21777,N_21343);
or U22189 (N_22189,N_21567,N_21709);
or U22190 (N_22190,N_21391,N_21466);
and U22191 (N_22191,N_21503,N_21335);
nor U22192 (N_22192,N_21616,N_21549);
and U22193 (N_22193,N_21353,N_21798);
nand U22194 (N_22194,N_21610,N_21362);
and U22195 (N_22195,N_21775,N_21688);
xnor U22196 (N_22196,N_21732,N_21848);
and U22197 (N_22197,N_21724,N_21311);
and U22198 (N_22198,N_21658,N_21817);
xor U22199 (N_22199,N_21657,N_21838);
xor U22200 (N_22200,N_21439,N_21256);
or U22201 (N_22201,N_21353,N_21808);
nor U22202 (N_22202,N_21839,N_21413);
nor U22203 (N_22203,N_21629,N_21663);
nor U22204 (N_22204,N_21315,N_21600);
nand U22205 (N_22205,N_21759,N_21785);
nor U22206 (N_22206,N_21276,N_21629);
nor U22207 (N_22207,N_21589,N_21612);
nor U22208 (N_22208,N_21345,N_21533);
and U22209 (N_22209,N_21607,N_21273);
xnor U22210 (N_22210,N_21428,N_21384);
or U22211 (N_22211,N_21301,N_21553);
or U22212 (N_22212,N_21431,N_21820);
or U22213 (N_22213,N_21260,N_21794);
nor U22214 (N_22214,N_21548,N_21415);
or U22215 (N_22215,N_21821,N_21361);
or U22216 (N_22216,N_21308,N_21632);
nor U22217 (N_22217,N_21780,N_21471);
nor U22218 (N_22218,N_21715,N_21333);
nor U22219 (N_22219,N_21305,N_21389);
or U22220 (N_22220,N_21774,N_21650);
nor U22221 (N_22221,N_21347,N_21310);
and U22222 (N_22222,N_21312,N_21275);
or U22223 (N_22223,N_21415,N_21343);
and U22224 (N_22224,N_21713,N_21650);
or U22225 (N_22225,N_21547,N_21437);
nand U22226 (N_22226,N_21424,N_21578);
and U22227 (N_22227,N_21818,N_21251);
or U22228 (N_22228,N_21532,N_21809);
nand U22229 (N_22229,N_21433,N_21302);
and U22230 (N_22230,N_21382,N_21756);
or U22231 (N_22231,N_21627,N_21653);
xor U22232 (N_22232,N_21549,N_21611);
nor U22233 (N_22233,N_21647,N_21683);
nor U22234 (N_22234,N_21699,N_21491);
and U22235 (N_22235,N_21350,N_21589);
nor U22236 (N_22236,N_21363,N_21767);
xor U22237 (N_22237,N_21791,N_21729);
xnor U22238 (N_22238,N_21531,N_21459);
nand U22239 (N_22239,N_21850,N_21626);
nor U22240 (N_22240,N_21506,N_21310);
nor U22241 (N_22241,N_21568,N_21796);
nand U22242 (N_22242,N_21487,N_21452);
xor U22243 (N_22243,N_21436,N_21625);
and U22244 (N_22244,N_21750,N_21481);
xor U22245 (N_22245,N_21359,N_21776);
and U22246 (N_22246,N_21353,N_21327);
nand U22247 (N_22247,N_21345,N_21699);
nand U22248 (N_22248,N_21516,N_21322);
and U22249 (N_22249,N_21632,N_21709);
and U22250 (N_22250,N_21565,N_21857);
nand U22251 (N_22251,N_21835,N_21673);
or U22252 (N_22252,N_21853,N_21706);
or U22253 (N_22253,N_21730,N_21401);
or U22254 (N_22254,N_21539,N_21400);
nand U22255 (N_22255,N_21401,N_21404);
nor U22256 (N_22256,N_21750,N_21633);
xor U22257 (N_22257,N_21447,N_21666);
xnor U22258 (N_22258,N_21297,N_21525);
or U22259 (N_22259,N_21526,N_21515);
nand U22260 (N_22260,N_21528,N_21448);
xnor U22261 (N_22261,N_21552,N_21315);
nand U22262 (N_22262,N_21856,N_21632);
or U22263 (N_22263,N_21770,N_21351);
and U22264 (N_22264,N_21487,N_21268);
or U22265 (N_22265,N_21715,N_21592);
nand U22266 (N_22266,N_21761,N_21538);
nor U22267 (N_22267,N_21783,N_21336);
nand U22268 (N_22268,N_21580,N_21446);
or U22269 (N_22269,N_21563,N_21529);
or U22270 (N_22270,N_21367,N_21354);
xnor U22271 (N_22271,N_21701,N_21268);
and U22272 (N_22272,N_21513,N_21692);
or U22273 (N_22273,N_21672,N_21337);
nor U22274 (N_22274,N_21628,N_21324);
nor U22275 (N_22275,N_21820,N_21762);
xnor U22276 (N_22276,N_21611,N_21264);
nand U22277 (N_22277,N_21391,N_21610);
and U22278 (N_22278,N_21633,N_21391);
or U22279 (N_22279,N_21663,N_21799);
nor U22280 (N_22280,N_21639,N_21389);
nor U22281 (N_22281,N_21805,N_21385);
and U22282 (N_22282,N_21453,N_21711);
nand U22283 (N_22283,N_21813,N_21514);
nor U22284 (N_22284,N_21870,N_21676);
nor U22285 (N_22285,N_21821,N_21261);
nor U22286 (N_22286,N_21562,N_21304);
nand U22287 (N_22287,N_21623,N_21493);
nand U22288 (N_22288,N_21358,N_21484);
or U22289 (N_22289,N_21459,N_21754);
or U22290 (N_22290,N_21659,N_21600);
or U22291 (N_22291,N_21811,N_21334);
or U22292 (N_22292,N_21437,N_21850);
and U22293 (N_22293,N_21497,N_21254);
nand U22294 (N_22294,N_21824,N_21678);
xor U22295 (N_22295,N_21484,N_21784);
nand U22296 (N_22296,N_21571,N_21530);
nor U22297 (N_22297,N_21732,N_21856);
xor U22298 (N_22298,N_21457,N_21854);
nor U22299 (N_22299,N_21865,N_21559);
and U22300 (N_22300,N_21325,N_21601);
nand U22301 (N_22301,N_21840,N_21520);
nand U22302 (N_22302,N_21278,N_21739);
nand U22303 (N_22303,N_21336,N_21605);
nand U22304 (N_22304,N_21369,N_21733);
nor U22305 (N_22305,N_21381,N_21869);
or U22306 (N_22306,N_21666,N_21449);
nand U22307 (N_22307,N_21555,N_21803);
or U22308 (N_22308,N_21608,N_21448);
and U22309 (N_22309,N_21407,N_21579);
nand U22310 (N_22310,N_21871,N_21519);
nand U22311 (N_22311,N_21474,N_21332);
nor U22312 (N_22312,N_21293,N_21593);
or U22313 (N_22313,N_21354,N_21834);
nand U22314 (N_22314,N_21861,N_21790);
nand U22315 (N_22315,N_21357,N_21668);
or U22316 (N_22316,N_21777,N_21395);
and U22317 (N_22317,N_21823,N_21518);
nor U22318 (N_22318,N_21316,N_21646);
nor U22319 (N_22319,N_21484,N_21619);
nor U22320 (N_22320,N_21789,N_21298);
or U22321 (N_22321,N_21266,N_21603);
or U22322 (N_22322,N_21666,N_21442);
nor U22323 (N_22323,N_21256,N_21633);
nor U22324 (N_22324,N_21255,N_21857);
nor U22325 (N_22325,N_21705,N_21399);
or U22326 (N_22326,N_21654,N_21782);
nor U22327 (N_22327,N_21642,N_21621);
or U22328 (N_22328,N_21849,N_21422);
and U22329 (N_22329,N_21689,N_21346);
and U22330 (N_22330,N_21856,N_21280);
nand U22331 (N_22331,N_21250,N_21417);
nor U22332 (N_22332,N_21357,N_21620);
and U22333 (N_22333,N_21366,N_21837);
and U22334 (N_22334,N_21796,N_21396);
or U22335 (N_22335,N_21268,N_21737);
and U22336 (N_22336,N_21741,N_21274);
or U22337 (N_22337,N_21794,N_21313);
nand U22338 (N_22338,N_21294,N_21788);
nand U22339 (N_22339,N_21379,N_21865);
xnor U22340 (N_22340,N_21474,N_21509);
nand U22341 (N_22341,N_21866,N_21591);
or U22342 (N_22342,N_21789,N_21399);
nor U22343 (N_22343,N_21738,N_21708);
nand U22344 (N_22344,N_21789,N_21802);
and U22345 (N_22345,N_21583,N_21700);
nand U22346 (N_22346,N_21301,N_21734);
or U22347 (N_22347,N_21663,N_21509);
or U22348 (N_22348,N_21793,N_21623);
nand U22349 (N_22349,N_21718,N_21577);
xnor U22350 (N_22350,N_21464,N_21324);
nor U22351 (N_22351,N_21506,N_21273);
nor U22352 (N_22352,N_21833,N_21273);
or U22353 (N_22353,N_21824,N_21550);
nand U22354 (N_22354,N_21390,N_21522);
xnor U22355 (N_22355,N_21843,N_21319);
xnor U22356 (N_22356,N_21372,N_21495);
nor U22357 (N_22357,N_21316,N_21434);
nand U22358 (N_22358,N_21550,N_21640);
nand U22359 (N_22359,N_21469,N_21628);
nand U22360 (N_22360,N_21615,N_21739);
nor U22361 (N_22361,N_21472,N_21338);
nand U22362 (N_22362,N_21533,N_21371);
and U22363 (N_22363,N_21713,N_21290);
xnor U22364 (N_22364,N_21354,N_21343);
and U22365 (N_22365,N_21546,N_21299);
nor U22366 (N_22366,N_21531,N_21386);
xor U22367 (N_22367,N_21608,N_21763);
or U22368 (N_22368,N_21271,N_21854);
nor U22369 (N_22369,N_21275,N_21397);
nor U22370 (N_22370,N_21820,N_21691);
xnor U22371 (N_22371,N_21727,N_21568);
and U22372 (N_22372,N_21479,N_21741);
and U22373 (N_22373,N_21725,N_21372);
and U22374 (N_22374,N_21836,N_21301);
and U22375 (N_22375,N_21581,N_21443);
xnor U22376 (N_22376,N_21509,N_21309);
and U22377 (N_22377,N_21811,N_21568);
nor U22378 (N_22378,N_21383,N_21830);
nor U22379 (N_22379,N_21439,N_21474);
nor U22380 (N_22380,N_21275,N_21837);
and U22381 (N_22381,N_21431,N_21859);
xnor U22382 (N_22382,N_21553,N_21504);
xor U22383 (N_22383,N_21475,N_21703);
or U22384 (N_22384,N_21562,N_21649);
nand U22385 (N_22385,N_21504,N_21760);
or U22386 (N_22386,N_21266,N_21530);
nor U22387 (N_22387,N_21675,N_21401);
nand U22388 (N_22388,N_21459,N_21742);
nor U22389 (N_22389,N_21799,N_21762);
and U22390 (N_22390,N_21610,N_21836);
and U22391 (N_22391,N_21873,N_21529);
nor U22392 (N_22392,N_21524,N_21404);
or U22393 (N_22393,N_21351,N_21423);
or U22394 (N_22394,N_21682,N_21256);
nand U22395 (N_22395,N_21471,N_21374);
nand U22396 (N_22396,N_21451,N_21412);
and U22397 (N_22397,N_21321,N_21647);
xor U22398 (N_22398,N_21802,N_21252);
or U22399 (N_22399,N_21821,N_21386);
xnor U22400 (N_22400,N_21539,N_21822);
nand U22401 (N_22401,N_21414,N_21821);
and U22402 (N_22402,N_21559,N_21368);
nand U22403 (N_22403,N_21265,N_21313);
xnor U22404 (N_22404,N_21747,N_21614);
nand U22405 (N_22405,N_21674,N_21268);
or U22406 (N_22406,N_21576,N_21598);
nand U22407 (N_22407,N_21791,N_21418);
or U22408 (N_22408,N_21736,N_21448);
nand U22409 (N_22409,N_21608,N_21612);
nand U22410 (N_22410,N_21346,N_21753);
or U22411 (N_22411,N_21862,N_21435);
xnor U22412 (N_22412,N_21707,N_21341);
xnor U22413 (N_22413,N_21594,N_21542);
or U22414 (N_22414,N_21753,N_21715);
nand U22415 (N_22415,N_21833,N_21694);
xor U22416 (N_22416,N_21829,N_21657);
or U22417 (N_22417,N_21357,N_21316);
or U22418 (N_22418,N_21281,N_21491);
or U22419 (N_22419,N_21413,N_21438);
nor U22420 (N_22420,N_21508,N_21871);
nand U22421 (N_22421,N_21610,N_21463);
and U22422 (N_22422,N_21599,N_21332);
nand U22423 (N_22423,N_21300,N_21459);
nor U22424 (N_22424,N_21792,N_21393);
xor U22425 (N_22425,N_21443,N_21377);
and U22426 (N_22426,N_21569,N_21683);
and U22427 (N_22427,N_21638,N_21390);
and U22428 (N_22428,N_21435,N_21551);
xnor U22429 (N_22429,N_21571,N_21828);
or U22430 (N_22430,N_21433,N_21430);
or U22431 (N_22431,N_21565,N_21373);
or U22432 (N_22432,N_21823,N_21868);
nor U22433 (N_22433,N_21715,N_21256);
xnor U22434 (N_22434,N_21738,N_21282);
nor U22435 (N_22435,N_21781,N_21273);
and U22436 (N_22436,N_21822,N_21417);
or U22437 (N_22437,N_21802,N_21267);
xnor U22438 (N_22438,N_21600,N_21329);
or U22439 (N_22439,N_21391,N_21371);
nor U22440 (N_22440,N_21286,N_21775);
nor U22441 (N_22441,N_21296,N_21841);
and U22442 (N_22442,N_21337,N_21353);
and U22443 (N_22443,N_21814,N_21817);
and U22444 (N_22444,N_21847,N_21863);
or U22445 (N_22445,N_21341,N_21789);
xor U22446 (N_22446,N_21346,N_21730);
xor U22447 (N_22447,N_21464,N_21535);
or U22448 (N_22448,N_21648,N_21400);
nand U22449 (N_22449,N_21862,N_21585);
nor U22450 (N_22450,N_21254,N_21615);
and U22451 (N_22451,N_21561,N_21592);
nand U22452 (N_22452,N_21690,N_21508);
and U22453 (N_22453,N_21867,N_21626);
nand U22454 (N_22454,N_21603,N_21366);
and U22455 (N_22455,N_21550,N_21478);
xnor U22456 (N_22456,N_21326,N_21325);
and U22457 (N_22457,N_21856,N_21396);
and U22458 (N_22458,N_21401,N_21659);
nand U22459 (N_22459,N_21439,N_21848);
xor U22460 (N_22460,N_21849,N_21796);
nand U22461 (N_22461,N_21837,N_21701);
and U22462 (N_22462,N_21802,N_21870);
or U22463 (N_22463,N_21795,N_21282);
nor U22464 (N_22464,N_21456,N_21738);
nor U22465 (N_22465,N_21516,N_21845);
or U22466 (N_22466,N_21340,N_21394);
and U22467 (N_22467,N_21316,N_21851);
xnor U22468 (N_22468,N_21763,N_21804);
nor U22469 (N_22469,N_21673,N_21820);
nor U22470 (N_22470,N_21755,N_21302);
or U22471 (N_22471,N_21744,N_21777);
or U22472 (N_22472,N_21870,N_21331);
or U22473 (N_22473,N_21770,N_21798);
xor U22474 (N_22474,N_21683,N_21813);
nor U22475 (N_22475,N_21355,N_21384);
or U22476 (N_22476,N_21551,N_21547);
or U22477 (N_22477,N_21690,N_21523);
xor U22478 (N_22478,N_21817,N_21806);
and U22479 (N_22479,N_21639,N_21567);
and U22480 (N_22480,N_21784,N_21593);
xor U22481 (N_22481,N_21273,N_21778);
and U22482 (N_22482,N_21835,N_21818);
nand U22483 (N_22483,N_21424,N_21432);
xor U22484 (N_22484,N_21267,N_21299);
or U22485 (N_22485,N_21778,N_21611);
and U22486 (N_22486,N_21845,N_21376);
nor U22487 (N_22487,N_21845,N_21858);
or U22488 (N_22488,N_21260,N_21254);
and U22489 (N_22489,N_21452,N_21441);
nand U22490 (N_22490,N_21791,N_21532);
nand U22491 (N_22491,N_21290,N_21717);
and U22492 (N_22492,N_21832,N_21356);
nand U22493 (N_22493,N_21774,N_21674);
nor U22494 (N_22494,N_21507,N_21697);
nor U22495 (N_22495,N_21340,N_21499);
or U22496 (N_22496,N_21538,N_21666);
nand U22497 (N_22497,N_21801,N_21715);
xor U22498 (N_22498,N_21297,N_21754);
nor U22499 (N_22499,N_21756,N_21759);
and U22500 (N_22500,N_22301,N_22336);
or U22501 (N_22501,N_21956,N_22078);
nand U22502 (N_22502,N_21903,N_21915);
nand U22503 (N_22503,N_21900,N_21986);
and U22504 (N_22504,N_22462,N_22353);
nand U22505 (N_22505,N_22213,N_22045);
xnor U22506 (N_22506,N_21934,N_22230);
nand U22507 (N_22507,N_22418,N_22089);
xor U22508 (N_22508,N_22240,N_22448);
nand U22509 (N_22509,N_22064,N_22383);
or U22510 (N_22510,N_22378,N_21924);
xor U22511 (N_22511,N_22478,N_22279);
or U22512 (N_22512,N_22063,N_22080);
nor U22513 (N_22513,N_21962,N_22485);
or U22514 (N_22514,N_22428,N_22390);
nor U22515 (N_22515,N_22342,N_22387);
xnor U22516 (N_22516,N_22169,N_22202);
or U22517 (N_22517,N_22103,N_21885);
nor U22518 (N_22518,N_21906,N_21899);
and U22519 (N_22519,N_22191,N_22211);
and U22520 (N_22520,N_22126,N_21960);
nand U22521 (N_22521,N_22246,N_22398);
nor U22522 (N_22522,N_21964,N_22059);
nand U22523 (N_22523,N_22312,N_22265);
nor U22524 (N_22524,N_21927,N_22134);
or U22525 (N_22525,N_22173,N_22360);
nor U22526 (N_22526,N_22273,N_22001);
xor U22527 (N_22527,N_21972,N_21910);
xor U22528 (N_22528,N_22074,N_22004);
xnor U22529 (N_22529,N_22395,N_22226);
xnor U22530 (N_22530,N_21938,N_22491);
nand U22531 (N_22531,N_22035,N_22164);
or U22532 (N_22532,N_22159,N_22350);
nand U22533 (N_22533,N_22236,N_22269);
nand U22534 (N_22534,N_22404,N_22371);
and U22535 (N_22535,N_21978,N_22010);
xnor U22536 (N_22536,N_22038,N_22490);
and U22537 (N_22537,N_22403,N_21957);
nand U22538 (N_22538,N_21913,N_22008);
nor U22539 (N_22539,N_21983,N_22188);
nor U22540 (N_22540,N_22100,N_22091);
or U22541 (N_22541,N_22281,N_21998);
xor U22542 (N_22542,N_22104,N_22168);
or U22543 (N_22543,N_21912,N_22186);
nor U22544 (N_22544,N_21961,N_22200);
or U22545 (N_22545,N_22361,N_22384);
and U22546 (N_22546,N_22304,N_22308);
and U22547 (N_22547,N_21932,N_21989);
and U22548 (N_22548,N_22155,N_22024);
or U22549 (N_22549,N_22254,N_22460);
xor U22550 (N_22550,N_22271,N_22461);
and U22551 (N_22551,N_22034,N_22095);
xor U22552 (N_22552,N_22058,N_21997);
nand U22553 (N_22553,N_22107,N_22499);
xnor U22554 (N_22554,N_22219,N_22454);
and U22555 (N_22555,N_22272,N_22175);
nand U22556 (N_22556,N_22036,N_22225);
and U22557 (N_22557,N_22380,N_22477);
xnor U22558 (N_22558,N_22305,N_22359);
and U22559 (N_22559,N_22425,N_22037);
xnor U22560 (N_22560,N_22182,N_22426);
or U22561 (N_22561,N_21968,N_22183);
or U22562 (N_22562,N_22190,N_22162);
and U22563 (N_22563,N_22363,N_22295);
xnor U22564 (N_22564,N_22357,N_22400);
nor U22565 (N_22565,N_22184,N_21917);
xor U22566 (N_22566,N_22451,N_22253);
nor U22567 (N_22567,N_22027,N_21902);
nor U22568 (N_22568,N_22278,N_22017);
and U22569 (N_22569,N_22094,N_22379);
xor U22570 (N_22570,N_22487,N_22386);
xor U22571 (N_22571,N_22423,N_22157);
and U22572 (N_22572,N_22204,N_22318);
and U22573 (N_22573,N_22430,N_22255);
nand U22574 (N_22574,N_21916,N_21930);
nand U22575 (N_22575,N_22261,N_22263);
and U22576 (N_22576,N_22181,N_22003);
or U22577 (N_22577,N_22026,N_22142);
nand U22578 (N_22578,N_21894,N_22054);
and U22579 (N_22579,N_21970,N_22450);
and U22580 (N_22580,N_22101,N_22405);
nor U22581 (N_22581,N_22009,N_22061);
nor U22582 (N_22582,N_21973,N_22042);
and U22583 (N_22583,N_22138,N_22432);
xor U22584 (N_22584,N_22023,N_22315);
or U22585 (N_22585,N_22081,N_22108);
nor U22586 (N_22586,N_22102,N_21919);
nand U22587 (N_22587,N_22049,N_22283);
nor U22588 (N_22588,N_22067,N_22497);
or U22589 (N_22589,N_22411,N_21942);
nor U22590 (N_22590,N_21939,N_21933);
nor U22591 (N_22591,N_22310,N_21991);
nor U22592 (N_22592,N_22251,N_22112);
and U22593 (N_22593,N_22466,N_22401);
nand U22594 (N_22594,N_22389,N_22135);
and U22595 (N_22595,N_22196,N_22114);
or U22596 (N_22596,N_22287,N_22046);
nor U22597 (N_22597,N_22198,N_22167);
and U22598 (N_22598,N_22439,N_22165);
nor U22599 (N_22599,N_21884,N_22148);
nand U22600 (N_22600,N_22307,N_22412);
nand U22601 (N_22601,N_22410,N_22105);
and U22602 (N_22602,N_22099,N_22006);
nand U22603 (N_22603,N_21996,N_21949);
or U22604 (N_22604,N_21891,N_22073);
xnor U22605 (N_22605,N_22249,N_22041);
xnor U22606 (N_22606,N_22179,N_22072);
nand U22607 (N_22607,N_22097,N_22195);
nand U22608 (N_22608,N_22120,N_22421);
nand U22609 (N_22609,N_22327,N_22048);
xor U22610 (N_22610,N_22416,N_22393);
xnor U22611 (N_22611,N_22446,N_22233);
nand U22612 (N_22612,N_22476,N_22364);
and U22613 (N_22613,N_22291,N_22370);
nor U22614 (N_22614,N_22109,N_22177);
nor U22615 (N_22615,N_21898,N_22119);
nor U22616 (N_22616,N_22333,N_22498);
xnor U22617 (N_22617,N_22481,N_22445);
nand U22618 (N_22618,N_22187,N_22438);
and U22619 (N_22619,N_21963,N_22325);
and U22620 (N_22620,N_22229,N_21897);
xnor U22621 (N_22621,N_22464,N_22194);
nand U22622 (N_22622,N_22040,N_21954);
nor U22623 (N_22623,N_22096,N_21880);
or U22624 (N_22624,N_22334,N_21953);
and U22625 (N_22625,N_22266,N_22051);
and U22626 (N_22626,N_22176,N_22115);
nor U22627 (N_22627,N_22372,N_22362);
or U22628 (N_22628,N_22178,N_22424);
or U22629 (N_22629,N_22419,N_22206);
or U22630 (N_22630,N_21907,N_21937);
nand U22631 (N_22631,N_22012,N_21935);
xor U22632 (N_22632,N_22302,N_21888);
nor U22633 (N_22633,N_22232,N_22156);
and U22634 (N_22634,N_22311,N_21995);
xor U22635 (N_22635,N_21908,N_21886);
and U22636 (N_22636,N_22039,N_22224);
or U22637 (N_22637,N_22303,N_22128);
nand U22638 (N_22638,N_22329,N_22057);
nand U22639 (N_22639,N_21901,N_22288);
and U22640 (N_22640,N_21987,N_22330);
or U22641 (N_22641,N_22276,N_22453);
nand U22642 (N_22642,N_22468,N_22152);
xor U22643 (N_22643,N_22479,N_22488);
nor U22644 (N_22644,N_22163,N_21890);
xnor U22645 (N_22645,N_22250,N_21909);
xor U22646 (N_22646,N_22293,N_21926);
xor U22647 (N_22647,N_22349,N_22223);
and U22648 (N_22648,N_22489,N_22174);
or U22649 (N_22649,N_22131,N_22133);
or U22650 (N_22650,N_22463,N_22215);
nor U22651 (N_22651,N_22221,N_22415);
or U22652 (N_22652,N_22227,N_22209);
nand U22653 (N_22653,N_21952,N_22354);
nor U22654 (N_22654,N_22217,N_22417);
and U22655 (N_22655,N_22079,N_21879);
nor U22656 (N_22656,N_22070,N_22331);
or U22657 (N_22657,N_22257,N_22340);
nand U22658 (N_22658,N_22406,N_22388);
nor U22659 (N_22659,N_22121,N_21974);
or U22660 (N_22660,N_22002,N_21911);
or U22661 (N_22661,N_22345,N_22033);
nor U22662 (N_22662,N_21945,N_21925);
nor U22663 (N_22663,N_22483,N_22234);
nor U22664 (N_22664,N_22116,N_22117);
and U22665 (N_22665,N_22306,N_22088);
or U22666 (N_22666,N_22455,N_22136);
or U22667 (N_22667,N_22321,N_22050);
nor U22668 (N_22668,N_22443,N_21967);
and U22669 (N_22669,N_22189,N_22025);
or U22670 (N_22670,N_22486,N_21959);
xor U22671 (N_22671,N_21951,N_22444);
xnor U22672 (N_22672,N_22141,N_21893);
xor U22673 (N_22673,N_22267,N_22077);
xor U22674 (N_22674,N_22032,N_22324);
nor U22675 (N_22675,N_22338,N_21992);
or U22676 (N_22676,N_21881,N_22084);
and U22677 (N_22677,N_22289,N_22474);
or U22678 (N_22678,N_22222,N_22347);
and U22679 (N_22679,N_22270,N_22343);
nand U22680 (N_22680,N_22207,N_22402);
or U22681 (N_22681,N_22129,N_22172);
nand U22682 (N_22682,N_22437,N_21966);
xor U22683 (N_22683,N_22212,N_22130);
and U22684 (N_22684,N_22268,N_21876);
nand U22685 (N_22685,N_22422,N_22391);
nand U22686 (N_22686,N_22434,N_22473);
nor U22687 (N_22687,N_22031,N_22205);
nand U22688 (N_22688,N_22373,N_22242);
and U22689 (N_22689,N_21905,N_22066);
nand U22690 (N_22690,N_22285,N_22409);
and U22691 (N_22691,N_22431,N_22139);
xnor U22692 (N_22692,N_21950,N_22013);
nand U22693 (N_22693,N_21931,N_22397);
xor U22694 (N_22694,N_22435,N_22220);
or U22695 (N_22695,N_22294,N_22256);
and U22696 (N_22696,N_22166,N_22309);
and U22697 (N_22697,N_21999,N_22344);
or U22698 (N_22698,N_22366,N_22071);
nand U22699 (N_22699,N_21896,N_22098);
and U22700 (N_22700,N_22018,N_21947);
xor U22701 (N_22701,N_22286,N_22252);
nand U22702 (N_22702,N_21943,N_22277);
nor U22703 (N_22703,N_21984,N_22106);
or U22704 (N_22704,N_22355,N_22282);
and U22705 (N_22705,N_22458,N_21923);
nand U22706 (N_22706,N_22180,N_22262);
nand U22707 (N_22707,N_22260,N_21990);
nand U22708 (N_22708,N_22146,N_22123);
and U22709 (N_22709,N_22158,N_22392);
nand U22710 (N_22710,N_22440,N_22016);
nand U22711 (N_22711,N_22385,N_22193);
xor U22712 (N_22712,N_21976,N_22029);
and U22713 (N_22713,N_22238,N_22472);
xnor U22714 (N_22714,N_22339,N_22203);
xnor U22715 (N_22715,N_21955,N_22456);
or U22716 (N_22716,N_22028,N_21940);
nand U22717 (N_22717,N_22171,N_22297);
nand U22718 (N_22718,N_22376,N_22442);
nor U22719 (N_22719,N_21988,N_22326);
and U22720 (N_22720,N_21875,N_21994);
nor U22721 (N_22721,N_22143,N_22085);
nor U22722 (N_22722,N_22110,N_21982);
nor U22723 (N_22723,N_22153,N_22300);
and U22724 (N_22724,N_22471,N_22145);
or U22725 (N_22725,N_22076,N_22197);
or U22726 (N_22726,N_22322,N_22496);
xnor U22727 (N_22727,N_22298,N_22069);
nor U22728 (N_22728,N_22290,N_22082);
nor U22729 (N_22729,N_22299,N_22151);
xor U22730 (N_22730,N_22280,N_22239);
and U22731 (N_22731,N_22030,N_22122);
xnor U22732 (N_22732,N_21914,N_21944);
and U22733 (N_22733,N_22356,N_21946);
nand U22734 (N_22734,N_22284,N_22043);
xor U22735 (N_22735,N_22137,N_22492);
nor U22736 (N_22736,N_21985,N_22436);
and U22737 (N_22737,N_22480,N_22332);
nor U22738 (N_22738,N_22317,N_22092);
nand U22739 (N_22739,N_22228,N_22368);
nand U22740 (N_22740,N_22068,N_22218);
xor U22741 (N_22741,N_22093,N_22259);
nor U22742 (N_22742,N_22382,N_22000);
xor U22743 (N_22743,N_22020,N_22365);
xor U22744 (N_22744,N_21936,N_22144);
and U22745 (N_22745,N_22475,N_22052);
or U22746 (N_22746,N_21921,N_22019);
nand U22747 (N_22747,N_22358,N_21892);
nor U22748 (N_22748,N_22248,N_22216);
and U22749 (N_22749,N_22320,N_22015);
nor U22750 (N_22750,N_22414,N_21979);
or U22751 (N_22751,N_22275,N_21977);
and U22752 (N_22752,N_21895,N_22335);
or U22753 (N_22753,N_21948,N_22408);
nor U22754 (N_22754,N_21971,N_22022);
nand U22755 (N_22755,N_21958,N_22007);
or U22756 (N_22756,N_22161,N_22449);
or U22757 (N_22757,N_21993,N_21918);
nand U22758 (N_22758,N_21878,N_22208);
xnor U22759 (N_22759,N_22274,N_22053);
and U22760 (N_22760,N_22494,N_22258);
and U22761 (N_22761,N_22447,N_22060);
xnor U22762 (N_22762,N_22090,N_22149);
nand U22763 (N_22763,N_22055,N_22065);
and U22764 (N_22764,N_21922,N_22044);
and U22765 (N_22765,N_21904,N_22328);
nor U22766 (N_22766,N_22292,N_22433);
xor U22767 (N_22767,N_22241,N_22132);
xnor U22768 (N_22768,N_21941,N_22369);
nor U22769 (N_22769,N_22235,N_21877);
or U22770 (N_22770,N_22264,N_22374);
nor U22771 (N_22771,N_22192,N_22459);
xnor U22772 (N_22772,N_22469,N_22482);
or U22773 (N_22773,N_22441,N_21882);
and U22774 (N_22774,N_22375,N_22185);
nor U22775 (N_22775,N_22351,N_22124);
nand U22776 (N_22776,N_22231,N_22470);
xnor U22777 (N_22777,N_22367,N_22493);
nand U22778 (N_22778,N_22316,N_21883);
and U22779 (N_22779,N_21980,N_22377);
nor U22780 (N_22780,N_21920,N_22237);
nor U22781 (N_22781,N_22313,N_22087);
or U22782 (N_22782,N_22111,N_22413);
or U22783 (N_22783,N_22160,N_22348);
nand U22784 (N_22784,N_22127,N_22062);
and U22785 (N_22785,N_22381,N_22319);
and U22786 (N_22786,N_21889,N_22210);
nor U22787 (N_22787,N_22113,N_22394);
or U22788 (N_22788,N_22457,N_22337);
and U22789 (N_22789,N_22247,N_22296);
nor U22790 (N_22790,N_22314,N_22465);
or U22791 (N_22791,N_22245,N_22352);
and U22792 (N_22792,N_21965,N_22399);
or U22793 (N_22793,N_22005,N_21975);
xor U22794 (N_22794,N_22170,N_22346);
xor U22795 (N_22795,N_22214,N_22021);
and U22796 (N_22796,N_22467,N_22150);
xnor U22797 (N_22797,N_22429,N_22125);
nor U22798 (N_22798,N_22047,N_22396);
nor U22799 (N_22799,N_22420,N_22083);
and U22800 (N_22800,N_22407,N_22452);
nand U22801 (N_22801,N_21969,N_22323);
and U22802 (N_22802,N_21928,N_22011);
and U22803 (N_22803,N_22244,N_21981);
xor U22804 (N_22804,N_22075,N_22201);
or U22805 (N_22805,N_22427,N_22484);
nor U22806 (N_22806,N_22495,N_21887);
nor U22807 (N_22807,N_22154,N_22056);
or U22808 (N_22808,N_21929,N_22147);
or U22809 (N_22809,N_22341,N_22199);
or U22810 (N_22810,N_22243,N_22086);
and U22811 (N_22811,N_22140,N_22014);
nor U22812 (N_22812,N_22118,N_22204);
and U22813 (N_22813,N_22190,N_22139);
nor U22814 (N_22814,N_22265,N_21934);
or U22815 (N_22815,N_22162,N_22178);
nand U22816 (N_22816,N_21933,N_22302);
nor U22817 (N_22817,N_22455,N_22330);
and U22818 (N_22818,N_22072,N_21907);
nand U22819 (N_22819,N_22038,N_22402);
xnor U22820 (N_22820,N_22290,N_21971);
xor U22821 (N_22821,N_21935,N_22071);
xor U22822 (N_22822,N_22176,N_22311);
nand U22823 (N_22823,N_22295,N_22073);
and U22824 (N_22824,N_22075,N_22375);
xnor U22825 (N_22825,N_22232,N_22119);
xnor U22826 (N_22826,N_22318,N_22396);
xor U22827 (N_22827,N_22137,N_22169);
xor U22828 (N_22828,N_22102,N_22365);
xor U22829 (N_22829,N_21885,N_21986);
nand U22830 (N_22830,N_22278,N_21994);
nor U22831 (N_22831,N_22179,N_22377);
nand U22832 (N_22832,N_22442,N_21911);
or U22833 (N_22833,N_22443,N_22440);
nand U22834 (N_22834,N_22038,N_22144);
and U22835 (N_22835,N_21914,N_22304);
nor U22836 (N_22836,N_22191,N_22065);
nand U22837 (N_22837,N_22190,N_22231);
xor U22838 (N_22838,N_22120,N_22307);
nand U22839 (N_22839,N_21938,N_22154);
nor U22840 (N_22840,N_22208,N_21891);
nand U22841 (N_22841,N_22273,N_22223);
xor U22842 (N_22842,N_22388,N_21936);
and U22843 (N_22843,N_22172,N_22437);
xor U22844 (N_22844,N_22450,N_21913);
nand U22845 (N_22845,N_22477,N_22048);
nor U22846 (N_22846,N_22122,N_22395);
nor U22847 (N_22847,N_22020,N_22436);
or U22848 (N_22848,N_22497,N_21997);
nor U22849 (N_22849,N_22312,N_22482);
nor U22850 (N_22850,N_22286,N_22082);
or U22851 (N_22851,N_22149,N_22331);
nor U22852 (N_22852,N_22223,N_22005);
xnor U22853 (N_22853,N_22349,N_22065);
nor U22854 (N_22854,N_21905,N_22101);
and U22855 (N_22855,N_22181,N_22026);
and U22856 (N_22856,N_22380,N_22316);
nor U22857 (N_22857,N_22160,N_22196);
nor U22858 (N_22858,N_22397,N_21975);
nand U22859 (N_22859,N_22066,N_22357);
nand U22860 (N_22860,N_22177,N_22092);
nand U22861 (N_22861,N_22107,N_22247);
nor U22862 (N_22862,N_22082,N_22001);
xor U22863 (N_22863,N_22170,N_22491);
xor U22864 (N_22864,N_22379,N_22406);
nor U22865 (N_22865,N_22302,N_22345);
or U22866 (N_22866,N_22021,N_22179);
xnor U22867 (N_22867,N_22339,N_22297);
or U22868 (N_22868,N_22132,N_22380);
and U22869 (N_22869,N_22360,N_22423);
nor U22870 (N_22870,N_22189,N_22272);
nor U22871 (N_22871,N_22368,N_22367);
nor U22872 (N_22872,N_22035,N_22196);
nor U22873 (N_22873,N_22309,N_22426);
nor U22874 (N_22874,N_22188,N_22270);
xor U22875 (N_22875,N_21968,N_22494);
nor U22876 (N_22876,N_22017,N_22310);
nand U22877 (N_22877,N_22050,N_22195);
and U22878 (N_22878,N_22232,N_22170);
nor U22879 (N_22879,N_21990,N_22258);
or U22880 (N_22880,N_22226,N_22277);
nor U22881 (N_22881,N_22389,N_22481);
nor U22882 (N_22882,N_22186,N_22053);
or U22883 (N_22883,N_22205,N_22415);
and U22884 (N_22884,N_22090,N_21969);
or U22885 (N_22885,N_22048,N_21959);
nor U22886 (N_22886,N_21994,N_21945);
xor U22887 (N_22887,N_22474,N_22275);
and U22888 (N_22888,N_22495,N_22335);
and U22889 (N_22889,N_22338,N_22110);
and U22890 (N_22890,N_21936,N_22403);
nand U22891 (N_22891,N_22296,N_22122);
nand U22892 (N_22892,N_22070,N_22374);
nand U22893 (N_22893,N_22158,N_21925);
nor U22894 (N_22894,N_22473,N_22289);
and U22895 (N_22895,N_22114,N_22141);
nor U22896 (N_22896,N_22018,N_21982);
xnor U22897 (N_22897,N_22494,N_22403);
or U22898 (N_22898,N_21930,N_22207);
nor U22899 (N_22899,N_22264,N_22406);
nand U22900 (N_22900,N_22016,N_22469);
xor U22901 (N_22901,N_22087,N_22462);
and U22902 (N_22902,N_21908,N_21970);
xnor U22903 (N_22903,N_22128,N_22120);
or U22904 (N_22904,N_22494,N_22070);
nor U22905 (N_22905,N_22336,N_22292);
xor U22906 (N_22906,N_22240,N_22097);
or U22907 (N_22907,N_22464,N_22024);
nand U22908 (N_22908,N_22354,N_22223);
xnor U22909 (N_22909,N_22491,N_21925);
nand U22910 (N_22910,N_22178,N_22394);
or U22911 (N_22911,N_22067,N_21943);
or U22912 (N_22912,N_22193,N_22085);
nor U22913 (N_22913,N_22325,N_22101);
nand U22914 (N_22914,N_21945,N_22430);
or U22915 (N_22915,N_22385,N_22471);
xnor U22916 (N_22916,N_21912,N_22221);
nor U22917 (N_22917,N_22194,N_22451);
nand U22918 (N_22918,N_22001,N_21998);
or U22919 (N_22919,N_22332,N_22328);
nand U22920 (N_22920,N_21983,N_22390);
xor U22921 (N_22921,N_22148,N_22406);
and U22922 (N_22922,N_21957,N_22265);
nor U22923 (N_22923,N_22265,N_21966);
and U22924 (N_22924,N_22105,N_21885);
nor U22925 (N_22925,N_22375,N_21982);
and U22926 (N_22926,N_22019,N_21918);
nand U22927 (N_22927,N_22220,N_22001);
and U22928 (N_22928,N_22202,N_22214);
nand U22929 (N_22929,N_21968,N_22040);
and U22930 (N_22930,N_22380,N_22054);
nor U22931 (N_22931,N_22019,N_21956);
nand U22932 (N_22932,N_22040,N_22436);
xnor U22933 (N_22933,N_21966,N_21900);
xnor U22934 (N_22934,N_21950,N_22187);
nand U22935 (N_22935,N_22074,N_22407);
and U22936 (N_22936,N_22453,N_22335);
nand U22937 (N_22937,N_22063,N_21940);
nor U22938 (N_22938,N_22168,N_22215);
nor U22939 (N_22939,N_22304,N_22263);
or U22940 (N_22940,N_22247,N_22257);
nand U22941 (N_22941,N_21998,N_22018);
or U22942 (N_22942,N_22179,N_22341);
and U22943 (N_22943,N_22463,N_22260);
xor U22944 (N_22944,N_21882,N_22319);
or U22945 (N_22945,N_22260,N_21985);
and U22946 (N_22946,N_22420,N_22320);
nor U22947 (N_22947,N_22249,N_22106);
nand U22948 (N_22948,N_22307,N_22025);
or U22949 (N_22949,N_22410,N_22312);
xnor U22950 (N_22950,N_22017,N_22208);
nor U22951 (N_22951,N_22318,N_22225);
xor U22952 (N_22952,N_22271,N_21936);
or U22953 (N_22953,N_22399,N_21923);
nand U22954 (N_22954,N_22009,N_22326);
xnor U22955 (N_22955,N_22143,N_22491);
and U22956 (N_22956,N_22196,N_22059);
nor U22957 (N_22957,N_22329,N_22071);
nor U22958 (N_22958,N_22152,N_22048);
xor U22959 (N_22959,N_22169,N_21963);
nor U22960 (N_22960,N_22489,N_22281);
xnor U22961 (N_22961,N_22384,N_22421);
and U22962 (N_22962,N_21901,N_22107);
nor U22963 (N_22963,N_22043,N_22248);
nor U22964 (N_22964,N_22090,N_22195);
and U22965 (N_22965,N_22173,N_22285);
nor U22966 (N_22966,N_22176,N_21934);
nand U22967 (N_22967,N_22323,N_21996);
or U22968 (N_22968,N_22088,N_22319);
and U22969 (N_22969,N_22495,N_22375);
xor U22970 (N_22970,N_22044,N_22411);
or U22971 (N_22971,N_22179,N_22197);
or U22972 (N_22972,N_22470,N_22494);
xnor U22973 (N_22973,N_22235,N_22012);
nand U22974 (N_22974,N_22088,N_22110);
xor U22975 (N_22975,N_22364,N_21933);
xor U22976 (N_22976,N_22497,N_22455);
and U22977 (N_22977,N_22071,N_22092);
nor U22978 (N_22978,N_22486,N_22274);
xnor U22979 (N_22979,N_22271,N_22316);
or U22980 (N_22980,N_21904,N_21939);
nand U22981 (N_22981,N_22046,N_21900);
xor U22982 (N_22982,N_22108,N_22485);
xor U22983 (N_22983,N_22106,N_22101);
nor U22984 (N_22984,N_22241,N_22343);
and U22985 (N_22985,N_21876,N_21961);
nand U22986 (N_22986,N_22019,N_22193);
nand U22987 (N_22987,N_22349,N_22056);
nor U22988 (N_22988,N_22333,N_22252);
or U22989 (N_22989,N_22340,N_22356);
nand U22990 (N_22990,N_22196,N_22475);
nand U22991 (N_22991,N_22133,N_22075);
and U22992 (N_22992,N_22088,N_22002);
and U22993 (N_22993,N_22207,N_22299);
xnor U22994 (N_22994,N_22356,N_21923);
xnor U22995 (N_22995,N_22365,N_21962);
nand U22996 (N_22996,N_22434,N_22303);
nor U22997 (N_22997,N_22207,N_21938);
nand U22998 (N_22998,N_22343,N_22309);
xor U22999 (N_22999,N_22074,N_22341);
xor U23000 (N_23000,N_22202,N_22147);
and U23001 (N_23001,N_21990,N_22215);
xnor U23002 (N_23002,N_22012,N_21967);
and U23003 (N_23003,N_22242,N_22365);
xnor U23004 (N_23004,N_22487,N_22030);
and U23005 (N_23005,N_22275,N_22139);
and U23006 (N_23006,N_22053,N_22243);
and U23007 (N_23007,N_22263,N_22194);
nand U23008 (N_23008,N_22008,N_22165);
nand U23009 (N_23009,N_22034,N_22392);
and U23010 (N_23010,N_22264,N_22388);
or U23011 (N_23011,N_22209,N_22061);
and U23012 (N_23012,N_22001,N_21982);
and U23013 (N_23013,N_22418,N_21879);
nand U23014 (N_23014,N_22308,N_22280);
and U23015 (N_23015,N_22339,N_22039);
xnor U23016 (N_23016,N_22425,N_21980);
nor U23017 (N_23017,N_22294,N_22492);
xor U23018 (N_23018,N_22359,N_22330);
nand U23019 (N_23019,N_22130,N_22027);
nand U23020 (N_23020,N_22394,N_22115);
xor U23021 (N_23021,N_21994,N_22045);
nand U23022 (N_23022,N_22479,N_21915);
or U23023 (N_23023,N_22034,N_21994);
and U23024 (N_23024,N_22055,N_22409);
nor U23025 (N_23025,N_22348,N_22236);
xnor U23026 (N_23026,N_22177,N_22294);
nor U23027 (N_23027,N_22286,N_22492);
and U23028 (N_23028,N_21958,N_22153);
and U23029 (N_23029,N_22149,N_21970);
nand U23030 (N_23030,N_22084,N_22313);
and U23031 (N_23031,N_22369,N_22237);
nor U23032 (N_23032,N_22442,N_22409);
and U23033 (N_23033,N_22446,N_22413);
nand U23034 (N_23034,N_22172,N_22089);
xnor U23035 (N_23035,N_21912,N_22286);
nand U23036 (N_23036,N_22330,N_22401);
and U23037 (N_23037,N_22266,N_22025);
nand U23038 (N_23038,N_22431,N_22067);
xor U23039 (N_23039,N_22356,N_22112);
nor U23040 (N_23040,N_22240,N_22266);
and U23041 (N_23041,N_22214,N_22303);
and U23042 (N_23042,N_22372,N_22136);
xnor U23043 (N_23043,N_22266,N_22308);
or U23044 (N_23044,N_22240,N_22075);
xor U23045 (N_23045,N_21987,N_22100);
nand U23046 (N_23046,N_22190,N_22160);
or U23047 (N_23047,N_22279,N_22044);
nand U23048 (N_23048,N_21948,N_22166);
xor U23049 (N_23049,N_22406,N_22336);
and U23050 (N_23050,N_22009,N_21906);
and U23051 (N_23051,N_22106,N_21939);
and U23052 (N_23052,N_21961,N_22141);
xnor U23053 (N_23053,N_22111,N_22476);
nand U23054 (N_23054,N_22408,N_22349);
and U23055 (N_23055,N_22406,N_22173);
nand U23056 (N_23056,N_21907,N_22422);
nand U23057 (N_23057,N_22003,N_22416);
or U23058 (N_23058,N_22281,N_22488);
xnor U23059 (N_23059,N_22335,N_22399);
nor U23060 (N_23060,N_22328,N_22439);
and U23061 (N_23061,N_22387,N_22110);
nand U23062 (N_23062,N_22238,N_22207);
or U23063 (N_23063,N_22369,N_22459);
xnor U23064 (N_23064,N_21961,N_22174);
xor U23065 (N_23065,N_22354,N_21972);
and U23066 (N_23066,N_21898,N_22443);
nand U23067 (N_23067,N_22478,N_22353);
and U23068 (N_23068,N_21911,N_22375);
xnor U23069 (N_23069,N_22301,N_22098);
xnor U23070 (N_23070,N_22085,N_22096);
nor U23071 (N_23071,N_22084,N_22062);
and U23072 (N_23072,N_22355,N_22237);
xor U23073 (N_23073,N_22234,N_22047);
or U23074 (N_23074,N_22306,N_22161);
nor U23075 (N_23075,N_22426,N_22250);
nor U23076 (N_23076,N_21999,N_21947);
and U23077 (N_23077,N_22402,N_22443);
xor U23078 (N_23078,N_22155,N_22309);
nor U23079 (N_23079,N_22322,N_22498);
xor U23080 (N_23080,N_21913,N_22317);
xnor U23081 (N_23081,N_22069,N_22138);
and U23082 (N_23082,N_21935,N_21989);
nand U23083 (N_23083,N_22233,N_22098);
and U23084 (N_23084,N_22052,N_22298);
and U23085 (N_23085,N_22118,N_21997);
nand U23086 (N_23086,N_22247,N_22044);
or U23087 (N_23087,N_22477,N_22115);
nand U23088 (N_23088,N_22472,N_22204);
nand U23089 (N_23089,N_22057,N_22152);
nor U23090 (N_23090,N_22472,N_22028);
xnor U23091 (N_23091,N_22203,N_22317);
nor U23092 (N_23092,N_22006,N_22147);
nor U23093 (N_23093,N_22047,N_22049);
xor U23094 (N_23094,N_22299,N_22290);
nor U23095 (N_23095,N_22030,N_22032);
nand U23096 (N_23096,N_22186,N_22471);
and U23097 (N_23097,N_22243,N_22483);
and U23098 (N_23098,N_21973,N_22457);
xnor U23099 (N_23099,N_22274,N_22014);
and U23100 (N_23100,N_22182,N_22452);
xor U23101 (N_23101,N_22087,N_22071);
nor U23102 (N_23102,N_21959,N_22123);
nor U23103 (N_23103,N_22108,N_22149);
nand U23104 (N_23104,N_22158,N_22402);
and U23105 (N_23105,N_22441,N_22445);
xor U23106 (N_23106,N_22486,N_22474);
and U23107 (N_23107,N_22304,N_22326);
and U23108 (N_23108,N_21921,N_22397);
or U23109 (N_23109,N_22120,N_22154);
and U23110 (N_23110,N_21988,N_22186);
and U23111 (N_23111,N_22243,N_22350);
and U23112 (N_23112,N_21903,N_21913);
nand U23113 (N_23113,N_21957,N_22487);
nor U23114 (N_23114,N_22165,N_22304);
xor U23115 (N_23115,N_22065,N_21997);
or U23116 (N_23116,N_22216,N_22479);
or U23117 (N_23117,N_21886,N_22395);
nand U23118 (N_23118,N_22204,N_21964);
and U23119 (N_23119,N_22417,N_22300);
xnor U23120 (N_23120,N_22416,N_22100);
nand U23121 (N_23121,N_22179,N_22198);
nand U23122 (N_23122,N_21946,N_22119);
xnor U23123 (N_23123,N_22357,N_22453);
nand U23124 (N_23124,N_22082,N_22284);
or U23125 (N_23125,N_22574,N_22548);
and U23126 (N_23126,N_22505,N_22781);
or U23127 (N_23127,N_22522,N_23035);
or U23128 (N_23128,N_22603,N_22747);
or U23129 (N_23129,N_22580,N_22982);
nor U23130 (N_23130,N_22838,N_22792);
and U23131 (N_23131,N_22585,N_23110);
or U23132 (N_23132,N_22993,N_23074);
nor U23133 (N_23133,N_22519,N_22961);
and U23134 (N_23134,N_23007,N_22782);
xnor U23135 (N_23135,N_22924,N_22698);
nor U23136 (N_23136,N_22570,N_22798);
and U23137 (N_23137,N_23099,N_22773);
and U23138 (N_23138,N_22926,N_22897);
or U23139 (N_23139,N_23045,N_22694);
nand U23140 (N_23140,N_23098,N_22659);
and U23141 (N_23141,N_22507,N_22651);
and U23142 (N_23142,N_22965,N_22801);
nor U23143 (N_23143,N_22776,N_23108);
or U23144 (N_23144,N_23012,N_22779);
xor U23145 (N_23145,N_22612,N_22707);
and U23146 (N_23146,N_22597,N_22606);
nor U23147 (N_23147,N_22885,N_22821);
xor U23148 (N_23148,N_23105,N_22508);
nor U23149 (N_23149,N_22509,N_22919);
nor U23150 (N_23150,N_22544,N_22980);
nand U23151 (N_23151,N_22736,N_22896);
and U23152 (N_23152,N_23075,N_23034);
nor U23153 (N_23153,N_22882,N_22725);
and U23154 (N_23154,N_22990,N_23070);
or U23155 (N_23155,N_22696,N_22527);
nand U23156 (N_23156,N_22648,N_23043);
xor U23157 (N_23157,N_22975,N_22667);
nand U23158 (N_23158,N_22640,N_22616);
and U23159 (N_23159,N_22869,N_22810);
nor U23160 (N_23160,N_23032,N_22905);
nor U23161 (N_23161,N_22845,N_22750);
xnor U23162 (N_23162,N_23063,N_23042);
nand U23163 (N_23163,N_22978,N_22786);
nand U23164 (N_23164,N_22662,N_22745);
and U23165 (N_23165,N_23083,N_22578);
nor U23166 (N_23166,N_22940,N_22976);
nand U23167 (N_23167,N_22774,N_22877);
or U23168 (N_23168,N_23091,N_22604);
or U23169 (N_23169,N_22681,N_22756);
or U23170 (N_23170,N_22683,N_22890);
and U23171 (N_23171,N_22692,N_22675);
nand U23172 (N_23172,N_22899,N_22611);
xnor U23173 (N_23173,N_22695,N_23020);
nand U23174 (N_23174,N_23031,N_22615);
nand U23175 (N_23175,N_22970,N_23018);
or U23176 (N_23176,N_22589,N_22793);
or U23177 (N_23177,N_22730,N_22534);
nand U23178 (N_23178,N_22533,N_22958);
nor U23179 (N_23179,N_22956,N_22992);
nor U23180 (N_23180,N_22904,N_22946);
and U23181 (N_23181,N_22920,N_22629);
and U23182 (N_23182,N_22915,N_22559);
nor U23183 (N_23183,N_23080,N_22962);
or U23184 (N_23184,N_22973,N_22518);
nand U23185 (N_23185,N_22858,N_23086);
nand U23186 (N_23186,N_22770,N_22727);
nand U23187 (N_23187,N_22828,N_23118);
nor U23188 (N_23188,N_22822,N_22647);
or U23189 (N_23189,N_23064,N_23071);
xor U23190 (N_23190,N_23005,N_22688);
nand U23191 (N_23191,N_22878,N_23114);
nand U23192 (N_23192,N_22985,N_23121);
nor U23193 (N_23193,N_22678,N_22861);
or U23194 (N_23194,N_22729,N_22785);
nand U23195 (N_23195,N_22656,N_22718);
nand U23196 (N_23196,N_22663,N_23019);
or U23197 (N_23197,N_22528,N_22853);
nor U23198 (N_23198,N_23077,N_23009);
or U23199 (N_23199,N_22733,N_23095);
xnor U23200 (N_23200,N_22637,N_23062);
xor U23201 (N_23201,N_22622,N_22842);
or U23202 (N_23202,N_22954,N_22598);
nor U23203 (N_23203,N_22847,N_22511);
xnor U23204 (N_23204,N_22969,N_22642);
or U23205 (N_23205,N_22816,N_22711);
and U23206 (N_23206,N_22631,N_22942);
nand U23207 (N_23207,N_22743,N_22766);
or U23208 (N_23208,N_22561,N_23106);
and U23209 (N_23209,N_22911,N_22800);
xnor U23210 (N_23210,N_22824,N_22555);
xor U23211 (N_23211,N_23021,N_22762);
or U23212 (N_23212,N_23119,N_23078);
nand U23213 (N_23213,N_22596,N_23059);
xnor U23214 (N_23214,N_22971,N_22901);
and U23215 (N_23215,N_22851,N_23017);
nor U23216 (N_23216,N_23092,N_22545);
nand U23217 (N_23217,N_22997,N_22796);
or U23218 (N_23218,N_22714,N_23085);
and U23219 (N_23219,N_22812,N_23015);
nand U23220 (N_23220,N_22660,N_22655);
or U23221 (N_23221,N_22516,N_23024);
or U23222 (N_23222,N_22863,N_22582);
nor U23223 (N_23223,N_22741,N_22968);
and U23224 (N_23224,N_23067,N_22934);
xor U23225 (N_23225,N_23057,N_23004);
nor U23226 (N_23226,N_22674,N_22679);
nor U23227 (N_23227,N_22617,N_22814);
or U23228 (N_23228,N_22862,N_22523);
xnor U23229 (N_23229,N_22778,N_22873);
xor U23230 (N_23230,N_22728,N_22805);
xor U23231 (N_23231,N_22979,N_22587);
or U23232 (N_23232,N_22795,N_23052);
nor U23233 (N_23233,N_22550,N_22610);
or U23234 (N_23234,N_22646,N_22753);
or U23235 (N_23235,N_22588,N_22564);
or U23236 (N_23236,N_22569,N_22953);
nand U23237 (N_23237,N_22907,N_22691);
and U23238 (N_23238,N_22825,N_22594);
nand U23239 (N_23239,N_22680,N_22676);
xnor U23240 (N_23240,N_22767,N_22602);
nor U23241 (N_23241,N_22830,N_23051);
and U23242 (N_23242,N_22951,N_22627);
nand U23243 (N_23243,N_22738,N_22556);
nor U23244 (N_23244,N_23088,N_23014);
nor U23245 (N_23245,N_23084,N_22558);
xnor U23246 (N_23246,N_22909,N_23011);
nand U23247 (N_23247,N_22826,N_22848);
xnor U23248 (N_23248,N_22775,N_23101);
or U23249 (N_23249,N_22618,N_23104);
or U23250 (N_23250,N_22697,N_22693);
nor U23251 (N_23251,N_22948,N_23022);
nand U23252 (N_23252,N_23029,N_22723);
nor U23253 (N_23253,N_22840,N_22880);
or U23254 (N_23254,N_22744,N_22576);
xnor U23255 (N_23255,N_22987,N_22687);
nand U23256 (N_23256,N_23093,N_22790);
xnor U23257 (N_23257,N_23033,N_22634);
or U23258 (N_23258,N_22554,N_23013);
nor U23259 (N_23259,N_23041,N_22866);
xor U23260 (N_23260,N_22945,N_22636);
and U23261 (N_23261,N_22963,N_22713);
nand U23262 (N_23262,N_22595,N_23037);
xnor U23263 (N_23263,N_22834,N_22553);
nor U23264 (N_23264,N_22964,N_23003);
nor U23265 (N_23265,N_22734,N_22807);
or U23266 (N_23266,N_22635,N_22868);
nor U23267 (N_23267,N_22758,N_22536);
or U23268 (N_23268,N_22630,N_23023);
xnor U23269 (N_23269,N_22565,N_22930);
nand U23270 (N_23270,N_22833,N_22887);
and U23271 (N_23271,N_22607,N_22669);
and U23272 (N_23272,N_22895,N_22923);
nand U23273 (N_23273,N_22571,N_22879);
or U23274 (N_23274,N_22567,N_23055);
nand U23275 (N_23275,N_22906,N_22941);
xor U23276 (N_23276,N_22531,N_22755);
xnor U23277 (N_23277,N_22925,N_23123);
nand U23278 (N_23278,N_23030,N_22540);
and U23279 (N_23279,N_22974,N_22552);
and U23280 (N_23280,N_23079,N_22850);
nor U23281 (N_23281,N_22699,N_22605);
xor U23282 (N_23282,N_22892,N_22715);
or U23283 (N_23283,N_22752,N_22966);
or U23284 (N_23284,N_22783,N_22939);
nor U23285 (N_23285,N_22721,N_22742);
nor U23286 (N_23286,N_22671,N_22996);
xor U23287 (N_23287,N_22638,N_22652);
nor U23288 (N_23288,N_23046,N_22520);
nand U23289 (N_23289,N_22893,N_23001);
and U23290 (N_23290,N_23025,N_22563);
xor U23291 (N_23291,N_22947,N_22658);
or U23292 (N_23292,N_23039,N_22936);
nor U23293 (N_23293,N_22836,N_22600);
nor U23294 (N_23294,N_22809,N_22802);
nor U23295 (N_23295,N_22900,N_22748);
and U23296 (N_23296,N_22746,N_22672);
xnor U23297 (N_23297,N_22938,N_23006);
nor U23298 (N_23298,N_22872,N_23087);
or U23299 (N_23299,N_22501,N_22759);
xnor U23300 (N_23300,N_22760,N_22855);
xnor U23301 (N_23301,N_22769,N_22922);
or U23302 (N_23302,N_23027,N_23040);
and U23303 (N_23303,N_22876,N_23036);
xor U23304 (N_23304,N_23120,N_22670);
or U23305 (N_23305,N_22989,N_22967);
xor U23306 (N_23306,N_23016,N_22619);
and U23307 (N_23307,N_22983,N_22804);
nand U23308 (N_23308,N_22535,N_22891);
nand U23309 (N_23309,N_22547,N_22739);
or U23310 (N_23310,N_22856,N_22846);
nand U23311 (N_23311,N_22806,N_22815);
xor U23312 (N_23312,N_22572,N_22543);
nor U23313 (N_23313,N_22628,N_22551);
nor U23314 (N_23314,N_22912,N_22959);
nor U23315 (N_23315,N_22706,N_23097);
xnor U23316 (N_23316,N_23026,N_22771);
and U23317 (N_23317,N_22705,N_22632);
nand U23318 (N_23318,N_22537,N_22532);
nand U23319 (N_23319,N_22949,N_22944);
and U23320 (N_23320,N_22590,N_23076);
nor U23321 (N_23321,N_22829,N_22910);
nand U23322 (N_23322,N_22735,N_22512);
nor U23323 (N_23323,N_22685,N_22813);
or U23324 (N_23324,N_22883,N_22720);
xor U23325 (N_23325,N_22633,N_22927);
xnor U23326 (N_23326,N_22562,N_22625);
nand U23327 (N_23327,N_22831,N_22521);
or U23328 (N_23328,N_22724,N_22981);
xor U23329 (N_23329,N_22881,N_23010);
or U23330 (N_23330,N_22654,N_23061);
nor U23331 (N_23331,N_22995,N_22599);
and U23332 (N_23332,N_22972,N_22665);
xor U23333 (N_23333,N_22731,N_23109);
nand U23334 (N_23334,N_22888,N_22668);
nor U23335 (N_23335,N_23102,N_22709);
nor U23336 (N_23336,N_22504,N_22579);
xnor U23337 (N_23337,N_22716,N_22864);
or U23338 (N_23338,N_22643,N_22898);
xor U23339 (N_23339,N_22539,N_23107);
xor U23340 (N_23340,N_22871,N_23038);
and U23341 (N_23341,N_22991,N_22870);
nand U23342 (N_23342,N_22933,N_22852);
or U23343 (N_23343,N_22772,N_22732);
or U23344 (N_23344,N_22921,N_22935);
nor U23345 (N_23345,N_22682,N_22614);
nor U23346 (N_23346,N_22803,N_23081);
or U23347 (N_23347,N_22583,N_22557);
xnor U23348 (N_23348,N_22722,N_23049);
or U23349 (N_23349,N_22797,N_23060);
and U23350 (N_23350,N_22649,N_23112);
xnor U23351 (N_23351,N_22977,N_22931);
nor U23352 (N_23352,N_22808,N_22929);
nand U23353 (N_23353,N_22524,N_22865);
or U23354 (N_23354,N_22513,N_22994);
or U23355 (N_23355,N_22684,N_22517);
and U23356 (N_23356,N_23044,N_22549);
or U23357 (N_23357,N_22839,N_23056);
or U23358 (N_23358,N_23072,N_22515);
and U23359 (N_23359,N_22650,N_22928);
or U23360 (N_23360,N_22609,N_23073);
and U23361 (N_23361,N_22820,N_23115);
or U23362 (N_23362,N_22529,N_22791);
nand U23363 (N_23363,N_22677,N_22624);
nor U23364 (N_23364,N_22999,N_22704);
and U23365 (N_23365,N_22884,N_23116);
xnor U23366 (N_23366,N_22584,N_22566);
nand U23367 (N_23367,N_23066,N_22844);
nand U23368 (N_23368,N_22560,N_22960);
nand U23369 (N_23369,N_22998,N_22641);
xor U23370 (N_23370,N_23096,N_22645);
xnor U23371 (N_23371,N_22768,N_22573);
nand U23372 (N_23372,N_22986,N_22894);
and U23373 (N_23373,N_22788,N_22726);
nor U23374 (N_23374,N_22908,N_22593);
nand U23375 (N_23375,N_22666,N_22859);
xor U23376 (N_23376,N_22937,N_22874);
xor U23377 (N_23377,N_22541,N_22754);
nand U23378 (N_23378,N_22827,N_22837);
and U23379 (N_23379,N_22689,N_22932);
nand U23380 (N_23380,N_22644,N_22765);
nor U23381 (N_23381,N_22854,N_22601);
nand U23382 (N_23382,N_22664,N_22917);
and U23383 (N_23383,N_22832,N_22613);
nor U23384 (N_23384,N_22957,N_22546);
or U23385 (N_23385,N_22712,N_22903);
xnor U23386 (N_23386,N_22591,N_22918);
xnor U23387 (N_23387,N_22860,N_22955);
nor U23388 (N_23388,N_23008,N_22787);
or U23389 (N_23389,N_22777,N_23090);
and U23390 (N_23390,N_22500,N_22620);
or U23391 (N_23391,N_22701,N_22503);
xnor U23392 (N_23392,N_22823,N_22538);
xor U23393 (N_23393,N_22526,N_22889);
nor U23394 (N_23394,N_23047,N_22690);
nand U23395 (N_23395,N_23053,N_22568);
nor U23396 (N_23396,N_22717,N_22510);
nand U23397 (N_23397,N_22525,N_22811);
nand U23398 (N_23398,N_22657,N_22703);
nand U23399 (N_23399,N_22626,N_23028);
nor U23400 (N_23400,N_22700,N_23065);
xnor U23401 (N_23401,N_22740,N_22621);
nand U23402 (N_23402,N_22849,N_22506);
nand U23403 (N_23403,N_23054,N_23068);
and U23404 (N_23404,N_23069,N_22902);
xor U23405 (N_23405,N_22708,N_22749);
or U23406 (N_23406,N_22780,N_23117);
and U23407 (N_23407,N_22794,N_22702);
xnor U23408 (N_23408,N_22914,N_22952);
nor U23409 (N_23409,N_22763,N_22719);
nor U23410 (N_23410,N_22784,N_22819);
nand U23411 (N_23411,N_22789,N_22514);
nand U23412 (N_23412,N_22661,N_23094);
xnor U23413 (N_23413,N_22913,N_22653);
nand U23414 (N_23414,N_22586,N_22751);
and U23415 (N_23415,N_22843,N_22799);
xnor U23416 (N_23416,N_22984,N_22950);
or U23417 (N_23417,N_23113,N_22673);
and U23418 (N_23418,N_22886,N_23122);
or U23419 (N_23419,N_22757,N_22502);
and U23420 (N_23420,N_23000,N_22867);
nand U23421 (N_23421,N_22623,N_22530);
nand U23422 (N_23422,N_22764,N_22943);
or U23423 (N_23423,N_22875,N_23089);
xor U23424 (N_23424,N_22592,N_22857);
nor U23425 (N_23425,N_22577,N_22710);
xnor U23426 (N_23426,N_22841,N_23100);
and U23427 (N_23427,N_22542,N_23050);
or U23428 (N_23428,N_23002,N_23111);
or U23429 (N_23429,N_22737,N_22761);
or U23430 (N_23430,N_23048,N_23058);
nor U23431 (N_23431,N_23124,N_23082);
and U23432 (N_23432,N_22988,N_22608);
and U23433 (N_23433,N_22916,N_23103);
xnor U23434 (N_23434,N_22818,N_22639);
and U23435 (N_23435,N_22686,N_22817);
nor U23436 (N_23436,N_22575,N_22581);
and U23437 (N_23437,N_22835,N_22896);
xor U23438 (N_23438,N_22947,N_22673);
and U23439 (N_23439,N_22663,N_22984);
or U23440 (N_23440,N_22740,N_22771);
or U23441 (N_23441,N_22594,N_22729);
xor U23442 (N_23442,N_22844,N_22921);
nor U23443 (N_23443,N_22635,N_22906);
xor U23444 (N_23444,N_22572,N_22758);
xnor U23445 (N_23445,N_22700,N_22565);
nand U23446 (N_23446,N_22777,N_22591);
and U23447 (N_23447,N_22760,N_22519);
nor U23448 (N_23448,N_22610,N_22695);
and U23449 (N_23449,N_23024,N_22792);
or U23450 (N_23450,N_22797,N_23041);
nand U23451 (N_23451,N_23017,N_22674);
nor U23452 (N_23452,N_22633,N_22769);
and U23453 (N_23453,N_22806,N_22860);
xnor U23454 (N_23454,N_22628,N_23037);
and U23455 (N_23455,N_22595,N_22627);
or U23456 (N_23456,N_22978,N_22994);
or U23457 (N_23457,N_22908,N_22995);
xnor U23458 (N_23458,N_22665,N_23057);
nor U23459 (N_23459,N_23091,N_22628);
xnor U23460 (N_23460,N_23047,N_22814);
nor U23461 (N_23461,N_22948,N_22597);
or U23462 (N_23462,N_22788,N_22622);
nor U23463 (N_23463,N_22796,N_22980);
or U23464 (N_23464,N_22994,N_22549);
or U23465 (N_23465,N_22582,N_22979);
nand U23466 (N_23466,N_23107,N_22759);
xor U23467 (N_23467,N_22743,N_22923);
nand U23468 (N_23468,N_23031,N_22869);
nor U23469 (N_23469,N_22925,N_22568);
nand U23470 (N_23470,N_22756,N_23097);
and U23471 (N_23471,N_22505,N_22999);
and U23472 (N_23472,N_22756,N_23017);
nor U23473 (N_23473,N_22771,N_22621);
nand U23474 (N_23474,N_22536,N_22541);
nand U23475 (N_23475,N_22849,N_23025);
and U23476 (N_23476,N_22844,N_23030);
and U23477 (N_23477,N_22648,N_22519);
nand U23478 (N_23478,N_22812,N_22774);
and U23479 (N_23479,N_23111,N_22922);
xnor U23480 (N_23480,N_22638,N_22700);
and U23481 (N_23481,N_22965,N_23098);
and U23482 (N_23482,N_22532,N_22714);
or U23483 (N_23483,N_22584,N_22773);
nor U23484 (N_23484,N_22510,N_22788);
xnor U23485 (N_23485,N_22699,N_22550);
nand U23486 (N_23486,N_23082,N_22967);
or U23487 (N_23487,N_22846,N_22808);
nor U23488 (N_23488,N_22769,N_23006);
or U23489 (N_23489,N_22558,N_22864);
and U23490 (N_23490,N_23056,N_22732);
and U23491 (N_23491,N_22585,N_22738);
nand U23492 (N_23492,N_22907,N_22668);
and U23493 (N_23493,N_23067,N_23006);
or U23494 (N_23494,N_22874,N_23084);
nor U23495 (N_23495,N_23044,N_22874);
or U23496 (N_23496,N_23041,N_23091);
nand U23497 (N_23497,N_22929,N_22588);
nor U23498 (N_23498,N_22915,N_22566);
and U23499 (N_23499,N_22601,N_22750);
and U23500 (N_23500,N_22664,N_22937);
nand U23501 (N_23501,N_22876,N_22867);
or U23502 (N_23502,N_22943,N_22748);
xor U23503 (N_23503,N_22938,N_22611);
or U23504 (N_23504,N_22606,N_22936);
xnor U23505 (N_23505,N_22570,N_22906);
or U23506 (N_23506,N_22788,N_23121);
and U23507 (N_23507,N_22805,N_22851);
xor U23508 (N_23508,N_23016,N_22746);
xor U23509 (N_23509,N_23011,N_22844);
nand U23510 (N_23510,N_23004,N_22958);
nand U23511 (N_23511,N_23056,N_22930);
nor U23512 (N_23512,N_23100,N_22941);
nand U23513 (N_23513,N_22905,N_22525);
and U23514 (N_23514,N_22597,N_22569);
nor U23515 (N_23515,N_22992,N_22513);
or U23516 (N_23516,N_22928,N_22929);
nor U23517 (N_23517,N_22675,N_22737);
nor U23518 (N_23518,N_23121,N_22944);
nor U23519 (N_23519,N_22806,N_22917);
xnor U23520 (N_23520,N_23067,N_22650);
xor U23521 (N_23521,N_22820,N_23111);
and U23522 (N_23522,N_23041,N_22655);
nor U23523 (N_23523,N_22843,N_22900);
or U23524 (N_23524,N_22759,N_22637);
xor U23525 (N_23525,N_22951,N_22516);
nor U23526 (N_23526,N_22603,N_22790);
nand U23527 (N_23527,N_22508,N_22527);
nor U23528 (N_23528,N_22534,N_22690);
and U23529 (N_23529,N_22635,N_22620);
nand U23530 (N_23530,N_22814,N_23032);
or U23531 (N_23531,N_23057,N_23026);
xor U23532 (N_23532,N_23039,N_23048);
nor U23533 (N_23533,N_22802,N_22689);
nor U23534 (N_23534,N_22841,N_22680);
and U23535 (N_23535,N_22848,N_23120);
xnor U23536 (N_23536,N_22726,N_23022);
or U23537 (N_23537,N_22996,N_22730);
and U23538 (N_23538,N_23039,N_22844);
and U23539 (N_23539,N_22595,N_22834);
nand U23540 (N_23540,N_23021,N_22974);
and U23541 (N_23541,N_22700,N_22557);
nand U23542 (N_23542,N_23011,N_22837);
xor U23543 (N_23543,N_22849,N_22991);
or U23544 (N_23544,N_23007,N_22647);
nand U23545 (N_23545,N_22515,N_22502);
or U23546 (N_23546,N_22813,N_22715);
nor U23547 (N_23547,N_23112,N_22592);
or U23548 (N_23548,N_23031,N_23001);
or U23549 (N_23549,N_22832,N_23055);
and U23550 (N_23550,N_22932,N_22806);
and U23551 (N_23551,N_22786,N_22661);
or U23552 (N_23552,N_22771,N_22748);
nand U23553 (N_23553,N_23007,N_22678);
and U23554 (N_23554,N_22988,N_22921);
or U23555 (N_23555,N_23108,N_22847);
and U23556 (N_23556,N_22878,N_22875);
nand U23557 (N_23557,N_22545,N_22975);
and U23558 (N_23558,N_22936,N_23078);
and U23559 (N_23559,N_23016,N_22979);
nand U23560 (N_23560,N_22941,N_23083);
and U23561 (N_23561,N_22585,N_22576);
nand U23562 (N_23562,N_22943,N_22845);
or U23563 (N_23563,N_22718,N_22845);
nor U23564 (N_23564,N_22820,N_22623);
nor U23565 (N_23565,N_22904,N_22678);
or U23566 (N_23566,N_22695,N_23076);
nand U23567 (N_23567,N_23114,N_22862);
nor U23568 (N_23568,N_22661,N_22524);
nand U23569 (N_23569,N_22582,N_23083);
or U23570 (N_23570,N_22617,N_22600);
and U23571 (N_23571,N_22764,N_22540);
nand U23572 (N_23572,N_23024,N_22692);
nand U23573 (N_23573,N_22740,N_22938);
xnor U23574 (N_23574,N_22785,N_23082);
or U23575 (N_23575,N_22645,N_22833);
nand U23576 (N_23576,N_22970,N_23037);
nand U23577 (N_23577,N_23041,N_22579);
nand U23578 (N_23578,N_23121,N_23008);
xnor U23579 (N_23579,N_22875,N_22962);
xor U23580 (N_23580,N_22963,N_23082);
nand U23581 (N_23581,N_23031,N_22723);
xor U23582 (N_23582,N_22558,N_23056);
nand U23583 (N_23583,N_22754,N_22863);
and U23584 (N_23584,N_22541,N_23070);
and U23585 (N_23585,N_22780,N_22847);
xor U23586 (N_23586,N_23030,N_22906);
or U23587 (N_23587,N_22887,N_22818);
xor U23588 (N_23588,N_22572,N_22640);
or U23589 (N_23589,N_22858,N_22763);
nor U23590 (N_23590,N_22699,N_22960);
nand U23591 (N_23591,N_22805,N_22708);
nor U23592 (N_23592,N_22960,N_22917);
or U23593 (N_23593,N_22900,N_22913);
nor U23594 (N_23594,N_22831,N_22557);
and U23595 (N_23595,N_22563,N_22787);
or U23596 (N_23596,N_22711,N_22955);
xor U23597 (N_23597,N_23103,N_22941);
nand U23598 (N_23598,N_23100,N_22627);
xnor U23599 (N_23599,N_22860,N_23067);
and U23600 (N_23600,N_22623,N_23033);
or U23601 (N_23601,N_22692,N_22846);
and U23602 (N_23602,N_22829,N_22580);
xor U23603 (N_23603,N_22591,N_22910);
nor U23604 (N_23604,N_22659,N_22606);
and U23605 (N_23605,N_22832,N_22884);
nor U23606 (N_23606,N_22874,N_23065);
xor U23607 (N_23607,N_22612,N_22701);
nor U23608 (N_23608,N_22608,N_22578);
nor U23609 (N_23609,N_23076,N_22852);
and U23610 (N_23610,N_22537,N_22728);
nor U23611 (N_23611,N_22763,N_22723);
nor U23612 (N_23612,N_22958,N_22621);
nand U23613 (N_23613,N_22808,N_22612);
or U23614 (N_23614,N_22976,N_22705);
xnor U23615 (N_23615,N_22625,N_22655);
or U23616 (N_23616,N_22815,N_22873);
or U23617 (N_23617,N_22949,N_22615);
xnor U23618 (N_23618,N_22741,N_22503);
and U23619 (N_23619,N_22833,N_23066);
nand U23620 (N_23620,N_23024,N_22582);
nand U23621 (N_23621,N_22541,N_22849);
or U23622 (N_23622,N_23069,N_22540);
and U23623 (N_23623,N_22501,N_22556);
nor U23624 (N_23624,N_22535,N_22789);
nor U23625 (N_23625,N_23059,N_22773);
or U23626 (N_23626,N_22524,N_22575);
nand U23627 (N_23627,N_23015,N_22856);
or U23628 (N_23628,N_22937,N_23072);
nand U23629 (N_23629,N_22639,N_22973);
xor U23630 (N_23630,N_22964,N_22547);
or U23631 (N_23631,N_23018,N_22815);
xor U23632 (N_23632,N_22557,N_22719);
xnor U23633 (N_23633,N_22682,N_22647);
nor U23634 (N_23634,N_23100,N_22866);
nand U23635 (N_23635,N_23069,N_22668);
nor U23636 (N_23636,N_22923,N_23027);
nand U23637 (N_23637,N_22519,N_22912);
xor U23638 (N_23638,N_22967,N_22532);
and U23639 (N_23639,N_23078,N_22821);
and U23640 (N_23640,N_22915,N_23073);
nand U23641 (N_23641,N_23047,N_23031);
nor U23642 (N_23642,N_23108,N_22976);
nand U23643 (N_23643,N_22554,N_22979);
nand U23644 (N_23644,N_22546,N_22644);
nand U23645 (N_23645,N_22689,N_22966);
nand U23646 (N_23646,N_22919,N_22887);
nor U23647 (N_23647,N_22520,N_22557);
nand U23648 (N_23648,N_22809,N_22976);
nand U23649 (N_23649,N_22696,N_22773);
nor U23650 (N_23650,N_22967,N_22647);
nor U23651 (N_23651,N_22967,N_22577);
xnor U23652 (N_23652,N_22520,N_22738);
nor U23653 (N_23653,N_22700,N_23118);
nand U23654 (N_23654,N_22721,N_22893);
or U23655 (N_23655,N_22605,N_23031);
nor U23656 (N_23656,N_22896,N_22612);
xor U23657 (N_23657,N_22721,N_22756);
nor U23658 (N_23658,N_23105,N_22757);
or U23659 (N_23659,N_22718,N_22996);
xor U23660 (N_23660,N_22722,N_22890);
nand U23661 (N_23661,N_22804,N_22584);
nand U23662 (N_23662,N_23016,N_22562);
nor U23663 (N_23663,N_22986,N_23034);
or U23664 (N_23664,N_22824,N_22785);
nand U23665 (N_23665,N_23005,N_22987);
and U23666 (N_23666,N_22658,N_23018);
nand U23667 (N_23667,N_23087,N_23014);
and U23668 (N_23668,N_22985,N_23043);
nor U23669 (N_23669,N_22506,N_23016);
or U23670 (N_23670,N_22856,N_22822);
xor U23671 (N_23671,N_23001,N_22522);
xor U23672 (N_23672,N_22774,N_22665);
xnor U23673 (N_23673,N_22602,N_22641);
xnor U23674 (N_23674,N_23088,N_22648);
nor U23675 (N_23675,N_22603,N_22538);
and U23676 (N_23676,N_22861,N_23024);
nor U23677 (N_23677,N_22508,N_23034);
nor U23678 (N_23678,N_22974,N_22710);
xor U23679 (N_23679,N_22509,N_22676);
nor U23680 (N_23680,N_22772,N_22540);
nor U23681 (N_23681,N_22896,N_22817);
nand U23682 (N_23682,N_23025,N_22659);
nor U23683 (N_23683,N_22528,N_22507);
nand U23684 (N_23684,N_22907,N_22798);
nor U23685 (N_23685,N_22527,N_23004);
nor U23686 (N_23686,N_22943,N_23013);
and U23687 (N_23687,N_22654,N_22863);
xnor U23688 (N_23688,N_23036,N_22605);
nand U23689 (N_23689,N_22514,N_22965);
nor U23690 (N_23690,N_22566,N_22881);
and U23691 (N_23691,N_22537,N_22619);
nand U23692 (N_23692,N_22925,N_22945);
nand U23693 (N_23693,N_22700,N_23045);
xnor U23694 (N_23694,N_22774,N_22718);
and U23695 (N_23695,N_22938,N_22739);
and U23696 (N_23696,N_23056,N_22508);
nand U23697 (N_23697,N_22530,N_22853);
xnor U23698 (N_23698,N_22706,N_22714);
nand U23699 (N_23699,N_22968,N_22871);
or U23700 (N_23700,N_22667,N_23051);
nand U23701 (N_23701,N_22700,N_22989);
nand U23702 (N_23702,N_22882,N_22734);
nand U23703 (N_23703,N_23036,N_22550);
nand U23704 (N_23704,N_22711,N_22794);
nor U23705 (N_23705,N_22991,N_22706);
or U23706 (N_23706,N_22894,N_22716);
nand U23707 (N_23707,N_22927,N_22949);
xor U23708 (N_23708,N_23016,N_23083);
nand U23709 (N_23709,N_22921,N_22500);
or U23710 (N_23710,N_22900,N_22502);
nand U23711 (N_23711,N_23027,N_23008);
nor U23712 (N_23712,N_22924,N_22674);
nand U23713 (N_23713,N_23010,N_23086);
or U23714 (N_23714,N_22785,N_22976);
and U23715 (N_23715,N_22870,N_22556);
and U23716 (N_23716,N_22596,N_23013);
nor U23717 (N_23717,N_23121,N_22717);
xnor U23718 (N_23718,N_22747,N_22707);
nor U23719 (N_23719,N_22906,N_22510);
and U23720 (N_23720,N_23123,N_22997);
nor U23721 (N_23721,N_22721,N_22582);
nor U23722 (N_23722,N_22655,N_22548);
xor U23723 (N_23723,N_22667,N_22839);
nor U23724 (N_23724,N_23039,N_22862);
nor U23725 (N_23725,N_22671,N_22667);
and U23726 (N_23726,N_22866,N_22650);
nand U23727 (N_23727,N_22919,N_22774);
nand U23728 (N_23728,N_22850,N_22925);
nor U23729 (N_23729,N_23011,N_23073);
nor U23730 (N_23730,N_22526,N_22936);
nor U23731 (N_23731,N_22705,N_23058);
xor U23732 (N_23732,N_22827,N_22770);
xnor U23733 (N_23733,N_22606,N_22535);
xnor U23734 (N_23734,N_22832,N_22720);
nand U23735 (N_23735,N_22819,N_23007);
or U23736 (N_23736,N_22614,N_22946);
xor U23737 (N_23737,N_22755,N_22655);
or U23738 (N_23738,N_23122,N_22921);
or U23739 (N_23739,N_22826,N_22997);
and U23740 (N_23740,N_22814,N_23113);
or U23741 (N_23741,N_23090,N_22950);
nor U23742 (N_23742,N_22744,N_22527);
or U23743 (N_23743,N_23046,N_23118);
xor U23744 (N_23744,N_22654,N_23003);
xnor U23745 (N_23745,N_23055,N_22706);
nor U23746 (N_23746,N_22888,N_22710);
and U23747 (N_23747,N_22765,N_22827);
or U23748 (N_23748,N_22565,N_22889);
nor U23749 (N_23749,N_22925,N_23031);
nor U23750 (N_23750,N_23165,N_23198);
nand U23751 (N_23751,N_23462,N_23534);
xnor U23752 (N_23752,N_23632,N_23514);
xnor U23753 (N_23753,N_23718,N_23522);
nand U23754 (N_23754,N_23188,N_23590);
nand U23755 (N_23755,N_23459,N_23730);
nand U23756 (N_23756,N_23136,N_23502);
nor U23757 (N_23757,N_23224,N_23129);
nand U23758 (N_23758,N_23394,N_23527);
xnor U23759 (N_23759,N_23339,N_23252);
nor U23760 (N_23760,N_23728,N_23386);
xor U23761 (N_23761,N_23137,N_23537);
xnor U23762 (N_23762,N_23285,N_23202);
or U23763 (N_23763,N_23161,N_23562);
nor U23764 (N_23764,N_23688,N_23709);
xnor U23765 (N_23765,N_23524,N_23154);
and U23766 (N_23766,N_23417,N_23210);
nand U23767 (N_23767,N_23215,N_23484);
and U23768 (N_23768,N_23146,N_23474);
xor U23769 (N_23769,N_23585,N_23563);
nor U23770 (N_23770,N_23613,N_23656);
nor U23771 (N_23771,N_23406,N_23240);
and U23772 (N_23772,N_23259,N_23282);
nand U23773 (N_23773,N_23148,N_23635);
xor U23774 (N_23774,N_23349,N_23598);
or U23775 (N_23775,N_23315,N_23445);
and U23776 (N_23776,N_23227,N_23615);
nor U23777 (N_23777,N_23361,N_23271);
or U23778 (N_23778,N_23389,N_23393);
nor U23779 (N_23779,N_23722,N_23267);
nand U23780 (N_23780,N_23644,N_23345);
nor U23781 (N_23781,N_23144,N_23147);
xnor U23782 (N_23782,N_23641,N_23281);
nor U23783 (N_23783,N_23263,N_23592);
or U23784 (N_23784,N_23143,N_23627);
or U23785 (N_23785,N_23492,N_23691);
xnor U23786 (N_23786,N_23335,N_23578);
nand U23787 (N_23787,N_23682,N_23533);
and U23788 (N_23788,N_23631,N_23253);
xor U23789 (N_23789,N_23211,N_23535);
or U23790 (N_23790,N_23642,N_23217);
or U23791 (N_23791,N_23337,N_23530);
and U23792 (N_23792,N_23643,N_23612);
nor U23793 (N_23793,N_23673,N_23197);
and U23794 (N_23794,N_23424,N_23246);
nand U23795 (N_23795,N_23347,N_23367);
or U23796 (N_23796,N_23748,N_23505);
or U23797 (N_23797,N_23658,N_23395);
xnor U23798 (N_23798,N_23307,N_23278);
nor U23799 (N_23799,N_23482,N_23304);
nor U23800 (N_23800,N_23152,N_23457);
and U23801 (N_23801,N_23571,N_23473);
nor U23802 (N_23802,N_23580,N_23561);
xnor U23803 (N_23803,N_23189,N_23584);
and U23804 (N_23804,N_23277,N_23579);
and U23805 (N_23805,N_23149,N_23471);
nor U23806 (N_23806,N_23170,N_23316);
and U23807 (N_23807,N_23412,N_23679);
xor U23808 (N_23808,N_23551,N_23242);
and U23809 (N_23809,N_23485,N_23498);
nand U23810 (N_23810,N_23195,N_23302);
or U23811 (N_23811,N_23477,N_23313);
nand U23812 (N_23812,N_23318,N_23626);
nor U23813 (N_23813,N_23439,N_23745);
nor U23814 (N_23814,N_23620,N_23531);
xnor U23815 (N_23815,N_23448,N_23697);
xnor U23816 (N_23816,N_23290,N_23454);
nor U23817 (N_23817,N_23734,N_23659);
or U23818 (N_23818,N_23173,N_23350);
and U23819 (N_23819,N_23279,N_23251);
nor U23820 (N_23820,N_23223,N_23645);
or U23821 (N_23821,N_23175,N_23408);
xor U23822 (N_23822,N_23449,N_23567);
and U23823 (N_23823,N_23131,N_23591);
and U23824 (N_23824,N_23651,N_23736);
nor U23825 (N_23825,N_23258,N_23291);
or U23826 (N_23826,N_23469,N_23637);
nor U23827 (N_23827,N_23132,N_23476);
xnor U23828 (N_23828,N_23690,N_23647);
nand U23829 (N_23829,N_23687,N_23622);
and U23830 (N_23830,N_23694,N_23625);
and U23831 (N_23831,N_23411,N_23300);
and U23832 (N_23832,N_23582,N_23128);
and U23833 (N_23833,N_23553,N_23397);
nand U23834 (N_23834,N_23159,N_23216);
nor U23835 (N_23835,N_23499,N_23487);
nor U23836 (N_23836,N_23497,N_23603);
nor U23837 (N_23837,N_23156,N_23639);
and U23838 (N_23838,N_23396,N_23362);
or U23839 (N_23839,N_23623,N_23155);
xnor U23840 (N_23840,N_23384,N_23207);
xnor U23841 (N_23841,N_23440,N_23569);
xor U23842 (N_23842,N_23648,N_23262);
and U23843 (N_23843,N_23385,N_23157);
nand U23844 (N_23844,N_23238,N_23606);
xnor U23845 (N_23845,N_23650,N_23244);
nor U23846 (N_23846,N_23407,N_23654);
and U23847 (N_23847,N_23272,N_23324);
and U23848 (N_23848,N_23593,N_23204);
and U23849 (N_23849,N_23741,N_23518);
nand U23850 (N_23850,N_23400,N_23556);
nand U23851 (N_23851,N_23544,N_23399);
nor U23852 (N_23852,N_23376,N_23275);
or U23853 (N_23853,N_23139,N_23700);
and U23854 (N_23854,N_23609,N_23452);
and U23855 (N_23855,N_23586,N_23415);
nand U23856 (N_23856,N_23312,N_23607);
xor U23857 (N_23857,N_23322,N_23746);
nor U23858 (N_23858,N_23245,N_23209);
and U23859 (N_23859,N_23604,N_23683);
nor U23860 (N_23860,N_23575,N_23359);
and U23861 (N_23861,N_23416,N_23176);
or U23862 (N_23862,N_23310,N_23343);
xor U23863 (N_23863,N_23243,N_23461);
or U23864 (N_23864,N_23696,N_23213);
xor U23865 (N_23865,N_23419,N_23541);
and U23866 (N_23866,N_23463,N_23409);
and U23867 (N_23867,N_23355,N_23430);
nor U23868 (N_23868,N_23301,N_23319);
xor U23869 (N_23869,N_23169,N_23305);
and U23870 (N_23870,N_23520,N_23619);
or U23871 (N_23871,N_23550,N_23163);
and U23872 (N_23872,N_23368,N_23135);
or U23873 (N_23873,N_23515,N_23719);
nor U23874 (N_23874,N_23235,N_23381);
and U23875 (N_23875,N_23234,N_23605);
nor U23876 (N_23876,N_23655,N_23164);
nand U23877 (N_23877,N_23250,N_23331);
nand U23878 (N_23878,N_23392,N_23460);
xnor U23879 (N_23879,N_23671,N_23543);
nor U23880 (N_23880,N_23652,N_23327);
or U23881 (N_23881,N_23516,N_23583);
nand U23882 (N_23882,N_23491,N_23695);
nand U23883 (N_23883,N_23186,N_23721);
and U23884 (N_23884,N_23510,N_23507);
and U23885 (N_23885,N_23353,N_23595);
nand U23886 (N_23886,N_23618,N_23184);
xor U23887 (N_23887,N_23701,N_23720);
nor U23888 (N_23888,N_23303,N_23239);
xnor U23889 (N_23889,N_23669,N_23443);
nand U23890 (N_23890,N_23723,N_23434);
and U23891 (N_23891,N_23321,N_23504);
nor U23892 (N_23892,N_23320,N_23735);
nor U23893 (N_23893,N_23269,N_23179);
or U23894 (N_23894,N_23711,N_23194);
and U23895 (N_23895,N_23542,N_23662);
nand U23896 (N_23896,N_23427,N_23540);
or U23897 (N_23897,N_23724,N_23503);
nand U23898 (N_23898,N_23340,N_23266);
nor U23899 (N_23899,N_23180,N_23475);
nor U23900 (N_23900,N_23255,N_23576);
xnor U23901 (N_23901,N_23570,N_23494);
xor U23902 (N_23902,N_23692,N_23675);
and U23903 (N_23903,N_23441,N_23532);
nand U23904 (N_23904,N_23309,N_23557);
nor U23905 (N_23905,N_23436,N_23420);
or U23906 (N_23906,N_23193,N_23704);
xor U23907 (N_23907,N_23493,N_23699);
and U23908 (N_23908,N_23465,N_23232);
and U23909 (N_23909,N_23382,N_23572);
and U23910 (N_23910,N_23629,N_23130);
xnor U23911 (N_23911,N_23729,N_23222);
and U23912 (N_23912,N_23481,N_23358);
and U23913 (N_23913,N_23546,N_23306);
and U23914 (N_23914,N_23744,N_23265);
nand U23915 (N_23915,N_23374,N_23332);
nand U23916 (N_23916,N_23190,N_23438);
and U23917 (N_23917,N_23698,N_23435);
or U23918 (N_23918,N_23141,N_23685);
xor U23919 (N_23919,N_23166,N_23366);
and U23920 (N_23920,N_23348,N_23596);
or U23921 (N_23921,N_23589,N_23205);
and U23922 (N_23922,N_23525,N_23421);
or U23923 (N_23923,N_23588,N_23292);
nand U23924 (N_23924,N_23418,N_23717);
xnor U23925 (N_23925,N_23628,N_23138);
nand U23926 (N_23926,N_23201,N_23167);
xor U23927 (N_23927,N_23383,N_23512);
and U23928 (N_23928,N_23431,N_23248);
nor U23929 (N_23929,N_23508,N_23422);
nand U23930 (N_23930,N_23681,N_23749);
and U23931 (N_23931,N_23702,N_23496);
and U23932 (N_23932,N_23428,N_23483);
nand U23933 (N_23933,N_23293,N_23334);
xor U23934 (N_23934,N_23268,N_23614);
or U23935 (N_23935,N_23280,N_23432);
or U23936 (N_23936,N_23653,N_23674);
xnor U23937 (N_23937,N_23287,N_23707);
and U23938 (N_23938,N_23495,N_23549);
or U23939 (N_23939,N_23464,N_23247);
nand U23940 (N_23940,N_23488,N_23231);
xor U23941 (N_23941,N_23182,N_23689);
or U23942 (N_23942,N_23547,N_23710);
nand U23943 (N_23943,N_23172,N_23731);
xnor U23944 (N_23944,N_23555,N_23727);
and U23945 (N_23945,N_23726,N_23450);
and U23946 (N_23946,N_23425,N_23325);
or U23947 (N_23947,N_23296,N_23196);
or U23948 (N_23948,N_23388,N_23684);
and U23949 (N_23949,N_23564,N_23183);
nand U23950 (N_23950,N_23375,N_23559);
xnor U23951 (N_23951,N_23528,N_23241);
nand U23952 (N_23952,N_23526,N_23733);
nor U23953 (N_23953,N_23162,N_23686);
nand U23954 (N_23954,N_23599,N_23470);
xor U23955 (N_23955,N_23703,N_23661);
nand U23956 (N_23956,N_23127,N_23600);
nand U23957 (N_23957,N_23380,N_23519);
and U23958 (N_23958,N_23742,N_23456);
or U23959 (N_23959,N_23725,N_23151);
or U23960 (N_23960,N_23714,N_23297);
xnor U23961 (N_23961,N_23732,N_23501);
nor U23962 (N_23962,N_23597,N_23150);
nand U23963 (N_23963,N_23705,N_23370);
or U23964 (N_23964,N_23708,N_23574);
xor U23965 (N_23965,N_23214,N_23333);
or U23966 (N_23966,N_23125,N_23354);
and U23967 (N_23967,N_23608,N_23636);
and U23968 (N_23968,N_23486,N_23640);
xor U23969 (N_23969,N_23565,N_23511);
or U23970 (N_23970,N_23678,N_23660);
nor U23971 (N_23971,N_23233,N_23577);
nand U23972 (N_23972,N_23284,N_23667);
and U23973 (N_23973,N_23185,N_23371);
nand U23974 (N_23974,N_23455,N_23621);
or U23975 (N_23975,N_23208,N_23447);
nand U23976 (N_23976,N_23341,N_23747);
nand U23977 (N_23977,N_23230,N_23405);
xor U23978 (N_23978,N_23587,N_23342);
or U23979 (N_23979,N_23126,N_23478);
xnor U23980 (N_23980,N_23369,N_23560);
and U23981 (N_23981,N_23372,N_23346);
or U23982 (N_23982,N_23221,N_23288);
or U23983 (N_23983,N_23554,N_23490);
nand U23984 (N_23984,N_23168,N_23295);
xor U23985 (N_23985,N_23308,N_23545);
nand U23986 (N_23986,N_23433,N_23633);
and U23987 (N_23987,N_23377,N_23446);
and U23988 (N_23988,N_23274,N_23552);
nand U23989 (N_23989,N_23594,N_23451);
and U23990 (N_23990,N_23472,N_23133);
or U23991 (N_23991,N_23276,N_23521);
nand U23992 (N_23992,N_23517,N_23624);
and U23993 (N_23993,N_23538,N_23712);
nand U23994 (N_23994,N_23298,N_23672);
xnor U23995 (N_23995,N_23153,N_23479);
and U23996 (N_23996,N_23352,N_23174);
nand U23997 (N_23997,N_23500,N_23509);
xor U23998 (N_23998,N_23328,N_23713);
or U23999 (N_23999,N_23261,N_23229);
and U24000 (N_24000,N_23680,N_23379);
or U24001 (N_24001,N_23668,N_23513);
or U24002 (N_24002,N_23203,N_23351);
or U24003 (N_24003,N_23260,N_23738);
nor U24004 (N_24004,N_23191,N_23299);
xnor U24005 (N_24005,N_23663,N_23160);
nand U24006 (N_24006,N_23715,N_23294);
xnor U24007 (N_24007,N_23429,N_23363);
and U24008 (N_24008,N_23364,N_23228);
nor U24009 (N_24009,N_23237,N_23390);
xnor U24010 (N_24010,N_23638,N_23192);
xor U24011 (N_24011,N_23666,N_23444);
or U24012 (N_24012,N_23387,N_23336);
xor U24013 (N_24013,N_23134,N_23617);
and U24014 (N_24014,N_23329,N_23317);
and U24015 (N_24015,N_23740,N_23311);
or U24016 (N_24016,N_23236,N_23737);
nand U24017 (N_24017,N_23330,N_23670);
and U24018 (N_24018,N_23356,N_23743);
xor U24019 (N_24019,N_23206,N_23283);
xor U24020 (N_24020,N_23338,N_23693);
and U24021 (N_24021,N_23529,N_23523);
xnor U24022 (N_24022,N_23466,N_23257);
or U24023 (N_24023,N_23676,N_23218);
and U24024 (N_24024,N_23458,N_23187);
nor U24025 (N_24025,N_23142,N_23426);
nor U24026 (N_24026,N_23378,N_23220);
or U24027 (N_24027,N_23716,N_23610);
or U24028 (N_24028,N_23664,N_23401);
nor U24029 (N_24029,N_23437,N_23611);
xnor U24030 (N_24030,N_23410,N_23140);
or U24031 (N_24031,N_23177,N_23414);
nor U24032 (N_24032,N_23558,N_23423);
nand U24033 (N_24033,N_23403,N_23657);
and U24034 (N_24034,N_23467,N_23468);
nor U24035 (N_24035,N_23539,N_23630);
or U24036 (N_24036,N_23649,N_23398);
nor U24037 (N_24037,N_23226,N_23413);
and U24038 (N_24038,N_23453,N_23646);
nor U24039 (N_24039,N_23171,N_23402);
nor U24040 (N_24040,N_23568,N_23536);
xor U24041 (N_24041,N_23289,N_23373);
and U24042 (N_24042,N_23573,N_23602);
xnor U24043 (N_24043,N_23256,N_23548);
and U24044 (N_24044,N_23739,N_23178);
nand U24045 (N_24045,N_23357,N_23442);
nand U24046 (N_24046,N_23634,N_23601);
nor U24047 (N_24047,N_23145,N_23489);
nand U24048 (N_24048,N_23323,N_23158);
nand U24049 (N_24049,N_23581,N_23199);
and U24050 (N_24050,N_23181,N_23480);
nand U24051 (N_24051,N_23314,N_23365);
xor U24052 (N_24052,N_23391,N_23665);
or U24053 (N_24053,N_23344,N_23273);
and U24054 (N_24054,N_23249,N_23225);
nand U24055 (N_24055,N_23200,N_23616);
and U24056 (N_24056,N_23326,N_23212);
nor U24057 (N_24057,N_23677,N_23286);
nor U24058 (N_24058,N_23270,N_23706);
nand U24059 (N_24059,N_23506,N_23264);
nand U24060 (N_24060,N_23566,N_23360);
nor U24061 (N_24061,N_23254,N_23404);
nor U24062 (N_24062,N_23219,N_23528);
xnor U24063 (N_24063,N_23679,N_23289);
or U24064 (N_24064,N_23726,N_23348);
nor U24065 (N_24065,N_23280,N_23381);
and U24066 (N_24066,N_23711,N_23286);
and U24067 (N_24067,N_23684,N_23227);
or U24068 (N_24068,N_23254,N_23216);
nand U24069 (N_24069,N_23275,N_23324);
nor U24070 (N_24070,N_23492,N_23730);
xnor U24071 (N_24071,N_23495,N_23228);
xor U24072 (N_24072,N_23259,N_23462);
nor U24073 (N_24073,N_23694,N_23644);
or U24074 (N_24074,N_23702,N_23523);
or U24075 (N_24075,N_23454,N_23396);
and U24076 (N_24076,N_23512,N_23158);
and U24077 (N_24077,N_23150,N_23585);
and U24078 (N_24078,N_23402,N_23391);
or U24079 (N_24079,N_23743,N_23563);
nand U24080 (N_24080,N_23166,N_23245);
and U24081 (N_24081,N_23702,N_23274);
nor U24082 (N_24082,N_23466,N_23182);
nor U24083 (N_24083,N_23644,N_23718);
and U24084 (N_24084,N_23193,N_23672);
and U24085 (N_24085,N_23399,N_23536);
or U24086 (N_24086,N_23197,N_23691);
and U24087 (N_24087,N_23553,N_23162);
xnor U24088 (N_24088,N_23253,N_23535);
nand U24089 (N_24089,N_23140,N_23695);
nand U24090 (N_24090,N_23462,N_23697);
and U24091 (N_24091,N_23550,N_23426);
or U24092 (N_24092,N_23317,N_23272);
xnor U24093 (N_24093,N_23260,N_23254);
xnor U24094 (N_24094,N_23659,N_23712);
nand U24095 (N_24095,N_23546,N_23347);
nor U24096 (N_24096,N_23589,N_23361);
xor U24097 (N_24097,N_23280,N_23166);
or U24098 (N_24098,N_23275,N_23175);
or U24099 (N_24099,N_23681,N_23741);
and U24100 (N_24100,N_23529,N_23424);
nand U24101 (N_24101,N_23377,N_23209);
nand U24102 (N_24102,N_23193,N_23694);
xnor U24103 (N_24103,N_23724,N_23193);
and U24104 (N_24104,N_23264,N_23168);
nand U24105 (N_24105,N_23240,N_23538);
or U24106 (N_24106,N_23651,N_23525);
and U24107 (N_24107,N_23615,N_23486);
nand U24108 (N_24108,N_23224,N_23388);
or U24109 (N_24109,N_23126,N_23414);
xor U24110 (N_24110,N_23268,N_23447);
xor U24111 (N_24111,N_23586,N_23134);
nor U24112 (N_24112,N_23310,N_23644);
nor U24113 (N_24113,N_23690,N_23592);
nand U24114 (N_24114,N_23550,N_23158);
nor U24115 (N_24115,N_23356,N_23692);
xor U24116 (N_24116,N_23132,N_23290);
xor U24117 (N_24117,N_23348,N_23547);
nand U24118 (N_24118,N_23745,N_23658);
nor U24119 (N_24119,N_23667,N_23296);
nor U24120 (N_24120,N_23178,N_23644);
nand U24121 (N_24121,N_23177,N_23666);
nor U24122 (N_24122,N_23582,N_23334);
and U24123 (N_24123,N_23713,N_23264);
nor U24124 (N_24124,N_23163,N_23742);
xor U24125 (N_24125,N_23318,N_23688);
and U24126 (N_24126,N_23137,N_23541);
nand U24127 (N_24127,N_23548,N_23314);
xnor U24128 (N_24128,N_23134,N_23251);
xor U24129 (N_24129,N_23548,N_23674);
or U24130 (N_24130,N_23173,N_23224);
nand U24131 (N_24131,N_23231,N_23277);
nand U24132 (N_24132,N_23341,N_23566);
and U24133 (N_24133,N_23476,N_23422);
nor U24134 (N_24134,N_23746,N_23516);
or U24135 (N_24135,N_23708,N_23566);
and U24136 (N_24136,N_23698,N_23504);
and U24137 (N_24137,N_23455,N_23250);
nand U24138 (N_24138,N_23389,N_23622);
or U24139 (N_24139,N_23553,N_23696);
or U24140 (N_24140,N_23485,N_23651);
and U24141 (N_24141,N_23300,N_23656);
xor U24142 (N_24142,N_23306,N_23143);
nor U24143 (N_24143,N_23710,N_23499);
xor U24144 (N_24144,N_23417,N_23184);
or U24145 (N_24145,N_23507,N_23139);
or U24146 (N_24146,N_23217,N_23626);
and U24147 (N_24147,N_23283,N_23702);
and U24148 (N_24148,N_23551,N_23576);
nor U24149 (N_24149,N_23356,N_23305);
or U24150 (N_24150,N_23404,N_23151);
or U24151 (N_24151,N_23320,N_23633);
xor U24152 (N_24152,N_23453,N_23246);
or U24153 (N_24153,N_23403,N_23678);
xnor U24154 (N_24154,N_23710,N_23684);
nor U24155 (N_24155,N_23395,N_23744);
and U24156 (N_24156,N_23258,N_23718);
and U24157 (N_24157,N_23280,N_23335);
nor U24158 (N_24158,N_23521,N_23625);
and U24159 (N_24159,N_23503,N_23193);
xor U24160 (N_24160,N_23372,N_23295);
and U24161 (N_24161,N_23705,N_23179);
and U24162 (N_24162,N_23187,N_23483);
or U24163 (N_24163,N_23320,N_23133);
nand U24164 (N_24164,N_23494,N_23530);
nand U24165 (N_24165,N_23246,N_23489);
or U24166 (N_24166,N_23190,N_23166);
xnor U24167 (N_24167,N_23612,N_23422);
nor U24168 (N_24168,N_23525,N_23142);
and U24169 (N_24169,N_23238,N_23471);
nand U24170 (N_24170,N_23641,N_23338);
or U24171 (N_24171,N_23162,N_23470);
nor U24172 (N_24172,N_23214,N_23223);
nor U24173 (N_24173,N_23159,N_23304);
and U24174 (N_24174,N_23516,N_23567);
or U24175 (N_24175,N_23291,N_23531);
and U24176 (N_24176,N_23184,N_23197);
and U24177 (N_24177,N_23722,N_23549);
or U24178 (N_24178,N_23680,N_23160);
nor U24179 (N_24179,N_23544,N_23638);
nand U24180 (N_24180,N_23232,N_23536);
nand U24181 (N_24181,N_23125,N_23234);
and U24182 (N_24182,N_23722,N_23418);
nor U24183 (N_24183,N_23676,N_23240);
and U24184 (N_24184,N_23412,N_23325);
and U24185 (N_24185,N_23596,N_23178);
or U24186 (N_24186,N_23405,N_23495);
or U24187 (N_24187,N_23741,N_23278);
xor U24188 (N_24188,N_23256,N_23713);
or U24189 (N_24189,N_23633,N_23515);
xnor U24190 (N_24190,N_23314,N_23374);
nor U24191 (N_24191,N_23746,N_23728);
or U24192 (N_24192,N_23156,N_23556);
or U24193 (N_24193,N_23549,N_23227);
nand U24194 (N_24194,N_23455,N_23361);
or U24195 (N_24195,N_23163,N_23200);
and U24196 (N_24196,N_23569,N_23468);
and U24197 (N_24197,N_23700,N_23150);
nand U24198 (N_24198,N_23164,N_23694);
xor U24199 (N_24199,N_23492,N_23362);
xnor U24200 (N_24200,N_23432,N_23417);
and U24201 (N_24201,N_23440,N_23441);
and U24202 (N_24202,N_23336,N_23127);
and U24203 (N_24203,N_23395,N_23399);
xor U24204 (N_24204,N_23497,N_23588);
nand U24205 (N_24205,N_23231,N_23563);
nand U24206 (N_24206,N_23517,N_23704);
and U24207 (N_24207,N_23268,N_23365);
xor U24208 (N_24208,N_23732,N_23430);
or U24209 (N_24209,N_23324,N_23280);
nand U24210 (N_24210,N_23739,N_23528);
or U24211 (N_24211,N_23455,N_23326);
xnor U24212 (N_24212,N_23645,N_23148);
nor U24213 (N_24213,N_23346,N_23580);
nand U24214 (N_24214,N_23132,N_23365);
nand U24215 (N_24215,N_23552,N_23403);
xnor U24216 (N_24216,N_23497,N_23635);
or U24217 (N_24217,N_23645,N_23394);
xnor U24218 (N_24218,N_23646,N_23696);
nand U24219 (N_24219,N_23511,N_23446);
or U24220 (N_24220,N_23442,N_23345);
nor U24221 (N_24221,N_23179,N_23407);
nor U24222 (N_24222,N_23165,N_23587);
and U24223 (N_24223,N_23352,N_23461);
or U24224 (N_24224,N_23262,N_23681);
and U24225 (N_24225,N_23448,N_23545);
nor U24226 (N_24226,N_23528,N_23625);
and U24227 (N_24227,N_23352,N_23316);
xor U24228 (N_24228,N_23355,N_23139);
nor U24229 (N_24229,N_23539,N_23182);
and U24230 (N_24230,N_23218,N_23512);
or U24231 (N_24231,N_23381,N_23454);
or U24232 (N_24232,N_23194,N_23348);
xor U24233 (N_24233,N_23217,N_23711);
nand U24234 (N_24234,N_23459,N_23576);
nor U24235 (N_24235,N_23646,N_23269);
xor U24236 (N_24236,N_23498,N_23434);
nand U24237 (N_24237,N_23567,N_23394);
or U24238 (N_24238,N_23497,N_23485);
nor U24239 (N_24239,N_23181,N_23725);
and U24240 (N_24240,N_23197,N_23738);
and U24241 (N_24241,N_23744,N_23334);
and U24242 (N_24242,N_23212,N_23126);
xor U24243 (N_24243,N_23601,N_23391);
nand U24244 (N_24244,N_23432,N_23689);
xnor U24245 (N_24245,N_23199,N_23436);
or U24246 (N_24246,N_23187,N_23257);
or U24247 (N_24247,N_23441,N_23529);
or U24248 (N_24248,N_23227,N_23726);
and U24249 (N_24249,N_23701,N_23703);
or U24250 (N_24250,N_23132,N_23246);
xnor U24251 (N_24251,N_23225,N_23154);
nand U24252 (N_24252,N_23358,N_23625);
and U24253 (N_24253,N_23227,N_23355);
nor U24254 (N_24254,N_23213,N_23384);
nor U24255 (N_24255,N_23285,N_23621);
nor U24256 (N_24256,N_23233,N_23333);
or U24257 (N_24257,N_23308,N_23718);
nand U24258 (N_24258,N_23729,N_23208);
nor U24259 (N_24259,N_23611,N_23262);
nor U24260 (N_24260,N_23356,N_23721);
and U24261 (N_24261,N_23743,N_23613);
and U24262 (N_24262,N_23625,N_23320);
and U24263 (N_24263,N_23427,N_23383);
nand U24264 (N_24264,N_23344,N_23401);
xor U24265 (N_24265,N_23371,N_23675);
nand U24266 (N_24266,N_23404,N_23672);
nor U24267 (N_24267,N_23482,N_23449);
xor U24268 (N_24268,N_23380,N_23500);
xnor U24269 (N_24269,N_23495,N_23474);
xor U24270 (N_24270,N_23550,N_23683);
nor U24271 (N_24271,N_23607,N_23661);
nand U24272 (N_24272,N_23389,N_23270);
or U24273 (N_24273,N_23376,N_23443);
xor U24274 (N_24274,N_23269,N_23285);
nor U24275 (N_24275,N_23141,N_23313);
and U24276 (N_24276,N_23502,N_23693);
and U24277 (N_24277,N_23211,N_23616);
nand U24278 (N_24278,N_23272,N_23389);
nor U24279 (N_24279,N_23135,N_23587);
or U24280 (N_24280,N_23569,N_23217);
nand U24281 (N_24281,N_23687,N_23204);
xor U24282 (N_24282,N_23241,N_23229);
xor U24283 (N_24283,N_23375,N_23609);
and U24284 (N_24284,N_23387,N_23322);
nand U24285 (N_24285,N_23187,N_23601);
or U24286 (N_24286,N_23138,N_23682);
and U24287 (N_24287,N_23561,N_23485);
and U24288 (N_24288,N_23226,N_23175);
nand U24289 (N_24289,N_23556,N_23199);
and U24290 (N_24290,N_23403,N_23599);
and U24291 (N_24291,N_23491,N_23559);
nor U24292 (N_24292,N_23244,N_23432);
nand U24293 (N_24293,N_23477,N_23276);
and U24294 (N_24294,N_23714,N_23716);
xor U24295 (N_24295,N_23226,N_23336);
nand U24296 (N_24296,N_23698,N_23439);
xnor U24297 (N_24297,N_23273,N_23491);
xnor U24298 (N_24298,N_23146,N_23304);
nand U24299 (N_24299,N_23205,N_23529);
nand U24300 (N_24300,N_23316,N_23428);
xor U24301 (N_24301,N_23634,N_23713);
or U24302 (N_24302,N_23741,N_23472);
or U24303 (N_24303,N_23473,N_23248);
and U24304 (N_24304,N_23746,N_23320);
or U24305 (N_24305,N_23587,N_23304);
xor U24306 (N_24306,N_23688,N_23523);
nor U24307 (N_24307,N_23358,N_23258);
and U24308 (N_24308,N_23231,N_23244);
xor U24309 (N_24309,N_23575,N_23365);
xnor U24310 (N_24310,N_23731,N_23447);
xor U24311 (N_24311,N_23345,N_23425);
or U24312 (N_24312,N_23243,N_23232);
nor U24313 (N_24313,N_23748,N_23696);
nor U24314 (N_24314,N_23712,N_23275);
nor U24315 (N_24315,N_23227,N_23461);
or U24316 (N_24316,N_23357,N_23163);
nand U24317 (N_24317,N_23581,N_23196);
nor U24318 (N_24318,N_23676,N_23454);
and U24319 (N_24319,N_23556,N_23609);
nor U24320 (N_24320,N_23131,N_23302);
nand U24321 (N_24321,N_23348,N_23233);
and U24322 (N_24322,N_23625,N_23382);
and U24323 (N_24323,N_23549,N_23174);
nand U24324 (N_24324,N_23326,N_23595);
nand U24325 (N_24325,N_23576,N_23614);
or U24326 (N_24326,N_23653,N_23702);
nand U24327 (N_24327,N_23619,N_23587);
or U24328 (N_24328,N_23195,N_23128);
xnor U24329 (N_24329,N_23196,N_23317);
nor U24330 (N_24330,N_23143,N_23694);
xor U24331 (N_24331,N_23268,N_23455);
nor U24332 (N_24332,N_23661,N_23499);
nor U24333 (N_24333,N_23145,N_23441);
nand U24334 (N_24334,N_23479,N_23430);
or U24335 (N_24335,N_23397,N_23506);
and U24336 (N_24336,N_23219,N_23673);
xor U24337 (N_24337,N_23210,N_23339);
nand U24338 (N_24338,N_23136,N_23241);
nand U24339 (N_24339,N_23478,N_23128);
xnor U24340 (N_24340,N_23545,N_23575);
or U24341 (N_24341,N_23292,N_23126);
nand U24342 (N_24342,N_23433,N_23652);
and U24343 (N_24343,N_23176,N_23525);
or U24344 (N_24344,N_23333,N_23511);
xor U24345 (N_24345,N_23582,N_23554);
and U24346 (N_24346,N_23385,N_23382);
xnor U24347 (N_24347,N_23223,N_23369);
xor U24348 (N_24348,N_23747,N_23557);
nand U24349 (N_24349,N_23396,N_23570);
nor U24350 (N_24350,N_23180,N_23343);
nand U24351 (N_24351,N_23693,N_23283);
nand U24352 (N_24352,N_23203,N_23481);
nor U24353 (N_24353,N_23128,N_23730);
xor U24354 (N_24354,N_23156,N_23254);
nand U24355 (N_24355,N_23462,N_23140);
nor U24356 (N_24356,N_23680,N_23499);
or U24357 (N_24357,N_23385,N_23572);
xnor U24358 (N_24358,N_23484,N_23635);
and U24359 (N_24359,N_23505,N_23363);
nand U24360 (N_24360,N_23249,N_23619);
and U24361 (N_24361,N_23394,N_23173);
xor U24362 (N_24362,N_23362,N_23524);
nor U24363 (N_24363,N_23722,N_23322);
or U24364 (N_24364,N_23387,N_23657);
and U24365 (N_24365,N_23438,N_23145);
nor U24366 (N_24366,N_23524,N_23363);
nor U24367 (N_24367,N_23575,N_23578);
or U24368 (N_24368,N_23197,N_23524);
and U24369 (N_24369,N_23742,N_23408);
or U24370 (N_24370,N_23163,N_23737);
and U24371 (N_24371,N_23438,N_23526);
nand U24372 (N_24372,N_23677,N_23410);
nand U24373 (N_24373,N_23461,N_23262);
nor U24374 (N_24374,N_23315,N_23422);
and U24375 (N_24375,N_24280,N_23973);
nor U24376 (N_24376,N_23818,N_24204);
xnor U24377 (N_24377,N_24327,N_23951);
xnor U24378 (N_24378,N_24372,N_24335);
nand U24379 (N_24379,N_24306,N_24126);
and U24380 (N_24380,N_24309,N_24239);
or U24381 (N_24381,N_23942,N_23809);
xor U24382 (N_24382,N_24277,N_24143);
and U24383 (N_24383,N_24300,N_24153);
xor U24384 (N_24384,N_24190,N_23947);
nand U24385 (N_24385,N_23926,N_24073);
xnor U24386 (N_24386,N_24332,N_24171);
nor U24387 (N_24387,N_24361,N_24047);
and U24388 (N_24388,N_23823,N_24340);
nand U24389 (N_24389,N_24178,N_24363);
xnor U24390 (N_24390,N_24181,N_23800);
and U24391 (N_24391,N_24356,N_23970);
nand U24392 (N_24392,N_23849,N_24247);
nand U24393 (N_24393,N_23794,N_24129);
nand U24394 (N_24394,N_24368,N_23874);
or U24395 (N_24395,N_24021,N_23835);
nor U24396 (N_24396,N_24227,N_24032);
xnor U24397 (N_24397,N_24015,N_24290);
xnor U24398 (N_24398,N_24148,N_24042);
and U24399 (N_24399,N_24080,N_23937);
nor U24400 (N_24400,N_23959,N_24139);
nor U24401 (N_24401,N_24326,N_23995);
or U24402 (N_24402,N_24268,N_24233);
nand U24403 (N_24403,N_23953,N_24331);
xor U24404 (N_24404,N_23936,N_24196);
xnor U24405 (N_24405,N_24296,N_24088);
nand U24406 (N_24406,N_23838,N_23994);
nor U24407 (N_24407,N_23762,N_24229);
xnor U24408 (N_24408,N_23887,N_24096);
and U24409 (N_24409,N_24157,N_23998);
or U24410 (N_24410,N_23979,N_23894);
and U24411 (N_24411,N_24018,N_23969);
nor U24412 (N_24412,N_23948,N_23939);
nor U24413 (N_24413,N_24367,N_24225);
nor U24414 (N_24414,N_23836,N_24098);
and U24415 (N_24415,N_24184,N_24298);
and U24416 (N_24416,N_23899,N_23949);
or U24417 (N_24417,N_23802,N_23805);
xnor U24418 (N_24418,N_24220,N_23917);
and U24419 (N_24419,N_24149,N_23993);
nand U24420 (N_24420,N_23812,N_23879);
xnor U24421 (N_24421,N_24329,N_24369);
xnor U24422 (N_24422,N_23754,N_23892);
xnor U24423 (N_24423,N_23943,N_24138);
nand U24424 (N_24424,N_23893,N_23932);
nor U24425 (N_24425,N_24286,N_24173);
or U24426 (N_24426,N_23964,N_24275);
nor U24427 (N_24427,N_23867,N_24037);
or U24428 (N_24428,N_24234,N_24059);
and U24429 (N_24429,N_23840,N_24094);
and U24430 (N_24430,N_23858,N_23767);
nor U24431 (N_24431,N_23961,N_23880);
or U24432 (N_24432,N_24311,N_24231);
xnor U24433 (N_24433,N_24034,N_24095);
nor U24434 (N_24434,N_24048,N_24353);
xor U24435 (N_24435,N_24272,N_24045);
nand U24436 (N_24436,N_24036,N_24270);
or U24437 (N_24437,N_23864,N_23989);
nand U24438 (N_24438,N_23793,N_24030);
or U24439 (N_24439,N_23848,N_23967);
nand U24440 (N_24440,N_24226,N_24349);
and U24441 (N_24441,N_24359,N_24102);
or U24442 (N_24442,N_23869,N_24221);
nand U24443 (N_24443,N_24373,N_24144);
and U24444 (N_24444,N_24135,N_23915);
nand U24445 (N_24445,N_24086,N_24141);
or U24446 (N_24446,N_24186,N_23859);
xor U24447 (N_24447,N_24057,N_23900);
or U24448 (N_24448,N_24371,N_24164);
nor U24449 (N_24449,N_23830,N_24206);
xnor U24450 (N_24450,N_24198,N_23775);
or U24451 (N_24451,N_23790,N_24180);
nor U24452 (N_24452,N_24110,N_23924);
or U24453 (N_24453,N_24000,N_24299);
nor U24454 (N_24454,N_23952,N_24028);
nand U24455 (N_24455,N_24039,N_24238);
or U24456 (N_24456,N_24266,N_24117);
nand U24457 (N_24457,N_24063,N_24177);
and U24458 (N_24458,N_23907,N_24162);
nand U24459 (N_24459,N_23984,N_24109);
nand U24460 (N_24460,N_24195,N_24172);
nand U24461 (N_24461,N_23860,N_24161);
nand U24462 (N_24462,N_23895,N_24145);
and U24463 (N_24463,N_23996,N_23934);
nand U24464 (N_24464,N_23914,N_23824);
and U24465 (N_24465,N_24274,N_24257);
xnor U24466 (N_24466,N_23911,N_24338);
and U24467 (N_24467,N_23884,N_24054);
nor U24468 (N_24468,N_24342,N_24154);
nor U24469 (N_24469,N_24362,N_23971);
and U24470 (N_24470,N_24011,N_24201);
or U24471 (N_24471,N_24093,N_23769);
xnor U24472 (N_24472,N_24041,N_23891);
and U24473 (N_24473,N_24320,N_24151);
nor U24474 (N_24474,N_24033,N_24228);
nand U24475 (N_24475,N_23902,N_24288);
and U24476 (N_24476,N_24169,N_24189);
nand U24477 (N_24477,N_23904,N_24293);
nand U24478 (N_24478,N_24118,N_23751);
xnor U24479 (N_24479,N_24366,N_24273);
xor U24480 (N_24480,N_23842,N_23828);
or U24481 (N_24481,N_24344,N_23787);
nand U24482 (N_24482,N_24014,N_24315);
xor U24483 (N_24483,N_24205,N_24026);
or U24484 (N_24484,N_24152,N_24324);
or U24485 (N_24485,N_24097,N_24200);
nor U24486 (N_24486,N_23963,N_24016);
xnor U24487 (N_24487,N_24020,N_24217);
nor U24488 (N_24488,N_24009,N_24082);
or U24489 (N_24489,N_23811,N_24174);
and U24490 (N_24490,N_24251,N_24255);
nor U24491 (N_24491,N_24343,N_24328);
xor U24492 (N_24492,N_24165,N_23856);
or U24493 (N_24493,N_24051,N_24113);
xnor U24494 (N_24494,N_23863,N_23763);
nand U24495 (N_24495,N_24022,N_23789);
xnor U24496 (N_24496,N_24208,N_24269);
or U24497 (N_24497,N_23757,N_24112);
nor U24498 (N_24498,N_24240,N_23983);
xor U24499 (N_24499,N_24121,N_24218);
or U24500 (N_24500,N_24219,N_24285);
nor U24501 (N_24501,N_24313,N_24199);
and U24502 (N_24502,N_24179,N_23846);
or U24503 (N_24503,N_23791,N_23821);
or U24504 (N_24504,N_24297,N_23777);
nand U24505 (N_24505,N_23765,N_24235);
nor U24506 (N_24506,N_24302,N_24318);
nand U24507 (N_24507,N_24262,N_23922);
nor U24508 (N_24508,N_24339,N_23779);
and U24509 (N_24509,N_24325,N_24008);
nor U24510 (N_24510,N_23819,N_24007);
xor U24511 (N_24511,N_23861,N_24115);
nand U24512 (N_24512,N_24207,N_23945);
xor U24513 (N_24513,N_24136,N_24078);
or U24514 (N_24514,N_23816,N_24346);
nand U24515 (N_24515,N_23966,N_24002);
and U24516 (N_24516,N_23978,N_23999);
nand U24517 (N_24517,N_24004,N_24081);
and U24518 (N_24518,N_24100,N_24237);
or U24519 (N_24519,N_24191,N_24128);
xnor U24520 (N_24520,N_23933,N_24337);
and U24521 (N_24521,N_24071,N_24243);
nand U24522 (N_24522,N_23834,N_24261);
or U24523 (N_24523,N_23847,N_24083);
nor U24524 (N_24524,N_24156,N_23972);
nand U24525 (N_24525,N_23938,N_23956);
nand U24526 (N_24526,N_23962,N_24216);
or U24527 (N_24527,N_23782,N_24307);
and U24528 (N_24528,N_24055,N_24314);
and U24529 (N_24529,N_24246,N_24347);
nor U24530 (N_24530,N_24127,N_24074);
nand U24531 (N_24531,N_24305,N_23981);
or U24532 (N_24532,N_24035,N_24140);
nand U24533 (N_24533,N_24374,N_24292);
nand U24534 (N_24534,N_24213,N_24276);
nor U24535 (N_24535,N_24222,N_23946);
or U24536 (N_24536,N_24301,N_24012);
and U24537 (N_24537,N_23844,N_23991);
nand U24538 (N_24538,N_24355,N_24170);
nor U24539 (N_24539,N_23882,N_23795);
nor U24540 (N_24540,N_23813,N_23905);
and U24541 (N_24541,N_23797,N_23968);
xor U24542 (N_24542,N_24230,N_24304);
nand U24543 (N_24543,N_24303,N_23808);
nand U24544 (N_24544,N_23822,N_24250);
or U24545 (N_24545,N_24267,N_23903);
and U24546 (N_24546,N_23921,N_24215);
xor U24547 (N_24547,N_24253,N_24038);
xnor U24548 (N_24548,N_23997,N_24209);
xnor U24549 (N_24549,N_23778,N_24289);
nand U24550 (N_24550,N_24049,N_24260);
xnor U24551 (N_24551,N_24350,N_24079);
and U24552 (N_24552,N_23771,N_24124);
and U24553 (N_24553,N_24120,N_24029);
nand U24554 (N_24554,N_23871,N_24271);
xnor U24555 (N_24555,N_23875,N_23940);
nor U24556 (N_24556,N_24244,N_24291);
and U24557 (N_24557,N_23885,N_24053);
or U24558 (N_24558,N_24077,N_24319);
nor U24559 (N_24559,N_23753,N_24168);
nand U24560 (N_24560,N_23803,N_23928);
nor U24561 (N_24561,N_23992,N_24197);
and U24562 (N_24562,N_24076,N_23785);
or U24563 (N_24563,N_24187,N_24060);
or U24564 (N_24564,N_23944,N_23873);
and U24565 (N_24565,N_24264,N_23855);
and U24566 (N_24566,N_24099,N_24122);
xor U24567 (N_24567,N_23886,N_24236);
or U24568 (N_24568,N_24142,N_23941);
or U24569 (N_24569,N_23825,N_24123);
and U24570 (N_24570,N_23768,N_23990);
or U24571 (N_24571,N_24160,N_24104);
nor U24572 (N_24572,N_24175,N_24336);
and U24573 (N_24573,N_24248,N_24323);
xnor U24574 (N_24574,N_24075,N_24017);
xnor U24575 (N_24575,N_24125,N_24058);
and U24576 (N_24576,N_24134,N_23857);
or U24577 (N_24577,N_23906,N_23845);
or U24578 (N_24578,N_23985,N_24210);
or U24579 (N_24579,N_24070,N_23833);
nand U24580 (N_24580,N_23852,N_24006);
nor U24581 (N_24581,N_24067,N_23872);
and U24582 (N_24582,N_24295,N_24040);
and U24583 (N_24583,N_24345,N_24294);
and U24584 (N_24584,N_24322,N_24259);
nand U24585 (N_24585,N_23896,N_23841);
or U24586 (N_24586,N_24066,N_24223);
nor U24587 (N_24587,N_23986,N_23756);
xnor U24588 (N_24588,N_24043,N_23866);
nor U24589 (N_24589,N_24072,N_24321);
nand U24590 (N_24590,N_23807,N_23832);
or U24591 (N_24591,N_23919,N_23774);
nand U24592 (N_24592,N_23881,N_23930);
and U24593 (N_24593,N_23815,N_23876);
or U24594 (N_24594,N_23854,N_24085);
or U24595 (N_24595,N_23764,N_24069);
or U24596 (N_24596,N_24050,N_23798);
xnor U24597 (N_24597,N_24116,N_23801);
nand U24598 (N_24598,N_24281,N_24013);
and U24599 (N_24599,N_24283,N_23976);
or U24600 (N_24600,N_24245,N_23890);
nor U24601 (N_24601,N_23780,N_23988);
or U24602 (N_24602,N_23752,N_23960);
nor U24603 (N_24603,N_23806,N_24108);
xnor U24604 (N_24604,N_24370,N_24119);
nand U24605 (N_24605,N_23839,N_23931);
nand U24606 (N_24606,N_23916,N_24258);
nand U24607 (N_24607,N_24224,N_24146);
xor U24608 (N_24608,N_24334,N_23792);
xnor U24609 (N_24609,N_24263,N_23755);
or U24610 (N_24610,N_23776,N_23810);
or U24611 (N_24611,N_23814,N_23831);
nand U24612 (N_24612,N_24284,N_24131);
xnor U24613 (N_24613,N_24155,N_24027);
and U24614 (N_24614,N_24333,N_24052);
nor U24615 (N_24615,N_24001,N_23850);
nor U24616 (N_24616,N_24357,N_24194);
or U24617 (N_24617,N_24166,N_23759);
xnor U24618 (N_24618,N_23950,N_24106);
and U24619 (N_24619,N_24025,N_24341);
or U24620 (N_24620,N_24358,N_24330);
nand U24621 (N_24621,N_23918,N_24316);
xnor U24622 (N_24622,N_23868,N_23909);
and U24623 (N_24623,N_24354,N_24202);
or U24624 (N_24624,N_23804,N_24265);
or U24625 (N_24625,N_23851,N_23910);
nor U24626 (N_24626,N_24130,N_23758);
xnor U24627 (N_24627,N_24061,N_24241);
nor U24628 (N_24628,N_24312,N_23974);
nor U24629 (N_24629,N_24150,N_23954);
and U24630 (N_24630,N_23799,N_23929);
nor U24631 (N_24631,N_24163,N_24090);
nand U24632 (N_24632,N_24091,N_23829);
and U24633 (N_24633,N_23772,N_24065);
xor U24634 (N_24634,N_24352,N_23957);
nor U24635 (N_24635,N_24056,N_24046);
nand U24636 (N_24636,N_23862,N_23980);
and U24637 (N_24637,N_23853,N_23766);
nor U24638 (N_24638,N_24254,N_23977);
or U24639 (N_24639,N_23788,N_23913);
xnor U24640 (N_24640,N_23897,N_24214);
and U24641 (N_24641,N_24192,N_24137);
and U24642 (N_24642,N_23870,N_23901);
nor U24643 (N_24643,N_24010,N_23958);
nor U24644 (N_24644,N_24203,N_24182);
xnor U24645 (N_24645,N_23927,N_23965);
xor U24646 (N_24646,N_23784,N_23843);
xnor U24647 (N_24647,N_23923,N_23796);
nand U24648 (N_24648,N_23889,N_24183);
or U24649 (N_24649,N_23955,N_24064);
nor U24650 (N_24650,N_24044,N_24232);
and U24651 (N_24651,N_23817,N_24212);
nand U24652 (N_24652,N_24211,N_24351);
and U24653 (N_24653,N_24114,N_24132);
nand U24654 (N_24654,N_24279,N_23925);
xnor U24655 (N_24655,N_23987,N_24133);
nand U24656 (N_24656,N_24252,N_23898);
or U24657 (N_24657,N_24031,N_24103);
nor U24658 (N_24658,N_23878,N_24176);
xor U24659 (N_24659,N_24003,N_24278);
and U24660 (N_24660,N_23877,N_23783);
nand U24661 (N_24661,N_24005,N_24348);
nor U24662 (N_24662,N_24101,N_23761);
and U24663 (N_24663,N_24193,N_24249);
and U24664 (N_24664,N_24062,N_24107);
xor U24665 (N_24665,N_24147,N_23920);
and U24666 (N_24666,N_23935,N_23912);
and U24667 (N_24667,N_23908,N_24084);
nor U24668 (N_24668,N_23837,N_24317);
xnor U24669 (N_24669,N_24167,N_23826);
and U24670 (N_24670,N_24364,N_24256);
or U24671 (N_24671,N_24360,N_24242);
nand U24672 (N_24672,N_23982,N_24282);
or U24673 (N_24673,N_23773,N_24023);
and U24674 (N_24674,N_24185,N_23820);
and U24675 (N_24675,N_23975,N_24111);
nand U24676 (N_24676,N_23781,N_24188);
xnor U24677 (N_24677,N_24365,N_23888);
nand U24678 (N_24678,N_24089,N_23760);
xnor U24679 (N_24679,N_23770,N_24019);
nand U24680 (N_24680,N_24308,N_24310);
nand U24681 (N_24681,N_24287,N_23827);
nor U24682 (N_24682,N_24024,N_24092);
xnor U24683 (N_24683,N_23750,N_24105);
nor U24684 (N_24684,N_23865,N_23883);
or U24685 (N_24685,N_24158,N_23786);
nor U24686 (N_24686,N_24159,N_24087);
nand U24687 (N_24687,N_24068,N_23770);
and U24688 (N_24688,N_24115,N_24052);
nand U24689 (N_24689,N_23798,N_24077);
or U24690 (N_24690,N_24240,N_24258);
nor U24691 (N_24691,N_24206,N_23829);
or U24692 (N_24692,N_24286,N_24207);
xor U24693 (N_24693,N_24001,N_24302);
xor U24694 (N_24694,N_23752,N_24002);
nand U24695 (N_24695,N_23935,N_24308);
nor U24696 (N_24696,N_23869,N_24347);
and U24697 (N_24697,N_24227,N_24010);
or U24698 (N_24698,N_24156,N_24231);
or U24699 (N_24699,N_23799,N_23790);
nand U24700 (N_24700,N_24039,N_24159);
nor U24701 (N_24701,N_23761,N_24052);
or U24702 (N_24702,N_24118,N_23974);
nor U24703 (N_24703,N_24098,N_24284);
nand U24704 (N_24704,N_23868,N_24267);
and U24705 (N_24705,N_24150,N_24135);
or U24706 (N_24706,N_24225,N_23945);
or U24707 (N_24707,N_23780,N_23965);
xor U24708 (N_24708,N_24334,N_24369);
xnor U24709 (N_24709,N_23849,N_24164);
or U24710 (N_24710,N_24326,N_23813);
and U24711 (N_24711,N_24018,N_23945);
nor U24712 (N_24712,N_24288,N_23864);
nor U24713 (N_24713,N_24190,N_24334);
and U24714 (N_24714,N_24210,N_23867);
xnor U24715 (N_24715,N_23978,N_24142);
or U24716 (N_24716,N_23967,N_24334);
nand U24717 (N_24717,N_24198,N_24204);
nand U24718 (N_24718,N_24009,N_23835);
xnor U24719 (N_24719,N_23962,N_23846);
and U24720 (N_24720,N_24325,N_24052);
nand U24721 (N_24721,N_23888,N_23966);
nor U24722 (N_24722,N_24308,N_24094);
nand U24723 (N_24723,N_24320,N_23839);
nand U24724 (N_24724,N_24182,N_23897);
nand U24725 (N_24725,N_23785,N_23885);
and U24726 (N_24726,N_24146,N_24093);
or U24727 (N_24727,N_23924,N_23796);
or U24728 (N_24728,N_24373,N_24208);
nor U24729 (N_24729,N_24173,N_24267);
nor U24730 (N_24730,N_23996,N_23931);
xnor U24731 (N_24731,N_23960,N_24332);
and U24732 (N_24732,N_23949,N_23793);
xnor U24733 (N_24733,N_23964,N_23753);
or U24734 (N_24734,N_23756,N_23847);
nand U24735 (N_24735,N_24175,N_23831);
nand U24736 (N_24736,N_23966,N_24079);
or U24737 (N_24737,N_23949,N_23987);
nand U24738 (N_24738,N_23776,N_24173);
and U24739 (N_24739,N_24156,N_24202);
nand U24740 (N_24740,N_23773,N_24039);
and U24741 (N_24741,N_23750,N_24284);
nand U24742 (N_24742,N_24178,N_24218);
nand U24743 (N_24743,N_23949,N_24194);
and U24744 (N_24744,N_24097,N_23849);
nor U24745 (N_24745,N_24009,N_24284);
xnor U24746 (N_24746,N_24165,N_23750);
xor U24747 (N_24747,N_23935,N_23926);
nor U24748 (N_24748,N_23864,N_23970);
or U24749 (N_24749,N_24248,N_24274);
and U24750 (N_24750,N_23766,N_23842);
or U24751 (N_24751,N_24357,N_23980);
nor U24752 (N_24752,N_23913,N_24011);
and U24753 (N_24753,N_23945,N_24056);
xnor U24754 (N_24754,N_24055,N_24020);
or U24755 (N_24755,N_24345,N_23903);
nand U24756 (N_24756,N_24176,N_24233);
nand U24757 (N_24757,N_24148,N_23905);
nor U24758 (N_24758,N_24247,N_24263);
nor U24759 (N_24759,N_24002,N_23924);
or U24760 (N_24760,N_24152,N_24060);
nand U24761 (N_24761,N_23815,N_23809);
xor U24762 (N_24762,N_23853,N_24038);
nand U24763 (N_24763,N_24191,N_24355);
nand U24764 (N_24764,N_23891,N_23954);
nand U24765 (N_24765,N_24235,N_23838);
or U24766 (N_24766,N_23925,N_23973);
or U24767 (N_24767,N_24169,N_23820);
xor U24768 (N_24768,N_23929,N_23914);
nand U24769 (N_24769,N_23830,N_24031);
nand U24770 (N_24770,N_24353,N_24336);
xnor U24771 (N_24771,N_24360,N_24059);
nor U24772 (N_24772,N_23799,N_24009);
xor U24773 (N_24773,N_23814,N_23956);
or U24774 (N_24774,N_24325,N_24236);
xnor U24775 (N_24775,N_24235,N_24158);
or U24776 (N_24776,N_23878,N_24135);
xnor U24777 (N_24777,N_24362,N_24263);
or U24778 (N_24778,N_24117,N_24241);
nand U24779 (N_24779,N_23803,N_24131);
nor U24780 (N_24780,N_23847,N_24025);
or U24781 (N_24781,N_24310,N_24366);
or U24782 (N_24782,N_23961,N_24211);
nor U24783 (N_24783,N_24049,N_23766);
xnor U24784 (N_24784,N_24248,N_24263);
nand U24785 (N_24785,N_24163,N_24070);
or U24786 (N_24786,N_24320,N_23917);
and U24787 (N_24787,N_24068,N_24180);
and U24788 (N_24788,N_23824,N_24029);
and U24789 (N_24789,N_24017,N_24063);
nor U24790 (N_24790,N_23759,N_23777);
xor U24791 (N_24791,N_24230,N_24039);
nor U24792 (N_24792,N_23936,N_23810);
xnor U24793 (N_24793,N_24002,N_23831);
or U24794 (N_24794,N_24067,N_23789);
xnor U24795 (N_24795,N_24053,N_24140);
or U24796 (N_24796,N_24039,N_23854);
xnor U24797 (N_24797,N_24365,N_24167);
nor U24798 (N_24798,N_24273,N_24210);
nor U24799 (N_24799,N_23775,N_24177);
xor U24800 (N_24800,N_23854,N_24016);
nand U24801 (N_24801,N_24025,N_23961);
nand U24802 (N_24802,N_24160,N_24200);
xor U24803 (N_24803,N_24278,N_24062);
or U24804 (N_24804,N_24356,N_24223);
nor U24805 (N_24805,N_24339,N_24138);
and U24806 (N_24806,N_23940,N_23924);
or U24807 (N_24807,N_23947,N_24218);
nor U24808 (N_24808,N_23891,N_23878);
nor U24809 (N_24809,N_24331,N_24081);
and U24810 (N_24810,N_23805,N_23751);
xnor U24811 (N_24811,N_23969,N_23754);
xor U24812 (N_24812,N_24160,N_23752);
xnor U24813 (N_24813,N_23751,N_24060);
nand U24814 (N_24814,N_23790,N_24003);
xnor U24815 (N_24815,N_23949,N_24064);
nand U24816 (N_24816,N_23919,N_23826);
nand U24817 (N_24817,N_23806,N_23850);
and U24818 (N_24818,N_24207,N_24213);
nor U24819 (N_24819,N_23998,N_24326);
nand U24820 (N_24820,N_24329,N_23786);
and U24821 (N_24821,N_24184,N_23801);
xor U24822 (N_24822,N_24149,N_24343);
or U24823 (N_24823,N_23977,N_24227);
nand U24824 (N_24824,N_24034,N_24146);
or U24825 (N_24825,N_24067,N_24190);
and U24826 (N_24826,N_23842,N_24150);
and U24827 (N_24827,N_24099,N_24277);
xnor U24828 (N_24828,N_24060,N_24264);
nand U24829 (N_24829,N_24112,N_23945);
nand U24830 (N_24830,N_23785,N_23890);
nor U24831 (N_24831,N_24012,N_24313);
nor U24832 (N_24832,N_24043,N_23802);
xor U24833 (N_24833,N_23776,N_24033);
and U24834 (N_24834,N_24216,N_24151);
and U24835 (N_24835,N_24261,N_24034);
nor U24836 (N_24836,N_24227,N_24059);
nor U24837 (N_24837,N_24141,N_23913);
xor U24838 (N_24838,N_24275,N_24136);
xnor U24839 (N_24839,N_24011,N_24034);
and U24840 (N_24840,N_24067,N_24096);
nand U24841 (N_24841,N_23872,N_23937);
and U24842 (N_24842,N_24108,N_24124);
or U24843 (N_24843,N_23790,N_23830);
and U24844 (N_24844,N_24368,N_24055);
nand U24845 (N_24845,N_24250,N_24070);
or U24846 (N_24846,N_23803,N_23819);
nor U24847 (N_24847,N_23751,N_23772);
xnor U24848 (N_24848,N_23943,N_24339);
and U24849 (N_24849,N_23936,N_23915);
xnor U24850 (N_24850,N_24007,N_24048);
nand U24851 (N_24851,N_24097,N_23919);
xnor U24852 (N_24852,N_23791,N_24332);
and U24853 (N_24853,N_24371,N_24327);
and U24854 (N_24854,N_24346,N_23829);
nor U24855 (N_24855,N_24293,N_23895);
nor U24856 (N_24856,N_24189,N_24281);
nor U24857 (N_24857,N_24224,N_23974);
nor U24858 (N_24858,N_23791,N_24085);
nand U24859 (N_24859,N_23828,N_24236);
nor U24860 (N_24860,N_24277,N_24103);
xor U24861 (N_24861,N_23910,N_24072);
xor U24862 (N_24862,N_23783,N_23855);
xor U24863 (N_24863,N_23873,N_24245);
and U24864 (N_24864,N_24221,N_23866);
nand U24865 (N_24865,N_24339,N_23935);
nand U24866 (N_24866,N_24353,N_23829);
or U24867 (N_24867,N_24295,N_24194);
xor U24868 (N_24868,N_24054,N_24301);
nor U24869 (N_24869,N_24127,N_24299);
nand U24870 (N_24870,N_24351,N_24103);
or U24871 (N_24871,N_23870,N_23996);
and U24872 (N_24872,N_24010,N_24311);
or U24873 (N_24873,N_23777,N_23776);
or U24874 (N_24874,N_24336,N_23980);
nand U24875 (N_24875,N_24293,N_24046);
and U24876 (N_24876,N_24279,N_23931);
xor U24877 (N_24877,N_23941,N_23969);
xnor U24878 (N_24878,N_23919,N_24125);
and U24879 (N_24879,N_24077,N_24255);
and U24880 (N_24880,N_24167,N_24141);
xor U24881 (N_24881,N_24326,N_23939);
or U24882 (N_24882,N_24052,N_24004);
nor U24883 (N_24883,N_23804,N_23794);
nand U24884 (N_24884,N_24059,N_23853);
xor U24885 (N_24885,N_23770,N_23966);
xor U24886 (N_24886,N_24354,N_24017);
nand U24887 (N_24887,N_23864,N_24330);
xnor U24888 (N_24888,N_23864,N_23946);
xnor U24889 (N_24889,N_23765,N_24123);
xnor U24890 (N_24890,N_24146,N_23887);
nand U24891 (N_24891,N_24165,N_24317);
xor U24892 (N_24892,N_24042,N_23862);
xnor U24893 (N_24893,N_23942,N_24090);
or U24894 (N_24894,N_24281,N_23864);
xnor U24895 (N_24895,N_24122,N_24037);
nor U24896 (N_24896,N_23891,N_24196);
nand U24897 (N_24897,N_23779,N_23979);
xnor U24898 (N_24898,N_23826,N_24000);
or U24899 (N_24899,N_23795,N_24032);
nor U24900 (N_24900,N_24012,N_23871);
and U24901 (N_24901,N_24071,N_23930);
nand U24902 (N_24902,N_23754,N_23926);
nand U24903 (N_24903,N_24133,N_24196);
and U24904 (N_24904,N_24055,N_24137);
xor U24905 (N_24905,N_23947,N_24200);
nand U24906 (N_24906,N_24321,N_23784);
and U24907 (N_24907,N_24297,N_24289);
xor U24908 (N_24908,N_24367,N_23822);
and U24909 (N_24909,N_24107,N_24146);
or U24910 (N_24910,N_24264,N_24034);
and U24911 (N_24911,N_23755,N_24209);
or U24912 (N_24912,N_23771,N_24347);
nor U24913 (N_24913,N_23926,N_24024);
xnor U24914 (N_24914,N_23941,N_24285);
xor U24915 (N_24915,N_23907,N_23771);
nor U24916 (N_24916,N_24303,N_24117);
and U24917 (N_24917,N_24081,N_23823);
nand U24918 (N_24918,N_23996,N_24305);
nor U24919 (N_24919,N_24033,N_23833);
xnor U24920 (N_24920,N_24055,N_24349);
and U24921 (N_24921,N_24017,N_24093);
or U24922 (N_24922,N_23915,N_24343);
and U24923 (N_24923,N_23875,N_24283);
nor U24924 (N_24924,N_23963,N_24038);
nor U24925 (N_24925,N_24177,N_23846);
or U24926 (N_24926,N_24329,N_23942);
nor U24927 (N_24927,N_24084,N_23802);
or U24928 (N_24928,N_23915,N_23904);
and U24929 (N_24929,N_23908,N_24217);
nand U24930 (N_24930,N_24344,N_24014);
and U24931 (N_24931,N_24041,N_23883);
and U24932 (N_24932,N_23932,N_23762);
nor U24933 (N_24933,N_24119,N_24002);
or U24934 (N_24934,N_24258,N_24281);
xor U24935 (N_24935,N_24065,N_23854);
xor U24936 (N_24936,N_24256,N_23811);
or U24937 (N_24937,N_23840,N_24054);
nor U24938 (N_24938,N_23940,N_24240);
or U24939 (N_24939,N_24000,N_23921);
and U24940 (N_24940,N_23967,N_24214);
xnor U24941 (N_24941,N_23801,N_24351);
and U24942 (N_24942,N_24092,N_23830);
xnor U24943 (N_24943,N_24135,N_24252);
xor U24944 (N_24944,N_24124,N_23981);
or U24945 (N_24945,N_24029,N_23752);
or U24946 (N_24946,N_24068,N_23883);
nand U24947 (N_24947,N_24051,N_24353);
and U24948 (N_24948,N_24043,N_24105);
nor U24949 (N_24949,N_24333,N_23874);
or U24950 (N_24950,N_23836,N_24273);
or U24951 (N_24951,N_24147,N_23958);
nand U24952 (N_24952,N_23954,N_23910);
nand U24953 (N_24953,N_23765,N_24112);
or U24954 (N_24954,N_24068,N_23827);
nand U24955 (N_24955,N_24351,N_24213);
xor U24956 (N_24956,N_24094,N_24099);
or U24957 (N_24957,N_24374,N_23910);
xor U24958 (N_24958,N_24153,N_23902);
and U24959 (N_24959,N_23870,N_23888);
nand U24960 (N_24960,N_24138,N_24169);
or U24961 (N_24961,N_23764,N_24297);
xnor U24962 (N_24962,N_24010,N_24281);
nand U24963 (N_24963,N_23869,N_23969);
nand U24964 (N_24964,N_24219,N_24267);
xnor U24965 (N_24965,N_23844,N_24304);
or U24966 (N_24966,N_23899,N_24023);
and U24967 (N_24967,N_24239,N_24318);
xnor U24968 (N_24968,N_23862,N_23990);
or U24969 (N_24969,N_24010,N_23808);
nand U24970 (N_24970,N_24265,N_23751);
and U24971 (N_24971,N_24227,N_24041);
nand U24972 (N_24972,N_24153,N_23968);
or U24973 (N_24973,N_23955,N_23865);
nor U24974 (N_24974,N_24053,N_24292);
and U24975 (N_24975,N_23812,N_24286);
nor U24976 (N_24976,N_24133,N_24330);
xor U24977 (N_24977,N_24205,N_23756);
nor U24978 (N_24978,N_24342,N_23941);
and U24979 (N_24979,N_24042,N_24052);
and U24980 (N_24980,N_23799,N_24264);
and U24981 (N_24981,N_24273,N_24109);
or U24982 (N_24982,N_23862,N_24046);
or U24983 (N_24983,N_24242,N_24369);
xor U24984 (N_24984,N_24260,N_23888);
or U24985 (N_24985,N_23840,N_24228);
nand U24986 (N_24986,N_23763,N_24221);
nand U24987 (N_24987,N_24268,N_23801);
and U24988 (N_24988,N_23827,N_23809);
nand U24989 (N_24989,N_23899,N_24211);
and U24990 (N_24990,N_23934,N_23769);
nor U24991 (N_24991,N_24034,N_24110);
and U24992 (N_24992,N_23956,N_23884);
and U24993 (N_24993,N_23991,N_23882);
or U24994 (N_24994,N_24071,N_23763);
and U24995 (N_24995,N_24057,N_23855);
nand U24996 (N_24996,N_24368,N_23988);
xnor U24997 (N_24997,N_24326,N_23792);
nor U24998 (N_24998,N_24039,N_23946);
and U24999 (N_24999,N_24052,N_23752);
nand UO_0 (O_0,N_24811,N_24760);
and UO_1 (O_1,N_24881,N_24829);
or UO_2 (O_2,N_24433,N_24609);
or UO_3 (O_3,N_24737,N_24721);
and UO_4 (O_4,N_24405,N_24919);
or UO_5 (O_5,N_24685,N_24482);
nor UO_6 (O_6,N_24741,N_24650);
xnor UO_7 (O_7,N_24610,N_24856);
or UO_8 (O_8,N_24630,N_24455);
nand UO_9 (O_9,N_24873,N_24532);
nor UO_10 (O_10,N_24801,N_24653);
nor UO_11 (O_11,N_24850,N_24605);
nor UO_12 (O_12,N_24812,N_24566);
or UO_13 (O_13,N_24646,N_24460);
xor UO_14 (O_14,N_24902,N_24839);
and UO_15 (O_15,N_24843,N_24485);
xnor UO_16 (O_16,N_24535,N_24662);
and UO_17 (O_17,N_24614,N_24979);
or UO_18 (O_18,N_24488,N_24794);
xnor UO_19 (O_19,N_24771,N_24861);
and UO_20 (O_20,N_24865,N_24389);
nand UO_21 (O_21,N_24793,N_24571);
and UO_22 (O_22,N_24710,N_24836);
and UO_23 (O_23,N_24501,N_24676);
or UO_24 (O_24,N_24738,N_24623);
xnor UO_25 (O_25,N_24742,N_24819);
nor UO_26 (O_26,N_24953,N_24489);
nand UO_27 (O_27,N_24820,N_24492);
or UO_28 (O_28,N_24845,N_24739);
and UO_29 (O_29,N_24642,N_24858);
and UO_30 (O_30,N_24773,N_24823);
nor UO_31 (O_31,N_24443,N_24709);
nand UO_32 (O_32,N_24669,N_24528);
nor UO_33 (O_33,N_24929,N_24853);
or UO_34 (O_34,N_24775,N_24519);
nor UO_35 (O_35,N_24424,N_24608);
xnor UO_36 (O_36,N_24831,N_24525);
nand UO_37 (O_37,N_24493,N_24395);
nor UO_38 (O_38,N_24931,N_24841);
nor UO_39 (O_39,N_24572,N_24783);
nand UO_40 (O_40,N_24756,N_24692);
or UO_41 (O_41,N_24683,N_24705);
xor UO_42 (O_42,N_24536,N_24557);
or UO_43 (O_43,N_24654,N_24997);
and UO_44 (O_44,N_24896,N_24416);
nand UO_45 (O_45,N_24449,N_24659);
nand UO_46 (O_46,N_24852,N_24963);
nor UO_47 (O_47,N_24833,N_24516);
nand UO_48 (O_48,N_24696,N_24437);
and UO_49 (O_49,N_24450,N_24988);
nor UO_50 (O_50,N_24989,N_24969);
nor UO_51 (O_51,N_24951,N_24457);
nor UO_52 (O_52,N_24549,N_24418);
or UO_53 (O_53,N_24984,N_24815);
or UO_54 (O_54,N_24407,N_24500);
nor UO_55 (O_55,N_24644,N_24784);
xnor UO_56 (O_56,N_24928,N_24452);
xor UO_57 (O_57,N_24638,N_24734);
nand UO_58 (O_58,N_24480,N_24907);
nand UO_59 (O_59,N_24874,N_24503);
nand UO_60 (O_60,N_24816,N_24621);
nand UO_61 (O_61,N_24666,N_24444);
and UO_62 (O_62,N_24466,N_24565);
and UO_63 (O_63,N_24386,N_24461);
nand UO_64 (O_64,N_24691,N_24906);
or UO_65 (O_65,N_24553,N_24592);
and UO_66 (O_66,N_24766,N_24712);
nand UO_67 (O_67,N_24419,N_24959);
or UO_68 (O_68,N_24952,N_24392);
nand UO_69 (O_69,N_24505,N_24777);
xor UO_70 (O_70,N_24656,N_24698);
nor UO_71 (O_71,N_24383,N_24755);
xnor UO_72 (O_72,N_24910,N_24596);
or UO_73 (O_73,N_24926,N_24660);
or UO_74 (O_74,N_24504,N_24417);
xnor UO_75 (O_75,N_24943,N_24795);
or UO_76 (O_76,N_24378,N_24991);
xor UO_77 (O_77,N_24432,N_24606);
nor UO_78 (O_78,N_24915,N_24972);
nor UO_79 (O_79,N_24474,N_24448);
nand UO_80 (O_80,N_24736,N_24765);
nor UO_81 (O_81,N_24479,N_24851);
and UO_82 (O_82,N_24796,N_24577);
or UO_83 (O_83,N_24636,N_24468);
or UO_84 (O_84,N_24593,N_24380);
and UO_85 (O_85,N_24904,N_24453);
and UO_86 (O_86,N_24661,N_24863);
or UO_87 (O_87,N_24764,N_24758);
and UO_88 (O_88,N_24379,N_24387);
nor UO_89 (O_89,N_24899,N_24888);
or UO_90 (O_90,N_24626,N_24859);
or UO_91 (O_91,N_24876,N_24537);
xnor UO_92 (O_92,N_24624,N_24703);
nor UO_93 (O_93,N_24599,N_24600);
or UO_94 (O_94,N_24940,N_24830);
and UO_95 (O_95,N_24442,N_24441);
and UO_96 (O_96,N_24866,N_24579);
and UO_97 (O_97,N_24552,N_24996);
and UO_98 (O_98,N_24607,N_24499);
and UO_99 (O_99,N_24540,N_24822);
or UO_100 (O_100,N_24745,N_24456);
nand UO_101 (O_101,N_24498,N_24923);
nand UO_102 (O_102,N_24806,N_24918);
and UO_103 (O_103,N_24744,N_24882);
xor UO_104 (O_104,N_24476,N_24983);
xnor UO_105 (O_105,N_24717,N_24458);
and UO_106 (O_106,N_24772,N_24768);
nand UO_107 (O_107,N_24469,N_24451);
and UO_108 (O_108,N_24770,N_24686);
nand UO_109 (O_109,N_24994,N_24697);
or UO_110 (O_110,N_24995,N_24639);
and UO_111 (O_111,N_24531,N_24990);
nor UO_112 (O_112,N_24564,N_24715);
xnor UO_113 (O_113,N_24590,N_24497);
nor UO_114 (O_114,N_24725,N_24687);
nand UO_115 (O_115,N_24518,N_24975);
and UO_116 (O_116,N_24522,N_24818);
or UO_117 (O_117,N_24999,N_24707);
and UO_118 (O_118,N_24948,N_24809);
nor UO_119 (O_119,N_24837,N_24581);
xnor UO_120 (O_120,N_24539,N_24484);
nor UO_121 (O_121,N_24509,N_24752);
or UO_122 (O_122,N_24932,N_24584);
nand UO_123 (O_123,N_24708,N_24748);
nand UO_124 (O_124,N_24619,N_24699);
xor UO_125 (O_125,N_24917,N_24547);
and UO_126 (O_126,N_24527,N_24568);
or UO_127 (O_127,N_24757,N_24862);
and UO_128 (O_128,N_24467,N_24575);
or UO_129 (O_129,N_24804,N_24916);
or UO_130 (O_130,N_24462,N_24560);
xor UO_131 (O_131,N_24496,N_24561);
nand UO_132 (O_132,N_24478,N_24486);
nand UO_133 (O_133,N_24641,N_24652);
xor UO_134 (O_134,N_24912,N_24515);
and UO_135 (O_135,N_24588,N_24582);
nor UO_136 (O_136,N_24648,N_24807);
nand UO_137 (O_137,N_24838,N_24594);
and UO_138 (O_138,N_24665,N_24941);
nand UO_139 (O_139,N_24724,N_24643);
nand UO_140 (O_140,N_24747,N_24473);
nand UO_141 (O_141,N_24601,N_24595);
and UO_142 (O_142,N_24423,N_24868);
nand UO_143 (O_143,N_24754,N_24589);
or UO_144 (O_144,N_24440,N_24897);
nand UO_145 (O_145,N_24787,N_24920);
and UO_146 (O_146,N_24938,N_24970);
or UO_147 (O_147,N_24978,N_24835);
nor UO_148 (O_148,N_24554,N_24631);
or UO_149 (O_149,N_24821,N_24889);
and UO_150 (O_150,N_24377,N_24393);
nor UO_151 (O_151,N_24690,N_24834);
or UO_152 (O_152,N_24569,N_24967);
xnor UO_153 (O_153,N_24810,N_24957);
nand UO_154 (O_154,N_24769,N_24583);
xor UO_155 (O_155,N_24847,N_24625);
nor UO_156 (O_156,N_24936,N_24640);
or UO_157 (O_157,N_24883,N_24628);
and UO_158 (O_158,N_24611,N_24517);
or UO_159 (O_159,N_24550,N_24799);
nand UO_160 (O_160,N_24586,N_24844);
nand UO_161 (O_161,N_24421,N_24827);
nor UO_162 (O_162,N_24732,N_24950);
and UO_163 (O_163,N_24622,N_24849);
nor UO_164 (O_164,N_24427,N_24723);
nor UO_165 (O_165,N_24733,N_24598);
nand UO_166 (O_166,N_24776,N_24558);
xnor UO_167 (O_167,N_24574,N_24805);
xnor UO_168 (O_168,N_24746,N_24792);
nand UO_169 (O_169,N_24958,N_24510);
and UO_170 (O_170,N_24426,N_24658);
and UO_171 (O_171,N_24502,N_24790);
xor UO_172 (O_172,N_24872,N_24743);
or UO_173 (O_173,N_24908,N_24487);
nand UO_174 (O_174,N_24924,N_24727);
nor UO_175 (O_175,N_24668,N_24587);
nand UO_176 (O_176,N_24616,N_24753);
and UO_177 (O_177,N_24693,N_24701);
nor UO_178 (O_178,N_24922,N_24892);
nand UO_179 (O_179,N_24731,N_24800);
nand UO_180 (O_180,N_24678,N_24927);
and UO_181 (O_181,N_24490,N_24947);
nand UO_182 (O_182,N_24645,N_24559);
and UO_183 (O_183,N_24375,N_24446);
nor UO_184 (O_184,N_24533,N_24785);
xnor UO_185 (O_185,N_24798,N_24620);
or UO_186 (O_186,N_24401,N_24411);
nand UO_187 (O_187,N_24680,N_24993);
nand UO_188 (O_188,N_24431,N_24781);
xor UO_189 (O_189,N_24671,N_24846);
or UO_190 (O_190,N_24454,N_24774);
nor UO_191 (O_191,N_24430,N_24730);
or UO_192 (O_192,N_24570,N_24871);
or UO_193 (O_193,N_24848,N_24942);
nand UO_194 (O_194,N_24397,N_24403);
xor UO_195 (O_195,N_24935,N_24543);
nor UO_196 (O_196,N_24885,N_24637);
nand UO_197 (O_197,N_24491,N_24961);
nand UO_198 (O_198,N_24546,N_24713);
or UO_199 (O_199,N_24428,N_24657);
nor UO_200 (O_200,N_24884,N_24962);
xor UO_201 (O_201,N_24376,N_24400);
and UO_202 (O_202,N_24728,N_24808);
nor UO_203 (O_203,N_24413,N_24706);
nand UO_204 (O_204,N_24782,N_24627);
and UO_205 (O_205,N_24985,N_24980);
or UO_206 (O_206,N_24726,N_24524);
and UO_207 (O_207,N_24946,N_24767);
nand UO_208 (O_208,N_24465,N_24870);
and UO_209 (O_209,N_24689,N_24722);
xnor UO_210 (O_210,N_24530,N_24711);
or UO_211 (O_211,N_24495,N_24463);
and UO_212 (O_212,N_24511,N_24679);
or UO_213 (O_213,N_24651,N_24634);
nor UO_214 (O_214,N_24973,N_24508);
xnor UO_215 (O_215,N_24933,N_24481);
nand UO_216 (O_216,N_24802,N_24420);
and UO_217 (O_217,N_24814,N_24551);
and UO_218 (O_218,N_24716,N_24635);
and UO_219 (O_219,N_24789,N_24780);
xnor UO_220 (O_220,N_24398,N_24410);
xor UO_221 (O_221,N_24471,N_24913);
or UO_222 (O_222,N_24966,N_24576);
xnor UO_223 (O_223,N_24740,N_24388);
nand UO_224 (O_224,N_24521,N_24415);
and UO_225 (O_225,N_24880,N_24826);
xnor UO_226 (O_226,N_24914,N_24877);
and UO_227 (O_227,N_24925,N_24677);
nor UO_228 (O_228,N_24391,N_24857);
and UO_229 (O_229,N_24944,N_24682);
nor UO_230 (O_230,N_24567,N_24475);
xnor UO_231 (O_231,N_24613,N_24893);
xnor UO_232 (O_232,N_24986,N_24887);
and UO_233 (O_233,N_24900,N_24750);
xor UO_234 (O_234,N_24384,N_24905);
nor UO_235 (O_235,N_24779,N_24681);
or UO_236 (O_236,N_24909,N_24464);
nand UO_237 (O_237,N_24992,N_24414);
nand UO_238 (O_238,N_24939,N_24976);
or UO_239 (O_239,N_24633,N_24506);
and UO_240 (O_240,N_24629,N_24408);
nor UO_241 (O_241,N_24674,N_24447);
or UO_242 (O_242,N_24720,N_24615);
or UO_243 (O_243,N_24921,N_24949);
and UO_244 (O_244,N_24672,N_24700);
xnor UO_245 (O_245,N_24761,N_24520);
nor UO_246 (O_246,N_24390,N_24612);
nand UO_247 (O_247,N_24429,N_24472);
or UO_248 (O_248,N_24751,N_24759);
nor UO_249 (O_249,N_24470,N_24507);
xor UO_250 (O_250,N_24667,N_24542);
nor UO_251 (O_251,N_24869,N_24459);
and UO_252 (O_252,N_24791,N_24578);
xnor UO_253 (O_253,N_24494,N_24523);
xnor UO_254 (O_254,N_24778,N_24675);
nand UO_255 (O_255,N_24512,N_24585);
and UO_256 (O_256,N_24937,N_24555);
nand UO_257 (O_257,N_24664,N_24435);
or UO_258 (O_258,N_24749,N_24824);
nand UO_259 (O_259,N_24832,N_24898);
or UO_260 (O_260,N_24903,N_24655);
xor UO_261 (O_261,N_24878,N_24409);
xor UO_262 (O_262,N_24434,N_24911);
nor UO_263 (O_263,N_24477,N_24597);
nor UO_264 (O_264,N_24573,N_24890);
nor UO_265 (O_265,N_24617,N_24875);
xor UO_266 (O_266,N_24860,N_24735);
xnor UO_267 (O_267,N_24945,N_24422);
or UO_268 (O_268,N_24385,N_24513);
and UO_269 (O_269,N_24394,N_24526);
nand UO_270 (O_270,N_24602,N_24894);
xnor UO_271 (O_271,N_24439,N_24649);
nor UO_272 (O_272,N_24534,N_24483);
or UO_273 (O_273,N_24563,N_24647);
or UO_274 (O_274,N_24854,N_24842);
and UO_275 (O_275,N_24406,N_24425);
nand UO_276 (O_276,N_24977,N_24436);
and UO_277 (O_277,N_24895,N_24545);
or UO_278 (O_278,N_24987,N_24688);
xor UO_279 (O_279,N_24718,N_24956);
nand UO_280 (O_280,N_24438,N_24381);
or UO_281 (O_281,N_24797,N_24673);
and UO_282 (O_282,N_24632,N_24603);
nand UO_283 (O_283,N_24901,N_24763);
nand UO_284 (O_284,N_24934,N_24840);
xnor UO_285 (O_285,N_24684,N_24982);
xnor UO_286 (O_286,N_24813,N_24412);
nor UO_287 (O_287,N_24930,N_24729);
or UO_288 (O_288,N_24719,N_24788);
xnor UO_289 (O_289,N_24954,N_24803);
and UO_290 (O_290,N_24762,N_24825);
nor UO_291 (O_291,N_24864,N_24541);
xor UO_292 (O_292,N_24404,N_24618);
nor UO_293 (O_293,N_24886,N_24694);
or UO_294 (O_294,N_24704,N_24879);
nand UO_295 (O_295,N_24971,N_24399);
or UO_296 (O_296,N_24663,N_24556);
and UO_297 (O_297,N_24960,N_24529);
nand UO_298 (O_298,N_24964,N_24855);
nor UO_299 (O_299,N_24695,N_24514);
and UO_300 (O_300,N_24544,N_24965);
nor UO_301 (O_301,N_24402,N_24538);
or UO_302 (O_302,N_24445,N_24548);
xnor UO_303 (O_303,N_24591,N_24670);
and UO_304 (O_304,N_24396,N_24867);
and UO_305 (O_305,N_24562,N_24714);
nor UO_306 (O_306,N_24968,N_24974);
nand UO_307 (O_307,N_24786,N_24891);
nor UO_308 (O_308,N_24955,N_24998);
and UO_309 (O_309,N_24580,N_24817);
and UO_310 (O_310,N_24828,N_24702);
xor UO_311 (O_311,N_24382,N_24604);
nand UO_312 (O_312,N_24981,N_24985);
nor UO_313 (O_313,N_24845,N_24431);
nor UO_314 (O_314,N_24733,N_24820);
nor UO_315 (O_315,N_24872,N_24830);
xnor UO_316 (O_316,N_24798,N_24528);
xnor UO_317 (O_317,N_24579,N_24389);
xor UO_318 (O_318,N_24805,N_24749);
xor UO_319 (O_319,N_24726,N_24899);
nand UO_320 (O_320,N_24567,N_24946);
xor UO_321 (O_321,N_24752,N_24960);
nand UO_322 (O_322,N_24454,N_24442);
nor UO_323 (O_323,N_24978,N_24429);
xor UO_324 (O_324,N_24933,N_24583);
or UO_325 (O_325,N_24688,N_24650);
nand UO_326 (O_326,N_24759,N_24774);
or UO_327 (O_327,N_24648,N_24502);
nand UO_328 (O_328,N_24825,N_24446);
nor UO_329 (O_329,N_24820,N_24896);
nand UO_330 (O_330,N_24583,N_24646);
and UO_331 (O_331,N_24982,N_24379);
xor UO_332 (O_332,N_24403,N_24885);
nor UO_333 (O_333,N_24379,N_24679);
nand UO_334 (O_334,N_24429,N_24559);
and UO_335 (O_335,N_24521,N_24472);
nor UO_336 (O_336,N_24614,N_24870);
xor UO_337 (O_337,N_24577,N_24926);
nand UO_338 (O_338,N_24519,N_24977);
xor UO_339 (O_339,N_24394,N_24459);
nor UO_340 (O_340,N_24435,N_24584);
and UO_341 (O_341,N_24405,N_24986);
and UO_342 (O_342,N_24497,N_24930);
or UO_343 (O_343,N_24743,N_24487);
nor UO_344 (O_344,N_24700,N_24840);
nand UO_345 (O_345,N_24375,N_24903);
or UO_346 (O_346,N_24711,N_24567);
xor UO_347 (O_347,N_24966,N_24833);
or UO_348 (O_348,N_24961,N_24588);
and UO_349 (O_349,N_24782,N_24484);
nor UO_350 (O_350,N_24453,N_24496);
and UO_351 (O_351,N_24380,N_24705);
xnor UO_352 (O_352,N_24886,N_24898);
or UO_353 (O_353,N_24545,N_24729);
nand UO_354 (O_354,N_24679,N_24978);
and UO_355 (O_355,N_24454,N_24768);
nand UO_356 (O_356,N_24943,N_24621);
nand UO_357 (O_357,N_24919,N_24981);
nand UO_358 (O_358,N_24922,N_24632);
xor UO_359 (O_359,N_24638,N_24680);
nor UO_360 (O_360,N_24546,N_24544);
xnor UO_361 (O_361,N_24688,N_24509);
nor UO_362 (O_362,N_24928,N_24988);
and UO_363 (O_363,N_24959,N_24492);
nor UO_364 (O_364,N_24634,N_24568);
xnor UO_365 (O_365,N_24442,N_24618);
and UO_366 (O_366,N_24705,N_24748);
nor UO_367 (O_367,N_24868,N_24999);
or UO_368 (O_368,N_24955,N_24553);
or UO_369 (O_369,N_24478,N_24698);
nand UO_370 (O_370,N_24653,N_24634);
and UO_371 (O_371,N_24654,N_24586);
and UO_372 (O_372,N_24477,N_24389);
nor UO_373 (O_373,N_24468,N_24517);
xnor UO_374 (O_374,N_24648,N_24819);
or UO_375 (O_375,N_24630,N_24708);
nor UO_376 (O_376,N_24949,N_24746);
nand UO_377 (O_377,N_24446,N_24813);
or UO_378 (O_378,N_24622,N_24477);
xnor UO_379 (O_379,N_24934,N_24492);
or UO_380 (O_380,N_24647,N_24535);
or UO_381 (O_381,N_24841,N_24522);
or UO_382 (O_382,N_24392,N_24457);
nor UO_383 (O_383,N_24496,N_24990);
or UO_384 (O_384,N_24645,N_24581);
nor UO_385 (O_385,N_24376,N_24488);
or UO_386 (O_386,N_24526,N_24511);
or UO_387 (O_387,N_24903,N_24398);
or UO_388 (O_388,N_24392,N_24887);
and UO_389 (O_389,N_24981,N_24711);
nand UO_390 (O_390,N_24448,N_24916);
and UO_391 (O_391,N_24707,N_24452);
or UO_392 (O_392,N_24953,N_24574);
xor UO_393 (O_393,N_24585,N_24750);
nand UO_394 (O_394,N_24561,N_24386);
xor UO_395 (O_395,N_24740,N_24465);
nand UO_396 (O_396,N_24867,N_24516);
and UO_397 (O_397,N_24572,N_24627);
nand UO_398 (O_398,N_24583,N_24880);
or UO_399 (O_399,N_24492,N_24587);
xor UO_400 (O_400,N_24780,N_24915);
xor UO_401 (O_401,N_24439,N_24938);
and UO_402 (O_402,N_24580,N_24724);
xnor UO_403 (O_403,N_24623,N_24932);
or UO_404 (O_404,N_24460,N_24541);
or UO_405 (O_405,N_24912,N_24678);
or UO_406 (O_406,N_24856,N_24600);
and UO_407 (O_407,N_24389,N_24709);
or UO_408 (O_408,N_24882,N_24910);
nor UO_409 (O_409,N_24593,N_24813);
nand UO_410 (O_410,N_24420,N_24988);
nor UO_411 (O_411,N_24723,N_24446);
and UO_412 (O_412,N_24500,N_24674);
nand UO_413 (O_413,N_24993,N_24441);
nand UO_414 (O_414,N_24880,N_24701);
or UO_415 (O_415,N_24563,N_24627);
xnor UO_416 (O_416,N_24723,N_24665);
nor UO_417 (O_417,N_24887,N_24705);
xor UO_418 (O_418,N_24456,N_24537);
nand UO_419 (O_419,N_24422,N_24449);
or UO_420 (O_420,N_24600,N_24577);
nor UO_421 (O_421,N_24444,N_24834);
xnor UO_422 (O_422,N_24642,N_24412);
nor UO_423 (O_423,N_24678,N_24588);
nand UO_424 (O_424,N_24478,N_24594);
xor UO_425 (O_425,N_24591,N_24796);
nor UO_426 (O_426,N_24941,N_24886);
and UO_427 (O_427,N_24771,N_24910);
nand UO_428 (O_428,N_24922,N_24407);
nor UO_429 (O_429,N_24879,N_24842);
or UO_430 (O_430,N_24878,N_24927);
and UO_431 (O_431,N_24904,N_24745);
nor UO_432 (O_432,N_24758,N_24445);
nor UO_433 (O_433,N_24526,N_24897);
and UO_434 (O_434,N_24555,N_24811);
and UO_435 (O_435,N_24999,N_24744);
and UO_436 (O_436,N_24537,N_24727);
xor UO_437 (O_437,N_24457,N_24448);
and UO_438 (O_438,N_24904,N_24726);
xnor UO_439 (O_439,N_24675,N_24739);
nor UO_440 (O_440,N_24693,N_24996);
or UO_441 (O_441,N_24639,N_24843);
nor UO_442 (O_442,N_24746,N_24822);
xor UO_443 (O_443,N_24887,N_24385);
nor UO_444 (O_444,N_24466,N_24548);
or UO_445 (O_445,N_24377,N_24811);
xnor UO_446 (O_446,N_24555,N_24759);
nand UO_447 (O_447,N_24818,N_24483);
or UO_448 (O_448,N_24484,N_24909);
or UO_449 (O_449,N_24646,N_24657);
or UO_450 (O_450,N_24884,N_24907);
xor UO_451 (O_451,N_24637,N_24500);
xnor UO_452 (O_452,N_24638,N_24403);
nand UO_453 (O_453,N_24521,N_24813);
or UO_454 (O_454,N_24948,N_24544);
and UO_455 (O_455,N_24780,N_24409);
xor UO_456 (O_456,N_24744,N_24521);
nand UO_457 (O_457,N_24766,N_24762);
nor UO_458 (O_458,N_24615,N_24704);
nor UO_459 (O_459,N_24919,N_24907);
xnor UO_460 (O_460,N_24398,N_24630);
nor UO_461 (O_461,N_24481,N_24672);
or UO_462 (O_462,N_24899,N_24488);
nor UO_463 (O_463,N_24440,N_24786);
nor UO_464 (O_464,N_24568,N_24936);
xor UO_465 (O_465,N_24639,N_24663);
or UO_466 (O_466,N_24893,N_24796);
or UO_467 (O_467,N_24885,N_24929);
nand UO_468 (O_468,N_24992,N_24771);
nand UO_469 (O_469,N_24455,N_24553);
and UO_470 (O_470,N_24916,N_24410);
xnor UO_471 (O_471,N_24719,N_24868);
nor UO_472 (O_472,N_24419,N_24410);
xnor UO_473 (O_473,N_24476,N_24812);
xor UO_474 (O_474,N_24929,N_24975);
xnor UO_475 (O_475,N_24972,N_24665);
nor UO_476 (O_476,N_24828,N_24956);
xor UO_477 (O_477,N_24906,N_24772);
nor UO_478 (O_478,N_24621,N_24458);
nor UO_479 (O_479,N_24812,N_24850);
xor UO_480 (O_480,N_24755,N_24449);
xnor UO_481 (O_481,N_24459,N_24559);
nand UO_482 (O_482,N_24987,N_24624);
xor UO_483 (O_483,N_24474,N_24582);
and UO_484 (O_484,N_24949,N_24510);
nor UO_485 (O_485,N_24425,N_24655);
or UO_486 (O_486,N_24789,N_24717);
nor UO_487 (O_487,N_24536,N_24767);
and UO_488 (O_488,N_24801,N_24541);
nor UO_489 (O_489,N_24818,N_24946);
nand UO_490 (O_490,N_24724,N_24428);
nand UO_491 (O_491,N_24882,N_24843);
and UO_492 (O_492,N_24696,N_24771);
nor UO_493 (O_493,N_24594,N_24906);
or UO_494 (O_494,N_24523,N_24786);
nor UO_495 (O_495,N_24460,N_24431);
xnor UO_496 (O_496,N_24714,N_24553);
or UO_497 (O_497,N_24748,N_24626);
xor UO_498 (O_498,N_24882,N_24504);
or UO_499 (O_499,N_24801,N_24774);
or UO_500 (O_500,N_24508,N_24783);
or UO_501 (O_501,N_24560,N_24851);
xnor UO_502 (O_502,N_24972,N_24427);
xor UO_503 (O_503,N_24840,N_24419);
nand UO_504 (O_504,N_24941,N_24692);
nand UO_505 (O_505,N_24608,N_24945);
nor UO_506 (O_506,N_24835,N_24379);
and UO_507 (O_507,N_24506,N_24834);
and UO_508 (O_508,N_24403,N_24553);
nand UO_509 (O_509,N_24733,N_24874);
or UO_510 (O_510,N_24651,N_24971);
nor UO_511 (O_511,N_24732,N_24832);
nand UO_512 (O_512,N_24827,N_24839);
or UO_513 (O_513,N_24453,N_24594);
xnor UO_514 (O_514,N_24593,N_24556);
or UO_515 (O_515,N_24615,N_24861);
nand UO_516 (O_516,N_24715,N_24409);
and UO_517 (O_517,N_24693,N_24535);
nand UO_518 (O_518,N_24816,N_24757);
or UO_519 (O_519,N_24396,N_24987);
or UO_520 (O_520,N_24818,N_24405);
or UO_521 (O_521,N_24580,N_24969);
and UO_522 (O_522,N_24695,N_24926);
or UO_523 (O_523,N_24762,N_24526);
and UO_524 (O_524,N_24677,N_24746);
or UO_525 (O_525,N_24625,N_24826);
xnor UO_526 (O_526,N_24577,N_24928);
nand UO_527 (O_527,N_24785,N_24896);
or UO_528 (O_528,N_24954,N_24926);
xnor UO_529 (O_529,N_24795,N_24924);
or UO_530 (O_530,N_24946,N_24920);
or UO_531 (O_531,N_24849,N_24389);
nand UO_532 (O_532,N_24603,N_24508);
xnor UO_533 (O_533,N_24710,N_24848);
xnor UO_534 (O_534,N_24540,N_24993);
xnor UO_535 (O_535,N_24483,N_24945);
nand UO_536 (O_536,N_24453,N_24471);
nor UO_537 (O_537,N_24553,N_24865);
or UO_538 (O_538,N_24377,N_24905);
and UO_539 (O_539,N_24463,N_24988);
nor UO_540 (O_540,N_24810,N_24704);
nand UO_541 (O_541,N_24671,N_24456);
or UO_542 (O_542,N_24634,N_24465);
and UO_543 (O_543,N_24874,N_24675);
or UO_544 (O_544,N_24767,N_24418);
nand UO_545 (O_545,N_24493,N_24423);
nand UO_546 (O_546,N_24793,N_24805);
and UO_547 (O_547,N_24621,N_24774);
and UO_548 (O_548,N_24495,N_24448);
nor UO_549 (O_549,N_24428,N_24850);
nor UO_550 (O_550,N_24603,N_24803);
nand UO_551 (O_551,N_24752,N_24700);
xnor UO_552 (O_552,N_24389,N_24815);
or UO_553 (O_553,N_24536,N_24850);
nand UO_554 (O_554,N_24742,N_24820);
nand UO_555 (O_555,N_24955,N_24903);
nor UO_556 (O_556,N_24494,N_24987);
xor UO_557 (O_557,N_24825,N_24552);
nand UO_558 (O_558,N_24711,N_24905);
nand UO_559 (O_559,N_24774,N_24583);
and UO_560 (O_560,N_24438,N_24672);
or UO_561 (O_561,N_24638,N_24855);
nand UO_562 (O_562,N_24598,N_24824);
or UO_563 (O_563,N_24791,N_24525);
and UO_564 (O_564,N_24890,N_24809);
and UO_565 (O_565,N_24799,N_24971);
nand UO_566 (O_566,N_24976,N_24803);
and UO_567 (O_567,N_24382,N_24541);
nand UO_568 (O_568,N_24465,N_24947);
and UO_569 (O_569,N_24412,N_24911);
xor UO_570 (O_570,N_24437,N_24931);
nor UO_571 (O_571,N_24379,N_24768);
nand UO_572 (O_572,N_24954,N_24543);
or UO_573 (O_573,N_24433,N_24943);
nor UO_574 (O_574,N_24681,N_24453);
nor UO_575 (O_575,N_24413,N_24522);
xor UO_576 (O_576,N_24477,N_24845);
nand UO_577 (O_577,N_24851,N_24806);
and UO_578 (O_578,N_24454,N_24890);
nor UO_579 (O_579,N_24377,N_24637);
nand UO_580 (O_580,N_24880,N_24854);
nor UO_581 (O_581,N_24524,N_24788);
or UO_582 (O_582,N_24553,N_24731);
and UO_583 (O_583,N_24512,N_24394);
xnor UO_584 (O_584,N_24792,N_24822);
or UO_585 (O_585,N_24603,N_24879);
and UO_586 (O_586,N_24559,N_24713);
nand UO_587 (O_587,N_24646,N_24654);
nand UO_588 (O_588,N_24943,N_24755);
nor UO_589 (O_589,N_24554,N_24847);
xor UO_590 (O_590,N_24684,N_24734);
and UO_591 (O_591,N_24729,N_24724);
nor UO_592 (O_592,N_24411,N_24560);
and UO_593 (O_593,N_24777,N_24449);
nor UO_594 (O_594,N_24737,N_24853);
and UO_595 (O_595,N_24464,N_24515);
and UO_596 (O_596,N_24663,N_24581);
nand UO_597 (O_597,N_24905,N_24498);
nand UO_598 (O_598,N_24659,N_24557);
and UO_599 (O_599,N_24445,N_24659);
nor UO_600 (O_600,N_24542,N_24636);
or UO_601 (O_601,N_24624,N_24566);
nor UO_602 (O_602,N_24985,N_24722);
xnor UO_603 (O_603,N_24865,N_24421);
nor UO_604 (O_604,N_24389,N_24707);
or UO_605 (O_605,N_24621,N_24593);
or UO_606 (O_606,N_24741,N_24591);
nand UO_607 (O_607,N_24813,N_24493);
and UO_608 (O_608,N_24880,N_24625);
and UO_609 (O_609,N_24692,N_24818);
and UO_610 (O_610,N_24838,N_24540);
xor UO_611 (O_611,N_24654,N_24474);
nor UO_612 (O_612,N_24545,N_24799);
xnor UO_613 (O_613,N_24798,N_24948);
or UO_614 (O_614,N_24505,N_24906);
xnor UO_615 (O_615,N_24806,N_24881);
xnor UO_616 (O_616,N_24731,N_24817);
and UO_617 (O_617,N_24893,N_24997);
or UO_618 (O_618,N_24598,N_24696);
or UO_619 (O_619,N_24676,N_24666);
xnor UO_620 (O_620,N_24976,N_24627);
or UO_621 (O_621,N_24914,N_24375);
xnor UO_622 (O_622,N_24792,N_24469);
xor UO_623 (O_623,N_24635,N_24849);
nand UO_624 (O_624,N_24692,N_24380);
or UO_625 (O_625,N_24629,N_24731);
nor UO_626 (O_626,N_24884,N_24565);
or UO_627 (O_627,N_24728,N_24679);
nand UO_628 (O_628,N_24527,N_24780);
and UO_629 (O_629,N_24895,N_24872);
nor UO_630 (O_630,N_24615,N_24975);
nand UO_631 (O_631,N_24525,N_24629);
or UO_632 (O_632,N_24907,N_24863);
nor UO_633 (O_633,N_24380,N_24490);
xnor UO_634 (O_634,N_24820,N_24524);
or UO_635 (O_635,N_24460,N_24754);
nor UO_636 (O_636,N_24957,N_24507);
nand UO_637 (O_637,N_24706,N_24666);
nand UO_638 (O_638,N_24681,N_24930);
nor UO_639 (O_639,N_24516,N_24762);
nand UO_640 (O_640,N_24673,N_24713);
nor UO_641 (O_641,N_24690,N_24537);
or UO_642 (O_642,N_24383,N_24505);
nand UO_643 (O_643,N_24391,N_24652);
nor UO_644 (O_644,N_24652,N_24477);
or UO_645 (O_645,N_24520,N_24858);
and UO_646 (O_646,N_24380,N_24387);
or UO_647 (O_647,N_24390,N_24910);
or UO_648 (O_648,N_24955,N_24383);
nand UO_649 (O_649,N_24586,N_24874);
nand UO_650 (O_650,N_24968,N_24685);
nand UO_651 (O_651,N_24641,N_24704);
or UO_652 (O_652,N_24413,N_24711);
and UO_653 (O_653,N_24471,N_24793);
nand UO_654 (O_654,N_24864,N_24887);
nor UO_655 (O_655,N_24967,N_24484);
or UO_656 (O_656,N_24489,N_24990);
xnor UO_657 (O_657,N_24803,N_24463);
xnor UO_658 (O_658,N_24419,N_24949);
and UO_659 (O_659,N_24725,N_24622);
and UO_660 (O_660,N_24751,N_24909);
nand UO_661 (O_661,N_24718,N_24770);
nor UO_662 (O_662,N_24656,N_24818);
xor UO_663 (O_663,N_24811,N_24651);
nand UO_664 (O_664,N_24607,N_24467);
or UO_665 (O_665,N_24605,N_24655);
nand UO_666 (O_666,N_24545,N_24817);
nand UO_667 (O_667,N_24669,N_24682);
nor UO_668 (O_668,N_24539,N_24923);
xnor UO_669 (O_669,N_24954,N_24392);
xor UO_670 (O_670,N_24811,N_24498);
or UO_671 (O_671,N_24659,N_24417);
nand UO_672 (O_672,N_24908,N_24927);
nand UO_673 (O_673,N_24583,N_24494);
xnor UO_674 (O_674,N_24823,N_24883);
or UO_675 (O_675,N_24772,N_24821);
nor UO_676 (O_676,N_24455,N_24592);
xnor UO_677 (O_677,N_24759,N_24848);
or UO_678 (O_678,N_24637,N_24977);
nor UO_679 (O_679,N_24539,N_24740);
or UO_680 (O_680,N_24548,N_24680);
nand UO_681 (O_681,N_24462,N_24677);
or UO_682 (O_682,N_24435,N_24724);
and UO_683 (O_683,N_24685,N_24547);
or UO_684 (O_684,N_24763,N_24615);
nand UO_685 (O_685,N_24727,N_24397);
or UO_686 (O_686,N_24588,N_24572);
nand UO_687 (O_687,N_24477,N_24608);
or UO_688 (O_688,N_24842,N_24474);
nor UO_689 (O_689,N_24570,N_24449);
nor UO_690 (O_690,N_24713,N_24671);
and UO_691 (O_691,N_24586,N_24549);
nor UO_692 (O_692,N_24909,N_24991);
xor UO_693 (O_693,N_24958,N_24613);
nor UO_694 (O_694,N_24569,N_24494);
xor UO_695 (O_695,N_24736,N_24591);
xor UO_696 (O_696,N_24972,N_24580);
xor UO_697 (O_697,N_24458,N_24630);
nor UO_698 (O_698,N_24650,N_24518);
nand UO_699 (O_699,N_24947,N_24715);
nor UO_700 (O_700,N_24867,N_24543);
and UO_701 (O_701,N_24721,N_24520);
and UO_702 (O_702,N_24614,N_24775);
nor UO_703 (O_703,N_24998,N_24460);
and UO_704 (O_704,N_24410,N_24764);
nand UO_705 (O_705,N_24990,N_24778);
and UO_706 (O_706,N_24995,N_24474);
and UO_707 (O_707,N_24613,N_24693);
or UO_708 (O_708,N_24773,N_24748);
or UO_709 (O_709,N_24956,N_24993);
and UO_710 (O_710,N_24673,N_24784);
nor UO_711 (O_711,N_24479,N_24934);
or UO_712 (O_712,N_24612,N_24650);
nor UO_713 (O_713,N_24719,N_24995);
or UO_714 (O_714,N_24458,N_24628);
nand UO_715 (O_715,N_24542,N_24478);
nand UO_716 (O_716,N_24852,N_24578);
or UO_717 (O_717,N_24632,N_24967);
nand UO_718 (O_718,N_24786,N_24969);
or UO_719 (O_719,N_24415,N_24686);
and UO_720 (O_720,N_24600,N_24471);
and UO_721 (O_721,N_24382,N_24862);
nor UO_722 (O_722,N_24509,N_24507);
nor UO_723 (O_723,N_24741,N_24467);
or UO_724 (O_724,N_24803,N_24601);
or UO_725 (O_725,N_24685,N_24415);
nor UO_726 (O_726,N_24601,N_24665);
nand UO_727 (O_727,N_24954,N_24473);
or UO_728 (O_728,N_24598,N_24793);
nand UO_729 (O_729,N_24923,N_24840);
and UO_730 (O_730,N_24462,N_24692);
nor UO_731 (O_731,N_24585,N_24903);
nor UO_732 (O_732,N_24898,N_24589);
or UO_733 (O_733,N_24981,N_24407);
or UO_734 (O_734,N_24455,N_24941);
nor UO_735 (O_735,N_24465,N_24571);
nand UO_736 (O_736,N_24644,N_24540);
nand UO_737 (O_737,N_24710,N_24595);
and UO_738 (O_738,N_24865,N_24705);
nor UO_739 (O_739,N_24531,N_24729);
nor UO_740 (O_740,N_24801,N_24424);
and UO_741 (O_741,N_24786,N_24540);
nand UO_742 (O_742,N_24996,N_24472);
or UO_743 (O_743,N_24485,N_24700);
nor UO_744 (O_744,N_24752,N_24889);
or UO_745 (O_745,N_24563,N_24752);
xor UO_746 (O_746,N_24524,N_24718);
nand UO_747 (O_747,N_24429,N_24747);
and UO_748 (O_748,N_24861,N_24416);
or UO_749 (O_749,N_24937,N_24389);
or UO_750 (O_750,N_24590,N_24577);
xnor UO_751 (O_751,N_24973,N_24517);
nor UO_752 (O_752,N_24853,N_24636);
nand UO_753 (O_753,N_24867,N_24645);
nand UO_754 (O_754,N_24679,N_24995);
nand UO_755 (O_755,N_24692,N_24440);
or UO_756 (O_756,N_24567,N_24473);
xnor UO_757 (O_757,N_24702,N_24674);
and UO_758 (O_758,N_24414,N_24919);
nor UO_759 (O_759,N_24521,N_24493);
and UO_760 (O_760,N_24574,N_24679);
and UO_761 (O_761,N_24715,N_24468);
or UO_762 (O_762,N_24849,N_24962);
nand UO_763 (O_763,N_24887,N_24612);
xnor UO_764 (O_764,N_24795,N_24503);
xnor UO_765 (O_765,N_24484,N_24686);
nor UO_766 (O_766,N_24590,N_24855);
xnor UO_767 (O_767,N_24872,N_24984);
nand UO_768 (O_768,N_24487,N_24617);
xor UO_769 (O_769,N_24988,N_24536);
xnor UO_770 (O_770,N_24828,N_24450);
nand UO_771 (O_771,N_24449,N_24698);
xnor UO_772 (O_772,N_24803,N_24517);
and UO_773 (O_773,N_24461,N_24483);
and UO_774 (O_774,N_24495,N_24710);
xnor UO_775 (O_775,N_24573,N_24495);
xnor UO_776 (O_776,N_24916,N_24722);
xnor UO_777 (O_777,N_24840,N_24490);
and UO_778 (O_778,N_24942,N_24438);
and UO_779 (O_779,N_24856,N_24722);
nor UO_780 (O_780,N_24887,N_24999);
or UO_781 (O_781,N_24433,N_24856);
nand UO_782 (O_782,N_24794,N_24914);
nor UO_783 (O_783,N_24877,N_24498);
and UO_784 (O_784,N_24383,N_24899);
nand UO_785 (O_785,N_24425,N_24824);
and UO_786 (O_786,N_24610,N_24817);
nand UO_787 (O_787,N_24766,N_24792);
and UO_788 (O_788,N_24544,N_24534);
nor UO_789 (O_789,N_24775,N_24642);
xnor UO_790 (O_790,N_24377,N_24891);
nor UO_791 (O_791,N_24701,N_24375);
and UO_792 (O_792,N_24886,N_24999);
or UO_793 (O_793,N_24493,N_24804);
xnor UO_794 (O_794,N_24874,N_24404);
or UO_795 (O_795,N_24544,N_24529);
nand UO_796 (O_796,N_24872,N_24845);
xnor UO_797 (O_797,N_24940,N_24931);
xnor UO_798 (O_798,N_24906,N_24522);
xnor UO_799 (O_799,N_24745,N_24866);
nor UO_800 (O_800,N_24909,N_24850);
nor UO_801 (O_801,N_24968,N_24616);
nand UO_802 (O_802,N_24920,N_24864);
nor UO_803 (O_803,N_24884,N_24476);
or UO_804 (O_804,N_24705,N_24879);
xor UO_805 (O_805,N_24386,N_24944);
and UO_806 (O_806,N_24855,N_24501);
and UO_807 (O_807,N_24732,N_24375);
nand UO_808 (O_808,N_24426,N_24754);
nor UO_809 (O_809,N_24880,N_24445);
nor UO_810 (O_810,N_24887,N_24573);
and UO_811 (O_811,N_24572,N_24581);
nor UO_812 (O_812,N_24864,N_24876);
nand UO_813 (O_813,N_24820,N_24696);
xnor UO_814 (O_814,N_24804,N_24715);
nand UO_815 (O_815,N_24820,N_24540);
and UO_816 (O_816,N_24843,N_24862);
xor UO_817 (O_817,N_24930,N_24997);
or UO_818 (O_818,N_24771,N_24661);
nor UO_819 (O_819,N_24684,N_24776);
xnor UO_820 (O_820,N_24971,N_24855);
or UO_821 (O_821,N_24480,N_24993);
xnor UO_822 (O_822,N_24596,N_24815);
and UO_823 (O_823,N_24656,N_24429);
and UO_824 (O_824,N_24956,N_24717);
and UO_825 (O_825,N_24640,N_24945);
or UO_826 (O_826,N_24396,N_24681);
or UO_827 (O_827,N_24946,N_24552);
or UO_828 (O_828,N_24553,N_24752);
and UO_829 (O_829,N_24704,N_24771);
or UO_830 (O_830,N_24964,N_24418);
nand UO_831 (O_831,N_24518,N_24450);
nand UO_832 (O_832,N_24628,N_24402);
or UO_833 (O_833,N_24748,N_24670);
or UO_834 (O_834,N_24819,N_24979);
or UO_835 (O_835,N_24898,N_24484);
nor UO_836 (O_836,N_24814,N_24603);
and UO_837 (O_837,N_24696,N_24736);
nor UO_838 (O_838,N_24636,N_24753);
nand UO_839 (O_839,N_24988,N_24952);
xor UO_840 (O_840,N_24615,N_24597);
and UO_841 (O_841,N_24902,N_24393);
nand UO_842 (O_842,N_24956,N_24768);
xor UO_843 (O_843,N_24587,N_24391);
xnor UO_844 (O_844,N_24518,N_24736);
and UO_845 (O_845,N_24552,N_24649);
and UO_846 (O_846,N_24602,N_24677);
nand UO_847 (O_847,N_24482,N_24622);
xor UO_848 (O_848,N_24804,N_24592);
nor UO_849 (O_849,N_24828,N_24703);
nand UO_850 (O_850,N_24674,N_24882);
nand UO_851 (O_851,N_24433,N_24494);
or UO_852 (O_852,N_24857,N_24382);
nand UO_853 (O_853,N_24518,N_24946);
nor UO_854 (O_854,N_24556,N_24901);
or UO_855 (O_855,N_24479,N_24772);
or UO_856 (O_856,N_24454,N_24758);
nand UO_857 (O_857,N_24706,N_24451);
and UO_858 (O_858,N_24430,N_24427);
nor UO_859 (O_859,N_24519,N_24509);
nand UO_860 (O_860,N_24594,N_24782);
and UO_861 (O_861,N_24899,N_24639);
nor UO_862 (O_862,N_24526,N_24485);
nand UO_863 (O_863,N_24474,N_24603);
or UO_864 (O_864,N_24562,N_24474);
xor UO_865 (O_865,N_24414,N_24438);
nor UO_866 (O_866,N_24885,N_24448);
or UO_867 (O_867,N_24629,N_24835);
xnor UO_868 (O_868,N_24799,N_24677);
nor UO_869 (O_869,N_24524,N_24993);
and UO_870 (O_870,N_24573,N_24486);
or UO_871 (O_871,N_24466,N_24527);
xor UO_872 (O_872,N_24838,N_24652);
nor UO_873 (O_873,N_24429,N_24778);
or UO_874 (O_874,N_24920,N_24745);
xnor UO_875 (O_875,N_24535,N_24685);
nor UO_876 (O_876,N_24795,N_24414);
xor UO_877 (O_877,N_24650,N_24541);
nand UO_878 (O_878,N_24554,N_24572);
or UO_879 (O_879,N_24780,N_24526);
and UO_880 (O_880,N_24892,N_24944);
and UO_881 (O_881,N_24414,N_24471);
xor UO_882 (O_882,N_24646,N_24820);
and UO_883 (O_883,N_24942,N_24480);
nand UO_884 (O_884,N_24945,N_24560);
and UO_885 (O_885,N_24789,N_24831);
or UO_886 (O_886,N_24498,N_24483);
xnor UO_887 (O_887,N_24843,N_24928);
and UO_888 (O_888,N_24412,N_24781);
nand UO_889 (O_889,N_24776,N_24849);
xnor UO_890 (O_890,N_24852,N_24394);
xnor UO_891 (O_891,N_24853,N_24523);
xor UO_892 (O_892,N_24642,N_24558);
nand UO_893 (O_893,N_24734,N_24508);
xnor UO_894 (O_894,N_24623,N_24718);
nor UO_895 (O_895,N_24394,N_24726);
nand UO_896 (O_896,N_24664,N_24752);
xor UO_897 (O_897,N_24487,N_24508);
xor UO_898 (O_898,N_24805,N_24539);
and UO_899 (O_899,N_24562,N_24875);
nand UO_900 (O_900,N_24916,N_24831);
xor UO_901 (O_901,N_24608,N_24472);
nor UO_902 (O_902,N_24972,N_24622);
and UO_903 (O_903,N_24933,N_24433);
nor UO_904 (O_904,N_24609,N_24424);
and UO_905 (O_905,N_24893,N_24524);
xor UO_906 (O_906,N_24641,N_24946);
or UO_907 (O_907,N_24601,N_24878);
nand UO_908 (O_908,N_24469,N_24892);
or UO_909 (O_909,N_24393,N_24708);
nand UO_910 (O_910,N_24554,N_24412);
and UO_911 (O_911,N_24537,N_24971);
xor UO_912 (O_912,N_24882,N_24473);
nand UO_913 (O_913,N_24580,N_24626);
nand UO_914 (O_914,N_24423,N_24629);
xnor UO_915 (O_915,N_24519,N_24489);
or UO_916 (O_916,N_24401,N_24565);
and UO_917 (O_917,N_24611,N_24401);
xnor UO_918 (O_918,N_24874,N_24800);
nor UO_919 (O_919,N_24408,N_24880);
xnor UO_920 (O_920,N_24722,N_24599);
and UO_921 (O_921,N_24614,N_24527);
xnor UO_922 (O_922,N_24378,N_24475);
xor UO_923 (O_923,N_24981,N_24583);
and UO_924 (O_924,N_24776,N_24702);
or UO_925 (O_925,N_24707,N_24683);
or UO_926 (O_926,N_24633,N_24833);
xor UO_927 (O_927,N_24811,N_24603);
xor UO_928 (O_928,N_24888,N_24395);
nand UO_929 (O_929,N_24692,N_24972);
nor UO_930 (O_930,N_24524,N_24438);
or UO_931 (O_931,N_24643,N_24859);
nand UO_932 (O_932,N_24448,N_24565);
nand UO_933 (O_933,N_24685,N_24798);
nand UO_934 (O_934,N_24727,N_24806);
nand UO_935 (O_935,N_24457,N_24637);
xnor UO_936 (O_936,N_24688,N_24642);
nand UO_937 (O_937,N_24468,N_24637);
or UO_938 (O_938,N_24838,N_24786);
nand UO_939 (O_939,N_24409,N_24385);
nand UO_940 (O_940,N_24592,N_24816);
xor UO_941 (O_941,N_24417,N_24565);
xor UO_942 (O_942,N_24816,N_24496);
or UO_943 (O_943,N_24747,N_24633);
nand UO_944 (O_944,N_24808,N_24949);
xnor UO_945 (O_945,N_24418,N_24945);
and UO_946 (O_946,N_24903,N_24626);
xnor UO_947 (O_947,N_24937,N_24970);
xor UO_948 (O_948,N_24403,N_24665);
or UO_949 (O_949,N_24441,N_24408);
and UO_950 (O_950,N_24990,N_24947);
or UO_951 (O_951,N_24811,N_24786);
nand UO_952 (O_952,N_24605,N_24946);
and UO_953 (O_953,N_24505,N_24803);
nor UO_954 (O_954,N_24698,N_24869);
xor UO_955 (O_955,N_24647,N_24907);
xor UO_956 (O_956,N_24645,N_24378);
and UO_957 (O_957,N_24947,N_24509);
nor UO_958 (O_958,N_24858,N_24612);
or UO_959 (O_959,N_24645,N_24623);
nand UO_960 (O_960,N_24740,N_24765);
and UO_961 (O_961,N_24551,N_24387);
or UO_962 (O_962,N_24426,N_24954);
nor UO_963 (O_963,N_24786,N_24686);
nor UO_964 (O_964,N_24731,N_24466);
xnor UO_965 (O_965,N_24862,N_24593);
or UO_966 (O_966,N_24775,N_24791);
or UO_967 (O_967,N_24691,N_24731);
and UO_968 (O_968,N_24377,N_24733);
nor UO_969 (O_969,N_24575,N_24826);
or UO_970 (O_970,N_24479,N_24961);
nor UO_971 (O_971,N_24421,N_24464);
or UO_972 (O_972,N_24594,N_24615);
nor UO_973 (O_973,N_24388,N_24984);
nand UO_974 (O_974,N_24966,N_24947);
and UO_975 (O_975,N_24603,N_24804);
nand UO_976 (O_976,N_24613,N_24766);
and UO_977 (O_977,N_24594,N_24882);
nor UO_978 (O_978,N_24486,N_24549);
nor UO_979 (O_979,N_24904,N_24852);
xnor UO_980 (O_980,N_24934,N_24430);
and UO_981 (O_981,N_24513,N_24934);
and UO_982 (O_982,N_24608,N_24884);
or UO_983 (O_983,N_24979,N_24619);
nand UO_984 (O_984,N_24991,N_24375);
xor UO_985 (O_985,N_24629,N_24474);
nand UO_986 (O_986,N_24942,N_24630);
and UO_987 (O_987,N_24422,N_24654);
or UO_988 (O_988,N_24402,N_24752);
or UO_989 (O_989,N_24754,N_24858);
nand UO_990 (O_990,N_24766,N_24503);
nand UO_991 (O_991,N_24683,N_24689);
xor UO_992 (O_992,N_24702,N_24939);
xor UO_993 (O_993,N_24632,N_24979);
or UO_994 (O_994,N_24583,N_24798);
or UO_995 (O_995,N_24397,N_24842);
or UO_996 (O_996,N_24604,N_24842);
and UO_997 (O_997,N_24585,N_24918);
nand UO_998 (O_998,N_24717,N_24840);
xor UO_999 (O_999,N_24809,N_24803);
and UO_1000 (O_1000,N_24985,N_24514);
and UO_1001 (O_1001,N_24993,N_24649);
and UO_1002 (O_1002,N_24401,N_24512);
xnor UO_1003 (O_1003,N_24415,N_24789);
xor UO_1004 (O_1004,N_24627,N_24565);
xor UO_1005 (O_1005,N_24662,N_24827);
or UO_1006 (O_1006,N_24426,N_24592);
xor UO_1007 (O_1007,N_24375,N_24864);
xnor UO_1008 (O_1008,N_24500,N_24979);
nand UO_1009 (O_1009,N_24984,N_24836);
nor UO_1010 (O_1010,N_24708,N_24538);
xor UO_1011 (O_1011,N_24618,N_24375);
xnor UO_1012 (O_1012,N_24500,N_24382);
or UO_1013 (O_1013,N_24893,N_24772);
nand UO_1014 (O_1014,N_24711,N_24638);
or UO_1015 (O_1015,N_24611,N_24853);
or UO_1016 (O_1016,N_24411,N_24415);
or UO_1017 (O_1017,N_24793,N_24997);
nand UO_1018 (O_1018,N_24927,N_24582);
and UO_1019 (O_1019,N_24693,N_24570);
nand UO_1020 (O_1020,N_24484,N_24637);
and UO_1021 (O_1021,N_24802,N_24597);
nand UO_1022 (O_1022,N_24747,N_24930);
xnor UO_1023 (O_1023,N_24759,N_24818);
nor UO_1024 (O_1024,N_24612,N_24835);
or UO_1025 (O_1025,N_24429,N_24466);
nor UO_1026 (O_1026,N_24913,N_24676);
xnor UO_1027 (O_1027,N_24735,N_24479);
nor UO_1028 (O_1028,N_24505,N_24945);
nand UO_1029 (O_1029,N_24476,N_24752);
or UO_1030 (O_1030,N_24671,N_24910);
xor UO_1031 (O_1031,N_24741,N_24489);
or UO_1032 (O_1032,N_24509,N_24923);
or UO_1033 (O_1033,N_24381,N_24697);
nand UO_1034 (O_1034,N_24765,N_24683);
xnor UO_1035 (O_1035,N_24434,N_24539);
and UO_1036 (O_1036,N_24905,N_24782);
and UO_1037 (O_1037,N_24424,N_24717);
or UO_1038 (O_1038,N_24533,N_24474);
or UO_1039 (O_1039,N_24418,N_24870);
xor UO_1040 (O_1040,N_24748,N_24712);
or UO_1041 (O_1041,N_24978,N_24516);
nor UO_1042 (O_1042,N_24828,N_24915);
or UO_1043 (O_1043,N_24931,N_24630);
or UO_1044 (O_1044,N_24711,N_24810);
xor UO_1045 (O_1045,N_24441,N_24798);
and UO_1046 (O_1046,N_24640,N_24404);
and UO_1047 (O_1047,N_24454,N_24408);
or UO_1048 (O_1048,N_24672,N_24405);
xor UO_1049 (O_1049,N_24870,N_24452);
nand UO_1050 (O_1050,N_24746,N_24532);
xor UO_1051 (O_1051,N_24695,N_24492);
nand UO_1052 (O_1052,N_24689,N_24866);
xnor UO_1053 (O_1053,N_24442,N_24497);
or UO_1054 (O_1054,N_24965,N_24597);
nand UO_1055 (O_1055,N_24920,N_24874);
and UO_1056 (O_1056,N_24751,N_24375);
xor UO_1057 (O_1057,N_24882,N_24696);
nand UO_1058 (O_1058,N_24888,N_24779);
or UO_1059 (O_1059,N_24831,N_24403);
and UO_1060 (O_1060,N_24677,N_24555);
and UO_1061 (O_1061,N_24837,N_24440);
and UO_1062 (O_1062,N_24978,N_24718);
and UO_1063 (O_1063,N_24544,N_24968);
xnor UO_1064 (O_1064,N_24852,N_24559);
or UO_1065 (O_1065,N_24716,N_24732);
nand UO_1066 (O_1066,N_24752,N_24917);
and UO_1067 (O_1067,N_24493,N_24615);
nor UO_1068 (O_1068,N_24625,N_24673);
nor UO_1069 (O_1069,N_24820,N_24853);
or UO_1070 (O_1070,N_24420,N_24837);
nor UO_1071 (O_1071,N_24919,N_24689);
and UO_1072 (O_1072,N_24650,N_24813);
nand UO_1073 (O_1073,N_24525,N_24541);
nand UO_1074 (O_1074,N_24645,N_24862);
nand UO_1075 (O_1075,N_24596,N_24793);
nand UO_1076 (O_1076,N_24724,N_24929);
and UO_1077 (O_1077,N_24441,N_24724);
or UO_1078 (O_1078,N_24581,N_24695);
nor UO_1079 (O_1079,N_24668,N_24549);
nand UO_1080 (O_1080,N_24968,N_24902);
nand UO_1081 (O_1081,N_24935,N_24792);
or UO_1082 (O_1082,N_24488,N_24970);
xor UO_1083 (O_1083,N_24650,N_24831);
nand UO_1084 (O_1084,N_24887,N_24401);
and UO_1085 (O_1085,N_24899,N_24864);
nand UO_1086 (O_1086,N_24445,N_24988);
xor UO_1087 (O_1087,N_24708,N_24968);
nand UO_1088 (O_1088,N_24981,N_24712);
nor UO_1089 (O_1089,N_24777,N_24411);
and UO_1090 (O_1090,N_24501,N_24585);
or UO_1091 (O_1091,N_24753,N_24601);
and UO_1092 (O_1092,N_24625,N_24968);
and UO_1093 (O_1093,N_24457,N_24730);
nor UO_1094 (O_1094,N_24424,N_24912);
nand UO_1095 (O_1095,N_24865,N_24890);
xnor UO_1096 (O_1096,N_24615,N_24781);
or UO_1097 (O_1097,N_24516,N_24810);
xnor UO_1098 (O_1098,N_24380,N_24887);
or UO_1099 (O_1099,N_24534,N_24621);
nand UO_1100 (O_1100,N_24604,N_24800);
and UO_1101 (O_1101,N_24985,N_24829);
nand UO_1102 (O_1102,N_24887,N_24395);
xor UO_1103 (O_1103,N_24764,N_24979);
or UO_1104 (O_1104,N_24713,N_24430);
or UO_1105 (O_1105,N_24468,N_24532);
or UO_1106 (O_1106,N_24763,N_24421);
or UO_1107 (O_1107,N_24727,N_24421);
nand UO_1108 (O_1108,N_24900,N_24990);
and UO_1109 (O_1109,N_24604,N_24705);
xor UO_1110 (O_1110,N_24417,N_24509);
nor UO_1111 (O_1111,N_24917,N_24781);
or UO_1112 (O_1112,N_24689,N_24841);
or UO_1113 (O_1113,N_24818,N_24801);
and UO_1114 (O_1114,N_24790,N_24495);
nor UO_1115 (O_1115,N_24497,N_24473);
xnor UO_1116 (O_1116,N_24895,N_24656);
xor UO_1117 (O_1117,N_24451,N_24610);
xor UO_1118 (O_1118,N_24573,N_24688);
nand UO_1119 (O_1119,N_24723,N_24871);
nand UO_1120 (O_1120,N_24719,N_24569);
xor UO_1121 (O_1121,N_24584,N_24904);
nor UO_1122 (O_1122,N_24947,N_24468);
nand UO_1123 (O_1123,N_24655,N_24705);
nor UO_1124 (O_1124,N_24490,N_24594);
xor UO_1125 (O_1125,N_24933,N_24707);
and UO_1126 (O_1126,N_24562,N_24624);
nand UO_1127 (O_1127,N_24581,N_24378);
nor UO_1128 (O_1128,N_24915,N_24553);
nor UO_1129 (O_1129,N_24683,N_24432);
nand UO_1130 (O_1130,N_24697,N_24541);
nand UO_1131 (O_1131,N_24568,N_24569);
or UO_1132 (O_1132,N_24627,N_24490);
and UO_1133 (O_1133,N_24887,N_24952);
and UO_1134 (O_1134,N_24868,N_24546);
nor UO_1135 (O_1135,N_24482,N_24902);
nand UO_1136 (O_1136,N_24796,N_24810);
and UO_1137 (O_1137,N_24392,N_24654);
or UO_1138 (O_1138,N_24907,N_24739);
nor UO_1139 (O_1139,N_24563,N_24955);
xor UO_1140 (O_1140,N_24452,N_24795);
and UO_1141 (O_1141,N_24633,N_24782);
or UO_1142 (O_1142,N_24627,N_24470);
xnor UO_1143 (O_1143,N_24640,N_24873);
xnor UO_1144 (O_1144,N_24568,N_24566);
and UO_1145 (O_1145,N_24599,N_24387);
nand UO_1146 (O_1146,N_24643,N_24783);
nand UO_1147 (O_1147,N_24985,N_24710);
and UO_1148 (O_1148,N_24508,N_24980);
and UO_1149 (O_1149,N_24881,N_24468);
xnor UO_1150 (O_1150,N_24891,N_24801);
xnor UO_1151 (O_1151,N_24806,N_24694);
nand UO_1152 (O_1152,N_24379,N_24545);
xnor UO_1153 (O_1153,N_24545,N_24514);
or UO_1154 (O_1154,N_24676,N_24514);
and UO_1155 (O_1155,N_24437,N_24665);
and UO_1156 (O_1156,N_24408,N_24491);
nand UO_1157 (O_1157,N_24841,N_24428);
xor UO_1158 (O_1158,N_24690,N_24902);
nand UO_1159 (O_1159,N_24803,N_24419);
nand UO_1160 (O_1160,N_24731,N_24827);
xnor UO_1161 (O_1161,N_24720,N_24551);
or UO_1162 (O_1162,N_24843,N_24848);
nand UO_1163 (O_1163,N_24926,N_24768);
and UO_1164 (O_1164,N_24801,N_24616);
xor UO_1165 (O_1165,N_24845,N_24505);
xor UO_1166 (O_1166,N_24473,N_24825);
and UO_1167 (O_1167,N_24953,N_24522);
nor UO_1168 (O_1168,N_24706,N_24973);
or UO_1169 (O_1169,N_24783,N_24740);
or UO_1170 (O_1170,N_24650,N_24495);
nor UO_1171 (O_1171,N_24469,N_24411);
nor UO_1172 (O_1172,N_24632,N_24500);
nand UO_1173 (O_1173,N_24924,N_24928);
nand UO_1174 (O_1174,N_24409,N_24597);
xor UO_1175 (O_1175,N_24923,N_24947);
nand UO_1176 (O_1176,N_24661,N_24967);
nor UO_1177 (O_1177,N_24862,N_24423);
xnor UO_1178 (O_1178,N_24970,N_24405);
or UO_1179 (O_1179,N_24762,N_24513);
nor UO_1180 (O_1180,N_24880,N_24775);
xnor UO_1181 (O_1181,N_24396,N_24636);
nor UO_1182 (O_1182,N_24903,N_24717);
nand UO_1183 (O_1183,N_24456,N_24518);
xor UO_1184 (O_1184,N_24865,N_24918);
nor UO_1185 (O_1185,N_24888,N_24638);
nor UO_1186 (O_1186,N_24887,N_24695);
nor UO_1187 (O_1187,N_24399,N_24508);
nor UO_1188 (O_1188,N_24821,N_24885);
nand UO_1189 (O_1189,N_24929,N_24404);
nand UO_1190 (O_1190,N_24799,N_24790);
xor UO_1191 (O_1191,N_24880,N_24457);
nand UO_1192 (O_1192,N_24487,N_24385);
nand UO_1193 (O_1193,N_24484,N_24442);
and UO_1194 (O_1194,N_24734,N_24548);
nand UO_1195 (O_1195,N_24572,N_24486);
nand UO_1196 (O_1196,N_24562,N_24742);
nor UO_1197 (O_1197,N_24623,N_24577);
and UO_1198 (O_1198,N_24487,N_24519);
and UO_1199 (O_1199,N_24684,N_24900);
xnor UO_1200 (O_1200,N_24435,N_24834);
nor UO_1201 (O_1201,N_24785,N_24786);
and UO_1202 (O_1202,N_24380,N_24395);
xnor UO_1203 (O_1203,N_24909,N_24972);
nand UO_1204 (O_1204,N_24617,N_24663);
and UO_1205 (O_1205,N_24929,N_24499);
xor UO_1206 (O_1206,N_24395,N_24482);
and UO_1207 (O_1207,N_24992,N_24847);
xnor UO_1208 (O_1208,N_24565,N_24507);
or UO_1209 (O_1209,N_24817,N_24880);
or UO_1210 (O_1210,N_24922,N_24564);
and UO_1211 (O_1211,N_24442,N_24676);
nor UO_1212 (O_1212,N_24423,N_24656);
and UO_1213 (O_1213,N_24411,N_24878);
xor UO_1214 (O_1214,N_24500,N_24523);
xor UO_1215 (O_1215,N_24443,N_24661);
nand UO_1216 (O_1216,N_24522,N_24809);
nand UO_1217 (O_1217,N_24490,N_24497);
xor UO_1218 (O_1218,N_24827,N_24376);
or UO_1219 (O_1219,N_24737,N_24539);
and UO_1220 (O_1220,N_24650,N_24721);
nor UO_1221 (O_1221,N_24378,N_24412);
nand UO_1222 (O_1222,N_24821,N_24450);
or UO_1223 (O_1223,N_24420,N_24782);
xnor UO_1224 (O_1224,N_24816,N_24952);
nor UO_1225 (O_1225,N_24962,N_24882);
xor UO_1226 (O_1226,N_24723,N_24412);
nand UO_1227 (O_1227,N_24601,N_24842);
or UO_1228 (O_1228,N_24847,N_24799);
or UO_1229 (O_1229,N_24499,N_24483);
nor UO_1230 (O_1230,N_24441,N_24640);
or UO_1231 (O_1231,N_24520,N_24855);
nor UO_1232 (O_1232,N_24891,N_24647);
nand UO_1233 (O_1233,N_24938,N_24509);
or UO_1234 (O_1234,N_24489,N_24797);
nor UO_1235 (O_1235,N_24817,N_24807);
xnor UO_1236 (O_1236,N_24909,N_24726);
nor UO_1237 (O_1237,N_24606,N_24821);
xor UO_1238 (O_1238,N_24865,N_24619);
and UO_1239 (O_1239,N_24911,N_24871);
nor UO_1240 (O_1240,N_24503,N_24575);
or UO_1241 (O_1241,N_24525,N_24691);
nand UO_1242 (O_1242,N_24885,N_24931);
and UO_1243 (O_1243,N_24908,N_24833);
nor UO_1244 (O_1244,N_24715,N_24767);
nand UO_1245 (O_1245,N_24917,N_24585);
or UO_1246 (O_1246,N_24508,N_24663);
nand UO_1247 (O_1247,N_24377,N_24722);
nor UO_1248 (O_1248,N_24988,N_24815);
xor UO_1249 (O_1249,N_24577,N_24732);
nor UO_1250 (O_1250,N_24996,N_24391);
nand UO_1251 (O_1251,N_24413,N_24850);
nand UO_1252 (O_1252,N_24454,N_24517);
xor UO_1253 (O_1253,N_24831,N_24385);
nand UO_1254 (O_1254,N_24722,N_24780);
xor UO_1255 (O_1255,N_24414,N_24673);
and UO_1256 (O_1256,N_24803,N_24975);
or UO_1257 (O_1257,N_24822,N_24747);
nor UO_1258 (O_1258,N_24885,N_24851);
nor UO_1259 (O_1259,N_24609,N_24818);
xnor UO_1260 (O_1260,N_24808,N_24640);
xnor UO_1261 (O_1261,N_24411,N_24488);
nand UO_1262 (O_1262,N_24827,N_24471);
and UO_1263 (O_1263,N_24748,N_24864);
xnor UO_1264 (O_1264,N_24746,N_24490);
nor UO_1265 (O_1265,N_24428,N_24468);
and UO_1266 (O_1266,N_24775,N_24589);
or UO_1267 (O_1267,N_24884,N_24650);
or UO_1268 (O_1268,N_24698,N_24582);
or UO_1269 (O_1269,N_24413,N_24379);
nand UO_1270 (O_1270,N_24953,N_24662);
nor UO_1271 (O_1271,N_24995,N_24559);
nand UO_1272 (O_1272,N_24785,N_24934);
nor UO_1273 (O_1273,N_24862,N_24883);
nand UO_1274 (O_1274,N_24611,N_24897);
and UO_1275 (O_1275,N_24810,N_24809);
nand UO_1276 (O_1276,N_24878,N_24958);
nor UO_1277 (O_1277,N_24787,N_24871);
nor UO_1278 (O_1278,N_24889,N_24724);
nor UO_1279 (O_1279,N_24851,N_24814);
xnor UO_1280 (O_1280,N_24529,N_24427);
or UO_1281 (O_1281,N_24628,N_24730);
and UO_1282 (O_1282,N_24479,N_24869);
nand UO_1283 (O_1283,N_24492,N_24938);
xor UO_1284 (O_1284,N_24964,N_24440);
nand UO_1285 (O_1285,N_24682,N_24899);
nor UO_1286 (O_1286,N_24931,N_24483);
xnor UO_1287 (O_1287,N_24688,N_24968);
xor UO_1288 (O_1288,N_24523,N_24705);
and UO_1289 (O_1289,N_24570,N_24486);
nor UO_1290 (O_1290,N_24701,N_24513);
and UO_1291 (O_1291,N_24531,N_24720);
and UO_1292 (O_1292,N_24969,N_24811);
and UO_1293 (O_1293,N_24560,N_24595);
nand UO_1294 (O_1294,N_24918,N_24662);
nand UO_1295 (O_1295,N_24631,N_24895);
or UO_1296 (O_1296,N_24980,N_24740);
nand UO_1297 (O_1297,N_24435,N_24894);
nor UO_1298 (O_1298,N_24634,N_24423);
nand UO_1299 (O_1299,N_24782,N_24966);
or UO_1300 (O_1300,N_24396,N_24497);
nor UO_1301 (O_1301,N_24659,N_24611);
and UO_1302 (O_1302,N_24775,N_24433);
nor UO_1303 (O_1303,N_24403,N_24724);
or UO_1304 (O_1304,N_24999,N_24775);
nor UO_1305 (O_1305,N_24820,N_24414);
xnor UO_1306 (O_1306,N_24934,N_24552);
xor UO_1307 (O_1307,N_24768,N_24896);
nand UO_1308 (O_1308,N_24647,N_24777);
nor UO_1309 (O_1309,N_24808,N_24889);
or UO_1310 (O_1310,N_24730,N_24912);
or UO_1311 (O_1311,N_24871,N_24955);
and UO_1312 (O_1312,N_24577,N_24678);
and UO_1313 (O_1313,N_24995,N_24429);
nor UO_1314 (O_1314,N_24879,N_24631);
or UO_1315 (O_1315,N_24701,N_24526);
nand UO_1316 (O_1316,N_24508,N_24469);
nor UO_1317 (O_1317,N_24554,N_24439);
xor UO_1318 (O_1318,N_24695,N_24609);
nor UO_1319 (O_1319,N_24510,N_24796);
nor UO_1320 (O_1320,N_24766,N_24519);
xnor UO_1321 (O_1321,N_24664,N_24974);
or UO_1322 (O_1322,N_24731,N_24867);
nand UO_1323 (O_1323,N_24487,N_24941);
nand UO_1324 (O_1324,N_24682,N_24860);
nand UO_1325 (O_1325,N_24998,N_24448);
xnor UO_1326 (O_1326,N_24717,N_24712);
nand UO_1327 (O_1327,N_24635,N_24681);
and UO_1328 (O_1328,N_24603,N_24925);
nand UO_1329 (O_1329,N_24390,N_24392);
nor UO_1330 (O_1330,N_24637,N_24577);
nand UO_1331 (O_1331,N_24388,N_24593);
nand UO_1332 (O_1332,N_24536,N_24602);
and UO_1333 (O_1333,N_24907,N_24745);
or UO_1334 (O_1334,N_24388,N_24983);
and UO_1335 (O_1335,N_24810,N_24477);
xnor UO_1336 (O_1336,N_24404,N_24968);
or UO_1337 (O_1337,N_24720,N_24702);
or UO_1338 (O_1338,N_24877,N_24607);
nand UO_1339 (O_1339,N_24526,N_24551);
xor UO_1340 (O_1340,N_24924,N_24453);
nand UO_1341 (O_1341,N_24901,N_24752);
nand UO_1342 (O_1342,N_24443,N_24510);
and UO_1343 (O_1343,N_24480,N_24755);
xnor UO_1344 (O_1344,N_24738,N_24467);
nand UO_1345 (O_1345,N_24610,N_24811);
nand UO_1346 (O_1346,N_24723,N_24853);
and UO_1347 (O_1347,N_24582,N_24585);
nand UO_1348 (O_1348,N_24879,N_24841);
nor UO_1349 (O_1349,N_24708,N_24851);
and UO_1350 (O_1350,N_24666,N_24730);
nand UO_1351 (O_1351,N_24897,N_24714);
nand UO_1352 (O_1352,N_24950,N_24574);
nand UO_1353 (O_1353,N_24716,N_24990);
or UO_1354 (O_1354,N_24827,N_24710);
xnor UO_1355 (O_1355,N_24956,N_24996);
nor UO_1356 (O_1356,N_24601,N_24589);
nand UO_1357 (O_1357,N_24620,N_24670);
nor UO_1358 (O_1358,N_24965,N_24468);
xor UO_1359 (O_1359,N_24410,N_24872);
nor UO_1360 (O_1360,N_24411,N_24483);
xor UO_1361 (O_1361,N_24540,N_24985);
nand UO_1362 (O_1362,N_24518,N_24854);
and UO_1363 (O_1363,N_24381,N_24775);
or UO_1364 (O_1364,N_24865,N_24759);
nor UO_1365 (O_1365,N_24854,N_24617);
or UO_1366 (O_1366,N_24604,N_24565);
xor UO_1367 (O_1367,N_24547,N_24635);
and UO_1368 (O_1368,N_24601,N_24677);
or UO_1369 (O_1369,N_24548,N_24866);
and UO_1370 (O_1370,N_24894,N_24664);
or UO_1371 (O_1371,N_24704,N_24964);
or UO_1372 (O_1372,N_24431,N_24375);
xor UO_1373 (O_1373,N_24788,N_24437);
nor UO_1374 (O_1374,N_24843,N_24914);
and UO_1375 (O_1375,N_24494,N_24385);
nor UO_1376 (O_1376,N_24481,N_24715);
or UO_1377 (O_1377,N_24858,N_24414);
nor UO_1378 (O_1378,N_24906,N_24417);
and UO_1379 (O_1379,N_24583,N_24899);
or UO_1380 (O_1380,N_24388,N_24728);
nor UO_1381 (O_1381,N_24883,N_24379);
or UO_1382 (O_1382,N_24772,N_24679);
nor UO_1383 (O_1383,N_24428,N_24640);
or UO_1384 (O_1384,N_24504,N_24426);
and UO_1385 (O_1385,N_24980,N_24829);
and UO_1386 (O_1386,N_24586,N_24474);
nor UO_1387 (O_1387,N_24613,N_24727);
or UO_1388 (O_1388,N_24759,N_24807);
xor UO_1389 (O_1389,N_24635,N_24969);
and UO_1390 (O_1390,N_24756,N_24546);
nor UO_1391 (O_1391,N_24990,N_24404);
xnor UO_1392 (O_1392,N_24432,N_24686);
nor UO_1393 (O_1393,N_24624,N_24947);
or UO_1394 (O_1394,N_24853,N_24615);
xor UO_1395 (O_1395,N_24861,N_24954);
nor UO_1396 (O_1396,N_24578,N_24719);
or UO_1397 (O_1397,N_24524,N_24715);
and UO_1398 (O_1398,N_24925,N_24528);
nor UO_1399 (O_1399,N_24418,N_24535);
nand UO_1400 (O_1400,N_24646,N_24383);
nor UO_1401 (O_1401,N_24582,N_24849);
and UO_1402 (O_1402,N_24606,N_24731);
or UO_1403 (O_1403,N_24961,N_24529);
or UO_1404 (O_1404,N_24545,N_24998);
nand UO_1405 (O_1405,N_24844,N_24690);
nor UO_1406 (O_1406,N_24613,N_24649);
nor UO_1407 (O_1407,N_24792,N_24991);
nand UO_1408 (O_1408,N_24528,N_24940);
nand UO_1409 (O_1409,N_24797,N_24865);
xnor UO_1410 (O_1410,N_24554,N_24991);
or UO_1411 (O_1411,N_24867,N_24478);
or UO_1412 (O_1412,N_24902,N_24761);
and UO_1413 (O_1413,N_24447,N_24605);
nand UO_1414 (O_1414,N_24638,N_24662);
nor UO_1415 (O_1415,N_24601,N_24866);
nand UO_1416 (O_1416,N_24527,N_24761);
and UO_1417 (O_1417,N_24743,N_24493);
or UO_1418 (O_1418,N_24385,N_24443);
xor UO_1419 (O_1419,N_24613,N_24927);
or UO_1420 (O_1420,N_24952,N_24831);
nor UO_1421 (O_1421,N_24605,N_24385);
or UO_1422 (O_1422,N_24786,N_24931);
or UO_1423 (O_1423,N_24481,N_24440);
or UO_1424 (O_1424,N_24580,N_24757);
or UO_1425 (O_1425,N_24638,N_24515);
nand UO_1426 (O_1426,N_24755,N_24512);
xor UO_1427 (O_1427,N_24490,N_24414);
nand UO_1428 (O_1428,N_24670,N_24704);
or UO_1429 (O_1429,N_24658,N_24387);
nand UO_1430 (O_1430,N_24925,N_24711);
nor UO_1431 (O_1431,N_24645,N_24982);
or UO_1432 (O_1432,N_24872,N_24443);
xor UO_1433 (O_1433,N_24657,N_24742);
nand UO_1434 (O_1434,N_24567,N_24460);
or UO_1435 (O_1435,N_24902,N_24423);
and UO_1436 (O_1436,N_24801,N_24957);
and UO_1437 (O_1437,N_24747,N_24981);
or UO_1438 (O_1438,N_24973,N_24459);
nand UO_1439 (O_1439,N_24804,N_24974);
and UO_1440 (O_1440,N_24680,N_24854);
and UO_1441 (O_1441,N_24480,N_24627);
and UO_1442 (O_1442,N_24765,N_24837);
and UO_1443 (O_1443,N_24823,N_24895);
or UO_1444 (O_1444,N_24976,N_24745);
nor UO_1445 (O_1445,N_24456,N_24907);
nand UO_1446 (O_1446,N_24588,N_24903);
xnor UO_1447 (O_1447,N_24942,N_24552);
nand UO_1448 (O_1448,N_24646,N_24843);
or UO_1449 (O_1449,N_24829,N_24684);
xnor UO_1450 (O_1450,N_24706,N_24708);
nor UO_1451 (O_1451,N_24740,N_24561);
or UO_1452 (O_1452,N_24909,N_24905);
nand UO_1453 (O_1453,N_24716,N_24992);
nand UO_1454 (O_1454,N_24869,N_24480);
nor UO_1455 (O_1455,N_24519,N_24730);
nor UO_1456 (O_1456,N_24755,N_24667);
nor UO_1457 (O_1457,N_24651,N_24929);
nand UO_1458 (O_1458,N_24941,N_24848);
nand UO_1459 (O_1459,N_24975,N_24950);
or UO_1460 (O_1460,N_24547,N_24732);
xor UO_1461 (O_1461,N_24405,N_24757);
nor UO_1462 (O_1462,N_24432,N_24632);
xnor UO_1463 (O_1463,N_24808,N_24603);
xnor UO_1464 (O_1464,N_24436,N_24848);
nand UO_1465 (O_1465,N_24498,N_24919);
xnor UO_1466 (O_1466,N_24940,N_24782);
nand UO_1467 (O_1467,N_24775,N_24645);
and UO_1468 (O_1468,N_24813,N_24450);
nand UO_1469 (O_1469,N_24887,N_24622);
and UO_1470 (O_1470,N_24527,N_24404);
and UO_1471 (O_1471,N_24637,N_24424);
xnor UO_1472 (O_1472,N_24698,N_24526);
xnor UO_1473 (O_1473,N_24396,N_24884);
and UO_1474 (O_1474,N_24528,N_24871);
nor UO_1475 (O_1475,N_24493,N_24710);
or UO_1476 (O_1476,N_24768,N_24401);
or UO_1477 (O_1477,N_24383,N_24879);
nor UO_1478 (O_1478,N_24429,N_24660);
or UO_1479 (O_1479,N_24679,N_24750);
nand UO_1480 (O_1480,N_24802,N_24539);
nor UO_1481 (O_1481,N_24932,N_24931);
nor UO_1482 (O_1482,N_24420,N_24833);
or UO_1483 (O_1483,N_24436,N_24725);
or UO_1484 (O_1484,N_24811,N_24587);
or UO_1485 (O_1485,N_24777,N_24816);
and UO_1486 (O_1486,N_24848,N_24687);
xor UO_1487 (O_1487,N_24507,N_24682);
and UO_1488 (O_1488,N_24797,N_24571);
nor UO_1489 (O_1489,N_24877,N_24662);
or UO_1490 (O_1490,N_24461,N_24999);
nor UO_1491 (O_1491,N_24925,N_24852);
and UO_1492 (O_1492,N_24732,N_24390);
nor UO_1493 (O_1493,N_24598,N_24847);
nor UO_1494 (O_1494,N_24480,N_24512);
and UO_1495 (O_1495,N_24409,N_24897);
or UO_1496 (O_1496,N_24952,N_24805);
or UO_1497 (O_1497,N_24868,N_24416);
nand UO_1498 (O_1498,N_24625,N_24517);
or UO_1499 (O_1499,N_24595,N_24989);
nand UO_1500 (O_1500,N_24708,N_24893);
nand UO_1501 (O_1501,N_24680,N_24793);
nand UO_1502 (O_1502,N_24900,N_24507);
xor UO_1503 (O_1503,N_24807,N_24895);
nor UO_1504 (O_1504,N_24766,N_24568);
nor UO_1505 (O_1505,N_24887,N_24871);
or UO_1506 (O_1506,N_24684,N_24499);
or UO_1507 (O_1507,N_24395,N_24853);
or UO_1508 (O_1508,N_24971,N_24707);
or UO_1509 (O_1509,N_24782,N_24727);
and UO_1510 (O_1510,N_24721,N_24590);
nand UO_1511 (O_1511,N_24564,N_24770);
nand UO_1512 (O_1512,N_24513,N_24913);
and UO_1513 (O_1513,N_24679,N_24643);
nor UO_1514 (O_1514,N_24429,N_24396);
and UO_1515 (O_1515,N_24860,N_24854);
nand UO_1516 (O_1516,N_24796,N_24553);
nor UO_1517 (O_1517,N_24856,N_24739);
xor UO_1518 (O_1518,N_24461,N_24944);
xnor UO_1519 (O_1519,N_24777,N_24799);
xor UO_1520 (O_1520,N_24780,N_24599);
or UO_1521 (O_1521,N_24946,N_24526);
xnor UO_1522 (O_1522,N_24685,N_24408);
nand UO_1523 (O_1523,N_24830,N_24850);
and UO_1524 (O_1524,N_24420,N_24661);
nand UO_1525 (O_1525,N_24737,N_24449);
or UO_1526 (O_1526,N_24840,N_24442);
and UO_1527 (O_1527,N_24732,N_24608);
nand UO_1528 (O_1528,N_24505,N_24614);
or UO_1529 (O_1529,N_24519,N_24508);
nor UO_1530 (O_1530,N_24577,N_24588);
or UO_1531 (O_1531,N_24990,N_24940);
nand UO_1532 (O_1532,N_24981,N_24598);
or UO_1533 (O_1533,N_24388,N_24592);
and UO_1534 (O_1534,N_24811,N_24805);
xor UO_1535 (O_1535,N_24717,N_24581);
or UO_1536 (O_1536,N_24977,N_24713);
and UO_1537 (O_1537,N_24687,N_24758);
or UO_1538 (O_1538,N_24505,N_24438);
nor UO_1539 (O_1539,N_24452,N_24771);
nor UO_1540 (O_1540,N_24536,N_24489);
xor UO_1541 (O_1541,N_24851,N_24975);
and UO_1542 (O_1542,N_24870,N_24878);
nand UO_1543 (O_1543,N_24908,N_24597);
nand UO_1544 (O_1544,N_24897,N_24523);
nand UO_1545 (O_1545,N_24416,N_24520);
nor UO_1546 (O_1546,N_24480,N_24667);
nor UO_1547 (O_1547,N_24896,N_24828);
or UO_1548 (O_1548,N_24602,N_24613);
and UO_1549 (O_1549,N_24456,N_24780);
xor UO_1550 (O_1550,N_24901,N_24804);
and UO_1551 (O_1551,N_24819,N_24784);
xnor UO_1552 (O_1552,N_24876,N_24534);
or UO_1553 (O_1553,N_24635,N_24944);
xnor UO_1554 (O_1554,N_24978,N_24588);
xor UO_1555 (O_1555,N_24382,N_24916);
nor UO_1556 (O_1556,N_24886,N_24853);
or UO_1557 (O_1557,N_24992,N_24878);
or UO_1558 (O_1558,N_24595,N_24575);
xor UO_1559 (O_1559,N_24856,N_24720);
and UO_1560 (O_1560,N_24839,N_24810);
xnor UO_1561 (O_1561,N_24753,N_24491);
xnor UO_1562 (O_1562,N_24428,N_24928);
nand UO_1563 (O_1563,N_24482,N_24403);
and UO_1564 (O_1564,N_24494,N_24435);
nand UO_1565 (O_1565,N_24420,N_24871);
xnor UO_1566 (O_1566,N_24887,N_24483);
nor UO_1567 (O_1567,N_24896,N_24566);
or UO_1568 (O_1568,N_24657,N_24542);
and UO_1569 (O_1569,N_24434,N_24946);
nor UO_1570 (O_1570,N_24793,N_24995);
nor UO_1571 (O_1571,N_24376,N_24604);
and UO_1572 (O_1572,N_24808,N_24997);
nor UO_1573 (O_1573,N_24714,N_24716);
or UO_1574 (O_1574,N_24825,N_24619);
xor UO_1575 (O_1575,N_24756,N_24867);
nand UO_1576 (O_1576,N_24910,N_24818);
nor UO_1577 (O_1577,N_24814,N_24744);
xnor UO_1578 (O_1578,N_24734,N_24752);
nor UO_1579 (O_1579,N_24680,N_24869);
nor UO_1580 (O_1580,N_24730,N_24458);
or UO_1581 (O_1581,N_24959,N_24768);
nor UO_1582 (O_1582,N_24724,N_24502);
and UO_1583 (O_1583,N_24769,N_24644);
or UO_1584 (O_1584,N_24415,N_24380);
xnor UO_1585 (O_1585,N_24681,N_24434);
and UO_1586 (O_1586,N_24808,N_24708);
nor UO_1587 (O_1587,N_24630,N_24603);
nand UO_1588 (O_1588,N_24603,N_24398);
nor UO_1589 (O_1589,N_24768,N_24637);
nor UO_1590 (O_1590,N_24662,N_24464);
or UO_1591 (O_1591,N_24952,N_24923);
xnor UO_1592 (O_1592,N_24527,N_24403);
nor UO_1593 (O_1593,N_24892,N_24757);
and UO_1594 (O_1594,N_24593,N_24665);
xor UO_1595 (O_1595,N_24850,N_24663);
and UO_1596 (O_1596,N_24550,N_24831);
nor UO_1597 (O_1597,N_24998,N_24948);
or UO_1598 (O_1598,N_24505,N_24566);
nand UO_1599 (O_1599,N_24975,N_24783);
or UO_1600 (O_1600,N_24416,N_24420);
nor UO_1601 (O_1601,N_24691,N_24375);
nor UO_1602 (O_1602,N_24973,N_24426);
and UO_1603 (O_1603,N_24793,N_24650);
xnor UO_1604 (O_1604,N_24496,N_24656);
or UO_1605 (O_1605,N_24647,N_24513);
nor UO_1606 (O_1606,N_24505,N_24888);
nand UO_1607 (O_1607,N_24488,N_24919);
nor UO_1608 (O_1608,N_24712,N_24554);
xnor UO_1609 (O_1609,N_24872,N_24905);
or UO_1610 (O_1610,N_24783,N_24755);
nor UO_1611 (O_1611,N_24905,N_24619);
nand UO_1612 (O_1612,N_24436,N_24586);
or UO_1613 (O_1613,N_24851,N_24829);
or UO_1614 (O_1614,N_24987,N_24504);
and UO_1615 (O_1615,N_24854,N_24415);
xnor UO_1616 (O_1616,N_24683,N_24456);
nand UO_1617 (O_1617,N_24446,N_24790);
xor UO_1618 (O_1618,N_24859,N_24914);
nor UO_1619 (O_1619,N_24669,N_24868);
nor UO_1620 (O_1620,N_24895,N_24842);
and UO_1621 (O_1621,N_24816,N_24603);
or UO_1622 (O_1622,N_24611,N_24644);
xor UO_1623 (O_1623,N_24813,N_24958);
and UO_1624 (O_1624,N_24859,N_24723);
nor UO_1625 (O_1625,N_24390,N_24411);
xnor UO_1626 (O_1626,N_24447,N_24612);
or UO_1627 (O_1627,N_24830,N_24401);
xnor UO_1628 (O_1628,N_24825,N_24535);
or UO_1629 (O_1629,N_24394,N_24381);
nor UO_1630 (O_1630,N_24519,N_24699);
nor UO_1631 (O_1631,N_24542,N_24858);
or UO_1632 (O_1632,N_24977,N_24520);
and UO_1633 (O_1633,N_24798,N_24910);
nor UO_1634 (O_1634,N_24397,N_24597);
xnor UO_1635 (O_1635,N_24867,N_24553);
nand UO_1636 (O_1636,N_24552,N_24683);
nor UO_1637 (O_1637,N_24977,N_24721);
xor UO_1638 (O_1638,N_24518,N_24762);
nor UO_1639 (O_1639,N_24654,N_24457);
xnor UO_1640 (O_1640,N_24725,N_24967);
xor UO_1641 (O_1641,N_24541,N_24592);
or UO_1642 (O_1642,N_24951,N_24725);
xnor UO_1643 (O_1643,N_24763,N_24594);
nand UO_1644 (O_1644,N_24627,N_24953);
or UO_1645 (O_1645,N_24687,N_24935);
nand UO_1646 (O_1646,N_24516,N_24927);
or UO_1647 (O_1647,N_24802,N_24958);
or UO_1648 (O_1648,N_24780,N_24825);
nor UO_1649 (O_1649,N_24637,N_24485);
or UO_1650 (O_1650,N_24653,N_24655);
or UO_1651 (O_1651,N_24874,N_24534);
or UO_1652 (O_1652,N_24903,N_24817);
and UO_1653 (O_1653,N_24678,N_24583);
nor UO_1654 (O_1654,N_24467,N_24495);
nand UO_1655 (O_1655,N_24750,N_24574);
nor UO_1656 (O_1656,N_24859,N_24713);
and UO_1657 (O_1657,N_24630,N_24900);
nand UO_1658 (O_1658,N_24639,N_24942);
xor UO_1659 (O_1659,N_24735,N_24842);
nor UO_1660 (O_1660,N_24858,N_24611);
and UO_1661 (O_1661,N_24734,N_24621);
nor UO_1662 (O_1662,N_24481,N_24637);
or UO_1663 (O_1663,N_24969,N_24574);
or UO_1664 (O_1664,N_24910,N_24473);
xnor UO_1665 (O_1665,N_24403,N_24695);
or UO_1666 (O_1666,N_24627,N_24669);
or UO_1667 (O_1667,N_24832,N_24477);
and UO_1668 (O_1668,N_24703,N_24595);
and UO_1669 (O_1669,N_24391,N_24664);
nand UO_1670 (O_1670,N_24705,N_24946);
or UO_1671 (O_1671,N_24829,N_24815);
and UO_1672 (O_1672,N_24928,N_24403);
nor UO_1673 (O_1673,N_24843,N_24735);
and UO_1674 (O_1674,N_24480,N_24861);
nor UO_1675 (O_1675,N_24486,N_24802);
or UO_1676 (O_1676,N_24650,N_24382);
and UO_1677 (O_1677,N_24936,N_24395);
and UO_1678 (O_1678,N_24967,N_24810);
nor UO_1679 (O_1679,N_24652,N_24687);
xnor UO_1680 (O_1680,N_24447,N_24422);
or UO_1681 (O_1681,N_24458,N_24847);
nor UO_1682 (O_1682,N_24467,N_24459);
nand UO_1683 (O_1683,N_24658,N_24722);
nor UO_1684 (O_1684,N_24718,N_24724);
xor UO_1685 (O_1685,N_24679,N_24936);
and UO_1686 (O_1686,N_24854,N_24852);
nor UO_1687 (O_1687,N_24954,N_24415);
and UO_1688 (O_1688,N_24583,N_24841);
xnor UO_1689 (O_1689,N_24669,N_24705);
or UO_1690 (O_1690,N_24544,N_24995);
and UO_1691 (O_1691,N_24770,N_24834);
nor UO_1692 (O_1692,N_24765,N_24522);
and UO_1693 (O_1693,N_24635,N_24956);
and UO_1694 (O_1694,N_24949,N_24960);
or UO_1695 (O_1695,N_24642,N_24871);
and UO_1696 (O_1696,N_24905,N_24888);
or UO_1697 (O_1697,N_24573,N_24469);
or UO_1698 (O_1698,N_24399,N_24567);
nor UO_1699 (O_1699,N_24389,N_24994);
xnor UO_1700 (O_1700,N_24932,N_24802);
and UO_1701 (O_1701,N_24670,N_24375);
nand UO_1702 (O_1702,N_24797,N_24811);
xnor UO_1703 (O_1703,N_24917,N_24996);
nor UO_1704 (O_1704,N_24950,N_24968);
nor UO_1705 (O_1705,N_24509,N_24660);
or UO_1706 (O_1706,N_24482,N_24983);
nand UO_1707 (O_1707,N_24737,N_24410);
and UO_1708 (O_1708,N_24720,N_24697);
nor UO_1709 (O_1709,N_24684,N_24755);
nor UO_1710 (O_1710,N_24432,N_24780);
nand UO_1711 (O_1711,N_24654,N_24978);
and UO_1712 (O_1712,N_24716,N_24888);
nand UO_1713 (O_1713,N_24846,N_24906);
nand UO_1714 (O_1714,N_24814,N_24421);
and UO_1715 (O_1715,N_24606,N_24389);
nand UO_1716 (O_1716,N_24863,N_24486);
nor UO_1717 (O_1717,N_24855,N_24904);
nor UO_1718 (O_1718,N_24701,N_24840);
or UO_1719 (O_1719,N_24836,N_24970);
xnor UO_1720 (O_1720,N_24528,N_24658);
nor UO_1721 (O_1721,N_24447,N_24978);
or UO_1722 (O_1722,N_24733,N_24680);
nand UO_1723 (O_1723,N_24796,N_24876);
nor UO_1724 (O_1724,N_24588,N_24525);
nor UO_1725 (O_1725,N_24405,N_24946);
or UO_1726 (O_1726,N_24935,N_24779);
nor UO_1727 (O_1727,N_24881,N_24977);
nand UO_1728 (O_1728,N_24647,N_24854);
xor UO_1729 (O_1729,N_24831,N_24615);
xnor UO_1730 (O_1730,N_24732,N_24899);
xnor UO_1731 (O_1731,N_24577,N_24425);
or UO_1732 (O_1732,N_24413,N_24677);
and UO_1733 (O_1733,N_24851,N_24845);
nand UO_1734 (O_1734,N_24899,N_24840);
nor UO_1735 (O_1735,N_24933,N_24544);
nand UO_1736 (O_1736,N_24439,N_24893);
nor UO_1737 (O_1737,N_24794,N_24703);
and UO_1738 (O_1738,N_24942,N_24873);
xnor UO_1739 (O_1739,N_24934,N_24698);
xor UO_1740 (O_1740,N_24494,N_24857);
nor UO_1741 (O_1741,N_24748,N_24958);
nand UO_1742 (O_1742,N_24852,N_24796);
nor UO_1743 (O_1743,N_24790,N_24954);
and UO_1744 (O_1744,N_24991,N_24766);
nor UO_1745 (O_1745,N_24596,N_24971);
nand UO_1746 (O_1746,N_24458,N_24396);
xnor UO_1747 (O_1747,N_24789,N_24875);
xor UO_1748 (O_1748,N_24802,N_24898);
xnor UO_1749 (O_1749,N_24958,N_24893);
or UO_1750 (O_1750,N_24489,N_24712);
or UO_1751 (O_1751,N_24981,N_24926);
nand UO_1752 (O_1752,N_24502,N_24870);
xnor UO_1753 (O_1753,N_24876,N_24705);
and UO_1754 (O_1754,N_24497,N_24759);
nand UO_1755 (O_1755,N_24871,N_24605);
nand UO_1756 (O_1756,N_24751,N_24565);
nor UO_1757 (O_1757,N_24695,N_24467);
nor UO_1758 (O_1758,N_24396,N_24718);
or UO_1759 (O_1759,N_24772,N_24472);
xor UO_1760 (O_1760,N_24737,N_24716);
xnor UO_1761 (O_1761,N_24547,N_24828);
or UO_1762 (O_1762,N_24572,N_24602);
nor UO_1763 (O_1763,N_24756,N_24705);
nand UO_1764 (O_1764,N_24910,N_24894);
and UO_1765 (O_1765,N_24983,N_24528);
and UO_1766 (O_1766,N_24595,N_24565);
xnor UO_1767 (O_1767,N_24703,N_24588);
or UO_1768 (O_1768,N_24713,N_24458);
or UO_1769 (O_1769,N_24591,N_24816);
nor UO_1770 (O_1770,N_24454,N_24938);
nand UO_1771 (O_1771,N_24641,N_24746);
nor UO_1772 (O_1772,N_24949,N_24647);
and UO_1773 (O_1773,N_24428,N_24392);
nand UO_1774 (O_1774,N_24914,N_24377);
xor UO_1775 (O_1775,N_24626,N_24730);
nand UO_1776 (O_1776,N_24574,N_24384);
or UO_1777 (O_1777,N_24599,N_24928);
nand UO_1778 (O_1778,N_24929,N_24552);
or UO_1779 (O_1779,N_24543,N_24778);
xor UO_1780 (O_1780,N_24677,N_24906);
xor UO_1781 (O_1781,N_24688,N_24445);
or UO_1782 (O_1782,N_24763,N_24993);
and UO_1783 (O_1783,N_24951,N_24739);
nor UO_1784 (O_1784,N_24467,N_24501);
or UO_1785 (O_1785,N_24614,N_24955);
nand UO_1786 (O_1786,N_24925,N_24896);
xor UO_1787 (O_1787,N_24645,N_24926);
nor UO_1788 (O_1788,N_24500,N_24831);
nor UO_1789 (O_1789,N_24521,N_24570);
nand UO_1790 (O_1790,N_24714,N_24391);
xnor UO_1791 (O_1791,N_24823,N_24446);
or UO_1792 (O_1792,N_24520,N_24698);
or UO_1793 (O_1793,N_24409,N_24431);
nand UO_1794 (O_1794,N_24995,N_24448);
and UO_1795 (O_1795,N_24717,N_24495);
nand UO_1796 (O_1796,N_24409,N_24447);
nor UO_1797 (O_1797,N_24884,N_24842);
nor UO_1798 (O_1798,N_24451,N_24820);
nor UO_1799 (O_1799,N_24501,N_24964);
nand UO_1800 (O_1800,N_24525,N_24658);
or UO_1801 (O_1801,N_24802,N_24817);
or UO_1802 (O_1802,N_24603,N_24739);
or UO_1803 (O_1803,N_24670,N_24567);
nor UO_1804 (O_1804,N_24475,N_24476);
nand UO_1805 (O_1805,N_24526,N_24458);
nand UO_1806 (O_1806,N_24905,N_24732);
xnor UO_1807 (O_1807,N_24587,N_24458);
nor UO_1808 (O_1808,N_24714,N_24930);
nand UO_1809 (O_1809,N_24495,N_24514);
and UO_1810 (O_1810,N_24802,N_24893);
nand UO_1811 (O_1811,N_24840,N_24972);
and UO_1812 (O_1812,N_24780,N_24603);
nor UO_1813 (O_1813,N_24612,N_24656);
and UO_1814 (O_1814,N_24797,N_24699);
xor UO_1815 (O_1815,N_24909,N_24497);
nor UO_1816 (O_1816,N_24815,N_24874);
and UO_1817 (O_1817,N_24887,N_24909);
xor UO_1818 (O_1818,N_24579,N_24914);
xnor UO_1819 (O_1819,N_24448,N_24631);
or UO_1820 (O_1820,N_24861,N_24993);
nand UO_1821 (O_1821,N_24749,N_24630);
and UO_1822 (O_1822,N_24396,N_24391);
and UO_1823 (O_1823,N_24794,N_24918);
and UO_1824 (O_1824,N_24813,N_24422);
nor UO_1825 (O_1825,N_24770,N_24694);
and UO_1826 (O_1826,N_24538,N_24552);
xor UO_1827 (O_1827,N_24470,N_24485);
nand UO_1828 (O_1828,N_24982,N_24722);
and UO_1829 (O_1829,N_24797,N_24815);
nor UO_1830 (O_1830,N_24847,N_24457);
or UO_1831 (O_1831,N_24908,N_24377);
xor UO_1832 (O_1832,N_24832,N_24573);
nor UO_1833 (O_1833,N_24570,N_24614);
nor UO_1834 (O_1834,N_24610,N_24573);
nand UO_1835 (O_1835,N_24411,N_24740);
xnor UO_1836 (O_1836,N_24990,N_24709);
nor UO_1837 (O_1837,N_24884,N_24952);
xor UO_1838 (O_1838,N_24511,N_24627);
xor UO_1839 (O_1839,N_24710,N_24602);
nor UO_1840 (O_1840,N_24906,N_24476);
or UO_1841 (O_1841,N_24385,N_24787);
nand UO_1842 (O_1842,N_24492,N_24914);
nand UO_1843 (O_1843,N_24384,N_24627);
xor UO_1844 (O_1844,N_24861,N_24908);
nand UO_1845 (O_1845,N_24952,N_24969);
nor UO_1846 (O_1846,N_24937,N_24429);
nand UO_1847 (O_1847,N_24992,N_24674);
xor UO_1848 (O_1848,N_24701,N_24659);
or UO_1849 (O_1849,N_24963,N_24964);
or UO_1850 (O_1850,N_24644,N_24741);
xor UO_1851 (O_1851,N_24855,N_24940);
nand UO_1852 (O_1852,N_24917,N_24472);
nand UO_1853 (O_1853,N_24596,N_24716);
nand UO_1854 (O_1854,N_24612,N_24446);
nand UO_1855 (O_1855,N_24571,N_24609);
nor UO_1856 (O_1856,N_24844,N_24492);
and UO_1857 (O_1857,N_24994,N_24906);
nand UO_1858 (O_1858,N_24402,N_24462);
and UO_1859 (O_1859,N_24985,N_24932);
xnor UO_1860 (O_1860,N_24984,N_24884);
nor UO_1861 (O_1861,N_24735,N_24679);
or UO_1862 (O_1862,N_24411,N_24441);
nor UO_1863 (O_1863,N_24844,N_24728);
or UO_1864 (O_1864,N_24524,N_24678);
nor UO_1865 (O_1865,N_24418,N_24830);
nor UO_1866 (O_1866,N_24564,N_24578);
nand UO_1867 (O_1867,N_24435,N_24965);
or UO_1868 (O_1868,N_24717,N_24617);
and UO_1869 (O_1869,N_24684,N_24613);
nor UO_1870 (O_1870,N_24422,N_24794);
nor UO_1871 (O_1871,N_24808,N_24672);
nand UO_1872 (O_1872,N_24711,N_24535);
nand UO_1873 (O_1873,N_24759,N_24569);
xnor UO_1874 (O_1874,N_24424,N_24636);
nand UO_1875 (O_1875,N_24541,N_24446);
nand UO_1876 (O_1876,N_24439,N_24917);
nor UO_1877 (O_1877,N_24745,N_24658);
xor UO_1878 (O_1878,N_24974,N_24464);
xnor UO_1879 (O_1879,N_24375,N_24813);
nor UO_1880 (O_1880,N_24957,N_24423);
or UO_1881 (O_1881,N_24712,N_24432);
nand UO_1882 (O_1882,N_24500,N_24982);
and UO_1883 (O_1883,N_24863,N_24516);
nor UO_1884 (O_1884,N_24681,N_24917);
nand UO_1885 (O_1885,N_24457,N_24663);
and UO_1886 (O_1886,N_24823,N_24962);
nor UO_1887 (O_1887,N_24646,N_24587);
or UO_1888 (O_1888,N_24882,N_24789);
nand UO_1889 (O_1889,N_24547,N_24545);
nor UO_1890 (O_1890,N_24609,N_24884);
xnor UO_1891 (O_1891,N_24607,N_24639);
or UO_1892 (O_1892,N_24685,N_24513);
nor UO_1893 (O_1893,N_24461,N_24553);
xnor UO_1894 (O_1894,N_24966,N_24429);
or UO_1895 (O_1895,N_24683,N_24709);
xnor UO_1896 (O_1896,N_24642,N_24753);
xnor UO_1897 (O_1897,N_24684,N_24554);
nor UO_1898 (O_1898,N_24685,N_24909);
and UO_1899 (O_1899,N_24557,N_24464);
xnor UO_1900 (O_1900,N_24384,N_24972);
nand UO_1901 (O_1901,N_24988,N_24523);
or UO_1902 (O_1902,N_24990,N_24398);
xnor UO_1903 (O_1903,N_24771,N_24415);
xor UO_1904 (O_1904,N_24825,N_24936);
nand UO_1905 (O_1905,N_24887,N_24616);
or UO_1906 (O_1906,N_24856,N_24744);
or UO_1907 (O_1907,N_24898,N_24451);
nor UO_1908 (O_1908,N_24627,N_24637);
nand UO_1909 (O_1909,N_24976,N_24680);
nor UO_1910 (O_1910,N_24675,N_24630);
nand UO_1911 (O_1911,N_24532,N_24703);
or UO_1912 (O_1912,N_24888,N_24756);
and UO_1913 (O_1913,N_24681,N_24548);
nor UO_1914 (O_1914,N_24576,N_24931);
and UO_1915 (O_1915,N_24757,N_24459);
nand UO_1916 (O_1916,N_24709,N_24547);
nor UO_1917 (O_1917,N_24699,N_24872);
and UO_1918 (O_1918,N_24739,N_24918);
or UO_1919 (O_1919,N_24859,N_24902);
and UO_1920 (O_1920,N_24779,N_24674);
xnor UO_1921 (O_1921,N_24738,N_24711);
nand UO_1922 (O_1922,N_24952,N_24676);
xor UO_1923 (O_1923,N_24483,N_24789);
nand UO_1924 (O_1924,N_24806,N_24943);
xnor UO_1925 (O_1925,N_24629,N_24628);
nor UO_1926 (O_1926,N_24633,N_24791);
nor UO_1927 (O_1927,N_24811,N_24378);
and UO_1928 (O_1928,N_24613,N_24612);
nor UO_1929 (O_1929,N_24735,N_24972);
nor UO_1930 (O_1930,N_24789,N_24610);
nand UO_1931 (O_1931,N_24716,N_24738);
and UO_1932 (O_1932,N_24951,N_24435);
or UO_1933 (O_1933,N_24461,N_24667);
or UO_1934 (O_1934,N_24861,N_24997);
xor UO_1935 (O_1935,N_24995,N_24545);
and UO_1936 (O_1936,N_24524,N_24926);
and UO_1937 (O_1937,N_24706,N_24518);
nor UO_1938 (O_1938,N_24995,N_24766);
or UO_1939 (O_1939,N_24414,N_24559);
nor UO_1940 (O_1940,N_24446,N_24443);
nor UO_1941 (O_1941,N_24601,N_24703);
nor UO_1942 (O_1942,N_24629,N_24786);
nand UO_1943 (O_1943,N_24981,N_24389);
or UO_1944 (O_1944,N_24380,N_24548);
xor UO_1945 (O_1945,N_24879,N_24688);
nor UO_1946 (O_1946,N_24922,N_24647);
nor UO_1947 (O_1947,N_24504,N_24395);
nand UO_1948 (O_1948,N_24632,N_24815);
xnor UO_1949 (O_1949,N_24917,N_24661);
or UO_1950 (O_1950,N_24801,N_24973);
xnor UO_1951 (O_1951,N_24919,N_24484);
nor UO_1952 (O_1952,N_24498,N_24481);
or UO_1953 (O_1953,N_24839,N_24885);
nor UO_1954 (O_1954,N_24431,N_24721);
nand UO_1955 (O_1955,N_24805,N_24679);
xor UO_1956 (O_1956,N_24634,N_24661);
xor UO_1957 (O_1957,N_24513,N_24923);
nor UO_1958 (O_1958,N_24475,N_24850);
or UO_1959 (O_1959,N_24595,N_24662);
nand UO_1960 (O_1960,N_24748,N_24816);
nand UO_1961 (O_1961,N_24853,N_24910);
nor UO_1962 (O_1962,N_24902,N_24819);
nor UO_1963 (O_1963,N_24736,N_24738);
or UO_1964 (O_1964,N_24462,N_24518);
and UO_1965 (O_1965,N_24547,N_24883);
nor UO_1966 (O_1966,N_24539,N_24841);
nor UO_1967 (O_1967,N_24600,N_24837);
nand UO_1968 (O_1968,N_24752,N_24526);
or UO_1969 (O_1969,N_24939,N_24670);
xnor UO_1970 (O_1970,N_24588,N_24398);
nor UO_1971 (O_1971,N_24522,N_24802);
or UO_1972 (O_1972,N_24930,N_24905);
xor UO_1973 (O_1973,N_24991,N_24887);
and UO_1974 (O_1974,N_24705,N_24431);
xor UO_1975 (O_1975,N_24794,N_24700);
or UO_1976 (O_1976,N_24789,N_24382);
and UO_1977 (O_1977,N_24885,N_24619);
xnor UO_1978 (O_1978,N_24668,N_24943);
xor UO_1979 (O_1979,N_24991,N_24790);
nor UO_1980 (O_1980,N_24767,N_24406);
and UO_1981 (O_1981,N_24532,N_24913);
and UO_1982 (O_1982,N_24521,N_24897);
and UO_1983 (O_1983,N_24729,N_24564);
xor UO_1984 (O_1984,N_24961,N_24749);
or UO_1985 (O_1985,N_24456,N_24540);
or UO_1986 (O_1986,N_24941,N_24919);
or UO_1987 (O_1987,N_24953,N_24661);
and UO_1988 (O_1988,N_24939,N_24828);
and UO_1989 (O_1989,N_24990,N_24639);
nand UO_1990 (O_1990,N_24942,N_24627);
nor UO_1991 (O_1991,N_24590,N_24555);
or UO_1992 (O_1992,N_24666,N_24930);
nor UO_1993 (O_1993,N_24386,N_24597);
nor UO_1994 (O_1994,N_24668,N_24997);
nor UO_1995 (O_1995,N_24984,N_24481);
nand UO_1996 (O_1996,N_24839,N_24520);
nand UO_1997 (O_1997,N_24521,N_24412);
nor UO_1998 (O_1998,N_24954,N_24587);
nor UO_1999 (O_1999,N_24994,N_24496);
nand UO_2000 (O_2000,N_24488,N_24799);
nand UO_2001 (O_2001,N_24870,N_24919);
nor UO_2002 (O_2002,N_24805,N_24481);
xnor UO_2003 (O_2003,N_24716,N_24541);
xnor UO_2004 (O_2004,N_24774,N_24946);
nand UO_2005 (O_2005,N_24394,N_24493);
xor UO_2006 (O_2006,N_24901,N_24801);
nor UO_2007 (O_2007,N_24882,N_24496);
nand UO_2008 (O_2008,N_24932,N_24731);
or UO_2009 (O_2009,N_24906,N_24917);
or UO_2010 (O_2010,N_24435,N_24817);
and UO_2011 (O_2011,N_24430,N_24388);
or UO_2012 (O_2012,N_24662,N_24965);
and UO_2013 (O_2013,N_24894,N_24941);
nand UO_2014 (O_2014,N_24753,N_24845);
nor UO_2015 (O_2015,N_24759,N_24381);
or UO_2016 (O_2016,N_24951,N_24578);
or UO_2017 (O_2017,N_24829,N_24921);
nor UO_2018 (O_2018,N_24663,N_24568);
or UO_2019 (O_2019,N_24482,N_24974);
xor UO_2020 (O_2020,N_24636,N_24674);
or UO_2021 (O_2021,N_24490,N_24718);
and UO_2022 (O_2022,N_24468,N_24488);
xnor UO_2023 (O_2023,N_24475,N_24853);
or UO_2024 (O_2024,N_24797,N_24774);
and UO_2025 (O_2025,N_24793,N_24706);
xor UO_2026 (O_2026,N_24817,N_24475);
nand UO_2027 (O_2027,N_24473,N_24885);
xor UO_2028 (O_2028,N_24788,N_24895);
xor UO_2029 (O_2029,N_24636,N_24956);
nor UO_2030 (O_2030,N_24512,N_24975);
xnor UO_2031 (O_2031,N_24867,N_24585);
and UO_2032 (O_2032,N_24801,N_24468);
nand UO_2033 (O_2033,N_24814,N_24795);
or UO_2034 (O_2034,N_24531,N_24921);
and UO_2035 (O_2035,N_24543,N_24852);
nand UO_2036 (O_2036,N_24483,N_24464);
or UO_2037 (O_2037,N_24978,N_24681);
or UO_2038 (O_2038,N_24807,N_24896);
and UO_2039 (O_2039,N_24560,N_24581);
or UO_2040 (O_2040,N_24429,N_24962);
or UO_2041 (O_2041,N_24883,N_24592);
xnor UO_2042 (O_2042,N_24570,N_24744);
nor UO_2043 (O_2043,N_24839,N_24542);
or UO_2044 (O_2044,N_24580,N_24959);
xor UO_2045 (O_2045,N_24935,N_24637);
nor UO_2046 (O_2046,N_24867,N_24576);
nand UO_2047 (O_2047,N_24447,N_24860);
and UO_2048 (O_2048,N_24606,N_24930);
and UO_2049 (O_2049,N_24772,N_24938);
and UO_2050 (O_2050,N_24408,N_24875);
nor UO_2051 (O_2051,N_24709,N_24526);
nand UO_2052 (O_2052,N_24681,N_24502);
or UO_2053 (O_2053,N_24844,N_24508);
and UO_2054 (O_2054,N_24978,N_24660);
or UO_2055 (O_2055,N_24421,N_24510);
and UO_2056 (O_2056,N_24496,N_24417);
nor UO_2057 (O_2057,N_24508,N_24377);
or UO_2058 (O_2058,N_24490,N_24995);
and UO_2059 (O_2059,N_24731,N_24927);
nor UO_2060 (O_2060,N_24849,N_24995);
and UO_2061 (O_2061,N_24444,N_24860);
and UO_2062 (O_2062,N_24610,N_24424);
and UO_2063 (O_2063,N_24476,N_24799);
and UO_2064 (O_2064,N_24709,N_24808);
or UO_2065 (O_2065,N_24573,N_24609);
nand UO_2066 (O_2066,N_24427,N_24987);
and UO_2067 (O_2067,N_24721,N_24896);
xor UO_2068 (O_2068,N_24800,N_24844);
nand UO_2069 (O_2069,N_24807,N_24569);
nor UO_2070 (O_2070,N_24938,N_24709);
xor UO_2071 (O_2071,N_24736,N_24502);
nand UO_2072 (O_2072,N_24534,N_24816);
and UO_2073 (O_2073,N_24401,N_24872);
nor UO_2074 (O_2074,N_24558,N_24466);
nor UO_2075 (O_2075,N_24677,N_24787);
nand UO_2076 (O_2076,N_24490,N_24485);
nand UO_2077 (O_2077,N_24551,N_24717);
and UO_2078 (O_2078,N_24830,N_24883);
nor UO_2079 (O_2079,N_24780,N_24851);
xor UO_2080 (O_2080,N_24928,N_24457);
or UO_2081 (O_2081,N_24432,N_24849);
or UO_2082 (O_2082,N_24897,N_24470);
nand UO_2083 (O_2083,N_24528,N_24797);
nand UO_2084 (O_2084,N_24695,N_24993);
and UO_2085 (O_2085,N_24500,N_24965);
and UO_2086 (O_2086,N_24419,N_24823);
nor UO_2087 (O_2087,N_24881,N_24614);
nand UO_2088 (O_2088,N_24513,N_24623);
or UO_2089 (O_2089,N_24760,N_24563);
nor UO_2090 (O_2090,N_24670,N_24783);
nor UO_2091 (O_2091,N_24436,N_24546);
and UO_2092 (O_2092,N_24561,N_24798);
and UO_2093 (O_2093,N_24999,N_24432);
nand UO_2094 (O_2094,N_24924,N_24697);
xnor UO_2095 (O_2095,N_24728,N_24420);
and UO_2096 (O_2096,N_24530,N_24928);
and UO_2097 (O_2097,N_24966,N_24679);
xnor UO_2098 (O_2098,N_24657,N_24958);
xor UO_2099 (O_2099,N_24794,N_24499);
and UO_2100 (O_2100,N_24423,N_24590);
nand UO_2101 (O_2101,N_24532,N_24530);
xor UO_2102 (O_2102,N_24909,N_24660);
or UO_2103 (O_2103,N_24998,N_24599);
and UO_2104 (O_2104,N_24402,N_24612);
xnor UO_2105 (O_2105,N_24766,N_24552);
nand UO_2106 (O_2106,N_24565,N_24383);
and UO_2107 (O_2107,N_24415,N_24986);
or UO_2108 (O_2108,N_24995,N_24428);
nand UO_2109 (O_2109,N_24656,N_24926);
nor UO_2110 (O_2110,N_24973,N_24889);
xnor UO_2111 (O_2111,N_24811,N_24847);
xor UO_2112 (O_2112,N_24904,N_24917);
nor UO_2113 (O_2113,N_24407,N_24998);
xor UO_2114 (O_2114,N_24813,N_24997);
and UO_2115 (O_2115,N_24582,N_24715);
or UO_2116 (O_2116,N_24543,N_24859);
xnor UO_2117 (O_2117,N_24840,N_24984);
and UO_2118 (O_2118,N_24445,N_24644);
or UO_2119 (O_2119,N_24908,N_24842);
nor UO_2120 (O_2120,N_24557,N_24514);
xnor UO_2121 (O_2121,N_24516,N_24426);
xor UO_2122 (O_2122,N_24529,N_24882);
and UO_2123 (O_2123,N_24519,N_24454);
xnor UO_2124 (O_2124,N_24561,N_24649);
xnor UO_2125 (O_2125,N_24733,N_24753);
nor UO_2126 (O_2126,N_24545,N_24662);
nand UO_2127 (O_2127,N_24505,N_24634);
and UO_2128 (O_2128,N_24678,N_24572);
nand UO_2129 (O_2129,N_24779,N_24673);
and UO_2130 (O_2130,N_24506,N_24661);
nand UO_2131 (O_2131,N_24587,N_24923);
nor UO_2132 (O_2132,N_24907,N_24388);
nor UO_2133 (O_2133,N_24686,N_24813);
and UO_2134 (O_2134,N_24461,N_24480);
and UO_2135 (O_2135,N_24884,N_24558);
nor UO_2136 (O_2136,N_24822,N_24503);
or UO_2137 (O_2137,N_24891,N_24826);
or UO_2138 (O_2138,N_24854,N_24877);
and UO_2139 (O_2139,N_24555,N_24913);
and UO_2140 (O_2140,N_24636,N_24582);
nor UO_2141 (O_2141,N_24498,N_24710);
xor UO_2142 (O_2142,N_24888,N_24982);
nor UO_2143 (O_2143,N_24530,N_24472);
or UO_2144 (O_2144,N_24887,N_24729);
or UO_2145 (O_2145,N_24970,N_24404);
or UO_2146 (O_2146,N_24408,N_24414);
nor UO_2147 (O_2147,N_24806,N_24995);
or UO_2148 (O_2148,N_24802,N_24833);
nand UO_2149 (O_2149,N_24491,N_24970);
nor UO_2150 (O_2150,N_24845,N_24726);
nor UO_2151 (O_2151,N_24741,N_24988);
and UO_2152 (O_2152,N_24582,N_24725);
nor UO_2153 (O_2153,N_24954,N_24887);
or UO_2154 (O_2154,N_24573,N_24738);
nand UO_2155 (O_2155,N_24524,N_24895);
and UO_2156 (O_2156,N_24929,N_24469);
or UO_2157 (O_2157,N_24607,N_24814);
or UO_2158 (O_2158,N_24405,N_24615);
or UO_2159 (O_2159,N_24807,N_24469);
xnor UO_2160 (O_2160,N_24955,N_24498);
nor UO_2161 (O_2161,N_24874,N_24737);
and UO_2162 (O_2162,N_24713,N_24556);
nand UO_2163 (O_2163,N_24754,N_24484);
or UO_2164 (O_2164,N_24889,N_24856);
or UO_2165 (O_2165,N_24975,N_24726);
nor UO_2166 (O_2166,N_24964,N_24668);
nand UO_2167 (O_2167,N_24978,N_24998);
nand UO_2168 (O_2168,N_24920,N_24929);
nor UO_2169 (O_2169,N_24967,N_24985);
nand UO_2170 (O_2170,N_24813,N_24880);
xnor UO_2171 (O_2171,N_24637,N_24376);
and UO_2172 (O_2172,N_24984,N_24696);
nand UO_2173 (O_2173,N_24438,N_24379);
nand UO_2174 (O_2174,N_24730,N_24598);
or UO_2175 (O_2175,N_24467,N_24698);
or UO_2176 (O_2176,N_24890,N_24696);
or UO_2177 (O_2177,N_24653,N_24424);
and UO_2178 (O_2178,N_24723,N_24686);
nand UO_2179 (O_2179,N_24703,N_24732);
nor UO_2180 (O_2180,N_24646,N_24409);
nor UO_2181 (O_2181,N_24593,N_24603);
nand UO_2182 (O_2182,N_24959,N_24857);
nand UO_2183 (O_2183,N_24948,N_24404);
nor UO_2184 (O_2184,N_24519,N_24975);
or UO_2185 (O_2185,N_24390,N_24878);
nand UO_2186 (O_2186,N_24593,N_24496);
nor UO_2187 (O_2187,N_24797,N_24772);
or UO_2188 (O_2188,N_24545,N_24898);
or UO_2189 (O_2189,N_24980,N_24753);
and UO_2190 (O_2190,N_24386,N_24754);
nand UO_2191 (O_2191,N_24821,N_24831);
and UO_2192 (O_2192,N_24566,N_24677);
xnor UO_2193 (O_2193,N_24427,N_24715);
nand UO_2194 (O_2194,N_24424,N_24430);
and UO_2195 (O_2195,N_24934,N_24998);
xnor UO_2196 (O_2196,N_24763,N_24764);
nor UO_2197 (O_2197,N_24708,N_24704);
and UO_2198 (O_2198,N_24967,N_24954);
or UO_2199 (O_2199,N_24902,N_24809);
xor UO_2200 (O_2200,N_24563,N_24718);
nand UO_2201 (O_2201,N_24994,N_24924);
nand UO_2202 (O_2202,N_24575,N_24718);
nand UO_2203 (O_2203,N_24635,N_24832);
and UO_2204 (O_2204,N_24426,N_24672);
nand UO_2205 (O_2205,N_24699,N_24651);
nand UO_2206 (O_2206,N_24780,N_24532);
nor UO_2207 (O_2207,N_24433,N_24501);
nand UO_2208 (O_2208,N_24874,N_24542);
nand UO_2209 (O_2209,N_24438,N_24578);
or UO_2210 (O_2210,N_24492,N_24497);
or UO_2211 (O_2211,N_24815,N_24814);
nor UO_2212 (O_2212,N_24442,N_24767);
xor UO_2213 (O_2213,N_24691,N_24847);
and UO_2214 (O_2214,N_24863,N_24903);
xor UO_2215 (O_2215,N_24594,N_24992);
nor UO_2216 (O_2216,N_24850,N_24725);
nand UO_2217 (O_2217,N_24400,N_24881);
and UO_2218 (O_2218,N_24773,N_24486);
and UO_2219 (O_2219,N_24958,N_24393);
nor UO_2220 (O_2220,N_24895,N_24547);
nor UO_2221 (O_2221,N_24643,N_24487);
or UO_2222 (O_2222,N_24719,N_24454);
or UO_2223 (O_2223,N_24676,N_24534);
and UO_2224 (O_2224,N_24912,N_24651);
nor UO_2225 (O_2225,N_24838,N_24531);
xnor UO_2226 (O_2226,N_24745,N_24537);
or UO_2227 (O_2227,N_24600,N_24860);
or UO_2228 (O_2228,N_24817,N_24900);
and UO_2229 (O_2229,N_24659,N_24626);
nor UO_2230 (O_2230,N_24435,N_24699);
nand UO_2231 (O_2231,N_24636,N_24623);
nand UO_2232 (O_2232,N_24984,N_24414);
nand UO_2233 (O_2233,N_24840,N_24721);
nor UO_2234 (O_2234,N_24892,N_24540);
nor UO_2235 (O_2235,N_24510,N_24861);
nor UO_2236 (O_2236,N_24461,N_24630);
and UO_2237 (O_2237,N_24806,N_24731);
or UO_2238 (O_2238,N_24789,N_24979);
and UO_2239 (O_2239,N_24595,N_24873);
or UO_2240 (O_2240,N_24613,N_24670);
or UO_2241 (O_2241,N_24652,N_24946);
or UO_2242 (O_2242,N_24905,N_24462);
xor UO_2243 (O_2243,N_24814,N_24785);
nor UO_2244 (O_2244,N_24820,N_24402);
or UO_2245 (O_2245,N_24700,N_24499);
nor UO_2246 (O_2246,N_24390,N_24819);
xnor UO_2247 (O_2247,N_24823,N_24744);
nand UO_2248 (O_2248,N_24956,N_24589);
nand UO_2249 (O_2249,N_24441,N_24739);
nor UO_2250 (O_2250,N_24407,N_24576);
or UO_2251 (O_2251,N_24479,N_24474);
xor UO_2252 (O_2252,N_24949,N_24645);
and UO_2253 (O_2253,N_24848,N_24972);
xor UO_2254 (O_2254,N_24793,N_24425);
and UO_2255 (O_2255,N_24645,N_24613);
nand UO_2256 (O_2256,N_24640,N_24914);
xor UO_2257 (O_2257,N_24696,N_24836);
and UO_2258 (O_2258,N_24954,N_24445);
nor UO_2259 (O_2259,N_24573,N_24928);
nor UO_2260 (O_2260,N_24556,N_24963);
nand UO_2261 (O_2261,N_24589,N_24854);
nor UO_2262 (O_2262,N_24689,N_24437);
xor UO_2263 (O_2263,N_24607,N_24960);
and UO_2264 (O_2264,N_24621,N_24791);
or UO_2265 (O_2265,N_24385,N_24863);
or UO_2266 (O_2266,N_24618,N_24421);
xor UO_2267 (O_2267,N_24574,N_24657);
nand UO_2268 (O_2268,N_24567,N_24511);
or UO_2269 (O_2269,N_24816,N_24401);
nand UO_2270 (O_2270,N_24533,N_24614);
xor UO_2271 (O_2271,N_24508,N_24607);
or UO_2272 (O_2272,N_24401,N_24916);
or UO_2273 (O_2273,N_24562,N_24543);
or UO_2274 (O_2274,N_24456,N_24522);
xnor UO_2275 (O_2275,N_24570,N_24491);
nor UO_2276 (O_2276,N_24908,N_24944);
nand UO_2277 (O_2277,N_24449,N_24856);
xor UO_2278 (O_2278,N_24974,N_24922);
and UO_2279 (O_2279,N_24443,N_24687);
nand UO_2280 (O_2280,N_24749,N_24716);
nand UO_2281 (O_2281,N_24595,N_24602);
or UO_2282 (O_2282,N_24699,N_24831);
nand UO_2283 (O_2283,N_24487,N_24443);
and UO_2284 (O_2284,N_24779,N_24857);
nor UO_2285 (O_2285,N_24709,N_24572);
xnor UO_2286 (O_2286,N_24385,N_24613);
nor UO_2287 (O_2287,N_24429,N_24994);
nor UO_2288 (O_2288,N_24525,N_24751);
and UO_2289 (O_2289,N_24674,N_24835);
and UO_2290 (O_2290,N_24497,N_24789);
nand UO_2291 (O_2291,N_24607,N_24902);
nor UO_2292 (O_2292,N_24743,N_24797);
xnor UO_2293 (O_2293,N_24651,N_24982);
or UO_2294 (O_2294,N_24784,N_24552);
nand UO_2295 (O_2295,N_24672,N_24750);
nor UO_2296 (O_2296,N_24769,N_24970);
nor UO_2297 (O_2297,N_24616,N_24923);
xnor UO_2298 (O_2298,N_24640,N_24854);
nand UO_2299 (O_2299,N_24869,N_24492);
nor UO_2300 (O_2300,N_24834,N_24479);
or UO_2301 (O_2301,N_24851,N_24517);
xnor UO_2302 (O_2302,N_24482,N_24916);
and UO_2303 (O_2303,N_24816,N_24722);
nand UO_2304 (O_2304,N_24601,N_24903);
nand UO_2305 (O_2305,N_24744,N_24826);
or UO_2306 (O_2306,N_24456,N_24970);
or UO_2307 (O_2307,N_24409,N_24630);
xnor UO_2308 (O_2308,N_24383,N_24758);
nor UO_2309 (O_2309,N_24488,N_24729);
nand UO_2310 (O_2310,N_24873,N_24676);
and UO_2311 (O_2311,N_24803,N_24674);
and UO_2312 (O_2312,N_24433,N_24944);
and UO_2313 (O_2313,N_24731,N_24646);
nand UO_2314 (O_2314,N_24519,N_24905);
or UO_2315 (O_2315,N_24867,N_24490);
or UO_2316 (O_2316,N_24666,N_24836);
xor UO_2317 (O_2317,N_24376,N_24651);
nand UO_2318 (O_2318,N_24735,N_24583);
and UO_2319 (O_2319,N_24762,N_24695);
or UO_2320 (O_2320,N_24805,N_24448);
nand UO_2321 (O_2321,N_24920,N_24626);
or UO_2322 (O_2322,N_24951,N_24884);
xor UO_2323 (O_2323,N_24819,N_24516);
xnor UO_2324 (O_2324,N_24406,N_24772);
nor UO_2325 (O_2325,N_24622,N_24449);
xnor UO_2326 (O_2326,N_24715,N_24491);
xnor UO_2327 (O_2327,N_24472,N_24468);
or UO_2328 (O_2328,N_24651,N_24555);
nor UO_2329 (O_2329,N_24736,N_24419);
xnor UO_2330 (O_2330,N_24393,N_24544);
or UO_2331 (O_2331,N_24777,N_24841);
nand UO_2332 (O_2332,N_24752,N_24494);
xnor UO_2333 (O_2333,N_24954,N_24976);
nand UO_2334 (O_2334,N_24656,N_24669);
nor UO_2335 (O_2335,N_24606,N_24705);
nand UO_2336 (O_2336,N_24536,N_24580);
xnor UO_2337 (O_2337,N_24787,N_24852);
nor UO_2338 (O_2338,N_24991,N_24931);
nand UO_2339 (O_2339,N_24738,N_24851);
or UO_2340 (O_2340,N_24404,N_24790);
xor UO_2341 (O_2341,N_24893,N_24799);
nand UO_2342 (O_2342,N_24735,N_24552);
or UO_2343 (O_2343,N_24591,N_24958);
and UO_2344 (O_2344,N_24852,N_24865);
xor UO_2345 (O_2345,N_24527,N_24432);
and UO_2346 (O_2346,N_24835,N_24664);
or UO_2347 (O_2347,N_24868,N_24710);
and UO_2348 (O_2348,N_24680,N_24964);
or UO_2349 (O_2349,N_24661,N_24701);
nand UO_2350 (O_2350,N_24624,N_24542);
nor UO_2351 (O_2351,N_24385,N_24518);
nor UO_2352 (O_2352,N_24802,N_24749);
xor UO_2353 (O_2353,N_24683,N_24821);
xnor UO_2354 (O_2354,N_24790,N_24747);
nand UO_2355 (O_2355,N_24726,N_24437);
nor UO_2356 (O_2356,N_24774,N_24936);
xnor UO_2357 (O_2357,N_24398,N_24845);
nand UO_2358 (O_2358,N_24437,N_24546);
and UO_2359 (O_2359,N_24890,N_24693);
or UO_2360 (O_2360,N_24497,N_24912);
nand UO_2361 (O_2361,N_24457,N_24999);
nor UO_2362 (O_2362,N_24769,N_24680);
nor UO_2363 (O_2363,N_24747,N_24474);
nand UO_2364 (O_2364,N_24574,N_24804);
and UO_2365 (O_2365,N_24778,N_24911);
nor UO_2366 (O_2366,N_24834,N_24676);
and UO_2367 (O_2367,N_24755,N_24837);
nor UO_2368 (O_2368,N_24824,N_24792);
xnor UO_2369 (O_2369,N_24945,N_24576);
and UO_2370 (O_2370,N_24405,N_24869);
nand UO_2371 (O_2371,N_24633,N_24375);
xnor UO_2372 (O_2372,N_24989,N_24787);
nand UO_2373 (O_2373,N_24928,N_24443);
nand UO_2374 (O_2374,N_24529,N_24591);
and UO_2375 (O_2375,N_24537,N_24620);
or UO_2376 (O_2376,N_24534,N_24411);
nor UO_2377 (O_2377,N_24860,N_24993);
nand UO_2378 (O_2378,N_24565,N_24818);
nor UO_2379 (O_2379,N_24454,N_24882);
nor UO_2380 (O_2380,N_24684,N_24968);
xnor UO_2381 (O_2381,N_24614,N_24830);
or UO_2382 (O_2382,N_24797,N_24633);
nand UO_2383 (O_2383,N_24436,N_24673);
and UO_2384 (O_2384,N_24702,N_24786);
and UO_2385 (O_2385,N_24454,N_24394);
xnor UO_2386 (O_2386,N_24972,N_24435);
xnor UO_2387 (O_2387,N_24491,N_24751);
nand UO_2388 (O_2388,N_24443,N_24377);
xnor UO_2389 (O_2389,N_24609,N_24549);
and UO_2390 (O_2390,N_24379,N_24711);
xnor UO_2391 (O_2391,N_24978,N_24980);
or UO_2392 (O_2392,N_24699,N_24620);
xnor UO_2393 (O_2393,N_24690,N_24817);
nor UO_2394 (O_2394,N_24696,N_24799);
or UO_2395 (O_2395,N_24926,N_24965);
and UO_2396 (O_2396,N_24701,N_24399);
nand UO_2397 (O_2397,N_24887,N_24535);
xnor UO_2398 (O_2398,N_24414,N_24948);
and UO_2399 (O_2399,N_24937,N_24579);
or UO_2400 (O_2400,N_24971,N_24555);
and UO_2401 (O_2401,N_24511,N_24861);
or UO_2402 (O_2402,N_24404,N_24746);
nand UO_2403 (O_2403,N_24948,N_24576);
or UO_2404 (O_2404,N_24926,N_24839);
nand UO_2405 (O_2405,N_24867,N_24892);
xor UO_2406 (O_2406,N_24427,N_24776);
xor UO_2407 (O_2407,N_24473,N_24905);
xnor UO_2408 (O_2408,N_24425,N_24795);
nand UO_2409 (O_2409,N_24741,N_24731);
xnor UO_2410 (O_2410,N_24721,N_24526);
xor UO_2411 (O_2411,N_24574,N_24454);
or UO_2412 (O_2412,N_24479,N_24427);
nor UO_2413 (O_2413,N_24545,N_24956);
nor UO_2414 (O_2414,N_24770,N_24774);
xor UO_2415 (O_2415,N_24739,N_24842);
nor UO_2416 (O_2416,N_24937,N_24983);
nand UO_2417 (O_2417,N_24964,N_24692);
xor UO_2418 (O_2418,N_24667,N_24469);
or UO_2419 (O_2419,N_24413,N_24505);
xnor UO_2420 (O_2420,N_24537,N_24678);
or UO_2421 (O_2421,N_24894,N_24965);
nor UO_2422 (O_2422,N_24682,N_24582);
and UO_2423 (O_2423,N_24809,N_24759);
and UO_2424 (O_2424,N_24981,N_24796);
nor UO_2425 (O_2425,N_24457,N_24391);
or UO_2426 (O_2426,N_24620,N_24943);
nor UO_2427 (O_2427,N_24594,N_24835);
and UO_2428 (O_2428,N_24497,N_24849);
nor UO_2429 (O_2429,N_24728,N_24919);
nand UO_2430 (O_2430,N_24466,N_24672);
and UO_2431 (O_2431,N_24565,N_24613);
or UO_2432 (O_2432,N_24697,N_24900);
xor UO_2433 (O_2433,N_24689,N_24926);
nand UO_2434 (O_2434,N_24422,N_24642);
nor UO_2435 (O_2435,N_24401,N_24706);
nand UO_2436 (O_2436,N_24827,N_24648);
xor UO_2437 (O_2437,N_24403,N_24902);
and UO_2438 (O_2438,N_24491,N_24877);
xnor UO_2439 (O_2439,N_24628,N_24910);
xor UO_2440 (O_2440,N_24922,N_24690);
nand UO_2441 (O_2441,N_24956,N_24417);
and UO_2442 (O_2442,N_24554,N_24601);
and UO_2443 (O_2443,N_24450,N_24738);
or UO_2444 (O_2444,N_24561,N_24591);
nand UO_2445 (O_2445,N_24607,N_24813);
nand UO_2446 (O_2446,N_24665,N_24778);
or UO_2447 (O_2447,N_24953,N_24990);
nor UO_2448 (O_2448,N_24529,N_24388);
nand UO_2449 (O_2449,N_24664,N_24453);
nand UO_2450 (O_2450,N_24704,N_24677);
and UO_2451 (O_2451,N_24864,N_24908);
xor UO_2452 (O_2452,N_24993,N_24805);
nand UO_2453 (O_2453,N_24822,N_24988);
xnor UO_2454 (O_2454,N_24450,N_24723);
xor UO_2455 (O_2455,N_24459,N_24535);
nor UO_2456 (O_2456,N_24503,N_24905);
and UO_2457 (O_2457,N_24910,N_24945);
nand UO_2458 (O_2458,N_24958,N_24742);
nor UO_2459 (O_2459,N_24678,N_24677);
nor UO_2460 (O_2460,N_24451,N_24495);
nand UO_2461 (O_2461,N_24504,N_24793);
or UO_2462 (O_2462,N_24985,N_24573);
or UO_2463 (O_2463,N_24721,N_24844);
and UO_2464 (O_2464,N_24691,N_24829);
nor UO_2465 (O_2465,N_24837,N_24607);
nor UO_2466 (O_2466,N_24835,N_24934);
and UO_2467 (O_2467,N_24393,N_24421);
and UO_2468 (O_2468,N_24565,N_24903);
or UO_2469 (O_2469,N_24763,N_24935);
nor UO_2470 (O_2470,N_24498,N_24894);
nand UO_2471 (O_2471,N_24402,N_24907);
nor UO_2472 (O_2472,N_24602,N_24451);
or UO_2473 (O_2473,N_24567,N_24737);
xor UO_2474 (O_2474,N_24627,N_24380);
nor UO_2475 (O_2475,N_24979,N_24984);
nor UO_2476 (O_2476,N_24702,N_24805);
nor UO_2477 (O_2477,N_24964,N_24984);
xor UO_2478 (O_2478,N_24515,N_24685);
or UO_2479 (O_2479,N_24606,N_24922);
xnor UO_2480 (O_2480,N_24537,N_24915);
xor UO_2481 (O_2481,N_24866,N_24825);
and UO_2482 (O_2482,N_24559,N_24448);
or UO_2483 (O_2483,N_24900,N_24546);
xnor UO_2484 (O_2484,N_24899,N_24524);
or UO_2485 (O_2485,N_24501,N_24504);
nand UO_2486 (O_2486,N_24768,N_24657);
and UO_2487 (O_2487,N_24570,N_24499);
nor UO_2488 (O_2488,N_24807,N_24406);
nand UO_2489 (O_2489,N_24907,N_24721);
nand UO_2490 (O_2490,N_24642,N_24424);
or UO_2491 (O_2491,N_24594,N_24625);
and UO_2492 (O_2492,N_24587,N_24590);
xor UO_2493 (O_2493,N_24826,N_24969);
and UO_2494 (O_2494,N_24770,N_24461);
and UO_2495 (O_2495,N_24753,N_24871);
nor UO_2496 (O_2496,N_24807,N_24917);
xor UO_2497 (O_2497,N_24740,N_24606);
nor UO_2498 (O_2498,N_24687,N_24877);
or UO_2499 (O_2499,N_24868,N_24887);
nand UO_2500 (O_2500,N_24813,N_24496);
or UO_2501 (O_2501,N_24786,N_24510);
xor UO_2502 (O_2502,N_24816,N_24626);
xnor UO_2503 (O_2503,N_24614,N_24423);
nor UO_2504 (O_2504,N_24572,N_24436);
and UO_2505 (O_2505,N_24547,N_24853);
nand UO_2506 (O_2506,N_24380,N_24750);
nor UO_2507 (O_2507,N_24724,N_24601);
nor UO_2508 (O_2508,N_24540,N_24554);
or UO_2509 (O_2509,N_24787,N_24954);
nand UO_2510 (O_2510,N_24965,N_24619);
and UO_2511 (O_2511,N_24515,N_24706);
xor UO_2512 (O_2512,N_24395,N_24438);
nand UO_2513 (O_2513,N_24401,N_24906);
nand UO_2514 (O_2514,N_24918,N_24824);
nand UO_2515 (O_2515,N_24863,N_24629);
nor UO_2516 (O_2516,N_24460,N_24731);
and UO_2517 (O_2517,N_24490,N_24487);
xor UO_2518 (O_2518,N_24594,N_24789);
nor UO_2519 (O_2519,N_24972,N_24942);
or UO_2520 (O_2520,N_24932,N_24550);
or UO_2521 (O_2521,N_24812,N_24806);
nor UO_2522 (O_2522,N_24412,N_24651);
nor UO_2523 (O_2523,N_24408,N_24798);
and UO_2524 (O_2524,N_24768,N_24709);
nor UO_2525 (O_2525,N_24955,N_24837);
nand UO_2526 (O_2526,N_24679,N_24592);
nand UO_2527 (O_2527,N_24653,N_24390);
xnor UO_2528 (O_2528,N_24606,N_24806);
or UO_2529 (O_2529,N_24632,N_24833);
and UO_2530 (O_2530,N_24660,N_24825);
nor UO_2531 (O_2531,N_24890,N_24532);
and UO_2532 (O_2532,N_24783,N_24767);
or UO_2533 (O_2533,N_24664,N_24906);
nor UO_2534 (O_2534,N_24994,N_24669);
or UO_2535 (O_2535,N_24527,N_24720);
or UO_2536 (O_2536,N_24564,N_24550);
and UO_2537 (O_2537,N_24582,N_24630);
and UO_2538 (O_2538,N_24874,N_24587);
nand UO_2539 (O_2539,N_24666,N_24494);
or UO_2540 (O_2540,N_24937,N_24610);
and UO_2541 (O_2541,N_24782,N_24731);
and UO_2542 (O_2542,N_24904,N_24832);
or UO_2543 (O_2543,N_24492,N_24644);
nor UO_2544 (O_2544,N_24896,N_24597);
nor UO_2545 (O_2545,N_24469,N_24438);
or UO_2546 (O_2546,N_24486,N_24462);
and UO_2547 (O_2547,N_24758,N_24679);
xnor UO_2548 (O_2548,N_24631,N_24936);
xor UO_2549 (O_2549,N_24579,N_24817);
xnor UO_2550 (O_2550,N_24877,N_24774);
nor UO_2551 (O_2551,N_24433,N_24805);
xor UO_2552 (O_2552,N_24634,N_24406);
xnor UO_2553 (O_2553,N_24563,N_24808);
nand UO_2554 (O_2554,N_24406,N_24765);
and UO_2555 (O_2555,N_24892,N_24585);
and UO_2556 (O_2556,N_24945,N_24808);
xnor UO_2557 (O_2557,N_24991,N_24379);
or UO_2558 (O_2558,N_24691,N_24891);
xnor UO_2559 (O_2559,N_24887,N_24446);
or UO_2560 (O_2560,N_24630,N_24468);
or UO_2561 (O_2561,N_24547,N_24450);
xor UO_2562 (O_2562,N_24533,N_24400);
nand UO_2563 (O_2563,N_24672,N_24611);
nor UO_2564 (O_2564,N_24538,N_24602);
nand UO_2565 (O_2565,N_24737,N_24524);
nor UO_2566 (O_2566,N_24516,N_24499);
nand UO_2567 (O_2567,N_24900,N_24875);
nor UO_2568 (O_2568,N_24612,N_24813);
nand UO_2569 (O_2569,N_24383,N_24406);
or UO_2570 (O_2570,N_24915,N_24629);
and UO_2571 (O_2571,N_24748,N_24993);
xor UO_2572 (O_2572,N_24800,N_24469);
xnor UO_2573 (O_2573,N_24483,N_24636);
nand UO_2574 (O_2574,N_24732,N_24973);
nor UO_2575 (O_2575,N_24821,N_24502);
nand UO_2576 (O_2576,N_24891,N_24936);
xor UO_2577 (O_2577,N_24651,N_24624);
nor UO_2578 (O_2578,N_24817,N_24569);
nor UO_2579 (O_2579,N_24632,N_24519);
and UO_2580 (O_2580,N_24924,N_24590);
and UO_2581 (O_2581,N_24631,N_24523);
nand UO_2582 (O_2582,N_24726,N_24755);
nand UO_2583 (O_2583,N_24466,N_24743);
or UO_2584 (O_2584,N_24680,N_24982);
or UO_2585 (O_2585,N_24466,N_24944);
nand UO_2586 (O_2586,N_24722,N_24462);
or UO_2587 (O_2587,N_24718,N_24628);
and UO_2588 (O_2588,N_24492,N_24467);
nand UO_2589 (O_2589,N_24587,N_24841);
nand UO_2590 (O_2590,N_24899,N_24924);
xor UO_2591 (O_2591,N_24455,N_24882);
nor UO_2592 (O_2592,N_24702,N_24721);
xnor UO_2593 (O_2593,N_24644,N_24946);
nand UO_2594 (O_2594,N_24848,N_24614);
or UO_2595 (O_2595,N_24987,N_24875);
nand UO_2596 (O_2596,N_24393,N_24755);
or UO_2597 (O_2597,N_24908,N_24850);
nand UO_2598 (O_2598,N_24748,N_24739);
or UO_2599 (O_2599,N_24719,N_24545);
and UO_2600 (O_2600,N_24556,N_24787);
nor UO_2601 (O_2601,N_24458,N_24689);
xnor UO_2602 (O_2602,N_24878,N_24546);
or UO_2603 (O_2603,N_24795,N_24554);
nor UO_2604 (O_2604,N_24690,N_24481);
nor UO_2605 (O_2605,N_24802,N_24552);
nand UO_2606 (O_2606,N_24824,N_24493);
and UO_2607 (O_2607,N_24691,N_24497);
and UO_2608 (O_2608,N_24535,N_24866);
or UO_2609 (O_2609,N_24609,N_24808);
or UO_2610 (O_2610,N_24451,N_24704);
nand UO_2611 (O_2611,N_24552,N_24693);
nor UO_2612 (O_2612,N_24858,N_24869);
and UO_2613 (O_2613,N_24552,N_24505);
nor UO_2614 (O_2614,N_24638,N_24426);
or UO_2615 (O_2615,N_24844,N_24887);
and UO_2616 (O_2616,N_24704,N_24976);
nand UO_2617 (O_2617,N_24883,N_24871);
and UO_2618 (O_2618,N_24670,N_24787);
or UO_2619 (O_2619,N_24865,N_24795);
and UO_2620 (O_2620,N_24950,N_24802);
nor UO_2621 (O_2621,N_24568,N_24755);
xor UO_2622 (O_2622,N_24581,N_24576);
xnor UO_2623 (O_2623,N_24750,N_24858);
nor UO_2624 (O_2624,N_24638,N_24495);
xor UO_2625 (O_2625,N_24870,N_24845);
nor UO_2626 (O_2626,N_24853,N_24431);
nand UO_2627 (O_2627,N_24991,N_24739);
or UO_2628 (O_2628,N_24708,N_24878);
nor UO_2629 (O_2629,N_24680,N_24849);
nor UO_2630 (O_2630,N_24441,N_24566);
xnor UO_2631 (O_2631,N_24485,N_24967);
nor UO_2632 (O_2632,N_24866,N_24502);
xnor UO_2633 (O_2633,N_24403,N_24984);
nand UO_2634 (O_2634,N_24878,N_24934);
xor UO_2635 (O_2635,N_24472,N_24431);
nand UO_2636 (O_2636,N_24712,N_24697);
and UO_2637 (O_2637,N_24629,N_24771);
and UO_2638 (O_2638,N_24526,N_24453);
nand UO_2639 (O_2639,N_24892,N_24975);
or UO_2640 (O_2640,N_24922,N_24864);
and UO_2641 (O_2641,N_24925,N_24673);
and UO_2642 (O_2642,N_24628,N_24869);
xnor UO_2643 (O_2643,N_24527,N_24743);
and UO_2644 (O_2644,N_24648,N_24871);
xnor UO_2645 (O_2645,N_24454,N_24603);
and UO_2646 (O_2646,N_24509,N_24734);
or UO_2647 (O_2647,N_24910,N_24879);
nor UO_2648 (O_2648,N_24559,N_24406);
nand UO_2649 (O_2649,N_24898,N_24452);
nor UO_2650 (O_2650,N_24629,N_24717);
xnor UO_2651 (O_2651,N_24867,N_24631);
and UO_2652 (O_2652,N_24704,N_24899);
xor UO_2653 (O_2653,N_24597,N_24489);
nand UO_2654 (O_2654,N_24799,N_24789);
or UO_2655 (O_2655,N_24384,N_24560);
and UO_2656 (O_2656,N_24929,N_24862);
xnor UO_2657 (O_2657,N_24519,N_24713);
or UO_2658 (O_2658,N_24639,N_24410);
nand UO_2659 (O_2659,N_24721,N_24823);
nor UO_2660 (O_2660,N_24896,N_24972);
or UO_2661 (O_2661,N_24595,N_24425);
nor UO_2662 (O_2662,N_24820,N_24979);
or UO_2663 (O_2663,N_24857,N_24926);
nor UO_2664 (O_2664,N_24380,N_24974);
xor UO_2665 (O_2665,N_24658,N_24706);
nand UO_2666 (O_2666,N_24730,N_24483);
xnor UO_2667 (O_2667,N_24436,N_24544);
and UO_2668 (O_2668,N_24442,N_24727);
and UO_2669 (O_2669,N_24712,N_24573);
or UO_2670 (O_2670,N_24899,N_24908);
or UO_2671 (O_2671,N_24911,N_24765);
nor UO_2672 (O_2672,N_24519,N_24939);
and UO_2673 (O_2673,N_24986,N_24792);
nand UO_2674 (O_2674,N_24668,N_24446);
or UO_2675 (O_2675,N_24407,N_24389);
nand UO_2676 (O_2676,N_24583,N_24561);
xor UO_2677 (O_2677,N_24636,N_24990);
nand UO_2678 (O_2678,N_24817,N_24562);
nor UO_2679 (O_2679,N_24872,N_24758);
nor UO_2680 (O_2680,N_24955,N_24621);
or UO_2681 (O_2681,N_24772,N_24687);
nor UO_2682 (O_2682,N_24824,N_24874);
nand UO_2683 (O_2683,N_24806,N_24699);
or UO_2684 (O_2684,N_24822,N_24423);
or UO_2685 (O_2685,N_24591,N_24579);
nand UO_2686 (O_2686,N_24398,N_24709);
nand UO_2687 (O_2687,N_24561,N_24794);
nor UO_2688 (O_2688,N_24405,N_24884);
xor UO_2689 (O_2689,N_24453,N_24685);
and UO_2690 (O_2690,N_24788,N_24626);
nor UO_2691 (O_2691,N_24985,N_24591);
nor UO_2692 (O_2692,N_24784,N_24816);
nand UO_2693 (O_2693,N_24700,N_24778);
and UO_2694 (O_2694,N_24461,N_24854);
nor UO_2695 (O_2695,N_24683,N_24648);
nor UO_2696 (O_2696,N_24381,N_24885);
and UO_2697 (O_2697,N_24566,N_24661);
nor UO_2698 (O_2698,N_24833,N_24385);
and UO_2699 (O_2699,N_24966,N_24758);
nand UO_2700 (O_2700,N_24715,N_24956);
and UO_2701 (O_2701,N_24399,N_24516);
or UO_2702 (O_2702,N_24823,N_24930);
nand UO_2703 (O_2703,N_24578,N_24562);
nor UO_2704 (O_2704,N_24490,N_24685);
and UO_2705 (O_2705,N_24796,N_24596);
nor UO_2706 (O_2706,N_24686,N_24481);
xor UO_2707 (O_2707,N_24746,N_24631);
or UO_2708 (O_2708,N_24611,N_24714);
or UO_2709 (O_2709,N_24586,N_24599);
nand UO_2710 (O_2710,N_24391,N_24594);
xnor UO_2711 (O_2711,N_24628,N_24407);
nor UO_2712 (O_2712,N_24800,N_24379);
xor UO_2713 (O_2713,N_24856,N_24665);
and UO_2714 (O_2714,N_24452,N_24929);
xor UO_2715 (O_2715,N_24816,N_24890);
xor UO_2716 (O_2716,N_24551,N_24820);
and UO_2717 (O_2717,N_24896,N_24767);
and UO_2718 (O_2718,N_24474,N_24854);
or UO_2719 (O_2719,N_24752,N_24500);
xor UO_2720 (O_2720,N_24875,N_24854);
nand UO_2721 (O_2721,N_24884,N_24474);
or UO_2722 (O_2722,N_24649,N_24899);
xor UO_2723 (O_2723,N_24832,N_24589);
nor UO_2724 (O_2724,N_24725,N_24763);
nand UO_2725 (O_2725,N_24597,N_24790);
nor UO_2726 (O_2726,N_24708,N_24534);
nor UO_2727 (O_2727,N_24699,N_24869);
xnor UO_2728 (O_2728,N_24605,N_24822);
and UO_2729 (O_2729,N_24410,N_24569);
xor UO_2730 (O_2730,N_24993,N_24892);
and UO_2731 (O_2731,N_24758,N_24487);
nand UO_2732 (O_2732,N_24818,N_24958);
and UO_2733 (O_2733,N_24854,N_24923);
xnor UO_2734 (O_2734,N_24981,N_24862);
or UO_2735 (O_2735,N_24382,N_24899);
nor UO_2736 (O_2736,N_24886,N_24577);
xor UO_2737 (O_2737,N_24937,N_24537);
xnor UO_2738 (O_2738,N_24405,N_24926);
nand UO_2739 (O_2739,N_24654,N_24634);
nand UO_2740 (O_2740,N_24661,N_24618);
or UO_2741 (O_2741,N_24696,N_24489);
nand UO_2742 (O_2742,N_24763,N_24527);
nand UO_2743 (O_2743,N_24477,N_24648);
and UO_2744 (O_2744,N_24453,N_24619);
or UO_2745 (O_2745,N_24864,N_24517);
and UO_2746 (O_2746,N_24973,N_24855);
and UO_2747 (O_2747,N_24445,N_24576);
and UO_2748 (O_2748,N_24607,N_24947);
and UO_2749 (O_2749,N_24888,N_24663);
nor UO_2750 (O_2750,N_24862,N_24805);
xor UO_2751 (O_2751,N_24601,N_24841);
nand UO_2752 (O_2752,N_24683,N_24972);
xnor UO_2753 (O_2753,N_24428,N_24969);
xor UO_2754 (O_2754,N_24382,N_24910);
nor UO_2755 (O_2755,N_24742,N_24968);
nor UO_2756 (O_2756,N_24693,N_24942);
xnor UO_2757 (O_2757,N_24433,N_24645);
xnor UO_2758 (O_2758,N_24609,N_24384);
or UO_2759 (O_2759,N_24689,N_24556);
nand UO_2760 (O_2760,N_24703,N_24645);
or UO_2761 (O_2761,N_24938,N_24478);
or UO_2762 (O_2762,N_24790,N_24584);
or UO_2763 (O_2763,N_24854,N_24612);
or UO_2764 (O_2764,N_24978,N_24735);
or UO_2765 (O_2765,N_24465,N_24764);
and UO_2766 (O_2766,N_24791,N_24861);
nor UO_2767 (O_2767,N_24692,N_24625);
and UO_2768 (O_2768,N_24546,N_24424);
nor UO_2769 (O_2769,N_24532,N_24740);
xnor UO_2770 (O_2770,N_24628,N_24500);
and UO_2771 (O_2771,N_24655,N_24612);
xnor UO_2772 (O_2772,N_24612,N_24667);
nor UO_2773 (O_2773,N_24471,N_24682);
nand UO_2774 (O_2774,N_24998,N_24641);
and UO_2775 (O_2775,N_24697,N_24874);
nand UO_2776 (O_2776,N_24380,N_24755);
nor UO_2777 (O_2777,N_24775,N_24583);
and UO_2778 (O_2778,N_24682,N_24661);
nand UO_2779 (O_2779,N_24620,N_24720);
nand UO_2780 (O_2780,N_24645,N_24583);
or UO_2781 (O_2781,N_24747,N_24965);
nand UO_2782 (O_2782,N_24532,N_24994);
or UO_2783 (O_2783,N_24559,N_24799);
xor UO_2784 (O_2784,N_24701,N_24465);
or UO_2785 (O_2785,N_24629,N_24722);
or UO_2786 (O_2786,N_24997,N_24994);
and UO_2787 (O_2787,N_24625,N_24519);
nand UO_2788 (O_2788,N_24657,N_24859);
nor UO_2789 (O_2789,N_24540,N_24424);
xnor UO_2790 (O_2790,N_24567,N_24518);
or UO_2791 (O_2791,N_24516,N_24808);
or UO_2792 (O_2792,N_24734,N_24397);
and UO_2793 (O_2793,N_24834,N_24674);
nor UO_2794 (O_2794,N_24678,N_24647);
and UO_2795 (O_2795,N_24587,N_24599);
or UO_2796 (O_2796,N_24758,N_24727);
or UO_2797 (O_2797,N_24604,N_24416);
and UO_2798 (O_2798,N_24607,N_24763);
and UO_2799 (O_2799,N_24709,N_24455);
nor UO_2800 (O_2800,N_24940,N_24723);
xnor UO_2801 (O_2801,N_24526,N_24729);
nor UO_2802 (O_2802,N_24456,N_24657);
xor UO_2803 (O_2803,N_24801,N_24549);
xnor UO_2804 (O_2804,N_24854,N_24754);
nand UO_2805 (O_2805,N_24982,N_24578);
nor UO_2806 (O_2806,N_24773,N_24667);
or UO_2807 (O_2807,N_24415,N_24638);
or UO_2808 (O_2808,N_24805,N_24521);
nand UO_2809 (O_2809,N_24888,N_24721);
and UO_2810 (O_2810,N_24819,N_24541);
nand UO_2811 (O_2811,N_24763,N_24921);
or UO_2812 (O_2812,N_24486,N_24489);
nand UO_2813 (O_2813,N_24707,N_24928);
nor UO_2814 (O_2814,N_24597,N_24764);
xnor UO_2815 (O_2815,N_24393,N_24722);
nor UO_2816 (O_2816,N_24884,N_24408);
nor UO_2817 (O_2817,N_24387,N_24546);
xnor UO_2818 (O_2818,N_24619,N_24415);
nand UO_2819 (O_2819,N_24686,N_24562);
or UO_2820 (O_2820,N_24553,N_24468);
or UO_2821 (O_2821,N_24762,N_24793);
nor UO_2822 (O_2822,N_24594,N_24690);
nor UO_2823 (O_2823,N_24781,N_24390);
and UO_2824 (O_2824,N_24467,N_24393);
xor UO_2825 (O_2825,N_24757,N_24404);
or UO_2826 (O_2826,N_24856,N_24976);
or UO_2827 (O_2827,N_24732,N_24718);
and UO_2828 (O_2828,N_24596,N_24409);
xor UO_2829 (O_2829,N_24540,N_24914);
and UO_2830 (O_2830,N_24932,N_24951);
xor UO_2831 (O_2831,N_24679,N_24411);
or UO_2832 (O_2832,N_24538,N_24834);
xnor UO_2833 (O_2833,N_24428,N_24690);
nor UO_2834 (O_2834,N_24515,N_24971);
or UO_2835 (O_2835,N_24601,N_24726);
and UO_2836 (O_2836,N_24582,N_24815);
or UO_2837 (O_2837,N_24532,N_24608);
and UO_2838 (O_2838,N_24818,N_24658);
nor UO_2839 (O_2839,N_24836,N_24681);
and UO_2840 (O_2840,N_24796,N_24787);
xnor UO_2841 (O_2841,N_24517,N_24393);
and UO_2842 (O_2842,N_24943,N_24704);
xor UO_2843 (O_2843,N_24769,N_24826);
nand UO_2844 (O_2844,N_24747,N_24441);
xor UO_2845 (O_2845,N_24861,N_24385);
or UO_2846 (O_2846,N_24623,N_24809);
nand UO_2847 (O_2847,N_24759,N_24978);
and UO_2848 (O_2848,N_24721,N_24959);
or UO_2849 (O_2849,N_24535,N_24517);
and UO_2850 (O_2850,N_24527,N_24740);
or UO_2851 (O_2851,N_24812,N_24636);
and UO_2852 (O_2852,N_24414,N_24812);
or UO_2853 (O_2853,N_24969,N_24979);
or UO_2854 (O_2854,N_24954,N_24618);
nand UO_2855 (O_2855,N_24962,N_24977);
nand UO_2856 (O_2856,N_24944,N_24961);
or UO_2857 (O_2857,N_24790,N_24837);
nand UO_2858 (O_2858,N_24759,N_24955);
nand UO_2859 (O_2859,N_24999,N_24601);
nor UO_2860 (O_2860,N_24824,N_24958);
or UO_2861 (O_2861,N_24429,N_24586);
xnor UO_2862 (O_2862,N_24987,N_24686);
xor UO_2863 (O_2863,N_24596,N_24710);
nand UO_2864 (O_2864,N_24782,N_24376);
nand UO_2865 (O_2865,N_24824,N_24682);
or UO_2866 (O_2866,N_24384,N_24406);
xor UO_2867 (O_2867,N_24608,N_24784);
or UO_2868 (O_2868,N_24905,N_24875);
and UO_2869 (O_2869,N_24534,N_24402);
nand UO_2870 (O_2870,N_24539,N_24632);
and UO_2871 (O_2871,N_24653,N_24715);
xnor UO_2872 (O_2872,N_24936,N_24502);
nand UO_2873 (O_2873,N_24449,N_24829);
nand UO_2874 (O_2874,N_24995,N_24554);
and UO_2875 (O_2875,N_24613,N_24988);
nand UO_2876 (O_2876,N_24741,N_24835);
xnor UO_2877 (O_2877,N_24725,N_24595);
nor UO_2878 (O_2878,N_24921,N_24481);
xor UO_2879 (O_2879,N_24894,N_24964);
or UO_2880 (O_2880,N_24976,N_24587);
and UO_2881 (O_2881,N_24974,N_24907);
nand UO_2882 (O_2882,N_24419,N_24430);
nand UO_2883 (O_2883,N_24659,N_24642);
xor UO_2884 (O_2884,N_24456,N_24735);
or UO_2885 (O_2885,N_24994,N_24847);
nand UO_2886 (O_2886,N_24878,N_24549);
xnor UO_2887 (O_2887,N_24790,N_24667);
xnor UO_2888 (O_2888,N_24864,N_24998);
or UO_2889 (O_2889,N_24871,N_24498);
and UO_2890 (O_2890,N_24554,N_24538);
or UO_2891 (O_2891,N_24945,N_24876);
nand UO_2892 (O_2892,N_24387,N_24988);
and UO_2893 (O_2893,N_24952,N_24709);
nand UO_2894 (O_2894,N_24780,N_24856);
nor UO_2895 (O_2895,N_24902,N_24555);
nand UO_2896 (O_2896,N_24894,N_24759);
nand UO_2897 (O_2897,N_24961,N_24608);
or UO_2898 (O_2898,N_24849,N_24590);
or UO_2899 (O_2899,N_24765,N_24518);
nand UO_2900 (O_2900,N_24703,N_24598);
or UO_2901 (O_2901,N_24617,N_24432);
xor UO_2902 (O_2902,N_24982,N_24493);
or UO_2903 (O_2903,N_24525,N_24627);
or UO_2904 (O_2904,N_24596,N_24921);
nand UO_2905 (O_2905,N_24696,N_24785);
xor UO_2906 (O_2906,N_24511,N_24656);
or UO_2907 (O_2907,N_24437,N_24511);
and UO_2908 (O_2908,N_24939,N_24905);
xnor UO_2909 (O_2909,N_24596,N_24566);
nand UO_2910 (O_2910,N_24405,N_24526);
and UO_2911 (O_2911,N_24908,N_24984);
xnor UO_2912 (O_2912,N_24578,N_24615);
and UO_2913 (O_2913,N_24506,N_24505);
xnor UO_2914 (O_2914,N_24518,N_24623);
or UO_2915 (O_2915,N_24459,N_24731);
and UO_2916 (O_2916,N_24540,N_24915);
nor UO_2917 (O_2917,N_24957,N_24523);
and UO_2918 (O_2918,N_24613,N_24698);
nor UO_2919 (O_2919,N_24432,N_24502);
and UO_2920 (O_2920,N_24834,N_24839);
and UO_2921 (O_2921,N_24620,N_24384);
or UO_2922 (O_2922,N_24785,N_24652);
or UO_2923 (O_2923,N_24716,N_24512);
or UO_2924 (O_2924,N_24996,N_24874);
nand UO_2925 (O_2925,N_24661,N_24996);
xnor UO_2926 (O_2926,N_24389,N_24564);
or UO_2927 (O_2927,N_24393,N_24602);
nand UO_2928 (O_2928,N_24635,N_24420);
or UO_2929 (O_2929,N_24901,N_24535);
or UO_2930 (O_2930,N_24881,N_24550);
xnor UO_2931 (O_2931,N_24603,N_24410);
nand UO_2932 (O_2932,N_24443,N_24416);
or UO_2933 (O_2933,N_24902,N_24581);
and UO_2934 (O_2934,N_24693,N_24765);
nor UO_2935 (O_2935,N_24845,N_24710);
nand UO_2936 (O_2936,N_24896,N_24791);
or UO_2937 (O_2937,N_24931,N_24659);
nor UO_2938 (O_2938,N_24915,N_24967);
and UO_2939 (O_2939,N_24619,N_24714);
nand UO_2940 (O_2940,N_24901,N_24642);
nor UO_2941 (O_2941,N_24985,N_24524);
nand UO_2942 (O_2942,N_24502,N_24956);
nand UO_2943 (O_2943,N_24802,N_24942);
nor UO_2944 (O_2944,N_24497,N_24459);
and UO_2945 (O_2945,N_24514,N_24631);
and UO_2946 (O_2946,N_24932,N_24399);
nand UO_2947 (O_2947,N_24670,N_24490);
nand UO_2948 (O_2948,N_24487,N_24472);
xor UO_2949 (O_2949,N_24993,N_24739);
or UO_2950 (O_2950,N_24474,N_24583);
xor UO_2951 (O_2951,N_24519,N_24630);
nor UO_2952 (O_2952,N_24378,N_24439);
nand UO_2953 (O_2953,N_24653,N_24377);
xor UO_2954 (O_2954,N_24541,N_24735);
xnor UO_2955 (O_2955,N_24473,N_24678);
or UO_2956 (O_2956,N_24849,N_24605);
or UO_2957 (O_2957,N_24384,N_24390);
nor UO_2958 (O_2958,N_24717,N_24979);
nand UO_2959 (O_2959,N_24998,N_24900);
nor UO_2960 (O_2960,N_24935,N_24553);
or UO_2961 (O_2961,N_24805,N_24530);
nor UO_2962 (O_2962,N_24599,N_24509);
or UO_2963 (O_2963,N_24974,N_24645);
or UO_2964 (O_2964,N_24419,N_24673);
nand UO_2965 (O_2965,N_24424,N_24771);
nand UO_2966 (O_2966,N_24581,N_24535);
and UO_2967 (O_2967,N_24766,N_24902);
and UO_2968 (O_2968,N_24866,N_24510);
xor UO_2969 (O_2969,N_24562,N_24636);
nor UO_2970 (O_2970,N_24396,N_24552);
nor UO_2971 (O_2971,N_24635,N_24829);
nand UO_2972 (O_2972,N_24759,N_24452);
nand UO_2973 (O_2973,N_24437,N_24888);
xor UO_2974 (O_2974,N_24549,N_24493);
nor UO_2975 (O_2975,N_24688,N_24602);
or UO_2976 (O_2976,N_24543,N_24718);
nand UO_2977 (O_2977,N_24889,N_24927);
nand UO_2978 (O_2978,N_24627,N_24558);
nor UO_2979 (O_2979,N_24540,N_24539);
nor UO_2980 (O_2980,N_24934,N_24421);
nor UO_2981 (O_2981,N_24640,N_24586);
nand UO_2982 (O_2982,N_24738,N_24927);
or UO_2983 (O_2983,N_24393,N_24466);
or UO_2984 (O_2984,N_24753,N_24607);
nand UO_2985 (O_2985,N_24644,N_24710);
or UO_2986 (O_2986,N_24937,N_24985);
and UO_2987 (O_2987,N_24587,N_24566);
nor UO_2988 (O_2988,N_24618,N_24541);
nor UO_2989 (O_2989,N_24719,N_24770);
nor UO_2990 (O_2990,N_24909,N_24424);
or UO_2991 (O_2991,N_24886,N_24998);
and UO_2992 (O_2992,N_24756,N_24505);
or UO_2993 (O_2993,N_24462,N_24636);
nor UO_2994 (O_2994,N_24925,N_24729);
or UO_2995 (O_2995,N_24825,N_24925);
nor UO_2996 (O_2996,N_24735,N_24611);
and UO_2997 (O_2997,N_24579,N_24506);
nand UO_2998 (O_2998,N_24713,N_24674);
xnor UO_2999 (O_2999,N_24597,N_24540);
endmodule