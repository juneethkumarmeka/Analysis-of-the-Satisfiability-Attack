module basic_5000_50000_5000_25_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_1913,In_3063);
nand U1 (N_1,In_3938,In_749);
and U2 (N_2,In_597,In_3706);
and U3 (N_3,In_1410,In_704);
and U4 (N_4,In_1645,In_846);
nand U5 (N_5,In_216,In_3034);
nand U6 (N_6,In_2553,In_3309);
nand U7 (N_7,In_2149,In_3766);
nand U8 (N_8,In_3590,In_4163);
and U9 (N_9,In_2727,In_1818);
and U10 (N_10,In_4180,In_1139);
or U11 (N_11,In_250,In_480);
and U12 (N_12,In_2249,In_4706);
and U13 (N_13,In_624,In_4078);
nor U14 (N_14,In_3612,In_1123);
nor U15 (N_15,In_1878,In_2737);
nor U16 (N_16,In_2011,In_3521);
or U17 (N_17,In_3893,In_1553);
or U18 (N_18,In_4900,In_3404);
or U19 (N_19,In_4841,In_2684);
and U20 (N_20,In_2225,In_3563);
nand U21 (N_21,In_2317,In_1971);
and U22 (N_22,In_877,In_1910);
and U23 (N_23,In_4452,In_3725);
nor U24 (N_24,In_765,In_2319);
nand U25 (N_25,In_809,In_3900);
nand U26 (N_26,In_4682,In_2241);
or U27 (N_27,In_806,In_4644);
nor U28 (N_28,In_3299,In_2117);
or U29 (N_29,In_3882,In_4342);
and U30 (N_30,In_4166,In_930);
or U31 (N_31,In_2924,In_581);
and U32 (N_32,In_4708,In_42);
nand U33 (N_33,In_2891,In_4361);
and U34 (N_34,In_4110,In_3949);
xor U35 (N_35,In_2393,In_1314);
nor U36 (N_36,In_4696,In_2356);
or U37 (N_37,In_131,In_570);
nand U38 (N_38,In_753,In_3175);
nand U39 (N_39,In_1790,In_3545);
and U40 (N_40,In_123,In_2299);
nand U41 (N_41,In_3977,In_2086);
or U42 (N_42,In_1125,In_3867);
or U43 (N_43,In_1666,In_4099);
or U44 (N_44,In_2640,In_650);
or U45 (N_45,In_226,In_4018);
nor U46 (N_46,In_4568,In_3961);
nor U47 (N_47,In_1531,In_4354);
or U48 (N_48,In_610,In_4924);
or U49 (N_49,In_155,In_3992);
nand U50 (N_50,In_1166,In_2040);
nor U51 (N_51,In_1954,In_4135);
and U52 (N_52,In_2108,In_3744);
or U53 (N_53,In_1029,In_2754);
nor U54 (N_54,In_4829,In_4407);
nor U55 (N_55,In_3380,In_3814);
or U56 (N_56,In_3671,In_455);
nand U57 (N_57,In_3476,In_4022);
nor U58 (N_58,In_1179,In_1220);
or U59 (N_59,In_1068,In_4273);
and U60 (N_60,In_447,In_834);
nand U61 (N_61,In_2302,In_3005);
or U62 (N_62,In_2632,In_4119);
xor U63 (N_63,In_4676,In_492);
nand U64 (N_64,In_2325,In_2758);
and U65 (N_65,In_1981,In_1821);
or U66 (N_66,In_1258,In_2238);
nor U67 (N_67,In_4126,In_456);
nor U68 (N_68,In_2017,In_4425);
and U69 (N_69,In_4510,In_3548);
or U70 (N_70,In_2267,In_4859);
nor U71 (N_71,In_3734,In_65);
nor U72 (N_72,In_1849,In_2967);
nor U73 (N_73,In_781,In_3733);
or U74 (N_74,In_2699,In_502);
nand U75 (N_75,In_2045,In_1902);
nand U76 (N_76,In_2196,In_4581);
xnor U77 (N_77,In_2500,In_2425);
nor U78 (N_78,In_4797,In_579);
and U79 (N_79,In_3060,In_4551);
and U80 (N_80,In_1988,In_1586);
xor U81 (N_81,In_4516,In_2839);
and U82 (N_82,In_2170,In_3057);
nand U83 (N_83,In_4220,In_2979);
nand U84 (N_84,In_1593,In_1338);
nand U85 (N_85,In_3362,In_3340);
nand U86 (N_86,In_490,In_3341);
nor U87 (N_87,In_1128,In_2601);
nand U88 (N_88,In_1377,In_3004);
nand U89 (N_89,In_184,In_3209);
nor U90 (N_90,In_1236,In_4184);
and U91 (N_91,In_3518,In_3071);
or U92 (N_92,In_1490,In_1566);
and U93 (N_93,In_2949,In_4803);
and U94 (N_94,In_1898,In_1329);
nor U95 (N_95,In_3845,In_4420);
and U96 (N_96,In_1004,In_2157);
nand U97 (N_97,In_1079,In_3604);
and U98 (N_98,In_4573,In_4497);
nor U99 (N_99,In_3651,In_754);
and U100 (N_100,In_2387,In_873);
nor U101 (N_101,In_305,In_3935);
and U102 (N_102,In_576,In_395);
or U103 (N_103,In_3931,In_3825);
or U104 (N_104,In_891,In_318);
or U105 (N_105,In_2687,In_2043);
nor U106 (N_106,In_1016,In_3033);
nand U107 (N_107,In_371,In_3278);
and U108 (N_108,In_2051,In_1134);
and U109 (N_109,In_4403,In_516);
and U110 (N_110,In_1609,In_4316);
and U111 (N_111,In_4123,In_1114);
or U112 (N_112,In_620,In_1056);
nor U113 (N_113,In_384,In_279);
and U114 (N_114,In_2852,In_427);
and U115 (N_115,In_2643,In_1729);
and U116 (N_116,In_828,In_4784);
or U117 (N_117,In_4097,In_565);
and U118 (N_118,In_2923,In_2571);
and U119 (N_119,In_980,In_1953);
and U120 (N_120,In_2012,In_3003);
nor U121 (N_121,In_2429,In_3121);
and U122 (N_122,In_888,In_3602);
xor U123 (N_123,In_605,In_908);
nand U124 (N_124,In_4824,In_3660);
or U125 (N_125,In_665,In_402);
and U126 (N_126,In_2840,In_1630);
or U127 (N_127,In_2811,In_721);
nor U128 (N_128,In_4592,In_2195);
nor U129 (N_129,In_3317,In_2194);
nor U130 (N_130,In_473,In_2123);
nor U131 (N_131,In_2185,In_2879);
and U132 (N_132,In_3874,In_2420);
nor U133 (N_133,In_2791,In_3011);
nand U134 (N_134,In_3617,In_1570);
or U135 (N_135,In_160,In_3286);
nand U136 (N_136,In_2728,In_4986);
or U137 (N_137,In_1170,In_3042);
nor U138 (N_138,In_643,In_990);
nor U139 (N_139,In_4225,In_14);
nand U140 (N_140,In_1028,In_4241);
nor U141 (N_141,In_3635,In_4256);
xor U142 (N_142,In_4515,In_946);
and U143 (N_143,In_1797,In_4002);
nand U144 (N_144,In_1775,In_4858);
or U145 (N_145,In_3141,In_2853);
nor U146 (N_146,In_4437,In_1538);
and U147 (N_147,In_1425,In_3124);
nand U148 (N_148,In_2039,In_2454);
nor U149 (N_149,In_2602,In_718);
and U150 (N_150,In_1023,In_334);
and U151 (N_151,In_989,In_3339);
nand U152 (N_152,In_1416,In_2898);
xor U153 (N_153,In_4338,In_2616);
or U154 (N_154,In_2714,In_4199);
nor U155 (N_155,In_4766,In_2071);
nand U156 (N_156,In_4650,In_4266);
and U157 (N_157,In_2162,In_4961);
nand U158 (N_158,In_4206,In_159);
and U159 (N_159,In_276,In_2237);
nand U160 (N_160,In_3843,In_3074);
nand U161 (N_161,In_2872,In_3085);
nor U162 (N_162,In_3271,In_2215);
and U163 (N_163,In_2802,In_1649);
nor U164 (N_164,In_3139,In_4976);
and U165 (N_165,In_3966,In_2257);
or U166 (N_166,In_3098,In_1861);
nand U167 (N_167,In_1247,In_3592);
nand U168 (N_168,In_4419,In_4202);
xor U169 (N_169,In_4536,In_4312);
and U170 (N_170,In_4805,In_2207);
nor U171 (N_171,In_2966,In_603);
nand U172 (N_172,In_1762,In_2513);
nor U173 (N_173,In_1640,In_4363);
nand U174 (N_174,In_763,In_2491);
nor U175 (N_175,In_2175,In_2389);
nor U176 (N_176,In_513,In_975);
nand U177 (N_177,In_1401,In_3081);
xor U178 (N_178,In_2764,In_4004);
and U179 (N_179,In_2540,In_1669);
nor U180 (N_180,In_4382,In_2153);
and U181 (N_181,In_1826,In_938);
nor U182 (N_182,In_1869,In_582);
nor U183 (N_183,In_4869,In_1443);
nor U184 (N_184,In_3409,In_774);
and U185 (N_185,In_1422,In_4728);
xor U186 (N_186,In_4144,In_769);
nor U187 (N_187,In_2470,In_2069);
xor U188 (N_188,In_274,In_429);
nor U189 (N_189,In_2573,In_3760);
nor U190 (N_190,In_3572,In_1646);
and U191 (N_191,In_3956,In_2329);
xor U192 (N_192,In_1486,In_3815);
nand U193 (N_193,In_2283,In_810);
xnor U194 (N_194,In_1169,In_1828);
and U195 (N_195,In_127,In_3386);
nor U196 (N_196,In_3586,In_2064);
nor U197 (N_197,In_375,In_2461);
and U198 (N_198,In_1096,In_3072);
nor U199 (N_199,In_1484,In_4449);
nor U200 (N_200,In_895,In_3125);
or U201 (N_201,In_3377,In_4946);
and U202 (N_202,In_2368,In_1381);
nor U203 (N_203,In_521,In_4128);
nor U204 (N_204,In_567,In_4814);
or U205 (N_205,In_4487,In_4084);
or U206 (N_206,In_4998,In_1000);
or U207 (N_207,In_2845,In_4461);
and U208 (N_208,In_923,In_3629);
or U209 (N_209,In_1834,In_4246);
and U210 (N_210,In_1843,In_2630);
nand U211 (N_211,In_3305,In_1058);
or U212 (N_212,In_2925,In_3359);
xnor U213 (N_213,In_1823,In_1944);
and U214 (N_214,In_709,In_4102);
nand U215 (N_215,In_147,In_3023);
nor U216 (N_216,In_4656,In_2280);
and U217 (N_217,In_3922,In_4029);
and U218 (N_218,In_4164,In_2200);
xor U219 (N_219,In_1983,In_3254);
nor U220 (N_220,In_333,In_1868);
nor U221 (N_221,In_1812,In_1810);
and U222 (N_222,In_3414,In_3390);
nor U223 (N_223,In_3801,In_3226);
and U224 (N_224,In_2413,In_3043);
and U225 (N_225,In_3749,In_2642);
or U226 (N_226,In_4271,In_3691);
nand U227 (N_227,In_4935,In_3566);
or U228 (N_228,In_437,In_547);
or U229 (N_229,In_601,In_573);
nand U230 (N_230,In_972,In_3864);
nor U231 (N_231,In_3995,In_525);
and U232 (N_232,In_1282,In_4741);
and U233 (N_233,In_3703,In_4721);
nand U234 (N_234,In_2761,In_3046);
and U235 (N_235,In_4735,In_1995);
and U236 (N_236,In_4776,In_3841);
nand U237 (N_237,In_1431,In_4325);
and U238 (N_238,In_345,In_2219);
or U239 (N_239,In_2530,In_2133);
or U240 (N_240,In_741,In_3649);
or U241 (N_241,In_1288,In_3147);
nor U242 (N_242,In_1697,In_2469);
and U243 (N_243,In_1848,In_4168);
or U244 (N_244,In_4103,In_4816);
nand U245 (N_245,In_3668,In_2965);
nand U246 (N_246,In_1200,In_3818);
nand U247 (N_247,In_1005,In_3120);
nand U248 (N_248,In_532,In_2772);
or U249 (N_249,In_3876,In_4218);
or U250 (N_250,In_4445,In_1514);
xor U251 (N_251,In_2386,In_2474);
nand U252 (N_252,In_2375,In_1477);
nor U253 (N_253,In_4229,In_2326);
or U254 (N_254,In_1842,In_3675);
nor U255 (N_255,In_2908,In_1735);
nor U256 (N_256,In_2910,In_1598);
or U257 (N_257,In_2999,In_1015);
or U258 (N_258,In_331,In_2574);
and U259 (N_259,In_1793,In_381);
nand U260 (N_260,In_2141,In_1487);
and U261 (N_261,In_4739,In_2255);
nand U262 (N_262,In_2460,In_352);
or U263 (N_263,In_1440,In_178);
or U264 (N_264,In_1672,In_4075);
nor U265 (N_265,In_4709,In_3556);
or U266 (N_266,In_1002,In_3947);
xnor U267 (N_267,In_394,In_454);
nor U268 (N_268,In_1458,In_1313);
or U269 (N_269,In_901,In_3806);
or U270 (N_270,In_2430,In_1689);
nor U271 (N_271,In_3086,In_2948);
or U272 (N_272,In_3245,In_315);
and U273 (N_273,In_4173,In_1625);
or U274 (N_274,In_684,In_974);
nand U275 (N_275,In_4379,In_2973);
or U276 (N_276,In_2408,In_4888);
and U277 (N_277,In_180,In_1069);
and U278 (N_278,In_4506,In_4092);
nor U279 (N_279,In_1081,In_3070);
nand U280 (N_280,In_118,In_778);
or U281 (N_281,In_4021,In_3415);
and U282 (N_282,In_1164,In_1695);
or U283 (N_283,In_947,In_1774);
and U284 (N_284,In_1523,In_1432);
nor U285 (N_285,In_365,In_3450);
nand U286 (N_286,In_2247,In_324);
nand U287 (N_287,In_3458,In_1363);
nand U288 (N_288,In_1582,In_319);
nor U289 (N_289,In_858,In_3579);
or U290 (N_290,In_3597,In_2639);
and U291 (N_291,In_418,In_4504);
nand U292 (N_292,In_2376,In_3988);
nand U293 (N_293,In_1732,In_146);
nor U294 (N_294,In_3007,In_692);
and U295 (N_295,In_3606,In_770);
or U296 (N_296,In_3804,In_1102);
nand U297 (N_297,In_2036,In_1393);
nor U298 (N_298,In_4606,In_3748);
and U299 (N_299,In_2310,In_4632);
and U300 (N_300,In_3029,In_3670);
or U301 (N_301,In_896,In_4386);
and U302 (N_302,In_3270,In_949);
or U303 (N_303,In_2349,In_3443);
nor U304 (N_304,In_4699,In_284);
xor U305 (N_305,In_840,In_585);
and U306 (N_306,In_2323,In_3395);
nor U307 (N_307,In_4687,In_3530);
or U308 (N_308,In_831,In_3625);
and U309 (N_309,In_4901,In_4547);
and U310 (N_310,In_3231,In_849);
nor U311 (N_311,In_4411,In_2077);
xnor U312 (N_312,In_54,In_4183);
and U313 (N_313,In_3354,In_1932);
or U314 (N_314,In_2937,In_1550);
and U315 (N_315,In_1891,In_2516);
nand U316 (N_316,In_4391,In_3439);
nand U317 (N_317,In_1442,In_3911);
or U318 (N_318,In_1737,In_4850);
nor U319 (N_319,In_3520,In_2277);
and U320 (N_320,In_2384,In_1070);
or U321 (N_321,In_1364,In_2385);
nor U322 (N_322,In_2066,In_2807);
nor U323 (N_323,In_4886,In_1623);
and U324 (N_324,In_4340,In_1294);
and U325 (N_325,In_1872,In_182);
or U326 (N_326,In_2997,In_618);
nand U327 (N_327,In_1936,In_2274);
or U328 (N_328,In_512,In_2677);
nand U329 (N_329,In_733,In_1610);
or U330 (N_330,In_2822,In_820);
and U331 (N_331,In_4619,In_2477);
nor U332 (N_332,In_3408,In_4100);
nand U333 (N_333,In_4681,In_385);
nand U334 (N_334,In_2832,In_3393);
or U335 (N_335,In_2855,In_1138);
and U336 (N_336,In_3092,In_481);
nor U337 (N_337,In_3713,In_3319);
and U338 (N_338,In_3097,In_57);
nand U339 (N_339,In_166,In_2498);
or U340 (N_340,In_2786,In_2662);
and U341 (N_341,In_784,In_2611);
or U342 (N_342,In_4618,In_1186);
and U343 (N_343,In_1827,In_4336);
nand U344 (N_344,In_4863,In_1307);
xor U345 (N_345,In_2447,In_3334);
or U346 (N_346,In_286,In_2109);
nand U347 (N_347,In_2971,In_4343);
and U348 (N_348,In_878,In_4137);
and U349 (N_349,In_4170,In_4518);
xnor U350 (N_350,In_4280,In_3819);
nand U351 (N_351,In_4413,In_4570);
nand U352 (N_352,In_1185,In_86);
and U353 (N_353,In_4447,In_2496);
nor U354 (N_354,In_4066,In_882);
nand U355 (N_355,In_2179,In_1305);
and U356 (N_356,In_4494,In_1112);
nand U357 (N_357,In_1092,In_3784);
or U358 (N_358,In_3182,In_674);
nor U359 (N_359,In_3083,In_1206);
xor U360 (N_360,In_3471,In_1730);
nor U361 (N_361,In_2111,In_1304);
nor U362 (N_362,In_920,In_1345);
and U363 (N_363,In_970,In_1342);
or U364 (N_364,In_3161,In_3907);
and U365 (N_365,In_4118,In_1783);
or U366 (N_366,In_1333,In_3179);
and U367 (N_367,In_4085,In_3901);
or U368 (N_368,In_804,In_2236);
and U369 (N_369,In_4615,In_3553);
nand U370 (N_370,In_1951,In_561);
or U371 (N_371,In_1309,In_986);
and U372 (N_372,In_392,In_3402);
or U373 (N_373,In_759,In_41);
nand U374 (N_374,In_2027,In_3381);
or U375 (N_375,In_4251,In_2691);
or U376 (N_376,In_4833,In_637);
nor U377 (N_377,In_737,In_4716);
nand U378 (N_378,In_4275,In_983);
and U379 (N_379,In_3378,In_3432);
nand U380 (N_380,In_2,In_808);
or U381 (N_381,In_4378,In_4553);
xnor U382 (N_382,In_3306,In_1573);
nand U383 (N_383,In_4769,In_3202);
nor U384 (N_384,In_1167,In_4595);
nand U385 (N_385,In_1038,In_1986);
and U386 (N_386,In_3879,In_4427);
nand U387 (N_387,In_4959,In_1963);
nor U388 (N_388,In_4471,In_3795);
nand U389 (N_389,In_3477,In_2768);
nor U390 (N_390,In_2667,In_641);
and U391 (N_391,In_836,In_1297);
nor U392 (N_392,In_3420,In_4952);
nor U393 (N_393,In_1779,In_4817);
nor U394 (N_394,In_2259,In_4056);
and U395 (N_395,In_1929,In_3412);
and U396 (N_396,In_706,In_1060);
or U397 (N_397,In_4559,In_4594);
and U398 (N_398,In_2294,In_4027);
nor U399 (N_399,In_1895,In_1500);
or U400 (N_400,In_224,In_1419);
or U401 (N_401,In_823,In_4300);
and U402 (N_402,In_4171,In_3037);
or U403 (N_403,In_4995,In_3573);
nor U404 (N_404,In_1962,In_2929);
nand U405 (N_405,In_3677,In_1133);
or U406 (N_406,In_3866,In_2909);
nand U407 (N_407,In_3564,In_803);
xor U408 (N_408,In_3054,In_3982);
nand U409 (N_409,In_664,In_571);
nor U410 (N_410,In_1360,In_3969);
and U411 (N_411,In_4867,In_4459);
or U412 (N_412,In_5,In_3908);
nand U413 (N_413,In_855,In_3383);
nor U414 (N_414,In_2140,In_1569);
and U415 (N_415,In_1160,In_4667);
or U416 (N_416,In_1720,In_1927);
nor U417 (N_417,In_3645,In_1077);
and U418 (N_418,In_4422,In_1466);
nand U419 (N_419,In_3773,In_3533);
nor U420 (N_420,In_4645,In_380);
nor U421 (N_421,In_2715,In_2799);
nor U422 (N_422,In_3075,In_97);
nor U423 (N_423,In_1704,In_4605);
nor U424 (N_424,In_4042,In_4418);
or U425 (N_425,In_241,In_4598);
xnor U426 (N_426,In_837,In_921);
or U427 (N_427,In_3160,In_4834);
nand U428 (N_428,In_4724,In_646);
and U429 (N_429,In_3561,In_711);
or U430 (N_430,In_2049,In_157);
nor U431 (N_431,In_2324,In_2865);
and U432 (N_432,In_3942,In_2483);
and U433 (N_433,In_648,In_2838);
nand U434 (N_434,In_4177,In_1187);
xnor U435 (N_435,In_1208,In_4450);
and U436 (N_436,In_2673,In_3392);
xor U437 (N_437,In_1350,In_4194);
or U438 (N_438,In_1674,In_3345);
or U439 (N_439,In_3536,In_2378);
and U440 (N_440,In_262,In_4302);
and U441 (N_441,In_3473,In_417);
nor U442 (N_442,In_3501,In_604);
nand U443 (N_443,In_2619,In_841);
and U444 (N_444,In_3376,In_1923);
or U445 (N_445,In_145,In_4521);
nor U446 (N_446,In_4691,In_4399);
or U447 (N_447,In_557,In_2345);
and U448 (N_448,In_232,In_2969);
and U449 (N_449,In_444,In_2655);
and U450 (N_450,In_944,In_1822);
and U451 (N_451,In_657,In_2856);
or U452 (N_452,In_1014,In_4830);
or U453 (N_453,In_2796,In_1462);
or U454 (N_454,In_296,In_3531);
or U455 (N_455,In_534,In_2980);
nor U456 (N_456,In_2636,In_277);
nand U457 (N_457,In_3246,In_3827);
or U458 (N_458,In_3877,In_2557);
nand U459 (N_459,In_669,In_1232);
nor U460 (N_460,In_2493,In_1745);
nor U461 (N_461,In_4713,In_3019);
or U462 (N_462,In_3756,In_1964);
nor U463 (N_463,In_3131,In_423);
nor U464 (N_464,In_4988,In_4496);
or U465 (N_465,In_3030,In_707);
or U466 (N_466,In_788,In_4941);
or U467 (N_467,In_1412,In_3541);
or U468 (N_468,In_1694,In_2016);
and U469 (N_469,In_4908,In_1990);
nand U470 (N_470,In_1652,In_504);
or U471 (N_471,In_796,In_676);
and U472 (N_472,In_71,In_2223);
and U473 (N_473,In_4428,In_1839);
nor U474 (N_474,In_971,In_4871);
nor U475 (N_475,In_2970,In_2455);
nor U476 (N_476,In_1676,In_4937);
nand U477 (N_477,In_144,In_863);
and U478 (N_478,In_3224,In_2962);
and U479 (N_479,In_967,In_3574);
nor U480 (N_480,In_2563,In_4893);
nor U481 (N_481,In_1083,In_3027);
and U482 (N_482,In_1103,In_2887);
nor U483 (N_483,In_3682,In_3021);
or U484 (N_484,In_4324,In_3335);
or U485 (N_485,In_1811,In_2180);
and U486 (N_486,In_63,In_2607);
and U487 (N_487,In_1271,In_2809);
and U488 (N_488,In_4083,In_716);
nand U489 (N_489,In_1966,In_1244);
nand U490 (N_490,In_2138,In_2777);
nor U491 (N_491,In_1925,In_730);
or U492 (N_492,In_2090,In_1300);
and U493 (N_493,In_11,In_1837);
or U494 (N_494,In_2927,In_4621);
or U495 (N_495,In_3616,In_2703);
or U496 (N_496,In_2047,In_2952);
xor U497 (N_497,In_1135,In_406);
nor U498 (N_498,In_4740,In_389);
and U499 (N_499,In_4050,In_1389);
or U500 (N_500,In_1568,In_461);
and U501 (N_501,In_2650,In_2148);
nand U502 (N_502,In_2188,In_4371);
nand U503 (N_503,In_3885,In_4195);
nand U504 (N_504,In_4370,In_2057);
or U505 (N_505,In_3109,In_1930);
nor U506 (N_506,In_2472,In_338);
and U507 (N_507,In_4744,In_1600);
nor U508 (N_508,In_1054,In_235);
nand U509 (N_509,In_386,In_48);
or U510 (N_510,In_4526,In_4252);
and U511 (N_511,In_1158,In_3314);
nand U512 (N_512,In_1259,In_963);
and U513 (N_513,In_1887,In_4082);
and U514 (N_514,In_2436,In_261);
or U515 (N_515,In_544,In_4658);
nor U516 (N_516,In_3106,In_2450);
nor U517 (N_517,In_3778,In_1948);
or U518 (N_518,In_2533,In_4971);
nand U519 (N_519,In_3599,In_2785);
nor U520 (N_520,In_4774,In_1620);
nor U521 (N_521,In_3078,In_961);
or U522 (N_522,In_2334,In_1603);
nand U523 (N_523,In_1888,In_619);
and U524 (N_524,In_8,In_2261);
or U525 (N_525,In_3687,In_1257);
or U526 (N_526,In_3761,In_1973);
nand U527 (N_527,In_4040,In_1606);
or U528 (N_528,In_1760,In_835);
and U529 (N_529,In_644,In_1883);
or U530 (N_530,In_1544,In_675);
nor U531 (N_531,In_1238,In_2549);
nand U532 (N_532,In_2102,In_1789);
nand U533 (N_533,In_1065,In_2348);
nor U534 (N_534,In_317,In_2921);
or U535 (N_535,In_2930,In_668);
or U536 (N_536,In_1939,In_1648);
nor U537 (N_537,In_4599,In_1773);
or U538 (N_538,In_4695,In_1701);
nand U539 (N_539,In_2217,In_3844);
nor U540 (N_540,In_4239,In_149);
or U541 (N_541,In_4561,In_1190);
nand U542 (N_542,In_397,In_3559);
nand U543 (N_543,In_1692,In_1153);
nor U544 (N_544,In_3379,In_660);
or U545 (N_545,In_3052,In_4485);
and U546 (N_546,In_4139,In_2441);
and U547 (N_547,In_3002,In_1332);
and U548 (N_548,In_526,In_3132);
nor U549 (N_549,In_3917,In_4393);
nand U550 (N_550,In_3688,In_4141);
nor U551 (N_551,In_3111,In_1243);
or U552 (N_552,In_1261,In_1835);
or U553 (N_553,In_4479,In_851);
or U554 (N_554,In_4512,In_3297);
and U555 (N_555,In_4567,In_4622);
nor U556 (N_556,In_1358,In_1520);
xnor U557 (N_557,In_2951,In_2362);
or U558 (N_558,In_459,In_3102);
nor U559 (N_559,In_3394,In_1357);
or U560 (N_560,In_2744,In_2333);
and U561 (N_561,In_3720,In_926);
or U562 (N_562,In_3350,In_3262);
nand U563 (N_563,In_2978,In_779);
and U564 (N_564,In_4910,In_3697);
or U565 (N_565,In_4238,In_4294);
and U566 (N_566,In_3483,In_4453);
and U567 (N_567,In_4023,In_2070);
nand U568 (N_568,In_1885,In_1859);
nand U569 (N_569,In_3562,In_4702);
xor U570 (N_570,In_1525,In_2269);
or U571 (N_571,In_4198,In_3594);
nand U572 (N_572,In_4074,In_2305);
and U573 (N_573,In_3035,In_4675);
or U574 (N_574,In_413,In_3049);
nand U575 (N_575,In_1050,In_4111);
or U576 (N_576,In_1146,In_1884);
nand U577 (N_577,In_3100,In_2087);
or U578 (N_578,In_1734,In_1693);
nor U579 (N_579,In_1998,In_4914);
nor U580 (N_580,In_283,In_3329);
or U581 (N_581,In_2000,In_2848);
and U582 (N_582,In_3516,In_1651);
and U583 (N_583,In_4410,In_1549);
nand U584 (N_584,In_2416,In_399);
and U585 (N_585,In_70,In_2186);
nand U586 (N_586,In_4764,In_1752);
and U587 (N_587,In_203,In_1177);
nand U588 (N_588,In_2230,In_1479);
nor U589 (N_589,In_213,In_3356);
and U590 (N_590,In_3837,In_3967);
and U591 (N_591,In_1503,In_4038);
nor U592 (N_592,In_1595,In_3462);
and U593 (N_593,In_422,In_1473);
and U594 (N_594,In_3515,In_2943);
xor U595 (N_595,In_3360,In_4307);
xor U596 (N_596,In_622,In_3847);
nor U597 (N_597,In_3899,In_121);
or U598 (N_598,In_1414,In_3852);
and U599 (N_599,In_1143,In_1560);
nand U600 (N_600,In_2263,In_4680);
nand U601 (N_601,In_3603,In_1162);
or U602 (N_602,In_4114,In_4781);
and U603 (N_603,In_1911,In_469);
nand U604 (N_604,In_4353,In_2287);
and U605 (N_605,In_1691,In_4319);
or U606 (N_606,In_77,In_4788);
nor U607 (N_607,In_4439,In_1088);
and U608 (N_608,In_4255,In_3783);
nand U609 (N_609,In_1742,In_4041);
nor U610 (N_610,In_1303,In_2944);
or U611 (N_611,In_2256,In_4243);
nand U612 (N_612,In_3767,In_398);
xnor U613 (N_613,In_3229,In_786);
and U614 (N_614,In_2189,In_4253);
nor U615 (N_615,In_3405,In_4);
xnor U616 (N_616,In_859,In_4013);
nand U617 (N_617,In_631,In_1537);
or U618 (N_618,In_3351,In_1295);
or U619 (N_619,In_3740,In_4564);
and U620 (N_620,In_2360,In_3282);
nor U621 (N_621,In_2351,In_4778);
nand U622 (N_622,In_2272,In_931);
nor U623 (N_623,In_24,In_2245);
and U624 (N_624,In_4943,In_1912);
or U625 (N_625,In_4854,In_4067);
and U626 (N_626,In_1421,In_2697);
nand U627 (N_627,In_4938,In_1008);
nand U628 (N_628,In_3940,In_25);
nand U629 (N_629,In_2605,In_498);
nor U630 (N_630,In_2812,In_4532);
or U631 (N_631,In_4355,In_4763);
nand U632 (N_632,In_1637,In_518);
nand U633 (N_633,In_3352,In_1627);
or U634 (N_634,In_2733,In_2331);
or U635 (N_635,In_2633,In_2851);
nor U636 (N_636,In_2358,In_114);
or U637 (N_637,In_440,In_4210);
nor U638 (N_638,In_1831,In_3508);
or U639 (N_639,In_1084,In_2866);
nand U640 (N_640,In_1985,In_2537);
and U641 (N_641,In_4899,In_2723);
or U642 (N_642,In_2289,In_3364);
nor U643 (N_643,In_690,In_2211);
and U644 (N_644,In_1063,In_826);
or U645 (N_645,In_916,In_4426);
nand U646 (N_646,In_3509,In_3156);
nor U647 (N_647,In_2284,In_4897);
nand U648 (N_648,In_2964,In_3872);
and U649 (N_649,In_3526,In_4727);
nor U650 (N_650,In_2410,In_81);
and U651 (N_651,In_4073,In_2320);
and U652 (N_652,In_4033,In_4604);
or U653 (N_653,In_1334,In_2411);
or U654 (N_654,In_3628,In_376);
nand U655 (N_655,In_4076,In_2176);
xnor U656 (N_656,In_409,In_1682);
or U657 (N_657,In_1508,In_542);
and U658 (N_658,In_1025,In_2880);
and U659 (N_659,In_1279,In_568);
or U660 (N_660,In_3895,In_2092);
nand U661 (N_661,In_2592,In_3567);
nand U662 (N_662,In_4907,In_4648);
nor U663 (N_663,In_3537,In_4558);
and U664 (N_664,In_3388,In_903);
nor U665 (N_665,In_2704,In_238);
and U666 (N_666,In_4654,In_2304);
nor U667 (N_667,In_4563,In_727);
nor U668 (N_668,In_2110,In_120);
nor U669 (N_669,In_2377,In_4096);
or U670 (N_670,In_3884,In_4969);
xnor U671 (N_671,In_2243,In_1534);
or U672 (N_672,In_4237,In_2395);
nand U673 (N_673,In_2452,In_647);
xnor U674 (N_674,In_3490,In_1631);
nor U675 (N_675,In_2649,In_3173);
nor U676 (N_676,In_2591,In_2318);
nor U677 (N_677,In_190,In_1);
nand U678 (N_678,In_1850,In_3241);
nand U679 (N_679,In_2020,In_1254);
or U680 (N_680,In_3644,In_2803);
nor U681 (N_681,In_3913,In_939);
nor U682 (N_682,In_2945,In_2264);
xor U683 (N_683,In_4326,In_230);
nand U684 (N_684,In_2757,In_1908);
and U685 (N_685,In_4468,In_1189);
nor U686 (N_686,In_3225,In_2747);
nand U687 (N_687,In_507,In_37);
nand U688 (N_688,In_549,In_875);
and U689 (N_689,In_2152,In_985);
and U690 (N_690,In_2031,In_134);
nand U691 (N_691,In_468,In_2023);
or U692 (N_692,In_4396,In_3674);
nand U693 (N_693,In_3145,In_252);
or U694 (N_694,In_2831,In_548);
or U695 (N_695,In_4875,In_2829);
nor U696 (N_696,In_595,In_171);
and U697 (N_697,In_3919,In_388);
nand U698 (N_698,In_1324,In_3803);
or U699 (N_699,In_2725,In_2850);
or U700 (N_700,In_1504,In_4647);
or U701 (N_701,In_752,In_4975);
or U702 (N_702,In_2403,In_2079);
nand U703 (N_703,In_2167,In_3860);
nand U704 (N_704,In_4322,In_3168);
nand U705 (N_705,In_2379,In_1352);
nor U706 (N_706,In_3717,In_1758);
and U707 (N_707,In_2212,In_2629);
xnor U708 (N_708,In_1563,In_4600);
nor U709 (N_709,In_1751,In_2499);
nand U710 (N_710,In_4154,In_3869);
and U711 (N_711,In_2506,In_3365);
and U712 (N_712,In_2844,In_2805);
and U713 (N_713,In_1235,In_2572);
nand U714 (N_714,In_819,In_2099);
or U715 (N_715,In_865,In_766);
nand U716 (N_716,In_9,In_3044);
nor U717 (N_717,In_1996,In_1870);
nand U718 (N_718,In_59,In_4248);
nand U719 (N_719,In_897,In_2801);
nor U720 (N_720,In_3730,In_4991);
nand U721 (N_721,In_950,In_2718);
nand U722 (N_722,In_4917,In_4134);
or U723 (N_723,In_2448,In_4513);
and U724 (N_724,In_3684,In_1914);
nand U725 (N_725,In_3082,In_3469);
nand U726 (N_726,In_535,In_4780);
or U727 (N_727,In_1857,In_4247);
and U728 (N_728,In_2372,In_2906);
or U729 (N_729,In_3252,In_4463);
nor U730 (N_730,In_4362,In_4809);
and U731 (N_731,In_3496,In_3708);
nand U732 (N_732,In_4531,In_4845);
nand U733 (N_733,In_1091,In_1249);
or U734 (N_734,In_2072,In_3172);
nand U735 (N_735,In_4523,In_948);
nand U736 (N_736,In_2489,In_4757);
and U737 (N_737,In_3024,In_3600);
and U738 (N_738,In_4348,In_2531);
nor U739 (N_739,In_4148,In_964);
or U740 (N_740,In_4839,In_3930);
nand U741 (N_741,In_2584,In_3608);
nor U742 (N_742,In_3332,In_3823);
and U743 (N_743,In_320,In_702);
nand U744 (N_744,In_3292,In_1740);
and U745 (N_745,In_3721,In_2975);
or U746 (N_746,In_4372,In_4989);
nor U747 (N_747,In_187,In_4431);
nand U748 (N_748,In_1053,In_3194);
nor U749 (N_749,In_201,In_720);
and U750 (N_750,In_2495,In_4457);
nor U751 (N_751,In_2564,In_3646);
nand U752 (N_752,In_636,In_1461);
and U753 (N_753,In_4978,In_2817);
or U754 (N_754,In_4015,In_4662);
or U755 (N_755,In_1997,In_4359);
nand U756 (N_756,In_3571,In_3249);
and U757 (N_757,In_2075,In_1782);
and U758 (N_758,In_2467,In_614);
or U759 (N_759,In_128,In_1931);
or U760 (N_760,In_1106,In_2776);
nor U761 (N_761,In_3087,In_3346);
nor U762 (N_762,In_434,In_4505);
nand U763 (N_763,In_4008,In_357);
nor U764 (N_764,In_4704,In_1574);
and U765 (N_765,In_546,In_186);
and U766 (N_766,In_4586,In_2634);
nor U767 (N_767,In_1596,In_910);
nor U768 (N_768,In_3781,In_237);
and U769 (N_769,In_4678,In_3486);
xnor U770 (N_770,In_3223,In_4936);
and U771 (N_771,In_4963,In_1284);
xnor U772 (N_772,In_3148,In_2275);
or U773 (N_773,In_3343,In_578);
and U774 (N_774,In_1552,In_1854);
and U775 (N_775,In_3543,In_46);
and U776 (N_776,In_3472,In_4543);
nor U777 (N_777,In_443,In_4827);
nor U778 (N_778,In_3861,In_2082);
or U779 (N_779,In_2670,In_374);
or U780 (N_780,In_4293,In_1744);
nand U781 (N_781,In_2804,In_2007);
and U782 (N_782,In_1163,In_2330);
and U783 (N_783,In_3833,In_3547);
or U784 (N_784,In_2588,In_1562);
and U785 (N_785,In_1478,In_2339);
or U786 (N_786,In_3308,In_4005);
xor U787 (N_787,In_906,In_29);
and U788 (N_788,In_2240,In_4377);
or U789 (N_789,In_227,In_3751);
nand U790 (N_790,In_3960,In_703);
and U791 (N_791,In_2061,In_3948);
nand U792 (N_792,In_3410,In_3971);
and U793 (N_793,In_4337,In_1862);
or U794 (N_794,In_4299,In_691);
or U795 (N_795,In_2359,In_3775);
nor U796 (N_796,In_2029,In_588);
nand U797 (N_797,In_4545,In_4714);
and U798 (N_798,In_3596,In_4643);
or U799 (N_799,In_3765,In_2524);
nor U800 (N_800,In_4019,In_4222);
and U801 (N_801,In_1604,In_617);
or U802 (N_802,In_812,In_1960);
and U803 (N_803,In_2625,In_4947);
nand U804 (N_804,In_537,In_3826);
or U805 (N_805,In_4782,In_4043);
or U806 (N_806,In_3197,In_2181);
or U807 (N_807,In_4804,In_635);
nand U808 (N_808,In_3088,In_4116);
and U809 (N_809,In_1396,In_2414);
and U810 (N_810,In_1037,In_1787);
nand U811 (N_811,In_3798,In_757);
and U812 (N_812,In_1400,In_1266);
nor U813 (N_813,In_2350,In_2873);
and U814 (N_814,In_2143,In_3822);
or U815 (N_815,In_2749,In_1575);
and U816 (N_816,In_4617,In_3240);
nand U817 (N_817,In_2145,In_3770);
nand U818 (N_818,In_4832,In_2695);
or U819 (N_819,In_2440,In_4759);
and U820 (N_820,In_3137,In_3710);
and U821 (N_821,In_2052,In_956);
or U822 (N_822,In_4486,In_1890);
nor U823 (N_823,In_2692,In_1120);
and U824 (N_824,In_126,In_1211);
and U825 (N_825,In_438,In_1240);
nor U826 (N_826,In_189,In_606);
nand U827 (N_827,In_4213,In_2867);
nor U828 (N_828,In_4649,In_4851);
nor U829 (N_829,In_4121,In_2439);
nand U830 (N_830,In_387,In_249);
or U831 (N_831,In_335,In_1241);
nand U832 (N_832,In_3891,In_2622);
and U833 (N_833,In_3889,In_2234);
nor U834 (N_834,In_3090,In_4725);
and U835 (N_835,In_2548,In_2078);
nand U836 (N_836,In_1435,In_915);
or U837 (N_837,In_2158,In_4748);
or U838 (N_838,In_4423,In_2752);
or U839 (N_839,In_164,In_2321);
or U840 (N_840,In_1116,In_4847);
and U841 (N_841,In_3871,In_2374);
xnor U842 (N_842,In_3946,In_3640);
nor U843 (N_843,In_1958,In_4292);
and U844 (N_844,In_3810,In_1984);
nor U845 (N_845,In_1115,In_2645);
nor U846 (N_846,In_3838,In_1430);
and U847 (N_847,In_2151,In_183);
nand U848 (N_848,In_2551,In_1647);
or U849 (N_849,In_2849,In_3436);
nor U850 (N_850,In_2415,In_3119);
nor U851 (N_851,In_1748,In_2438);
or U852 (N_852,In_4566,In_2760);
and U853 (N_853,In_701,In_2419);
nand U854 (N_854,In_1717,In_1384);
nand U855 (N_855,In_1546,In_4488);
or U856 (N_856,In_430,In_1055);
nor U857 (N_857,In_4758,In_1230);
or U858 (N_858,In_1777,In_2056);
and U859 (N_859,In_3981,In_1950);
nor U860 (N_860,In_822,In_3222);
or U861 (N_861,In_4470,In_862);
nand U862 (N_862,In_1856,In_1959);
or U863 (N_863,In_1450,In_3774);
or U864 (N_864,In_2546,In_4973);
nand U865 (N_865,In_3511,In_3923);
or U866 (N_866,In_4852,In_3422);
and U867 (N_867,In_255,In_3073);
nor U868 (N_868,In_1899,In_4906);
or U869 (N_869,In_2171,In_1721);
nor U870 (N_870,In_2627,In_94);
or U871 (N_871,In_3146,In_1445);
nand U872 (N_872,In_2216,In_152);
or U873 (N_873,In_3061,In_87);
nand U874 (N_874,In_1965,In_2886);
nor U875 (N_875,In_1653,In_2732);
nor U876 (N_876,In_4993,In_968);
nand U877 (N_877,In_2600,In_3583);
xor U878 (N_878,In_4375,In_2621);
nand U879 (N_879,In_4972,In_1003);
nor U880 (N_880,In_2783,In_4367);
nand U881 (N_881,In_3250,In_1876);
and U882 (N_882,In_3551,In_2683);
and U883 (N_883,In_4345,In_368);
nor U884 (N_884,In_2093,In_3945);
nor U885 (N_885,In_3149,In_4483);
nor U886 (N_886,In_695,In_2631);
nand U887 (N_887,In_1087,In_452);
and U888 (N_888,In_1800,In_1203);
nor U889 (N_889,In_4277,In_2755);
or U890 (N_890,In_1719,In_1351);
or U891 (N_891,In_4873,In_3449);
xnor U892 (N_892,In_4270,In_2183);
or U893 (N_893,In_2570,In_4003);
nand U894 (N_894,In_2335,In_545);
or U895 (N_895,In_4591,In_1308);
nor U896 (N_896,In_2130,In_3627);
nor U897 (N_897,In_1205,In_725);
nor U898 (N_898,In_4208,In_1763);
or U899 (N_899,In_188,In_1299);
nand U900 (N_900,In_514,In_3493);
and U901 (N_901,In_1397,In_2782);
or U902 (N_902,In_3424,In_192);
xnor U903 (N_903,In_4138,In_4230);
and U904 (N_904,In_4499,In_4254);
or U905 (N_905,In_3812,In_1052);
nand U906 (N_906,In_1204,In_3746);
and U907 (N_907,In_3239,In_4446);
or U908 (N_908,In_2823,In_1471);
or U909 (N_909,In_2712,In_3598);
nand U910 (N_910,In_3817,In_566);
nor U911 (N_911,In_1532,In_524);
nand U912 (N_912,In_3479,In_4065);
or U913 (N_913,In_132,In_1654);
nand U914 (N_914,In_1476,In_1237);
nand U915 (N_915,In_267,In_240);
and U916 (N_916,In_3164,In_3366);
and U917 (N_917,In_3210,In_2373);
nand U918 (N_918,In_3679,In_686);
and U919 (N_919,In_3127,In_3655);
nor U920 (N_920,In_4221,In_3535);
nand U921 (N_921,In_876,In_2935);
xnor U922 (N_922,In_4894,In_1977);
nand U923 (N_923,In_1370,In_470);
or U924 (N_924,In_1889,In_100);
nor U925 (N_925,In_659,In_4984);
nand U926 (N_926,In_510,In_3743);
and U927 (N_927,In_4808,In_2527);
or U928 (N_928,In_130,In_1034);
xnor U929 (N_929,In_1577,In_2672);
nand U930 (N_930,In_4705,In_367);
or U931 (N_931,In_2746,In_4383);
nor U932 (N_932,In_4068,In_829);
nor U933 (N_933,In_1772,In_3578);
and U934 (N_934,In_3633,In_2300);
or U935 (N_935,In_999,In_3089);
nor U936 (N_936,In_3455,In_1331);
nand U937 (N_937,In_933,In_2126);
or U938 (N_938,In_3028,In_4638);
and U939 (N_939,In_4673,In_3676);
or U940 (N_940,In_3821,In_2202);
nor U941 (N_941,In_3134,In_111);
nand U942 (N_942,In_3921,In_2222);
and U943 (N_943,In_3058,In_520);
or U944 (N_944,In_1033,In_1624);
nor U945 (N_945,In_1860,In_4051);
and U946 (N_946,In_3474,In_2154);
nand U947 (N_947,In_2094,In_2566);
nand U948 (N_948,In_2242,In_3316);
and U949 (N_949,In_4528,In_2340);
and U950 (N_950,In_4957,In_2355);
or U951 (N_951,In_2120,In_3155);
nand U952 (N_952,In_2899,In_3217);
and U953 (N_953,In_1330,In_4263);
or U954 (N_954,In_1010,In_3138);
and U955 (N_955,In_4000,In_294);
and U956 (N_956,In_3371,In_1132);
and U957 (N_957,In_2828,In_1804);
nor U958 (N_958,In_3802,In_4311);
and U959 (N_959,In_2443,In_4282);
nor U960 (N_960,In_310,In_4105);
and U961 (N_961,In_1226,In_1943);
and U962 (N_962,In_2596,In_4562);
or U963 (N_963,In_4288,In_211);
or U964 (N_964,In_2080,In_3242);
nor U965 (N_965,In_3357,In_3470);
nor U966 (N_966,In_2229,In_1664);
nor U967 (N_967,In_4820,In_638);
nand U968 (N_968,In_3944,In_1343);
and U969 (N_969,In_1650,In_1753);
and U970 (N_970,In_150,In_4200);
nor U971 (N_971,In_1246,In_2717);
xor U972 (N_972,In_2678,In_27);
nor U973 (N_973,In_2038,In_2544);
and U974 (N_974,In_2905,In_401);
nand U975 (N_975,In_4369,In_1727);
nand U976 (N_976,In_866,In_3456);
nor U977 (N_977,In_4926,In_3772);
nand U978 (N_978,In_1356,In_681);
and U979 (N_979,In_1941,In_16);
nor U980 (N_980,In_3096,In_4223);
nand U981 (N_981,In_746,In_2308);
and U982 (N_982,In_1641,In_2518);
or U983 (N_983,In_4970,In_4717);
and U984 (N_984,In_1072,In_2998);
nand U985 (N_985,In_3206,In_1579);
nor U986 (N_986,In_3663,In_3048);
nor U987 (N_987,In_3274,In_421);
and U988 (N_988,In_2382,In_2048);
or U989 (N_989,In_1961,In_84);
and U990 (N_990,In_3636,In_4094);
nor U991 (N_991,In_2390,In_4583);
or U992 (N_992,In_2475,In_4686);
or U993 (N_993,In_1252,In_2567);
nor U994 (N_994,In_3650,In_449);
or U995 (N_995,In_905,In_3232);
nand U996 (N_996,In_3965,In_776);
nand U997 (N_997,In_2554,In_3401);
nand U998 (N_998,In_4500,In_1733);
nand U999 (N_999,In_3998,In_4131);
or U1000 (N_1000,In_1046,In_1127);
or U1001 (N_1001,In_3178,In_4133);
and U1002 (N_1002,In_2221,In_3926);
or U1003 (N_1003,In_1349,In_787);
or U1004 (N_1004,In_49,In_3642);
nor U1005 (N_1005,In_4069,In_1453);
and U1006 (N_1006,In_2144,In_1838);
or U1007 (N_1007,In_1585,In_299);
nand U1008 (N_1008,In_4753,In_1771);
or U1009 (N_1009,In_2492,In_2895);
nor U1010 (N_1010,In_4576,In_4495);
or U1011 (N_1011,In_3142,In_1690);
or U1012 (N_1012,In_4142,In_3514);
nor U1013 (N_1013,In_2113,In_3315);
nor U1014 (N_1014,In_2004,In_2690);
nand U1015 (N_1015,In_1043,In_4460);
or U1016 (N_1016,In_72,In_1619);
nand U1017 (N_1017,In_3170,In_1794);
or U1018 (N_1018,In_2821,In_4290);
and U1019 (N_1019,In_2647,In_4732);
nand U1020 (N_1020,In_1274,In_2955);
or U1021 (N_1021,In_4489,In_4169);
nor U1022 (N_1022,In_1180,In_4408);
or U1023 (N_1023,In_2191,In_2820);
and U1024 (N_1024,In_2664,In_3909);
and U1025 (N_1025,In_1880,In_2291);
and U1026 (N_1026,In_562,In_4889);
and U1027 (N_1027,In_3326,In_2515);
or U1028 (N_1028,In_867,In_3958);
nand U1029 (N_1029,In_3333,In_1875);
nor U1030 (N_1030,In_1601,In_2462);
and U1031 (N_1031,In_161,In_308);
and U1032 (N_1032,In_40,In_2301);
and U1033 (N_1033,In_2706,In_3742);
or U1034 (N_1034,In_1897,In_2105);
and U1035 (N_1035,In_4157,In_3718);
nand U1036 (N_1036,In_4831,In_372);
or U1037 (N_1037,In_621,In_1667);
nor U1038 (N_1038,In_3295,In_2025);
and U1039 (N_1039,In_988,In_3322);
or U1040 (N_1040,In_4376,In_2613);
and U1041 (N_1041,In_515,In_4779);
or U1042 (N_1042,In_1946,In_1615);
or U1043 (N_1043,In_3183,In_2604);
or U1044 (N_1044,In_4866,In_102);
nor U1045 (N_1045,In_1390,In_4178);
and U1046 (N_1046,In_1864,In_1426);
nand U1047 (N_1047,In_864,In_732);
nand U1048 (N_1048,In_4692,In_4818);
or U1049 (N_1049,In_2597,In_541);
nor U1050 (N_1050,In_23,In_3609);
and U1051 (N_1051,In_4580,In_4152);
or U1052 (N_1052,In_1272,In_3489);
nand U1053 (N_1053,In_4730,In_2437);
nor U1054 (N_1054,In_4542,In_1346);
nand U1055 (N_1055,In_563,In_1918);
nand U1056 (N_1056,In_4454,In_4109);
nand U1057 (N_1057,In_2453,In_2401);
or U1058 (N_1058,In_4707,In_3367);
and U1059 (N_1059,In_4077,In_4555);
nand U1060 (N_1060,In_2874,In_2134);
and U1061 (N_1061,In_3777,In_4731);
or U1062 (N_1062,In_3745,In_4982);
nand U1063 (N_1063,In_4939,In_3672);
or U1064 (N_1064,In_3059,In_1089);
nand U1065 (N_1065,In_2581,In_599);
nand U1066 (N_1066,In_4274,In_1590);
or U1067 (N_1067,In_3585,In_1480);
nand U1068 (N_1068,In_3176,In_4942);
nand U1069 (N_1069,In_2590,In_1256);
nand U1070 (N_1070,In_1281,In_3428);
and U1071 (N_1071,In_1298,In_3);
nand U1072 (N_1072,In_4979,In_3220);
nand U1073 (N_1073,In_3595,In_1093);
nand U1074 (N_1074,In_2173,In_33);
nand U1075 (N_1075,In_2653,In_2819);
nand U1076 (N_1076,In_1150,In_2076);
nand U1077 (N_1077,In_1635,In_1181);
or U1078 (N_1078,In_2426,In_1592);
nor U1079 (N_1079,In_1852,In_3009);
or U1080 (N_1080,In_4801,In_4368);
nor U1081 (N_1081,In_3523,In_2476);
nand U1082 (N_1082,In_2994,In_4887);
nor U1083 (N_1083,In_1101,In_4059);
and U1084 (N_1084,In_4722,In_4242);
nand U1085 (N_1085,In_4197,In_3391);
and U1086 (N_1086,In_3244,In_174);
or U1087 (N_1087,In_1209,In_3116);
nor U1088 (N_1088,In_3186,In_17);
nor U1089 (N_1089,In_1212,In_3227);
nand U1090 (N_1090,In_3280,In_693);
nand U1091 (N_1091,In_2399,In_4106);
nor U1092 (N_1092,In_3091,In_245);
nand U1093 (N_1093,In_3135,In_3039);
and U1094 (N_1094,In_2599,In_1798);
and U1095 (N_1095,In_4233,In_4268);
nand U1096 (N_1096,In_3208,In_4258);
xnor U1097 (N_1097,In_3328,In_816);
nor U1098 (N_1098,In_1866,In_2535);
or U1099 (N_1099,In_3972,In_2459);
nor U1100 (N_1100,In_957,In_1636);
nor U1101 (N_1101,In_4329,In_3512);
and U1102 (N_1102,In_890,In_272);
and U1103 (N_1103,In_2941,In_4994);
nor U1104 (N_1104,In_1706,In_3692);
nand U1105 (N_1105,In_3214,In_4344);
and U1106 (N_1106,In_487,In_4473);
nand U1107 (N_1107,In_758,In_3062);
nand U1108 (N_1108,In_1449,In_928);
or U1109 (N_1109,In_4752,In_3950);
and U1110 (N_1110,In_167,In_2987);
and U1111 (N_1111,In_667,In_3053);
nor U1112 (N_1112,In_2088,In_56);
nand U1113 (N_1113,In_3184,In_4602);
nand U1114 (N_1114,In_3936,In_4665);
nand U1115 (N_1115,In_50,In_2116);
and U1116 (N_1116,In_3790,In_663);
and U1117 (N_1117,In_1591,In_2790);
nand U1118 (N_1118,In_4214,In_405);
or U1119 (N_1119,In_282,In_266);
or U1120 (N_1120,In_3591,In_4761);
nor U1121 (N_1121,In_4577,In_3056);
nand U1122 (N_1122,In_2220,In_4544);
or U1123 (N_1123,In_297,In_3506);
and U1124 (N_1124,In_2569,In_3534);
nand U1125 (N_1125,In_4874,In_1974);
and U1126 (N_1126,In_101,In_36);
and U1127 (N_1127,In_4287,In_3166);
nand U1128 (N_1128,In_3355,In_4480);
nor U1129 (N_1129,In_1947,In_1795);
or U1130 (N_1130,In_4385,In_794);
or U1131 (N_1131,In_2309,In_4397);
nand U1132 (N_1132,In_844,In_4286);
nand U1133 (N_1133,In_729,In_2198);
and U1134 (N_1134,In_3398,In_2556);
nand U1135 (N_1135,In_4265,In_3979);
nand U1136 (N_1136,In_3959,In_2465);
nor U1137 (N_1137,In_4552,In_2694);
nor U1138 (N_1138,In_1201,In_3494);
nor U1139 (N_1139,In_1696,In_493);
nand U1140 (N_1140,In_1059,In_4304);
nor U1141 (N_1141,In_1519,In_2503);
or U1142 (N_1142,In_1260,In_4295);
nor U1143 (N_1143,In_158,In_1722);
nor U1144 (N_1144,In_2813,In_3434);
nor U1145 (N_1145,In_1877,In_1225);
or U1146 (N_1146,In_959,In_1554);
nand U1147 (N_1147,In_4127,In_807);
nand U1148 (N_1148,In_228,In_1467);
nand U1149 (N_1149,In_2912,In_2361);
nor U1150 (N_1150,In_3177,In_712);
and U1151 (N_1151,In_4527,In_1754);
nor U1152 (N_1152,In_3933,In_3465);
or U1153 (N_1153,In_2860,In_4228);
and U1154 (N_1154,In_1741,In_3107);
or U1155 (N_1155,In_4582,In_1207);
nor U1156 (N_1156,In_1969,In_1380);
and U1157 (N_1157,In_2128,In_1468);
and U1158 (N_1158,In_856,In_3338);
nor U1159 (N_1159,In_1154,In_3193);
nand U1160 (N_1160,In_3495,In_3752);
nor U1161 (N_1161,In_3731,In_3990);
or U1162 (N_1162,In_775,In_3108);
or U1163 (N_1163,In_1799,In_3207);
nor U1164 (N_1164,In_1219,In_1684);
nor U1165 (N_1165,In_347,In_886);
or U1166 (N_1166,In_4456,In_4794);
or U1167 (N_1167,In_500,In_4633);
or U1168 (N_1168,In_1766,In_307);
nand U1169 (N_1169,In_3957,In_4088);
nand U1170 (N_1170,In_441,In_3832);
nand U1171 (N_1171,In_4357,In_2434);
nor U1172 (N_1172,In_1340,In_2010);
nor U1173 (N_1173,In_2490,In_488);
nand U1174 (N_1174,In_1459,In_847);
nand U1175 (N_1175,In_1255,In_107);
or U1176 (N_1176,In_478,In_3187);
nand U1177 (N_1177,In_3457,In_3794);
and U1178 (N_1178,In_3503,In_4857);
nand U1179 (N_1179,In_4291,In_4113);
nand U1180 (N_1180,In_1144,In_2903);
and U1181 (N_1181,In_4918,In_2800);
or U1182 (N_1182,In_2095,In_590);
or U1183 (N_1183,In_1916,In_3896);
nand U1184 (N_1184,In_3786,In_223);
or U1185 (N_1185,In_1223,In_699);
or U1186 (N_1186,In_3051,In_2915);
nor U1187 (N_1187,In_2296,In_1506);
nand U1188 (N_1188,In_1949,In_1681);
nor U1189 (N_1189,In_1535,In_1900);
and U1190 (N_1190,In_4215,In_4985);
nand U1191 (N_1191,In_3375,In_2868);
nand U1192 (N_1192,In_3964,In_349);
and U1193 (N_1193,In_2406,In_3549);
nand U1194 (N_1194,In_4283,In_424);
nand U1195 (N_1195,In_2357,In_3522);
and U1196 (N_1196,In_2265,In_4124);
and U1197 (N_1197,In_1276,In_4356);
xnor U1198 (N_1198,In_1289,In_3859);
nor U1199 (N_1199,In_962,In_3620);
or U1200 (N_1200,In_3327,In_1685);
nor U1201 (N_1201,In_3807,In_1457);
nand U1202 (N_1202,In_4091,In_322);
xnor U1203 (N_1203,In_3912,In_1788);
nor U1204 (N_1204,In_364,In_4822);
nand U1205 (N_1205,In_1141,In_4151);
nor U1206 (N_1206,In_4465,In_2950);
nor U1207 (N_1207,In_3669,In_143);
or U1208 (N_1208,In_3219,In_463);
and U1209 (N_1209,In_3481,In_92);
or U1210 (N_1210,In_627,In_67);
or U1211 (N_1211,In_2794,In_1121);
and U1212 (N_1212,In_3324,In_894);
nor U1213 (N_1213,In_1472,In_1836);
nand U1214 (N_1214,In_4310,In_1409);
or U1215 (N_1215,In_3667,In_2096);
nand U1216 (N_1216,In_1216,In_4792);
nand U1217 (N_1217,In_3565,In_4467);
nor U1218 (N_1218,In_1767,In_1938);
nor U1219 (N_1219,In_4185,In_984);
nor U1220 (N_1220,In_4671,In_2101);
or U1221 (N_1221,In_2341,In_30);
or U1222 (N_1222,In_1175,In_3716);
nand U1223 (N_1223,In_208,In_1621);
or U1224 (N_1224,In_2651,In_353);
or U1225 (N_1225,In_3898,In_2423);
or U1226 (N_1226,In_580,In_4806);
or U1227 (N_1227,In_4079,In_2316);
and U1228 (N_1228,In_410,In_1080);
or U1229 (N_1229,In_4578,In_4932);
nand U1230 (N_1230,In_3656,In_4064);
and U1231 (N_1231,In_2182,In_805);
and U1232 (N_1232,In_2342,In_2960);
or U1233 (N_1233,In_4219,In_3272);
or U1234 (N_1234,In_1935,In_572);
or U1235 (N_1235,In_1530,In_3411);
nand U1236 (N_1236,In_3301,In_1540);
nor U1237 (N_1237,In_2295,In_4490);
nor U1238 (N_1238,In_1658,In_832);
and U1239 (N_1239,In_3610,In_243);
or U1240 (N_1240,In_1100,In_3368);
or U1241 (N_1241,In_656,In_1670);
or U1242 (N_1242,In_472,In_3431);
nand U1243 (N_1243,In_1991,In_362);
and U1244 (N_1244,In_2926,In_1817);
and U1245 (N_1245,In_2589,In_475);
or U1246 (N_1246,In_1022,In_586);
nand U1247 (N_1247,In_3887,In_2055);
nand U1248 (N_1248,In_4011,In_4655);
nor U1249 (N_1249,In_2446,In_2543);
nor U1250 (N_1250,In_1444,In_4334);
nor U1251 (N_1251,In_509,In_4508);
nor U1252 (N_1252,In_4203,In_2239);
and U1253 (N_1253,In_2232,In_652);
nand U1254 (N_1254,In_1551,In_613);
nor U1255 (N_1255,In_2913,In_1178);
or U1256 (N_1256,In_3702,In_4754);
nand U1257 (N_1257,In_2394,In_1919);
nor U1258 (N_1258,In_3269,In_2480);
nand U1259 (N_1259,In_1526,In_793);
and U1260 (N_1260,In_2132,In_292);
and U1261 (N_1261,In_185,In_4262);
or U1262 (N_1262,In_687,In_458);
and U1263 (N_1263,In_4036,In_2352);
and U1264 (N_1264,In_1073,In_4158);
or U1265 (N_1265,In_879,In_2209);
nor U1266 (N_1266,In_4030,In_62);
and U1267 (N_1267,In_902,In_361);
nor U1268 (N_1268,In_3069,In_1736);
or U1269 (N_1269,In_1527,In_3369);
or U1270 (N_1270,In_3630,In_3829);
nand U1271 (N_1271,In_4176,In_1979);
nand U1272 (N_1272,In_360,In_3055);
nand U1273 (N_1273,In_2696,In_4318);
or U1274 (N_1274,In_1594,In_3851);
nor U1275 (N_1275,In_2160,In_2824);
nor U1276 (N_1276,In_1040,In_428);
nor U1277 (N_1277,In_3927,In_1920);
and U1278 (N_1278,In_4269,In_2745);
and U1279 (N_1279,In_4700,In_3260);
or U1280 (N_1280,In_4796,In_1813);
and U1281 (N_1281,In_4679,In_3619);
nand U1282 (N_1282,In_3204,In_125);
or U1283 (N_1283,In_4045,In_3873);
or U1284 (N_1284,In_4862,In_745);
nand U1285 (N_1285,In_658,In_2497);
or U1286 (N_1286,In_4314,In_138);
nand U1287 (N_1287,In_273,In_738);
nor U1288 (N_1288,In_4366,In_3130);
and U1289 (N_1289,In_4861,In_1587);
xnor U1290 (N_1290,In_1761,In_38);
nor U1291 (N_1291,In_1614,In_1316);
nand U1292 (N_1292,In_4501,In_4575);
nor U1293 (N_1293,In_3468,In_4589);
or U1294 (N_1294,In_163,In_2235);
or U1295 (N_1295,In_3010,In_673);
and U1296 (N_1296,In_20,In_1485);
or U1297 (N_1297,In_1711,In_2003);
nor U1298 (N_1298,In_4236,In_743);
nor U1299 (N_1299,In_3546,In_3888);
and U1300 (N_1300,In_2681,In_960);
or U1301 (N_1301,In_852,In_979);
and U1302 (N_1302,In_3349,In_4235);
and U1303 (N_1303,In_1928,In_3830);
nand U1304 (N_1304,In_552,In_176);
or U1305 (N_1305,In_4205,In_2902);
or U1306 (N_1306,In_3705,In_2290);
nor U1307 (N_1307,In_4107,In_2091);
or U1308 (N_1308,In_2968,In_919);
and U1309 (N_1309,In_3118,In_1978);
nand U1310 (N_1310,In_3975,In_4201);
and U1311 (N_1311,In_2641,In_4944);
and U1312 (N_1312,In_814,In_1291);
or U1313 (N_1313,In_4652,In_2485);
nand U1314 (N_1314,In_529,In_1321);
and U1315 (N_1315,In_1161,In_3293);
and U1316 (N_1316,In_76,In_2190);
nor U1317 (N_1317,In_3425,In_1064);
nor U1318 (N_1318,In_1893,In_53);
or U1319 (N_1319,In_4216,In_683);
and U1320 (N_1320,In_124,In_550);
or U1321 (N_1321,In_1404,In_4057);
and U1322 (N_1322,In_2748,In_2169);
nand U1323 (N_1323,In_4017,In_4856);
and U1324 (N_1324,In_1660,In_3129);
nor U1325 (N_1325,In_3221,In_1511);
nor U1326 (N_1326,In_4749,In_2054);
or U1327 (N_1327,In_4996,In_3196);
and U1328 (N_1328,In_2644,In_4684);
and U1329 (N_1329,In_4967,In_655);
nor U1330 (N_1330,In_3902,In_3932);
or U1331 (N_1331,In_133,In_3484);
nor U1332 (N_1332,In_4087,In_922);
nor U1333 (N_1333,In_340,In_1904);
nand U1334 (N_1334,In_801,In_3846);
and U1335 (N_1335,In_996,In_2526);
nand U1336 (N_1336,In_3216,In_271);
nor U1337 (N_1337,In_4278,In_1677);
and U1338 (N_1338,In_2666,In_1915);
or U1339 (N_1339,In_540,In_680);
nand U1340 (N_1340,In_2336,In_2083);
or U1341 (N_1341,In_3491,In_2504);
or U1342 (N_1342,In_4187,In_4795);
and U1343 (N_1343,In_1738,In_1702);
nand U1344 (N_1344,In_1796,In_719);
nand U1345 (N_1345,In_1417,In_4443);
nor U1346 (N_1346,In_4204,In_4855);
nor U1347 (N_1347,In_1841,In_2559);
xnor U1348 (N_1348,In_1510,In_1217);
nor U1349 (N_1349,In_4651,In_2022);
nand U1350 (N_1350,In_1151,In_2614);
or U1351 (N_1351,In_4032,In_4037);
nor U1352 (N_1352,In_2593,In_44);
or U1353 (N_1353,In_1881,In_1157);
or U1354 (N_1354,In_2046,In_2197);
nand U1355 (N_1355,In_3588,In_942);
and U1356 (N_1356,In_2314,In_3985);
nor U1357 (N_1357,In_369,In_3849);
or U1358 (N_1358,In_3433,In_4746);
nor U1359 (N_1359,In_3886,In_1820);
and U1360 (N_1360,In_3426,In_3813);
and U1361 (N_1361,In_4890,In_4767);
and U1362 (N_1362,In_1769,In_4250);
nor U1363 (N_1363,In_3769,In_3453);
nand U1364 (N_1364,In_791,In_4609);
or U1365 (N_1365,In_3621,In_4534);
and U1366 (N_1366,In_3162,In_4472);
nand U1367 (N_1367,In_2488,In_3558);
and U1368 (N_1368,In_1262,In_193);
nor U1369 (N_1369,In_2468,In_3312);
xor U1370 (N_1370,In_4666,In_2192);
and U1371 (N_1371,In_2073,In_4677);
nor U1372 (N_1372,In_1287,In_726);
nor U1373 (N_1373,In_4049,In_4999);
or U1374 (N_1374,In_4309,In_4537);
nand U1375 (N_1375,In_419,In_4608);
and U1376 (N_1376,In_1972,In_3693);
and U1377 (N_1377,In_4160,In_404);
and U1378 (N_1378,In_2458,In_2857);
or U1379 (N_1379,In_3978,In_724);
or U1380 (N_1380,In_1903,In_2561);
and U1381 (N_1381,In_3920,In_2178);
or U1382 (N_1382,In_2934,In_1269);
and U1383 (N_1383,In_1545,In_4538);
nor U1384 (N_1384,In_3256,In_1781);
nor U1385 (N_1385,In_4878,In_2936);
and U1386 (N_1386,In_3389,In_1383);
or U1387 (N_1387,In_1633,In_4172);
nand U1388 (N_1388,In_2322,In_4791);
xnor U1389 (N_1389,In_78,In_3525);
and U1390 (N_1390,In_519,In_2738);
and U1391 (N_1391,In_448,In_4836);
nor U1392 (N_1392,In_3290,In_485);
and U1393 (N_1393,In_3704,In_3994);
and U1394 (N_1394,In_3031,In_156);
xnor U1395 (N_1395,In_2626,In_2293);
nor U1396 (N_1396,In_3529,In_4150);
nor U1397 (N_1397,In_2991,In_4698);
or U1398 (N_1398,In_4948,In_3892);
nand U1399 (N_1399,In_3283,In_136);
and U1400 (N_1400,In_2933,In_2635);
and U1401 (N_1401,In_0,In_2270);
nor U1402 (N_1402,In_3681,In_172);
nand U1403 (N_1403,In_503,In_1521);
nand U1404 (N_1404,In_4777,In_1611);
and U1405 (N_1405,In_135,In_4571);
and U1406 (N_1406,In_3444,In_64);
xnor U1407 (N_1407,In_4601,In_3510);
nand U1408 (N_1408,In_3737,In_2675);
or U1409 (N_1409,In_2818,In_2890);
nor U1410 (N_1410,In_1325,In_80);
nor U1411 (N_1411,In_4798,In_4052);
and U1412 (N_1412,In_1310,In_2528);
or U1413 (N_1413,In_2550,In_4317);
nand U1414 (N_1414,In_1147,In_247);
nor U1415 (N_1415,In_1536,In_2122);
and U1416 (N_1416,In_1366,In_2525);
nand U1417 (N_1417,In_2542,In_3205);
xor U1418 (N_1418,In_2481,In_1668);
xnor U1419 (N_1419,In_3273,In_2996);
and U1420 (N_1420,In_2201,In_1375);
and U1421 (N_1421,In_3550,In_976);
or U1422 (N_1422,In_642,In_4819);
or U1423 (N_1423,In_3914,In_3180);
nor U1424 (N_1424,In_314,In_269);
and U1425 (N_1425,In_1940,In_3430);
nand U1426 (N_1426,In_4303,In_2552);
and U1427 (N_1427,In_789,In_2877);
and U1428 (N_1428,In_2871,In_407);
nand U1429 (N_1429,In_1844,In_3188);
and U1430 (N_1430,In_3384,In_3538);
nand U1431 (N_1431,In_1253,In_4719);
and U1432 (N_1432,In_747,In_3664);
and U1433 (N_1433,In_2775,In_4261);
nand U1434 (N_1434,In_3904,In_1495);
and U1435 (N_1435,In_511,In_4607);
nor U1436 (N_1436,In_4417,In_4159);
nand U1437 (N_1437,In_2773,In_3934);
and U1438 (N_1438,In_21,In_4024);
xnor U1439 (N_1439,In_2435,In_4958);
and U1440 (N_1440,In_551,In_633);
nand U1441 (N_1441,In_1830,In_1802);
or U1442 (N_1442,In_446,In_2565);
or U1443 (N_1443,In_1195,In_4653);
and U1444 (N_1444,In_1952,In_3192);
nor U1445 (N_1445,In_761,In_662);
and U1446 (N_1446,In_220,In_1716);
nor U1447 (N_1447,In_2412,In_1159);
and U1448 (N_1448,In_1296,In_3158);
nor U1449 (N_1449,In_2206,In_4421);
or U1450 (N_1450,In_884,In_3446);
or U1451 (N_1451,In_4898,In_3662);
nand U1452 (N_1452,In_2231,In_426);
and U1453 (N_1453,In_2532,In_3014);
or U1454 (N_1454,In_2663,In_1441);
nand U1455 (N_1455,In_303,In_467);
and U1456 (N_1456,In_4149,In_453);
and U1457 (N_1457,In_907,In_2946);
nor U1458 (N_1458,In_293,In_4828);
and U1459 (N_1459,In_1199,In_1140);
nor U1460 (N_1460,In_992,In_2332);
and U1461 (N_1461,In_739,In_1335);
nand U1462 (N_1462,In_3711,In_1855);
or U1463 (N_1463,In_4909,In_734);
and U1464 (N_1464,In_3291,In_3984);
nand U1465 (N_1465,In_2187,In_2901);
and U1466 (N_1466,In_396,In_2992);
nand U1467 (N_1467,In_3459,In_3122);
or U1468 (N_1468,In_4697,In_1516);
nand U1469 (N_1469,In_2463,In_302);
and U1470 (N_1470,In_1090,In_4895);
nand U1471 (N_1471,In_1293,In_1778);
and U1472 (N_1472,In_4773,In_1725);
or U1473 (N_1473,In_4628,In_4881);
or U1474 (N_1474,In_3918,In_3785);
nand U1475 (N_1475,In_2702,In_3868);
or U1476 (N_1476,In_1045,In_1290);
or U1477 (N_1477,In_505,In_1286);
and U1478 (N_1478,In_2797,In_2942);
nor U1479 (N_1479,In_3714,In_898);
or U1480 (N_1480,In_3463,In_2560);
and U1481 (N_1481,In_531,In_2606);
or U1482 (N_1482,In_2251,In_1094);
nand U1483 (N_1483,In_4414,In_2806);
and U1484 (N_1484,In_22,In_3517);
or U1485 (N_1485,In_2510,In_257);
nor U1486 (N_1486,In_2520,In_4720);
nand U1487 (N_1487,In_4145,In_764);
nor U1488 (N_1488,In_3857,In_3213);
and U1489 (N_1489,In_4249,In_1196);
and U1490 (N_1490,In_2451,In_484);
or U1491 (N_1491,In_1218,In_3189);
or U1492 (N_1492,In_1191,In_2939);
or U1493 (N_1493,In_1388,In_43);
nand U1494 (N_1494,In_4381,In_4865);
nor U1495 (N_1495,In_499,In_1663);
nand U1496 (N_1496,In_4629,In_982);
or U1497 (N_1497,In_4143,In_1184);
or U1498 (N_1498,In_3811,In_119);
nor U1499 (N_1499,In_1867,In_4191);
nor U1500 (N_1500,In_1415,In_689);
and U1501 (N_1501,In_722,In_4533);
and U1502 (N_1502,In_3165,In_2661);
nor U1503 (N_1503,In_3416,In_1434);
xor U1504 (N_1504,In_4902,In_4025);
nor U1505 (N_1505,In_251,In_411);
and U1506 (N_1506,In_3251,In_373);
nor U1507 (N_1507,In_139,In_3302);
or U1508 (N_1508,In_2716,In_1712);
xor U1509 (N_1509,In_1703,In_4953);
nand U1510 (N_1510,In_2464,In_4224);
and U1511 (N_1511,In_1108,In_3277);
nand U1512 (N_1512,In_1456,In_3980);
nor U1513 (N_1513,In_1792,In_2843);
or U1514 (N_1514,In_4793,In_2756);
nor U1515 (N_1515,In_1743,In_3685);
or U1516 (N_1516,In_3824,In_4012);
nor U1517 (N_1517,In_3722,In_2125);
and U1518 (N_1518,In_1759,In_1024);
and U1519 (N_1519,In_3754,In_2623);
nor U1520 (N_1520,In_3077,In_755);
nand U1521 (N_1521,In_508,In_3279);
or U1522 (N_1522,In_142,In_4474);
and U1523 (N_1523,In_2798,In_4913);
nor U1524 (N_1524,In_306,In_4556);
nand U1525 (N_1525,In_2628,In_1347);
nor U1526 (N_1526,In_3480,In_3951);
nor U1527 (N_1527,In_952,In_4188);
or U1528 (N_1528,In_2137,In_1661);
nor U1529 (N_1529,In_2536,In_2993);
nor U1530 (N_1530,In_495,In_52);
nor U1531 (N_1531,In_1776,In_4789);
nor U1532 (N_1532,In_1814,In_3638);
or U1533 (N_1533,In_1049,In_4086);
nor U1534 (N_1534,In_981,In_3228);
and U1535 (N_1535,In_4737,In_3372);
nor U1536 (N_1536,In_3626,In_612);
and U1537 (N_1537,In_4415,In_2112);
or U1538 (N_1538,In_363,In_260);
and U1539 (N_1539,In_4911,In_685);
nor U1540 (N_1540,In_4389,In_4346);
and U1541 (N_1541,In_327,In_3438);
and U1542 (N_1542,In_955,In_4209);
or U1543 (N_1543,In_3429,In_12);
and U1544 (N_1544,In_698,In_2788);
nor U1545 (N_1545,In_2583,In_3406);
nand U1546 (N_1546,In_217,In_2961);
nor U1547 (N_1547,In_2624,In_1679);
nor U1548 (N_1548,In_2210,In_723);
nand U1549 (N_1549,In_99,In_1705);
and U1550 (N_1550,In_1197,In_1392);
nand U1551 (N_1551,In_4949,In_2159);
and U1552 (N_1552,In_3735,In_760);
and U1553 (N_1553,In_3435,In_3513);
or U1554 (N_1554,In_1428,In_4892);
nor U1555 (N_1555,In_2147,In_2456);
or U1556 (N_1556,In_4786,In_4507);
or U1557 (N_1557,In_207,In_1368);
xnor U1558 (N_1558,In_1605,In_2713);
and U1559 (N_1559,In_1497,In_1433);
nand U1560 (N_1560,In_2767,In_925);
and U1561 (N_1561,In_1909,In_2142);
nand U1562 (N_1562,In_4098,In_2118);
or U1563 (N_1563,In_1439,In_2397);
and U1564 (N_1564,In_108,In_3235);
nor U1565 (N_1565,In_3560,In_3485);
or U1566 (N_1566,In_291,In_2177);
or U1567 (N_1567,In_1320,In_2705);
nand U1568 (N_1568,In_2407,In_2168);
and U1569 (N_1569,In_2730,In_790);
nor U1570 (N_1570,In_2013,In_4660);
nor U1571 (N_1571,In_1301,In_654);
and U1572 (N_1572,In_3045,In_451);
nand U1573 (N_1573,In_1488,In_2507);
nand U1574 (N_1574,In_4674,In_3797);
nor U1575 (N_1575,In_3593,In_4320);
and U1576 (N_1576,In_91,In_4438);
or U1577 (N_1577,In_802,In_2711);
nand U1578 (N_1578,In_2598,In_1149);
nor U1579 (N_1579,In_1757,In_4734);
or U1580 (N_1580,In_4339,In_3577);
or U1581 (N_1581,In_818,In_1418);
xor U1582 (N_1582,In_3268,In_1354);
and U1583 (N_1583,In_2582,In_2244);
or U1584 (N_1584,In_2501,In_1394);
nand U1585 (N_1585,In_1643,In_4155);
nand U1586 (N_1586,In_3112,In_4535);
nand U1587 (N_1587,In_1026,In_1847);
nand U1588 (N_1588,In_522,In_194);
and U1589 (N_1589,In_911,In_1395);
nor U1590 (N_1590,In_4864,In_1829);
nor U1591 (N_1591,In_3318,In_2058);
nand U1592 (N_1592,In_1242,In_4125);
nand U1593 (N_1593,In_4047,In_4760);
nor U1594 (N_1594,In_2279,In_4435);
or U1595 (N_1595,In_2608,In_3587);
and U1596 (N_1596,In_4398,In_670);
and U1597 (N_1597,In_4683,In_1280);
nand U1598 (N_1598,In_2067,In_4081);
nor U1599 (N_1599,In_1067,In_2019);
and U1600 (N_1600,In_3154,In_1687);
or U1601 (N_1601,In_2587,In_2700);
nand U1602 (N_1602,In_28,In_4365);
nor U1603 (N_1603,In_918,In_198);
nor U1604 (N_1604,In_1097,In_412);
and U1605 (N_1605,In_4635,In_3248);
and U1606 (N_1606,In_1464,In_311);
or U1607 (N_1607,In_4055,In_4095);
or U1608 (N_1608,In_1853,In_3816);
nor U1609 (N_1609,In_2896,In_3601);
and U1610 (N_1610,In_2224,In_2312);
nor U1611 (N_1611,In_850,In_871);
nand U1612 (N_1612,In_3686,In_596);
or U1613 (N_1613,In_3881,In_2068);
nand U1614 (N_1614,In_653,In_270);
and U1615 (N_1615,In_4039,In_1264);
nand U1616 (N_1616,In_2825,In_4882);
and U1617 (N_1617,In_3255,In_4404);
or U1618 (N_1618,In_2618,In_4192);
nand U1619 (N_1619,In_4584,In_1589);
and U1620 (N_1620,In_2539,In_842);
nor U1621 (N_1621,In_2482,In_3294);
nor U1622 (N_1622,In_1558,In_1565);
or U1623 (N_1623,In_4823,In_3732);
or U1624 (N_1624,In_1539,In_1882);
nand U1625 (N_1625,In_2983,In_1580);
and U1626 (N_1626,In_1786,In_4983);
nand U1627 (N_1627,In_206,In_390);
or U1628 (N_1628,In_1017,In_2427);
nor U1629 (N_1629,In_1117,In_2826);
or U1630 (N_1630,In_1095,In_821);
and U1631 (N_1631,In_4458,In_3374);
and U1632 (N_1632,In_4016,In_1714);
nand U1633 (N_1633,In_2445,In_3953);
nand U1634 (N_1634,In_2595,In_221);
nor U1635 (N_1635,In_3589,In_3296);
nand U1636 (N_1636,In_4196,In_3101);
and U1637 (N_1637,In_88,In_1131);
nand U1638 (N_1638,In_2953,In_196);
nor U1639 (N_1639,In_4891,In_527);
or U1640 (N_1640,In_344,In_3257);
and U1641 (N_1641,In_4588,In_3032);
and U1642 (N_1642,In_1612,In_1407);
nand U1643 (N_1643,In_2578,In_4896);
nor U1644 (N_1644,In_4140,In_2365);
or U1645 (N_1645,In_3974,In_940);
or U1646 (N_1646,In_4464,In_1483);
nand U1647 (N_1647,In_140,In_2977);
and U1648 (N_1648,In_994,In_833);
and U1649 (N_1649,In_4257,In_4530);
xor U1650 (N_1650,In_2278,In_1723);
nor U1651 (N_1651,In_3678,In_2100);
xor U1652 (N_1652,In_225,In_2956);
or U1653 (N_1653,In_4990,In_313);
nand U1654 (N_1654,In_168,In_3200);
xnor U1655 (N_1655,In_2473,In_2617);
nor U1656 (N_1656,In_756,In_2371);
nand U1657 (N_1657,In_2433,In_2226);
or U1658 (N_1658,In_1638,In_1515);
or U1659 (N_1659,In_4388,In_462);
and U1660 (N_1660,In_2252,In_415);
nor U1661 (N_1661,In_1815,In_3285);
nor U1662 (N_1662,In_4821,In_2833);
nor U1663 (N_1663,In_4350,In_1512);
or U1664 (N_1664,In_2947,In_4181);
or U1665 (N_1665,In_1937,In_4800);
or U1666 (N_1666,In_4689,In_2928);
and U1667 (N_1667,In_2884,In_4080);
nand U1668 (N_1668,In_1341,In_1122);
nor U1669 (N_1669,In_4429,In_688);
xnor U1670 (N_1670,In_2808,In_103);
nor U1671 (N_1671,In_4751,In_482);
and U1672 (N_1672,In_1999,In_3461);
nor U1673 (N_1673,In_4330,In_4966);
or U1674 (N_1674,In_3038,In_2233);
nand U1675 (N_1675,In_2958,In_609);
or U1676 (N_1676,In_1007,In_3008);
nor U1677 (N_1677,In_1036,In_2479);
nand U1678 (N_1678,In_1399,In_3937);
nor U1679 (N_1679,In_1221,In_45);
or U1680 (N_1680,In_2421,In_615);
nand U1681 (N_1681,In_4475,In_1011);
nor U1682 (N_1682,In_3906,In_4612);
and U1683 (N_1683,In_4364,In_2610);
nor U1684 (N_1684,In_2018,In_104);
and U1685 (N_1685,In_3418,In_1228);
or U1686 (N_1686,In_2028,In_1968);
xor U1687 (N_1687,In_4560,In_1268);
and U1688 (N_1688,In_2575,In_229);
and U1689 (N_1689,In_3605,In_2163);
or U1690 (N_1690,In_2919,In_3460);
nor U1691 (N_1691,In_4860,In_4923);
and U1692 (N_1692,In_3080,In_678);
or U1693 (N_1693,In_1344,In_450);
nand U1694 (N_1694,In_1470,In_3298);
nor U1695 (N_1695,In_74,In_2396);
nor U1696 (N_1696,In_951,In_4498);
or U1697 (N_1697,In_2281,In_162);
or U1698 (N_1698,In_4374,In_1413);
or U1699 (N_1699,In_2981,In_4812);
or U1700 (N_1700,In_3622,In_4616);
or U1701 (N_1701,In_1805,In_1644);
and U1702 (N_1702,In_3025,In_3613);
nand U1703 (N_1703,In_3488,In_4384);
nand U1704 (N_1704,In_3555,In_1076);
nand U1705 (N_1705,In_115,In_3657);
nand U1706 (N_1706,In_3539,In_4227);
nand U1707 (N_1707,In_4659,In_3421);
xnor U1708 (N_1708,In_4341,In_3288);
or U1709 (N_1709,In_4590,In_4539);
xnor U1710 (N_1710,In_4844,In_708);
nand U1711 (N_1711,In_2720,In_1718);
nor U1712 (N_1712,In_4104,In_2369);
nor U1713 (N_1713,In_3519,In_4101);
nor U1714 (N_1714,In_4627,In_215);
nor U1715 (N_1715,In_2098,In_4916);
nor U1716 (N_1716,In_783,In_1557);
nand U1717 (N_1717,In_4048,In_3666);
nand U1718 (N_1718,In_3065,In_3954);
and U1719 (N_1719,In_1326,In_210);
nand U1720 (N_1720,In_1337,In_3699);
or U1721 (N_1721,In_2124,In_2576);
or U1722 (N_1722,In_2298,In_1807);
and U1723 (N_1723,In_4688,In_2894);
and U1724 (N_1724,In_2041,In_1378);
nand U1725 (N_1725,In_1571,In_205);
or U1726 (N_1726,In_3174,In_4646);
or U1727 (N_1727,In_339,In_4642);
nand U1728 (N_1728,In_3854,In_1583);
nor U1729 (N_1729,In_1047,In_1513);
or U1730 (N_1730,In_1429,In_1227);
nand U1731 (N_1731,In_137,In_2005);
and U1732 (N_1732,In_2888,In_696);
or U1733 (N_1733,In_3199,In_4060);
nand U1734 (N_1734,In_4451,In_751);
or U1735 (N_1735,In_61,In_1907);
and U1736 (N_1736,In_2139,In_932);
nand U1737 (N_1737,In_1840,In_4492);
and U1738 (N_1738,In_2327,In_1657);
and U1739 (N_1739,In_1234,In_945);
and U1740 (N_1740,In_4750,In_845);
or U1741 (N_1741,In_3647,In_181);
or U1742 (N_1742,In_3258,In_1543);
nor U1743 (N_1743,In_383,In_3999);
xor U1744 (N_1744,In_2030,In_2103);
nand U1745 (N_1745,In_3143,In_4541);
nand U1746 (N_1746,In_506,In_1806);
or U1747 (N_1747,In_69,In_3850);
or U1748 (N_1748,In_1780,In_4876);
and U1749 (N_1749,In_378,In_941);
and U1750 (N_1750,In_2743,In_432);
nand U1751 (N_1751,In_1976,In_403);
or U1752 (N_1752,In_2759,In_2739);
and U1753 (N_1753,In_4569,In_1499);
nand U1754 (N_1754,In_1750,In_1492);
nand U1755 (N_1755,In_2193,In_1386);
or U1756 (N_1756,In_2579,In_3719);
nor U1757 (N_1757,In_2511,In_4436);
nor U1758 (N_1758,In_4787,In_564);
nor U1759 (N_1759,In_3639,In_3159);
nand U1760 (N_1760,In_2534,In_4548);
xor U1761 (N_1761,In_4550,In_2957);
and U1762 (N_1762,In_843,In_3729);
or U1763 (N_1763,In_4785,In_170);
nand U1764 (N_1764,In_95,In_3344);
or U1765 (N_1765,In_3963,In_18);
or U1766 (N_1766,In_1229,In_2815);
or U1767 (N_1767,In_3800,In_2859);
and U1768 (N_1768,In_3310,In_4825);
nor U1769 (N_1769,In_593,In_4259);
nor U1770 (N_1770,In_792,In_666);
and U1771 (N_1771,In_1322,In_3683);
nor U1772 (N_1772,In_1982,In_2741);
and U1773 (N_1773,In_195,In_4603);
and U1774 (N_1774,In_4264,In_3307);
and U1775 (N_1775,In_3659,In_1768);
nand U1776 (N_1776,In_4925,In_4641);
xnor U1777 (N_1777,In_4373,In_442);
nor U1778 (N_1778,In_474,In_4557);
and U1779 (N_1779,In_3928,In_3789);
and U1780 (N_1780,In_2074,In_3212);
nand U1781 (N_1781,In_329,In_4718);
nand U1782 (N_1782,In_3808,In_4026);
or U1783 (N_1783,In_4955,In_998);
nand U1784 (N_1784,In_3259,In_2218);
nand U1785 (N_1785,In_256,In_817);
or U1786 (N_1786,In_1602,In_3022);
nand U1787 (N_1787,In_558,In_3916);
or U1788 (N_1788,In_83,In_4053);
nand U1789 (N_1789,In_583,In_594);
and U1790 (N_1790,In_2863,In_1816);
or U1791 (N_1791,In_1505,In_4046);
nor U1792 (N_1792,In_2671,In_2286);
or U1793 (N_1793,In_2972,In_2721);
and U1794 (N_1794,In_602,In_3528);
nand U1795 (N_1795,In_1086,In_2701);
or U1796 (N_1796,In_4661,In_89);
nor U1797 (N_1797,In_93,In_200);
or U1798 (N_1798,In_3487,In_2545);
and U1799 (N_1799,In_2315,In_2347);
or U1800 (N_1800,In_354,In_3614);
nand U1801 (N_1801,In_2878,In_2769);
nand U1802 (N_1802,In_391,In_4631);
or U1803 (N_1803,In_1956,In_735);
nand U1804 (N_1804,In_1292,In_2974);
and U1805 (N_1805,In_4711,In_1362);
and U1806 (N_1806,In_4115,In_3726);
nor U1807 (N_1807,In_1183,In_1475);
or U1808 (N_1808,In_3557,In_1567);
nand U1809 (N_1809,In_4061,In_4433);
nor U1810 (N_1810,In_4444,In_767);
nand U1811 (N_1811,In_4434,In_2431);
and U1812 (N_1812,In_2205,In_1285);
xor U1813 (N_1813,In_2722,In_3264);
nand U1814 (N_1814,In_4960,In_3820);
and U1815 (N_1815,In_3026,In_2724);
nor U1816 (N_1816,In_3787,In_3582);
nand U1817 (N_1817,In_1698,In_1845);
nand U1818 (N_1818,In_109,In_1994);
nand U1819 (N_1819,In_58,In_1756);
and U1820 (N_1820,In_4462,In_1283);
nand U1821 (N_1821,In_90,In_465);
nor U1822 (N_1822,In_1224,In_4179);
nor U1823 (N_1823,In_533,In_1359);
and U1824 (N_1824,In_1374,In_1239);
and U1825 (N_1825,In_4903,In_870);
xnor U1826 (N_1826,In_742,In_3013);
and U1827 (N_1827,In_1013,In_173);
xor U1828 (N_1828,In_4409,In_530);
or U1829 (N_1829,In_148,In_913);
nor U1830 (N_1830,In_1662,In_2816);
and U1831 (N_1831,In_4493,In_3505);
nor U1832 (N_1832,In_2885,In_4574);
nor U1833 (N_1833,In_4885,In_2558);
nor U1834 (N_1834,In_3584,In_4639);
nand U1835 (N_1835,In_4284,In_2876);
and U1836 (N_1836,In_2989,In_3413);
nor U1837 (N_1837,In_4933,In_1085);
nor U1838 (N_1838,In_4950,In_66);
or U1839 (N_1839,In_539,In_2882);
or U1840 (N_1840,In_3342,In_2780);
nor U1841 (N_1841,In_1728,In_4175);
xnor U1842 (N_1842,In_3169,In_4442);
or U1843 (N_1843,In_3284,In_1107);
or U1844 (N_1844,In_1041,In_827);
and U1845 (N_1845,In_3079,In_1424);
nand U1846 (N_1846,In_2719,In_4430);
nor U1847 (N_1847,In_4182,In_2652);
nand U1848 (N_1848,In_3736,In_1906);
nor U1849 (N_1849,In_4211,In_4811);
and U1850 (N_1850,In_2837,In_3370);
nand U1851 (N_1851,In_4122,In_4775);
or U1852 (N_1852,In_1934,In_4296);
and U1853 (N_1853,In_4843,In_591);
and U1854 (N_1854,In_1030,In_2904);
nor U1855 (N_1855,In_1369,In_4001);
and U1856 (N_1856,In_1411,In_268);
xnor U1857 (N_1857,In_4401,In_2354);
nand U1858 (N_1858,In_929,In_661);
or U1859 (N_1859,In_258,In_912);
nand U1860 (N_1860,In_4620,In_4174);
nand U1861 (N_1861,In_4014,In_154);
nand U1862 (N_1862,In_1509,In_1746);
and U1863 (N_1863,In_1613,In_4849);
nor U1864 (N_1864,In_2409,In_4826);
or U1865 (N_1865,In_4153,In_3658);
and U1866 (N_1866,In_3353,In_3738);
or U1867 (N_1867,In_1656,In_113);
nor U1868 (N_1868,In_3943,In_1710);
nand U1869 (N_1869,In_1210,In_1376);
nor U1870 (N_1870,In_4405,In_1152);
nand U1871 (N_1871,In_4217,In_772);
nand U1872 (N_1872,In_1454,In_869);
nand U1873 (N_1873,In_3238,In_3634);
or U1874 (N_1874,In_4226,In_3237);
or U1875 (N_1875,In_4070,In_445);
nand U1876 (N_1876,In_4929,In_3715);
nor U1877 (N_1877,In_3680,In_4987);
or U1878 (N_1878,In_1263,In_3105);
or U1879 (N_1879,In_1098,In_479);
nand U1880 (N_1880,In_3865,In_4962);
nand U1881 (N_1881,In_1104,In_3151);
nor U1882 (N_1882,In_3780,In_3724);
or U1883 (N_1883,In_4919,In_2114);
or U1884 (N_1884,In_3880,In_4883);
or U1885 (N_1885,In_1408,In_924);
nor U1886 (N_1886,In_3747,In_4625);
nand U1887 (N_1887,In_1031,In_861);
xor U1888 (N_1888,In_1311,In_96);
or U1889 (N_1889,In_263,In_848);
nand U1890 (N_1890,In_1957,In_3126);
nand U1891 (N_1891,In_1215,In_218);
and U1892 (N_1892,In_1113,In_2282);
or U1893 (N_1893,In_4305,In_2015);
and U1894 (N_1894,In_4062,In_3040);
or U1895 (N_1895,In_4044,In_1353);
nor U1896 (N_1896,In_973,In_3753);
nor U1897 (N_1897,In_2555,In_2659);
xnor U1898 (N_1898,In_4332,In_3191);
or U1899 (N_1899,In_2985,In_1109);
nor U1900 (N_1900,In_2063,In_3791);
xnor U1901 (N_1901,In_1129,In_943);
nor U1902 (N_1902,In_4476,In_1371);
or U1903 (N_1903,In_290,In_3643);
and U1904 (N_1904,In_2731,In_3201);
or U1905 (N_1905,In_1791,In_3451);
or U1906 (N_1906,In_4921,In_231);
nand U1907 (N_1907,In_3524,In_4668);
nand U1908 (N_1908,In_1328,In_1111);
and U1909 (N_1909,In_2449,In_3447);
and U1910 (N_1910,In_4840,In_3776);
nor U1911 (N_1911,In_2827,In_2680);
or U1912 (N_1912,In_3997,In_1423);
nand U1913 (N_1913,In_1541,In_4610);
and U1914 (N_1914,In_2346,In_3015);
or U1915 (N_1915,In_1452,In_598);
and U1916 (N_1916,In_1809,In_3397);
or U1917 (N_1917,In_4790,In_3648);
or U1918 (N_1918,In_3500,In_1933);
and U1919 (N_1919,In_4321,In_151);
and U1920 (N_1920,In_2106,In_19);
nor U1921 (N_1921,In_4387,In_32);
and U1922 (N_1922,In_4922,In_4509);
and U1923 (N_1923,In_1027,In_248);
nor U1924 (N_1924,In_3230,In_3110);
nand U1925 (N_1925,In_82,In_2059);
nand U1926 (N_1926,In_872,In_4009);
and U1927 (N_1927,In_3632,In_4402);
or U1928 (N_1928,In_3321,In_1078);
and U1929 (N_1929,In_1482,In_1989);
xor U1930 (N_1930,In_3799,In_2920);
nor U1931 (N_1931,In_799,In_1385);
or U1932 (N_1932,In_3445,In_1970);
or U1933 (N_1933,In_4815,In_4931);
or U1934 (N_1934,In_4189,In_2568);
and U1935 (N_1935,In_3796,In_2155);
nand U1936 (N_1936,In_3437,In_497);
nand U1937 (N_1937,In_1749,In_4352);
nand U1938 (N_1938,In_934,In_857);
or U1939 (N_1939,In_2693,In_811);
nand U1940 (N_1940,In_1446,In_1680);
nand U1941 (N_1941,In_1901,In_4129);
nor U1942 (N_1942,In_3163,In_73);
nor U1943 (N_1943,In_4484,In_2986);
or U1944 (N_1944,In_630,In_4930);
nand U1945 (N_1945,In_239,In_3939);
nand U1946 (N_1946,In_408,In_3399);
or U1947 (N_1947,In_2869,In_280);
xnor U1948 (N_1948,In_4156,In_2097);
nor U1949 (N_1949,In_285,In_3993);
nor U1950 (N_1950,In_4260,In_4522);
nand U1951 (N_1951,In_2502,In_4723);
nand U1952 (N_1952,In_1922,In_3701);
or U1953 (N_1953,In_2707,In_117);
nor U1954 (N_1954,In_2002,In_3203);
nor U1955 (N_1955,In_1764,In_476);
and U1956 (N_1956,In_2612,In_3289);
nand U1957 (N_1957,In_3336,In_3153);
and U1958 (N_1958,In_2364,In_4482);
and U1959 (N_1959,In_3618,In_1455);
nor U1960 (N_1960,In_1987,In_1542);
nand U1961 (N_1961,In_2026,In_2136);
nand U1962 (N_1962,In_3839,In_1373);
nand U1963 (N_1963,In_4980,In_1597);
or U1964 (N_1964,In_3924,In_3417);
and U1965 (N_1965,In_3128,In_3863);
nand U1966 (N_1966,In_165,In_3723);
nor U1967 (N_1967,In_4783,In_2900);
and U1968 (N_1968,In_346,In_553);
nor U1969 (N_1969,In_2391,In_4212);
nand U1970 (N_1970,In_416,In_351);
and U1971 (N_1971,In_1174,In_4231);
nor U1972 (N_1972,In_3970,In_649);
nor U1973 (N_1973,In_1231,In_3499);
and U1974 (N_1974,In_1372,In_1755);
nor U1975 (N_1975,In_700,In_3758);
or U1976 (N_1976,In_4670,In_325);
nand U1977 (N_1977,In_2784,In_4694);
nor U1978 (N_1978,In_2009,In_4813);
or U1979 (N_1979,In_740,In_4745);
nor U1980 (N_1980,In_892,In_4848);
and U1981 (N_1981,In_4327,In_4035);
nor U1982 (N_1982,In_2487,In_298);
or U1983 (N_1983,In_332,In_1967);
or U1984 (N_1984,In_3115,In_2609);
nor U1985 (N_1985,In_2127,In_2679);
and U1986 (N_1986,In_4054,In_4031);
nor U1987 (N_1987,In_3929,In_4715);
or U1988 (N_1988,In_3673,In_710);
and U1989 (N_1989,In_3104,In_358);
or U1990 (N_1990,In_1071,In_2916);
or U1991 (N_1991,In_2367,In_2001);
nand U1992 (N_1992,In_4146,In_1193);
and U1993 (N_1993,In_2172,In_433);
nor U1994 (N_1994,In_2008,In_1273);
nand U1995 (N_1995,In_1496,In_3764);
nand U1996 (N_1996,In_559,In_259);
nor U1997 (N_1997,In_1172,In_4281);
or U1998 (N_1998,In_2914,In_954);
and U1999 (N_1999,In_253,In_2508);
and U2000 (N_2000,N_1664,N_294);
or U2001 (N_2001,N_775,N_971);
or U2002 (N_2002,N_801,N_452);
nand U2003 (N_2003,N_1275,N_1366);
and U2004 (N_2004,N_826,In_2006);
nand U2005 (N_2005,N_904,N_1018);
nor U2006 (N_2006,N_148,In_629);
xor U2007 (N_2007,N_1623,N_43);
nor U2008 (N_2008,N_1154,In_1465);
and U2009 (N_2009,N_828,In_1616);
nand U2010 (N_2010,In_2688,N_1435);
and U2011 (N_2011,In_4915,In_222);
and U2012 (N_2012,N_1989,N_1469);
nor U2013 (N_2013,In_2404,N_170);
or U2014 (N_2014,In_1451,N_1607);
nor U2015 (N_2015,In_3848,N_264);
or U2016 (N_2016,In_4799,N_1026);
and U2017 (N_2017,N_479,N_974);
nor U2018 (N_2018,N_1001,In_1707);
or U2019 (N_2019,In_110,N_1629);
or U2020 (N_2020,N_1178,N_134);
or U2021 (N_2021,N_933,In_3313);
or U2022 (N_2022,In_464,N_131);
and U2023 (N_2023,In_3325,In_1642);
or U2024 (N_2024,N_768,N_144);
or U2025 (N_2025,N_1619,N_1176);
nand U2026 (N_2026,N_1819,In_584);
or U2027 (N_2027,N_389,N_310);
nor U2028 (N_2028,N_1695,In_4587);
and U2029 (N_2029,In_3000,In_177);
nor U2030 (N_2030,N_1875,N_525);
and U2031 (N_2031,N_1080,N_1155);
nor U2032 (N_2032,N_313,In_997);
and U2033 (N_2033,In_2512,N_1381);
and U2034 (N_2034,N_1598,N_1966);
nand U2035 (N_2035,N_1417,N_100);
and U2036 (N_2036,In_3788,In_3006);
nor U2037 (N_2037,N_1064,In_2762);
or U2038 (N_2038,N_318,N_1347);
or U2039 (N_2039,In_3047,N_488);
and U2040 (N_2040,N_1065,N_1451);
nand U2041 (N_2041,In_489,N_1864);
nor U2042 (N_2042,N_1359,In_2726);
or U2043 (N_2043,N_684,N_33);
and U2044 (N_2044,N_1218,N_1765);
or U2045 (N_2045,N_1112,N_1811);
and U2046 (N_2046,N_1676,N_965);
and U2047 (N_2047,N_633,In_3448);
nand U2048 (N_2048,N_512,In_1406);
and U2049 (N_2049,N_699,N_917);
or U2050 (N_2050,In_4190,N_436);
and U2051 (N_2051,N_618,N_1004);
or U2052 (N_2052,In_4020,N_1999);
nand U2053 (N_2053,N_1661,N_1358);
and U2054 (N_2054,N_231,N_1401);
and U2055 (N_2055,N_1856,N_1471);
nand U2056 (N_2056,In_3653,In_1673);
nand U2057 (N_2057,In_2428,N_1956);
nand U2058 (N_2058,N_276,N_1195);
nor U2059 (N_2059,N_1171,In_1171);
or U2060 (N_2060,In_4640,In_2146);
nor U2061 (N_2061,N_1031,In_2907);
or U2062 (N_2062,In_3552,N_536);
xnor U2063 (N_2063,In_2750,N_161);
nand U2064 (N_2064,N_1774,N_173);
nand U2065 (N_2065,N_261,In_2050);
nor U2066 (N_2066,N_157,In_3637);
and U2067 (N_2067,N_493,In_491);
and U2068 (N_2068,N_1878,N_766);
xnor U2069 (N_2069,N_1759,In_1202);
and U2070 (N_2070,N_1149,In_425);
nand U2071 (N_2071,In_2248,N_1115);
nand U2072 (N_2072,N_785,In_414);
and U2073 (N_2073,In_350,N_1309);
xor U2074 (N_2074,In_1318,N_657);
nand U2075 (N_2075,In_1865,N_1260);
nand U2076 (N_2076,N_915,N_353);
nand U2077 (N_2077,N_196,N_870);
and U2078 (N_2078,N_335,N_1280);
and U2079 (N_2079,In_10,In_4657);
nor U2080 (N_2080,In_4968,In_1075);
or U2081 (N_2081,N_150,N_991);
and U2082 (N_2082,In_2380,N_1543);
nor U2083 (N_2083,N_1046,N_172);
xnor U2084 (N_2084,In_2213,In_1137);
nand U2085 (N_2085,N_1750,N_1407);
and U2086 (N_2086,In_4347,In_4323);
or U2087 (N_2087,In_623,N_1785);
nand U2088 (N_2088,N_645,In_1222);
and U2089 (N_2089,N_1749,N_1170);
and U2090 (N_2090,N_485,N_760);
nand U2091 (N_2091,N_8,N_1457);
nand U2092 (N_2092,N_1207,In_1726);
and U2093 (N_2093,In_694,N_1893);
nor U2094 (N_2094,In_1700,N_1715);
nand U2095 (N_2095,N_115,N_797);
and U2096 (N_2096,N_985,N_240);
nand U2097 (N_2097,N_1644,N_0);
nor U2098 (N_2098,N_1883,N_1040);
and U2099 (N_2099,N_1116,N_1194);
nor U2100 (N_2100,N_1191,In_3782);
nand U2101 (N_2101,N_486,N_1498);
nand U2102 (N_2102,In_1622,N_1432);
nor U2103 (N_2103,In_328,N_1888);
nor U2104 (N_2104,N_234,N_1865);
nor U2105 (N_2105,N_95,N_1698);
nand U2106 (N_2106,N_208,In_179);
nor U2107 (N_2107,N_117,N_1125);
and U2108 (N_2108,N_959,N_204);
or U2109 (N_2109,N_1914,N_1775);
or U2110 (N_2110,N_783,N_744);
and U2111 (N_2111,N_1187,N_1078);
nand U2112 (N_2112,In_3234,In_348);
and U2113 (N_2113,N_725,In_2842);
nand U2114 (N_2114,In_2085,In_2161);
or U2115 (N_2115,N_96,In_2615);
xor U2116 (N_2116,N_1494,N_1103);
or U2117 (N_2117,N_1468,N_1434);
and U2118 (N_2118,N_219,In_1427);
and U2119 (N_2119,In_2514,In_2889);
nand U2120 (N_2120,N_1320,N_1674);
or U2121 (N_2121,In_1192,N_1671);
or U2122 (N_2122,N_1074,N_862);
or U2123 (N_2123,In_1581,N_1919);
or U2124 (N_2124,N_709,N_260);
nor U2125 (N_2125,In_854,In_717);
nor U2126 (N_2126,In_3925,N_542);
nand U2127 (N_2127,N_1660,In_1009);
nand U2128 (N_2128,In_4884,In_4733);
or U2129 (N_2129,N_563,In_927);
nand U2130 (N_2130,In_1176,N_1537);
xnor U2131 (N_2131,N_659,N_1473);
or U2132 (N_2132,In_2062,In_233);
nand U2133 (N_2133,In_4965,N_37);
nand U2134 (N_2134,In_3805,In_4549);
nor U2135 (N_2135,N_1860,In_3755);
or U2136 (N_2136,N_1076,In_1245);
nand U2137 (N_2137,N_327,N_1834);
and U2138 (N_2138,N_1995,In_575);
nor U2139 (N_2139,In_2976,N_742);
or U2140 (N_2140,N_564,N_1525);
xor U2141 (N_2141,N_1981,N_1464);
and U2142 (N_2142,N_1615,N_1997);
or U2143 (N_2143,In_677,In_3870);
nor U2144 (N_2144,N_1102,N_1789);
nor U2145 (N_2145,N_494,In_1547);
nand U2146 (N_2146,N_1497,In_987);
or U2147 (N_2147,In_917,N_65);
and U2148 (N_2148,N_1073,In_2258);
nor U2149 (N_2149,N_500,N_1418);
or U2150 (N_2150,N_929,N_325);
or U2151 (N_2151,N_859,In_1057);
nand U2152 (N_2152,N_805,N_1573);
or U2153 (N_2153,N_1005,N_832);
nor U2154 (N_2154,N_1262,N_1304);
and U2155 (N_2155,N_387,N_139);
and U2156 (N_2156,N_1727,N_1089);
nor U2157 (N_2157,N_1814,In_4297);
and U2158 (N_2158,N_1612,In_4478);
nand U2159 (N_2159,N_545,N_1202);
and U2160 (N_2160,N_395,N_1797);
nand U2161 (N_2161,N_995,N_1441);
and U2162 (N_2162,N_504,N_118);
nand U2163 (N_2163,N_601,N_1386);
and U2164 (N_2164,N_1265,In_2024);
or U2165 (N_2165,In_3878,N_943);
or U2166 (N_2166,In_3452,In_2307);
nand U2167 (N_2167,N_1662,In_1006);
nand U2168 (N_2168,In_3020,N_1338);
nor U2169 (N_2169,N_1458,N_1523);
or U2170 (N_2170,N_1688,N_1459);
nand U2171 (N_2171,N_1375,N_1571);
and U2172 (N_2172,In_1437,N_1602);
nor U2173 (N_2173,N_873,N_1060);
nor U2174 (N_2174,N_1673,N_60);
or U2175 (N_2175,In_1198,N_508);
and U2176 (N_2176,N_1857,In_4672);
and U2177 (N_2177,In_2834,N_390);
and U2178 (N_2178,N_680,In_3095);
nor U2179 (N_2179,N_1736,N_619);
nand U2180 (N_2180,N_632,N_171);
and U2181 (N_2181,In_342,N_1649);
nand U2182 (N_2182,In_853,N_228);
nor U2183 (N_2183,N_1693,In_1785);
or U2184 (N_2184,In_1323,In_3570);
or U2185 (N_2185,N_1488,N_582);
or U2186 (N_2186,N_872,N_654);
nor U2187 (N_2187,N_1861,In_4872);
or U2188 (N_2188,N_45,N_1740);
nand U2189 (N_2189,N_592,N_370);
nor U2190 (N_2190,N_286,N_954);
and U2191 (N_2191,N_1420,N_1166);
and U2192 (N_2192,In_4285,In_4992);
nor U2193 (N_2193,N_371,N_896);
or U2194 (N_2194,N_1576,N_356);
or U2195 (N_2195,N_1315,N_573);
or U2196 (N_2196,N_983,N_1217);
and U2197 (N_2197,In_2580,In_4663);
and U2198 (N_2198,In_3768,N_503);
xor U2199 (N_2199,N_1447,N_412);
nor U2200 (N_2200,N_1561,N_1354);
nor U2201 (N_2201,N_1540,In_2084);
nand U2202 (N_2202,N_738,In_2932);
nand U2203 (N_2203,N_1820,In_2486);
nor U2204 (N_2204,N_1762,N_1290);
or U2205 (N_2205,N_1609,In_3263);
nand U2206 (N_2206,N_185,N_112);
xnor U2207 (N_2207,In_4108,In_1731);
and U2208 (N_2208,N_711,N_1744);
and U2209 (N_2209,N_1419,In_3707);
or U2210 (N_2210,N_1379,In_477);
and U2211 (N_2211,In_2424,N_1168);
nand U2212 (N_2212,N_1737,N_346);
nand U2213 (N_2213,N_987,In_3348);
and U2214 (N_2214,N_558,In_2042);
and U2215 (N_2215,N_396,N_1097);
nor U2216 (N_2216,In_4349,N_723);
nor U2217 (N_2217,N_795,In_4112);
or U2218 (N_2218,N_763,N_1985);
or U2219 (N_2219,N_380,N_1397);
xor U2220 (N_2220,N_1872,In_2228);
or U2221 (N_2221,N_1533,N_679);
or U2222 (N_2222,In_60,N_1110);
and U2223 (N_2223,In_1365,In_3581);
and U2224 (N_2224,N_63,N_799);
nor U2225 (N_2225,N_74,N_1686);
nor U2226 (N_2226,N_1146,N_595);
nor U2227 (N_2227,N_569,N_774);
nand U2228 (N_2228,In_671,N_1958);
or U2229 (N_2229,In_1634,N_1942);
or U2230 (N_2230,In_2665,In_1688);
nand U2231 (N_2231,N_1901,N_1274);
nand U2232 (N_2232,In_3152,N_641);
and U2233 (N_2233,In_3991,N_1405);
xor U2234 (N_2234,N_574,In_4954);
nor U2235 (N_2235,In_3396,N_1306);
nor U2236 (N_2236,N_2,N_1563);
nand U2237 (N_2237,N_468,N_1236);
or U2238 (N_2238,N_1200,In_3303);
or U2239 (N_2239,N_379,In_1042);
nand U2240 (N_2240,N_658,N_702);
or U2241 (N_2241,N_1180,N_879);
nor U2242 (N_2242,In_2422,N_1617);
or U2243 (N_2243,In_3373,N_743);
and U2244 (N_2244,In_4147,N_919);
nand U2245 (N_2245,In_785,In_1871);
and U2246 (N_2246,In_3968,N_1164);
nand U2247 (N_2247,N_239,In_4807);
or U2248 (N_2248,N_451,N_1926);
xnor U2249 (N_2249,N_1099,N_938);
nand U2250 (N_2250,In_112,In_773);
nor U2251 (N_2251,In_3623,N_1302);
nor U2252 (N_2252,N_782,N_210);
xor U2253 (N_2253,In_288,In_1858);
and U2254 (N_2254,N_1951,N_1769);
nor U2255 (N_2255,N_643,In_1770);
or U2256 (N_2256,N_1998,N_871);
and U2257 (N_2257,N_806,In_3387);
nand U2258 (N_2258,N_439,N_928);
nor U2259 (N_2259,N_1550,N_693);
and U2260 (N_2260,N_1532,In_3093);
xnor U2261 (N_2261,N_179,N_526);
nor U2262 (N_2262,N_749,N_1931);
nand U2263 (N_2263,N_1876,N_976);
or U2264 (N_2264,N_1029,N_724);
or U2265 (N_2265,N_21,N_1467);
nand U2266 (N_2266,N_850,N_1545);
and U2267 (N_2267,In_3243,In_640);
xnor U2268 (N_2268,N_578,N_1424);
nor U2269 (N_2269,In_1808,N_858);
nor U2270 (N_2270,N_1719,N_302);
and U2271 (N_2271,N_445,N_391);
nand U2272 (N_2272,In_1398,N_233);
nor U2273 (N_2273,N_524,N_469);
nor U2274 (N_2274,In_3905,In_885);
nand U2275 (N_2275,N_1491,N_1758);
xnor U2276 (N_2276,N_275,N_24);
and U2277 (N_2277,In_1584,In_4313);
nand U2278 (N_2278,N_213,In_3527);
nor U2279 (N_2279,N_1882,N_1472);
nor U2280 (N_2280,N_1038,N_1826);
and U2281 (N_2281,N_85,In_3361);
nand U2282 (N_2282,N_577,In_4712);
or U2283 (N_2283,N_258,N_1082);
or U2284 (N_2284,N_540,N_250);
and U2285 (N_2285,N_1433,In_3114);
or U2286 (N_2286,N_1659,N_124);
nand U2287 (N_2287,In_2328,N_175);
and U2288 (N_2288,In_3103,N_1599);
nand U2289 (N_2289,N_72,N_4);
nand U2290 (N_2290,N_1140,In_1173);
nor U2291 (N_2291,N_714,N_423);
and U2292 (N_2292,N_649,N_1530);
xor U2293 (N_2293,N_1224,In_2121);
nand U2294 (N_2294,In_3331,N_565);
nor U2295 (N_2295,N_514,N_813);
and U2296 (N_2296,In_715,N_230);
or U2297 (N_2297,N_1984,N_430);
or U2298 (N_2298,N_1141,N_1173);
and U2299 (N_2299,N_53,N_1792);
and U2300 (N_2300,N_1212,N_77);
and U2301 (N_2301,N_1098,N_1802);
or U2302 (N_2302,In_2918,In_2793);
and U2303 (N_2303,N_424,N_664);
nor U2304 (N_2304,In_1438,N_1753);
or U2305 (N_2305,N_626,N_402);
nor U2306 (N_2306,In_457,N_587);
nand U2307 (N_2307,N_1847,N_1705);
or U2308 (N_2308,In_645,N_793);
and U2309 (N_2309,N_1585,In_1846);
nor U2310 (N_2310,In_4693,N_1186);
and U2311 (N_2311,In_1126,In_202);
nor U2312 (N_2312,In_75,In_1659);
or U2313 (N_2313,In_1118,N_1692);
or U2314 (N_2314,In_1405,In_705);
or U2315 (N_2315,N_1135,N_1685);
or U2316 (N_2316,N_579,N_555);
nand U2317 (N_2317,N_205,In_4432);
or U2318 (N_2318,In_1448,In_4455);
or U2319 (N_2319,In_2708,N_1591);
nand U2320 (N_2320,In_471,N_1292);
nor U2321 (N_2321,In_3580,N_1161);
and U2322 (N_2322,N_1221,N_981);
xnor U2323 (N_2323,In_4928,In_2585);
and U2324 (N_2324,N_94,N_1600);
or U2325 (N_2325,N_413,N_278);
or U2326 (N_2326,In_3050,N_128);
or U2327 (N_2327,In_969,N_613);
and U2328 (N_2328,N_238,N_151);
or U2329 (N_2329,In_2405,In_2637);
xnor U2330 (N_2330,N_481,In_1559);
and U2331 (N_2331,In_2119,N_638);
nor U2332 (N_2332,N_1858,In_2254);
or U2333 (N_2333,In_246,In_2521);
nand U2334 (N_2334,N_820,In_4392);
xnor U2335 (N_2335,N_366,N_67);
nor U2336 (N_2336,N_265,In_2789);
and U2337 (N_2337,In_4058,In_34);
nand U2338 (N_2338,N_1908,N_1158);
and U2339 (N_2339,N_1487,N_1970);
nand U2340 (N_2340,N_1798,In_2081);
nor U2341 (N_2341,In_4685,N_897);
nand U2342 (N_2342,N_1106,N_1936);
and U2343 (N_2343,In_3492,N_1075);
or U2344 (N_2344,In_4981,In_4380);
or U2345 (N_2345,N_1474,In_824);
nor U2346 (N_2346,In_1355,In_4879);
nand U2347 (N_2347,N_1070,N_1336);
and U2348 (N_2348,N_1890,In_589);
and U2349 (N_2349,N_952,N_947);
and U2350 (N_2350,N_843,N_1638);
nor U2351 (N_2351,In_2392,In_4997);
and U2352 (N_2352,N_1949,In_3962);
and U2353 (N_2353,N_596,N_89);
or U2354 (N_2354,N_1244,N_1559);
nand U2355 (N_2355,N_1138,N_1365);
nor U2356 (N_2356,N_1527,In_1317);
nand U2357 (N_2357,N_102,In_3709);
nand U2358 (N_2358,N_1203,N_378);
and U2359 (N_2359,In_3067,N_1809);
and U2360 (N_2360,N_1081,N_245);
and U2361 (N_2361,N_1059,In_2306);
nand U2362 (N_2362,N_308,N_369);
or U2363 (N_2363,In_2381,N_141);
or U2364 (N_2364,In_1576,N_1852);
or U2365 (N_2365,In_1502,N_283);
nand U2366 (N_2366,In_209,N_1581);
or U2367 (N_2367,In_51,N_1162);
or U2368 (N_2368,N_1894,N_1339);
or U2369 (N_2369,In_330,In_4880);
or U2370 (N_2370,In_1165,N_672);
nand U2371 (N_2371,N_660,In_169);
or U2372 (N_2372,In_3897,In_2792);
and U2373 (N_2373,N_908,In_1251);
nor U2374 (N_2374,In_1001,In_798);
and U2375 (N_2375,In_1074,N_1341);
or U2376 (N_2376,N_1514,In_697);
and U2377 (N_2377,In_3987,N_1206);
nor U2378 (N_2378,In_275,N_1622);
nor U2379 (N_2379,N_750,In_4596);
and U2380 (N_2380,In_2742,N_644);
and U2381 (N_2381,N_1509,N_1840);
and U2382 (N_2382,N_968,N_1185);
nand U2383 (N_2383,N_1730,N_681);
nand U2384 (N_2384,N_1625,In_2931);
nand U2385 (N_2385,N_999,In_1051);
nor U2386 (N_2386,N_47,N_1993);
nor U2387 (N_2387,N_31,N_1614);
nand U2388 (N_2388,N_823,N_1223);
nor U2389 (N_2389,In_4358,N_1558);
nand U2390 (N_2390,In_2689,N_602);
and U2391 (N_2391,N_361,N_110);
nand U2392 (N_2392,N_1606,N_155);
nand U2393 (N_2393,In_2660,N_1324);
or U2394 (N_2394,In_3690,N_1836);
or U2395 (N_2395,In_1233,N_492);
and U2396 (N_2396,N_317,N_1278);
and U2397 (N_2397,N_989,In_3862);
or U2398 (N_2398,In_2686,In_3757);
nand U2399 (N_2399,In_2751,N_336);
or U2400 (N_2400,In_3190,N_1553);
or U2401 (N_2401,In_815,In_556);
nand U2402 (N_2402,N_1144,N_1153);
nor U2403 (N_2403,In_4089,In_4810);
nand U2404 (N_2404,N_1681,In_1062);
and U2405 (N_2405,N_1416,N_937);
and U2406 (N_2406,N_463,N_1725);
nor U2407 (N_2407,N_1283,N_729);
nand U2408 (N_2408,In_2654,In_2292);
or U2409 (N_2409,N_352,In_4755);
nand U2410 (N_2410,N_1868,N_1770);
or U2411 (N_2411,In_2417,N_28);
and U2412 (N_2412,N_792,In_1436);
and U2413 (N_2413,N_1947,In_4768);
or U2414 (N_2414,N_97,N_1630);
nand U2415 (N_2415,N_1008,N_109);
and U2416 (N_2416,In_3631,In_3195);
and U2417 (N_2417,In_2343,In_1491);
and U2418 (N_2418,N_49,In_341);
or U2419 (N_2419,N_1699,N_1975);
nand U2420 (N_2420,N_1368,N_14);
and U2421 (N_2421,In_98,N_59);
or U2422 (N_2422,N_1470,N_1541);
nand U2423 (N_2423,In_1474,N_1850);
nand U2424 (N_2424,N_889,In_517);
or U2425 (N_2425,N_598,N_1163);
nand U2426 (N_2426,N_331,N_470);
and U2427 (N_2427,In_1213,N_1526);
or U2428 (N_2428,N_694,N_1702);
and U2429 (N_2429,N_851,N_136);
and U2430 (N_2430,N_1351,N_1729);
and U2431 (N_2431,In_2484,N_1377);
nand U2432 (N_2432,N_1621,N_1767);
nor U2433 (N_2433,N_1049,In_1501);
nand U2434 (N_2434,In_289,N_652);
nand U2435 (N_2435,In_2402,N_1979);
nand U2436 (N_2436,N_1738,N_127);
nor U2437 (N_2437,In_3576,N_1133);
nor U2438 (N_2438,N_87,N_1516);
nand U2439 (N_2439,In_1926,N_1904);
nor U2440 (N_2440,N_425,In_4360);
nand U2441 (N_2441,N_125,N_1519);
and U2442 (N_2442,N_1387,N_287);
and U2443 (N_2443,N_609,In_978);
nor U2444 (N_2444,N_1590,N_257);
nor U2445 (N_2445,N_1718,In_2836);
nor U2446 (N_2446,N_1788,In_3018);
and U2447 (N_2447,N_1314,N_1330);
nand U2448 (N_2448,N_1480,In_4328);
and U2449 (N_2449,N_1799,N_1954);
and U2450 (N_2450,In_4006,In_4267);
or U2451 (N_2451,N_1873,In_400);
and U2452 (N_2452,N_1717,N_55);
nor U2453 (N_2453,N_1579,N_1240);
nor U2454 (N_2454,N_36,N_1680);
nor U2455 (N_2455,N_82,In_3771);
nand U2456 (N_2456,In_4276,N_1228);
nor U2457 (N_2457,N_905,In_4770);
or U2458 (N_2458,N_1298,N_1192);
or U2459 (N_2459,In_899,In_4063);
or U2460 (N_2460,N_1911,N_416);
and U2461 (N_2461,In_3739,N_20);
xnor U2462 (N_2462,N_557,N_1395);
nor U2463 (N_2463,In_2847,In_3419);
and U2464 (N_2464,N_1264,N_66);
or U2465 (N_2465,N_1286,N_1577);
and U2466 (N_2466,N_203,N_498);
nor U2467 (N_2467,In_1021,N_1849);
or U2468 (N_2468,N_1829,In_4964);
or U2469 (N_2469,N_773,N_1215);
and U2470 (N_2470,N_612,N_1334);
and U2471 (N_2471,N_39,N_455);
or U2472 (N_2472,N_576,N_1136);
nor U2473 (N_2473,In_1578,N_863);
and U2474 (N_2474,N_400,In_3652);
and U2475 (N_2475,N_1022,In_543);
and U2476 (N_2476,N_314,In_1678);
or U2477 (N_2477,N_1483,N_875);
nand U2478 (N_2478,N_1437,N_1560);
nor U2479 (N_2479,N_1841,In_1665);
nand U2480 (N_2480,N_676,N_1079);
nand U2481 (N_2481,N_855,In_1801);
or U2482 (N_2482,N_878,In_466);
or U2483 (N_2483,In_1724,N_1524);
nand U2484 (N_2484,In_900,N_472);
and U2485 (N_2485,In_2954,In_2735);
or U2486 (N_2486,N_1597,N_1791);
and U2487 (N_2487,In_4406,N_1279);
and U2488 (N_2488,In_4007,In_2841);
nor U2489 (N_2489,N_883,In_2766);
xnor U2490 (N_2490,In_2523,N_1983);
nand U2491 (N_2491,N_1373,N_218);
and U2492 (N_2492,N_1874,N_708);
nor U2493 (N_2493,In_287,In_3267);
nor U2494 (N_2494,N_807,N_12);
and U2495 (N_2495,N_263,N_1915);
nor U2496 (N_2496,N_841,In_4636);
nor U2497 (N_2497,N_195,In_4132);
and U2498 (N_2498,N_748,In_3099);
xor U2499 (N_2499,N_556,N_1036);
or U2500 (N_2500,N_914,N_838);
nor U2501 (N_2501,In_2892,N_1455);
or U2502 (N_2502,N_1807,N_874);
or U2503 (N_2503,In_1671,N_1356);
nand U2504 (N_2504,N_1707,N_1077);
nor U2505 (N_2505,N_1086,In_4193);
or U2506 (N_2506,N_625,N_244);
nor U2507 (N_2507,N_372,N_716);
or U2508 (N_2508,N_712,N_1657);
nor U2509 (N_2509,N_1160,In_3809);
or U2510 (N_2510,In_860,N_794);
nor U2511 (N_2511,N_280,N_1731);
and U2512 (N_2512,N_519,N_891);
nand U2513 (N_2513,N_713,N_1613);
or U2514 (N_2514,N_784,N_1090);
and U2515 (N_2515,N_1549,In_2875);
nor U2516 (N_2516,N_502,In_3287);
nand U2517 (N_2517,N_1406,N_422);
or U2518 (N_2518,In_1066,In_1629);
nand U2519 (N_2519,In_35,N_130);
nor U2520 (N_2520,N_769,N_1723);
or U2521 (N_2521,N_1123,N_1250);
xnor U2522 (N_2522,N_1020,N_956);
nand U2523 (N_2523,N_1119,In_1275);
and U2524 (N_2524,In_2156,In_2710);
or U2525 (N_2525,N_1636,N_622);
and U2526 (N_2526,N_251,N_934);
or U2527 (N_2527,N_827,N_415);
and U2528 (N_2528,In_1061,N_50);
and U2529 (N_2529,N_786,N_1111);
or U2530 (N_2530,N_516,N_1547);
or U2531 (N_2531,N_191,N_1960);
and U2532 (N_2532,N_467,N_477);
nand U2533 (N_2533,N_437,N_1069);
or U2534 (N_2534,N_1353,In_359);
and U2535 (N_2535,N_1335,In_2053);
or U2536 (N_2536,N_922,N_674);
nand U2537 (N_2537,N_79,N_199);
nand U2538 (N_2538,N_836,In_2250);
or U2539 (N_2539,In_4572,N_814);
nand U2540 (N_2540,N_1974,In_1248);
or U2541 (N_2541,In_4090,N_886);
and U2542 (N_2542,N_861,In_748);
nor U2543 (N_2543,N_202,In_3502);
nand U2544 (N_2544,N_1242,N_696);
nand U2545 (N_2545,In_496,In_2522);
nor U2546 (N_2546,N_726,N_1114);
nand U2547 (N_2547,N_689,In_4772);
xnor U2548 (N_2548,N_1520,N_1107);
nor U2549 (N_2549,N_246,N_1535);
or U2550 (N_2550,N_1624,In_528);
and U2551 (N_2551,N_1461,N_994);
and U2552 (N_2552,N_950,In_1494);
or U2553 (N_2553,N_1151,In_4927);
nor U2554 (N_2554,In_1447,In_4272);
nand U2555 (N_2555,N_1087,N_521);
or U2556 (N_2556,N_1177,N_206);
or U2557 (N_2557,N_1877,N_1027);
and U2558 (N_2558,N_527,N_1404);
and U2559 (N_2559,In_887,N_1085);
nor U2560 (N_2560,In_2753,In_4424);
or U2561 (N_2561,N_1235,In_777);
nand U2562 (N_2562,N_1010,N_1297);
or U2563 (N_2563,In_1572,N_307);
and U2564 (N_2564,In_4351,N_733);
nand U2565 (N_2565,N_1805,N_129);
nand U2566 (N_2566,N_1982,N_253);
nand U2567 (N_2567,In_4630,N_1226);
nor U2568 (N_2568,N_1967,In_4771);
nand U2569 (N_2569,In_3320,In_2337);
or U2570 (N_2570,N_393,In_3694);
nand U2571 (N_2571,In_3712,N_930);
or U2572 (N_2572,In_2262,N_166);
nand U2573 (N_2573,In_321,In_780);
and U2574 (N_2574,In_2400,In_3497);
and U2575 (N_2575,N_1804,In_2037);
nor U2576 (N_2576,N_1068,N_1779);
nand U2577 (N_2577,In_2810,In_3853);
nor U2578 (N_2578,N_998,N_1646);
nor U2579 (N_2579,N_1887,In_3466);
and U2580 (N_2580,In_536,N_227);
nand U2581 (N_2581,N_215,N_355);
nand U2582 (N_2582,N_1101,N_692);
nand U2583 (N_2583,N_1542,N_1361);
nor U2584 (N_2584,N_93,N_1656);
nor U2585 (N_2585,N_964,In_3300);
nor U2586 (N_2586,N_337,In_1019);
xor U2587 (N_2587,N_1871,N_162);
nand U2588 (N_2588,N_41,In_3698);
nand U2589 (N_2589,N_1844,N_211);
nand U2590 (N_2590,In_1327,N_176);
and U2591 (N_2591,N_816,In_1699);
nor U2592 (N_2592,In_4951,In_4072);
nand U2593 (N_2593,In_3779,In_1819);
and U2594 (N_2594,N_1793,N_761);
and U2595 (N_2595,N_907,N_1724);
and U2596 (N_2596,N_163,N_1977);
or U2597 (N_2597,In_2787,N_1456);
or U2598 (N_2598,In_2288,N_1783);
nand U2599 (N_2599,N_1821,N_1551);
nand U2600 (N_2600,N_145,In_1463);
nor U2601 (N_2601,In_626,In_214);
or U2602 (N_2602,N_159,N_1083);
nor U2603 (N_2603,In_1879,N_1129);
or U2604 (N_2604,In_15,N_410);
or U2605 (N_2605,N_703,N_1117);
nand U2606 (N_2606,N_1100,N_1832);
and U2607 (N_2607,N_1616,N_473);
and U2608 (N_2608,N_818,N_686);
nand U2609 (N_2609,In_4634,In_1498);
and U2610 (N_2610,N_1534,N_538);
and U2611 (N_2611,N_1370,In_4742);
nand U2612 (N_2612,N_1992,N_614);
nor U2613 (N_2613,N_482,N_583);
and U2614 (N_2614,N_1654,N_1764);
or U2615 (N_2615,N_392,N_5);
or U2616 (N_2616,N_411,N_688);
nor U2617 (N_2617,N_1578,In_1739);
or U2618 (N_2618,N_25,In_3728);
or U2619 (N_2619,N_603,N_375);
and U2620 (N_2620,N_484,N_1327);
nor U2621 (N_2621,N_1500,In_3400);
or U2622 (N_2622,N_15,N_1916);
nand U2623 (N_2623,In_2995,N_320);
or U2624 (N_2624,In_4289,N_1300);
and U2625 (N_2625,N_248,In_953);
and U2626 (N_2626,In_4301,N_305);
nor U2627 (N_2627,N_1391,In_3661);
and U2628 (N_2628,N_553,N_295);
and U2629 (N_2629,In_2988,In_830);
nand U2630 (N_2630,N_121,In_355);
nand U2631 (N_2631,N_7,N_408);
nor U2632 (N_2632,In_2669,In_3996);
nand U2633 (N_2633,N_1881,In_2676);
or U2634 (N_2634,N_75,In_2893);
nand U2635 (N_2635,N_1583,N_456);
nand U2636 (N_2636,N_900,N_1481);
and U2637 (N_2637,In_4207,N_315);
nand U2638 (N_2638,N_303,N_912);
or U2639 (N_2639,In_1136,N_406);
nand U2640 (N_2640,In_175,In_1675);
and U2641 (N_2641,N_1167,In_4034);
nand U2642 (N_2642,N_247,In_1469);
or U2643 (N_2643,In_1825,In_1130);
and U2644 (N_2644,N_1045,In_4511);
and U2645 (N_2645,N_1209,N_894);
xnor U2646 (N_2646,In_574,N_1428);
and U2647 (N_2647,In_4161,N_429);
or U2648 (N_2648,N_1828,N_1854);
nor U2649 (N_2649,N_1735,N_433);
nand U2650 (N_2650,N_212,In_4412);
nor U2651 (N_2651,N_1667,In_1548);
nand U2652 (N_2652,N_385,In_3323);
xnor U2653 (N_2653,N_194,N_1384);
nand U2654 (N_2654,N_441,N_1452);
or U2655 (N_2655,N_363,N_1092);
or U2656 (N_2656,N_483,N_359);
nand U2657 (N_2657,N_547,In_560);
and U2658 (N_2658,In_3482,N_201);
nor U2659 (N_2659,N_158,In_782);
or U2660 (N_2660,In_2795,N_34);
nor U2661 (N_2661,In_1403,N_1493);
or U2662 (N_2662,N_1390,N_1042);
or U2663 (N_2663,N_207,In_2603);
nand U2664 (N_2664,In_958,N_1028);
or U2665 (N_2665,N_960,In_304);
nand U2666 (N_2666,N_1399,N_183);
nand U2667 (N_2667,N_256,N_1072);
nand U2668 (N_2668,N_899,N_791);
xnor U2669 (N_2669,N_1818,N_1760);
nand U2670 (N_2670,N_1900,N_1610);
nand U2671 (N_2671,N_719,N_734);
or U2672 (N_2672,N_330,N_497);
or U2673 (N_2673,N_1972,N_399);
nand U2674 (N_2674,In_1250,N_1608);
nand U2675 (N_2675,In_2729,N_1462);
or U2676 (N_2676,N_1238,N_1678);
or U2677 (N_2677,N_839,N_865);
and U2678 (N_2678,N_71,N_438);
nand U2679 (N_2679,In_2268,In_4400);
xor U2680 (N_2680,In_2620,N_1987);
nand U2681 (N_2681,N_491,In_993);
nor U2682 (N_2682,N_177,N_322);
and U2683 (N_2683,N_254,N_446);
and U2684 (N_2684,N_546,N_1756);
or U2685 (N_2685,N_197,N_99);
nor U2686 (N_2686,In_3117,In_2260);
nand U2687 (N_2687,N_665,N_1895);
nor U2688 (N_2688,In_797,N_409);
and U2689 (N_2689,In_1018,N_1174);
nand U2690 (N_2690,N_1198,N_731);
or U2691 (N_2691,N_1747,N_1287);
nand U2692 (N_2692,In_893,N_1003);
nand U2693 (N_2693,N_927,N_847);
or U2694 (N_2694,N_1007,N_435);
nor U2695 (N_2695,In_1032,In_4743);
and U2696 (N_2696,N_1439,N_46);
nand U2697 (N_2697,N_581,In_301);
nand U2698 (N_2698,In_4520,In_4416);
or U2699 (N_2699,N_225,In_2883);
or U2700 (N_2700,N_1586,N_394);
and U2701 (N_2701,In_3427,N_299);
or U2702 (N_2702,N_1927,N_137);
nor U2703 (N_2703,In_4315,N_1145);
or U2704 (N_2704,N_1522,N_1870);
or U2705 (N_2705,N_1910,In_3253);
nor U2706 (N_2706,In_937,N_1973);
and U2707 (N_2707,In_2115,N_1454);
or U2708 (N_2708,N_1012,In_3542);
nor U2709 (N_2709,N_1357,N_854);
and U2710 (N_2710,N_1130,N_1787);
or U2711 (N_2711,In_3211,N_1943);
nand U2712 (N_2712,N_1216,N_1352);
xnor U2713 (N_2713,In_2509,N_1641);
nand U2714 (N_2714,N_844,N_1786);
nor U2715 (N_2715,N_1751,N_1485);
xor U2716 (N_2716,In_555,N_1701);
and U2717 (N_2717,In_4611,N_1421);
nand U2718 (N_2718,In_3544,N_382);
or U2719 (N_2719,N_572,N_1842);
nand U2720 (N_2720,N_1658,N_103);
xnor U2721 (N_2721,N_639,N_1988);
nand U2722 (N_2722,N_1694,N_62);
nand U2723 (N_2723,In_2586,N_656);
and U2724 (N_2724,N_1584,N_671);
xor U2725 (N_2725,In_2246,In_2021);
nor U2726 (N_2726,N_1710,N_1831);
xor U2727 (N_2727,N_635,N_1157);
and U2728 (N_2728,N_610,In_1873);
nand U2729 (N_2729,N_132,In_122);
nand U2730 (N_2730,N_604,N_1466);
nor U2731 (N_2731,In_3989,In_1607);
xor U2732 (N_2732,N_1499,N_1968);
and U2733 (N_2733,N_1367,N_1448);
and U2734 (N_2734,In_672,N_91);
nor U2735 (N_2735,In_3689,N_19);
or U2736 (N_2736,In_995,N_1210);
or U2737 (N_2737,N_1372,N_1213);
nand U2738 (N_2738,N_1502,In_914);
nor U2739 (N_2739,N_1147,N_374);
nand U2740 (N_2740,N_274,N_1963);
nand U2741 (N_2741,In_3883,N_728);
nand U2742 (N_2742,N_1231,N_842);
nor U2743 (N_2743,N_1503,N_1030);
nand U2744 (N_2744,N_591,In_3855);
nand U2745 (N_2745,In_1336,N_1108);
nand U2746 (N_2746,N_1342,In_3068);
nand U2747 (N_2747,In_3171,In_3858);
nand U2748 (N_2748,N_328,N_825);
nor U2749 (N_2749,In_1267,N_1632);
nand U2750 (N_2750,N_1392,N_292);
or U2751 (N_2751,N_267,N_1679);
and U2752 (N_2752,N_584,In_1522);
or U2753 (N_2753,N_1477,N_266);
and U2754 (N_2754,In_4519,In_1391);
or U2755 (N_2755,N_1504,In_1529);
nor U2756 (N_2756,N_262,N_923);
or U2757 (N_2757,In_4010,N_397);
nor U2758 (N_2758,N_224,N_362);
nand U2759 (N_2759,In_3454,N_111);
or U2760 (N_2760,N_1969,N_364);
or U2761 (N_2761,N_1057,N_608);
and U2762 (N_2762,In_3569,In_3407);
nor U2763 (N_2763,N_637,In_265);
or U2764 (N_2764,N_38,In_736);
nand U2765 (N_2765,N_285,In_4481);
nand U2766 (N_2766,N_1971,In_2771);
xor U2767 (N_2767,In_1533,In_2709);
xor U2768 (N_2768,In_880,In_281);
nor U2769 (N_2769,In_1803,In_366);
nor U2770 (N_2770,In_2129,N_1);
and U2771 (N_2771,N_518,N_893);
or U2772 (N_2772,In_1528,N_539);
and U2773 (N_2773,N_1321,N_1095);
and U2774 (N_2774,N_701,In_1119);
xor U2775 (N_2775,N_168,In_3064);
nand U2776 (N_2776,N_386,N_977);
xor U2777 (N_2777,N_290,N_885);
nor U2778 (N_2778,In_1886,In_4904);
and U2779 (N_2779,N_1294,N_1415);
or U2780 (N_2780,N_368,In_3215);
nor U2781 (N_2781,N_880,In_838);
or U2782 (N_2782,N_1175,In_3792);
or U2783 (N_2783,N_1267,N_1071);
or U2784 (N_2784,N_1907,N_1595);
or U2785 (N_2785,N_510,N_944);
nand U2786 (N_2786,In_382,In_2032);
nand U2787 (N_2787,N_487,N_388);
nand U2788 (N_2788,N_323,N_720);
or U2789 (N_2789,N_68,N_142);
nor U2790 (N_2790,N_846,N_1272);
nand U2791 (N_2791,N_1815,N_1271);
nor U2792 (N_2792,N_1257,N_740);
nor U2793 (N_2793,N_1538,N_1869);
or U2794 (N_2794,N_350,In_731);
and U2795 (N_2795,N_1444,N_297);
nor U2796 (N_2796,N_17,N_1056);
and U2797 (N_2797,In_2044,N_1249);
or U2798 (N_2798,In_3233,N_687);
and U2799 (N_2799,N_106,In_2781);
nor U2800 (N_2800,N_1016,N_182);
and U2801 (N_2801,N_585,N_705);
and U2802 (N_2802,N_682,In_3382);
or U2803 (N_2803,N_1795,N_457);
or U2804 (N_2804,N_1867,N_1490);
and U2805 (N_2805,In_2444,N_1886);
nand U2806 (N_2806,N_187,In_2835);
or U2807 (N_2807,In_3611,In_3976);
nand U2808 (N_2808,N_114,N_848);
nand U2809 (N_2809,N_931,N_1891);
nor U2810 (N_2810,N_42,N_804);
xnor U2811 (N_2811,N_1190,N_718);
or U2812 (N_2812,In_3654,N_1229);
or U2813 (N_2813,N_961,N_529);
nand U2814 (N_2814,In_1556,In_3442);
or U2815 (N_2815,In_1975,N_108);
and U2816 (N_2816,In_2311,N_1385);
and U2817 (N_2817,N_296,In_2990);
or U2818 (N_2818,In_85,N_1643);
nand U2819 (N_2819,N_48,In_3759);
or U2820 (N_2820,In_4240,In_592);
and U2821 (N_2821,N_1440,In_1148);
nand U2822 (N_2822,N_963,N_697);
nand U2823 (N_2823,N_1941,In_2854);
nand U2824 (N_2824,In_2734,In_3076);
or U2825 (N_2825,In_312,N_69);
and U2826 (N_2826,N_1964,N_222);
nor U2827 (N_2827,In_1214,In_105);
and U2828 (N_2828,N_1402,N_464);
nor U2829 (N_2829,N_462,N_1055);
and U2830 (N_2830,N_935,N_1757);
or U2831 (N_2831,N_571,N_1562);
nor U2832 (N_2832,N_868,In_1564);
or U2833 (N_2833,N_1851,N_1587);
nor U2834 (N_2834,N_1225,N_509);
xor U2835 (N_2835,N_1000,In_4940);
nand U2836 (N_2836,In_538,N_1442);
nand U2837 (N_2837,N_1096,In_2471);
nand U2838 (N_2838,N_984,N_1343);
nor U2839 (N_2839,N_978,N_860);
nand U2840 (N_2840,In_2984,N_465);
nand U2841 (N_2841,In_4306,N_339);
nand U2842 (N_2842,N_252,N_119);
or U2843 (N_2843,In_1493,In_129);
or U2844 (N_2844,N_1768,In_2864);
nor U2845 (N_2845,N_448,N_1843);
nor U2846 (N_2846,N_1634,N_193);
or U2847 (N_2847,N_550,In_4186);
nand U2848 (N_2848,N_376,In_2184);
or U2849 (N_2849,N_1478,N_16);
and U2850 (N_2850,In_3157,In_3498);
and U2851 (N_2851,In_2285,N_675);
nand U2852 (N_2852,N_1690,N_1810);
and U2853 (N_2853,N_647,In_651);
nor U2854 (N_2854,In_3983,N_887);
nand U2855 (N_2855,N_1159,N_623);
nor U2856 (N_2856,In_611,N_1714);
nand U2857 (N_2857,N_1034,N_541);
nor U2858 (N_2858,N_663,N_837);
or U2859 (N_2859,N_1410,N_630);
nand U2860 (N_2860,N_520,N_300);
and U2861 (N_2861,N_475,In_242);
or U2862 (N_2862,N_1626,N_1884);
nor U2863 (N_2863,N_1839,N_1425);
and U2864 (N_2864,N_1726,N_903);
and U2865 (N_2865,N_812,N_815);
or U2866 (N_2866,In_68,In_4028);
or U2867 (N_2867,N_532,In_1306);
nand U2868 (N_2868,In_3337,N_242);
nor U2869 (N_2869,N_1918,In_2740);
or U2870 (N_2870,N_58,N_133);
nand U2871 (N_2871,In_3441,N_454);
nor U2872 (N_2872,In_2911,In_3986);
nand U2873 (N_2873,In_3532,N_217);
or U2874 (N_2874,N_1258,In_4974);
and U2875 (N_2875,N_1251,N_334);
or U2876 (N_2876,In_4868,N_329);
or U2877 (N_2877,N_1855,N_1991);
nor U2878 (N_2878,N_1812,N_351);
and U2879 (N_2879,N_471,In_295);
nand U2880 (N_2880,N_420,N_1938);
and U2881 (N_2881,In_1894,N_869);
or U2882 (N_2882,In_3903,In_393);
or U2883 (N_2883,N_648,N_566);
and U2884 (N_2884,N_523,N_113);
and U2885 (N_2885,N_924,N_272);
nor U2886 (N_2886,In_4912,N_1109);
nor U2887 (N_2887,In_4308,In_2203);
nor U2888 (N_2888,N_70,In_2881);
and U2889 (N_2889,N_770,N_824);
nor U2890 (N_2890,N_431,In_3218);
and U2891 (N_2891,In_2338,N_752);
xor U2892 (N_2892,In_1715,In_4623);
nand U2893 (N_2893,In_2638,N_1824);
or U2894 (N_2894,In_39,N_1496);
nor U2895 (N_2895,In_4466,In_4136);
and U2896 (N_2896,N_1708,N_1771);
and U2897 (N_2897,N_434,In_3198);
or U2898 (N_2898,In_679,In_4637);
nor U2899 (N_2899,In_3831,In_3017);
nand U2900 (N_2900,In_1765,N_1222);
or U2901 (N_2901,N_1976,N_324);
nor U2902 (N_2902,In_3265,N_1227);
nor U2903 (N_2903,N_1239,N_1255);
and U2904 (N_2904,N_901,N_1961);
and U2905 (N_2905,In_4802,N_1733);
nor U2906 (N_2906,N_1642,N_624);
or U2907 (N_2907,N_754,N_747);
nand U2908 (N_2908,N_1946,In_3423);
or U2909 (N_2909,In_1145,In_2529);
nor U2910 (N_2910,In_106,N_549);
and U2911 (N_2911,In_4747,In_889);
or U2912 (N_2912,In_1628,N_64);
nor U2913 (N_2913,N_1329,N_1722);
nor U2914 (N_2914,In_2276,N_273);
nor U2915 (N_2915,N_241,N_365);
nand U2916 (N_2916,N_617,N_840);
or U2917 (N_2917,In_1924,N_1552);
and U2918 (N_2918,N_1965,In_4838);
nor U2919 (N_2919,N_511,N_1669);
or U2920 (N_2920,N_1326,N_1067);
nand U2921 (N_2921,In_3554,N_636);
nor U2922 (N_2922,N_1363,In_2166);
or U2923 (N_2923,N_629,N_348);
nor U2924 (N_2924,In_3181,N_1665);
nor U2925 (N_2925,In_1348,In_1608);
nand U2926 (N_2926,N_1940,N_668);
nor U2927 (N_2927,N_1124,N_1214);
nand U2928 (N_2928,N_781,N_1755);
and U2929 (N_2929,N_40,In_4503);
and U2930 (N_2930,N_544,In_1099);
and U2931 (N_2931,N_1648,In_713);
or U2932 (N_2932,In_4690,N_1645);
or U2933 (N_2933,N_833,N_1555);
or U2934 (N_2934,In_4736,N_1037);
and U2935 (N_2935,N_1746,N_1959);
nand U2936 (N_2936,N_1396,N_683);
or U2937 (N_2937,In_2658,N_221);
nand U2938 (N_2938,N_1044,In_1874);
nand U2939 (N_2939,N_104,N_988);
and U2940 (N_2940,N_990,N_1909);
nand U2941 (N_2941,In_1713,N_236);
nor U2942 (N_2942,In_1124,N_957);
or U2943 (N_2943,In_3094,N_1521);
nor U2944 (N_2944,In_2648,N_1588);
nor U2945 (N_2945,N_338,N_1449);
and U2946 (N_2946,N_1618,In_883);
nand U2947 (N_2947,N_401,In_264);
and U2948 (N_2948,N_700,N_867);
nor U2949 (N_2949,N_149,N_810);
and U2950 (N_2950,N_92,N_570);
xnor U2951 (N_2951,In_3575,N_1806);
and U2952 (N_2952,N_1827,N_876);
nor U2953 (N_2953,In_2432,N_1047);
or U2954 (N_2954,N_51,N_1061);
and U2955 (N_2955,N_1403,In_323);
or U2956 (N_2956,In_682,N_1393);
nor U2957 (N_2957,N_1696,N_478);
nor U2958 (N_2958,N_1132,N_1501);
nand U2959 (N_2959,In_4614,N_1713);
or U2960 (N_2960,In_2214,N_1939);
nor U2961 (N_2961,N_495,N_319);
or U2962 (N_2962,N_936,In_4977);
or U2963 (N_2963,N_98,N_642);
xor U2964 (N_2964,N_1233,N_188);
nor U2965 (N_2965,N_948,N_381);
xor U2966 (N_2966,In_2034,N_809);
or U2967 (N_2967,In_2846,N_779);
nand U2968 (N_2968,N_403,In_219);
nor U2969 (N_2969,N_1319,N_1782);
xnor U2970 (N_2970,N_762,N_1019);
and U2971 (N_2971,N_1205,N_271);
nand U2972 (N_2972,In_4837,In_2541);
nand U2973 (N_2973,N_890,In_1892);
nand U2974 (N_2974,N_450,N_86);
or U2975 (N_2975,N_562,In_3066);
nand U2976 (N_2976,In_4597,In_2060);
xor U2977 (N_2977,N_1301,N_1460);
nor U2978 (N_2978,N_1482,N_249);
nor U2979 (N_2979,N_803,N_220);
nand U2980 (N_2980,In_2383,In_3875);
nor U2981 (N_2981,N_1021,In_3358);
and U2982 (N_2982,N_1880,N_1122);
or U2983 (N_2983,N_561,N_1801);
or U2984 (N_2984,N_1739,In_1188);
or U2985 (N_2985,N_1039,N_653);
or U2986 (N_2986,In_6,N_1593);
nor U2987 (N_2987,N_164,N_925);
and U2988 (N_2988,N_1344,N_1712);
nor U2989 (N_2989,In_4234,N_277);
nor U2990 (N_2990,N_669,N_289);
nand U2991 (N_2991,N_1345,In_2736);
nand U2992 (N_2992,N_1043,In_1420);
nand U2993 (N_2993,N_895,N_1990);
or U2994 (N_2994,N_235,In_4877);
and U2995 (N_2995,In_1686,In_3840);
or U2996 (N_2996,In_4469,In_1277);
or U2997 (N_2997,In_7,N_1137);
nand U2998 (N_2998,N_342,In_1708);
nand U2999 (N_2999,N_1364,In_244);
or U3000 (N_3000,N_120,In_4664);
nand U3001 (N_3001,N_1013,In_3261);
and U3002 (N_3002,N_970,N_126);
nand U3003 (N_3003,N_551,N_496);
nor U3004 (N_3004,In_1361,N_1650);
nand U3005 (N_3005,N_1033,In_234);
nand U3006 (N_3006,N_1528,N_1389);
nand U3007 (N_3007,In_1012,N_449);
and U3008 (N_3008,N_165,In_4502);
or U3009 (N_3009,In_3665,N_1017);
xor U3010 (N_3010,N_1199,In_4441);
and U3011 (N_3011,In_1319,In_1156);
nor U3012 (N_3012,N_1094,N_480);
or U3013 (N_3013,In_439,N_1349);
nor U3014 (N_3014,N_156,N_1284);
and U3015 (N_3015,N_1193,N_1113);
nor U3016 (N_3016,N_107,N_304);
nand U3017 (N_3017,N_780,N_1546);
xnor U3018 (N_3018,In_2164,N_1929);
nand U3019 (N_3019,In_1110,In_2959);
and U3020 (N_3020,N_830,In_4491);
or U3021 (N_3021,N_1261,N_1310);
nor U3022 (N_3022,In_4846,N_1299);
and U3023 (N_3023,In_4525,N_777);
or U3024 (N_3024,N_1293,In_4920);
or U3025 (N_3025,In_1507,N_1935);
nand U3026 (N_3026,N_834,N_1371);
and U3027 (N_3027,N_1230,N_537);
nor U3028 (N_3028,In_2313,N_360);
nand U3029 (N_3029,In_2814,N_606);
nand U3030 (N_3030,N_1281,N_1996);
nor U3031 (N_3031,N_1752,N_1570);
or U3032 (N_3032,In_3311,In_4956);
nor U3033 (N_3033,N_1436,N_1569);
nor U3034 (N_3034,In_1315,In_3330);
or U3035 (N_3035,In_3150,In_1402);
or U3036 (N_3036,N_1429,N_288);
or U3037 (N_3037,N_1510,N_1196);
and U3038 (N_3038,N_1903,N_1316);
nor U3039 (N_3039,In_1517,N_1346);
nor U3040 (N_3040,N_888,In_1626);
xnor U3041 (N_3041,N_83,In_1082);
nor U3042 (N_3042,In_881,N_1716);
or U3043 (N_3043,N_1378,N_404);
nor U3044 (N_3044,In_2517,N_1923);
or U3045 (N_3045,N_76,N_1476);
xor U3046 (N_3046,In_3266,In_3741);
nor U3047 (N_3047,In_2861,In_2253);
nand U3048 (N_3048,In_2519,In_2685);
xor U3049 (N_3049,N_1928,N_1628);
and U3050 (N_3050,N_505,N_962);
or U3051 (N_3051,N_1104,N_1889);
and U3052 (N_3052,N_1835,In_600);
nor U3053 (N_3053,N_1400,In_3696);
and U3054 (N_3054,N_1201,N_1655);
or U3055 (N_3055,In_3624,In_2199);
or U3056 (N_3056,In_813,N_1058);
nor U3057 (N_3057,N_829,In_2594);
nand U3058 (N_3058,N_1009,In_3890);
and U3059 (N_3059,In_3440,N_229);
or U3060 (N_3060,N_6,N_1181);
nor U3061 (N_3061,In_3403,N_1930);
or U3062 (N_3062,N_357,N_1002);
or U3063 (N_3063,N_1266,In_4440);
or U3064 (N_3064,N_946,N_1592);
and U3065 (N_3065,N_534,In_2774);
nand U3066 (N_3066,In_3836,In_2466);
or U3067 (N_3067,In_4762,In_212);
xor U3068 (N_3068,In_3123,In_356);
nand U3069 (N_3069,N_789,N_736);
and U3070 (N_3070,N_1677,N_1611);
and U3071 (N_3071,N_1620,In_4701);
and U3072 (N_3072,In_1489,N_513);
or U3073 (N_3073,N_421,In_1561);
or U3074 (N_3074,In_3236,N_18);
and U3075 (N_3075,N_1398,N_1035);
nand U3076 (N_3076,In_2370,N_1253);
nor U3077 (N_3077,N_552,N_1848);
nand U3078 (N_3078,N_306,N_662);
nor U3079 (N_3079,In_1387,N_1273);
or U3080 (N_3080,In_909,N_906);
xor U3081 (N_3081,N_214,N_243);
or U3082 (N_3082,In_3475,In_483);
or U3083 (N_3083,N_1409,N_1761);
and U3084 (N_3084,N_367,N_427);
nor U3085 (N_3085,N_1603,N_1957);
and U3086 (N_3086,N_1817,N_1663);
nor U3087 (N_3087,N_143,In_1044);
nor U3088 (N_3088,In_1747,N_1778);
or U3089 (N_3089,N_1311,N_458);
nand U3090 (N_3090,N_1475,N_1268);
and U3091 (N_3091,In_343,In_523);
and U3092 (N_3092,In_460,In_625);
nor U3093 (N_3093,N_628,In_309);
and U3094 (N_3094,In_2938,N_522);
nor U3095 (N_3095,In_435,N_1766);
and U3096 (N_3096,In_4167,N_651);
and U3097 (N_3097,In_2065,N_710);
and U3098 (N_3098,N_698,N_1803);
and U3099 (N_3099,N_1438,N_459);
nand U3100 (N_3100,N_1052,N_757);
or U3101 (N_3101,In_2770,N_1188);
nand U3102 (N_3102,N_1897,N_1539);
and U3103 (N_3103,In_2982,In_1194);
and U3104 (N_3104,In_1142,N_88);
nor U3105 (N_3105,In_4905,In_2353);
and U3106 (N_3106,N_268,N_44);
or U3107 (N_3107,In_1278,In_795);
nand U3108 (N_3108,In_4669,N_722);
nor U3109 (N_3109,N_1781,N_543);
nor U3110 (N_3110,N_32,In_116);
and U3111 (N_3111,N_650,N_1492);
or U3112 (N_3112,N_1128,N_1463);
or U3113 (N_3113,In_904,N_232);
nor U3114 (N_3114,In_4298,N_1859);
nand U3115 (N_3115,N_1572,N_1536);
nor U3116 (N_3116,In_2917,N_1945);
or U3117 (N_3117,In_2150,N_1277);
and U3118 (N_3118,N_1604,N_1484);
nand U3119 (N_3119,In_4842,N_640);
nor U3120 (N_3120,N_1728,N_605);
and U3121 (N_3121,N_1374,N_670);
or U3122 (N_3122,N_1978,N_1863);
nand U3123 (N_3123,N_1687,N_1784);
or U3124 (N_3124,In_2656,N_1024);
and U3125 (N_3125,N_160,N_344);
and U3126 (N_3126,In_1896,N_1340);
nor U3127 (N_3127,In_2208,In_4624);
nand U3128 (N_3128,N_405,N_1639);
nor U3129 (N_3129,N_1246,N_666);
and U3130 (N_3130,N_146,N_1312);
nand U3131 (N_3131,N_1380,In_4703);
nand U3132 (N_3132,N_758,N_29);
nor U3133 (N_3133,In_4585,N_154);
and U3134 (N_3134,In_4245,In_3834);
or U3135 (N_3135,In_1105,N_22);
nor U3136 (N_3136,N_426,In_199);
nand U3137 (N_3137,N_1912,N_1014);
nor U3138 (N_3138,N_1879,N_597);
or U3139 (N_3139,N_661,In_3385);
and U3140 (N_3140,N_1898,In_316);
or U3141 (N_3141,N_209,N_735);
nor U3142 (N_3142,N_1635,N_864);
and U3143 (N_3143,N_1450,N_237);
nand U3144 (N_3144,N_1507,N_1369);
nor U3145 (N_3145,N_593,In_1035);
nand U3146 (N_3146,In_3478,In_3363);
and U3147 (N_3147,In_2135,N_298);
or U3148 (N_3148,N_444,N_10);
and U3149 (N_3149,N_808,In_2388);
or U3150 (N_3150,N_1489,N_1208);
or U3151 (N_3151,In_4613,N_1800);
nand U3152 (N_3152,In_1655,N_975);
xnor U3153 (N_3153,In_3113,In_2538);
or U3154 (N_3154,N_1700,N_259);
nand U3155 (N_3155,In_4395,N_996);
or U3156 (N_3156,N_706,N_1732);
and U3157 (N_3157,N_341,N_1120);
nor U3158 (N_3158,In_4729,In_965);
and U3159 (N_3159,N_600,N_1913);
and U3160 (N_3160,N_1777,N_616);
or U3161 (N_3161,In_714,In_254);
nor U3162 (N_3162,N_730,In_4394);
nand U3163 (N_3163,N_717,In_4514);
nor U3164 (N_3164,N_1254,N_759);
nand U3165 (N_3165,In_3016,N_461);
and U3166 (N_3166,In_1980,In_4279);
xnor U3167 (N_3167,N_1270,N_138);
and U3168 (N_3168,N_690,N_1548);
xnor U3169 (N_3169,N_30,N_940);
and U3170 (N_3170,In_3952,N_1427);
or U3171 (N_3171,N_1962,In_1921);
nor U3172 (N_3172,N_1953,In_634);
and U3173 (N_3173,N_1948,N_1866);
and U3174 (N_3174,N_1564,N_1139);
nand U3175 (N_3175,N_490,N_1248);
nand U3176 (N_3176,N_1303,N_819);
and U3177 (N_3177,N_745,In_1917);
nand U3178 (N_3178,In_1833,In_379);
or U3179 (N_3179,In_4626,N_122);
and U3180 (N_3180,N_1143,In_607);
or U3181 (N_3181,In_1992,N_1443);
and U3182 (N_3182,N_1219,N_691);
nand U3183 (N_3183,N_326,N_1189);
or U3184 (N_3184,In_750,In_55);
and U3185 (N_3185,N_778,N_1921);
and U3186 (N_3186,N_153,In_3140);
and U3187 (N_3187,N_190,In_728);
or U3188 (N_3188,N_1142,N_52);
and U3189 (N_3189,N_1709,N_1220);
nand U3190 (N_3190,N_1323,In_4934);
or U3191 (N_3191,N_282,In_577);
nand U3192 (N_3192,N_419,N_1015);
or U3193 (N_3193,N_1823,In_839);
nand U3194 (N_3194,N_1743,N_737);
and U3195 (N_3195,N_685,In_4540);
nand U3196 (N_3196,In_204,N_178);
nand U3197 (N_3197,N_1933,In_2922);
or U3198 (N_3198,N_898,N_1062);
and U3199 (N_3199,N_321,N_772);
and U3200 (N_3200,N_972,N_1118);
and U3201 (N_3201,N_1651,N_1838);
nor U3202 (N_3202,N_852,In_4554);
and U3203 (N_3203,N_1691,N_620);
and U3204 (N_3204,N_81,In_3894);
xor U3205 (N_3205,N_1091,N_958);
nand U3206 (N_3206,N_223,In_4390);
nor U3207 (N_3207,In_3036,In_2478);
and U3208 (N_3208,N_751,N_1048);
and U3209 (N_3209,N_1704,N_312);
xor U3210 (N_3210,In_47,In_4756);
nor U3211 (N_3211,N_1413,N_721);
nor U3212 (N_3212,N_1259,N_1862);
and U3213 (N_3213,N_1465,N_1105);
nand U3214 (N_3214,N_1670,N_764);
nand U3215 (N_3215,N_1937,N_1601);
nor U3216 (N_3216,N_301,In_1993);
or U3217 (N_3217,N_73,N_1376);
nand U3218 (N_3218,In_2227,In_2765);
nand U3219 (N_3219,In_1339,N_902);
nand U3220 (N_3220,N_269,N_882);
or U3221 (N_3221,N_548,N_1822);
xor U3222 (N_3222,In_608,N_466);
and U3223 (N_3223,In_1618,N_909);
nand U3224 (N_3224,N_1247,In_2858);
nand U3225 (N_3225,N_1518,N_715);
or U3226 (N_3226,N_1830,In_2505);
or U3227 (N_3227,In_3041,N_1980);
nand U3228 (N_3228,In_431,In_1518);
and U3229 (N_3229,N_343,N_1653);
and U3230 (N_3230,In_2366,In_3276);
nor U3231 (N_3231,N_1121,N_560);
nor U3232 (N_3232,N_945,N_1084);
or U3233 (N_3233,N_817,N_575);
nor U3234 (N_3234,In_1632,In_436);
nor U3235 (N_3235,N_345,In_1039);
nand U3236 (N_3236,N_1846,N_1845);
or U3237 (N_3237,N_1675,N_1445);
or U3238 (N_3238,N_1412,N_634);
nor U3239 (N_3239,N_1816,N_1318);
nor U3240 (N_3240,N_140,In_874);
nand U3241 (N_3241,N_677,In_1784);
and U3242 (N_3242,In_4071,N_23);
nor U3243 (N_3243,N_1362,In_3763);
nand U3244 (N_3244,N_152,N_856);
nor U3245 (N_3245,N_967,N_200);
nand U3246 (N_3246,N_1023,In_191);
nand U3247 (N_3247,N_1833,N_1776);
xor U3248 (N_3248,In_370,N_1156);
nor U3249 (N_3249,N_530,In_2442);
or U3250 (N_3250,N_588,In_3275);
nand U3251 (N_3251,In_2963,In_300);
xor U3252 (N_3252,In_1379,In_3615);
or U3253 (N_3253,N_216,N_279);
and U3254 (N_3254,N_123,N_1204);
nor U3255 (N_3255,N_918,N_116);
or U3256 (N_3256,N_798,N_1066);
or U3257 (N_3257,N_1652,N_1355);
xnor U3258 (N_3258,N_84,N_982);
or U3259 (N_3259,In_3001,N_1032);
nand U3260 (N_3260,N_1322,N_1672);
or U3261 (N_3261,N_417,N_501);
nor U3262 (N_3262,In_337,In_197);
or U3263 (N_3263,N_695,N_1295);
or U3264 (N_3264,N_767,N_489);
or U3265 (N_3265,N_1183,N_1925);
nor U3266 (N_3266,N_1431,N_1252);
nor U3267 (N_3267,N_1703,N_198);
nand U3268 (N_3268,N_1408,N_1917);
or U3269 (N_3269,N_1922,In_1942);
nor U3270 (N_3270,In_3464,In_4546);
nor U3271 (N_3271,In_3467,In_2830);
nor U3272 (N_3272,N_174,N_447);
and U3273 (N_3273,In_2297,N_1296);
nor U3274 (N_3274,N_1896,N_169);
and U3275 (N_3275,In_3347,In_1555);
xnor U3276 (N_3276,In_800,N_1063);
xnor U3277 (N_3277,In_825,In_4726);
and U3278 (N_3278,N_1332,In_420);
nor U3279 (N_3279,In_26,In_1832);
nor U3280 (N_3280,In_1824,In_278);
nor U3281 (N_3281,In_4565,N_590);
and U3282 (N_3282,N_1394,N_1906);
or U3283 (N_3283,N_1232,N_507);
or U3284 (N_3284,In_4870,N_3);
and U3285 (N_3285,N_1631,N_340);
nand U3286 (N_3286,N_732,N_1041);
and U3287 (N_3287,N_255,N_1575);
and U3288 (N_3288,N_1165,In_2646);
and U3289 (N_3289,In_1683,In_4130);
nor U3290 (N_3290,N_1184,N_607);
xor U3291 (N_3291,N_771,In_1945);
xor U3292 (N_3292,N_11,N_1574);
or U3293 (N_3293,N_1813,In_31);
nand U3294 (N_3294,In_2418,N_1902);
and U3295 (N_3295,N_755,N_1172);
nor U3296 (N_3296,N_849,N_1025);
nor U3297 (N_3297,N_1134,N_776);
nor U3298 (N_3298,N_1932,In_1265);
nand U3299 (N_3299,N_57,N_383);
nor U3300 (N_3300,N_1150,In_3695);
and U3301 (N_3301,In_1367,N_1505);
nand U3302 (N_3302,N_739,N_1666);
nand U3303 (N_3303,In_2107,N_1256);
or U3304 (N_3304,In_4335,N_1360);
and U3305 (N_3305,N_167,N_1567);
nand U3306 (N_3306,N_1582,In_3793);
nand U3307 (N_3307,N_1772,N_398);
nor U3308 (N_3308,N_291,In_236);
and U3309 (N_3309,N_428,N_586);
or U3310 (N_3310,In_4524,N_506);
nand U3311 (N_3311,In_3185,In_1155);
and U3312 (N_3312,In_2303,N_293);
or U3313 (N_3313,N_1197,In_4333);
nor U3314 (N_3314,In_3641,N_916);
and U3315 (N_3315,N_1423,N_1263);
nand U3316 (N_3316,N_135,In_2494);
nor U3317 (N_3317,N_418,N_453);
or U3318 (N_3318,N_646,N_979);
nand U3319 (N_3319,N_921,N_753);
and U3320 (N_3320,N_281,N_78);
nand U3321 (N_3321,N_1414,N_1512);
nand U3322 (N_3322,N_1513,In_2104);
nor U3323 (N_3323,N_1808,N_1934);
nand U3324 (N_3324,N_1388,In_2547);
and U3325 (N_3325,In_935,In_4593);
nand U3326 (N_3326,In_1851,In_2035);
nand U3327 (N_3327,N_631,N_741);
and U3328 (N_3328,N_1711,In_3012);
nand U3329 (N_3329,N_1245,In_616);
and U3330 (N_3330,In_3835,N_309);
and U3331 (N_3331,N_567,In_3750);
and U3332 (N_3332,N_1289,N_589);
nand U3333 (N_3333,N_568,In_2682);
or U3334 (N_3334,N_1994,In_868);
nor U3335 (N_3335,N_1637,N_822);
nand U3336 (N_3336,N_407,In_2763);
or U3337 (N_3337,N_1291,In_3540);
nor U3338 (N_3338,N_800,N_476);
nand U3339 (N_3339,N_881,In_3167);
and U3340 (N_3340,N_877,N_1986);
and U3341 (N_3341,N_1446,N_27);
and U3342 (N_3342,N_1568,In_1020);
nor U3343 (N_3343,In_771,N_1350);
or U3344 (N_3344,N_1837,N_1697);
or U3345 (N_3345,N_1011,In_4529);
and U3346 (N_3346,N_1288,In_3084);
nand U3347 (N_3347,N_1565,N_845);
nor U3348 (N_3348,N_1308,N_1689);
and U3349 (N_3349,In_3247,N_284);
nor U3350 (N_3350,N_1950,N_1269);
nor U3351 (N_3351,N_1088,N_1955);
or U3352 (N_3352,N_673,In_1599);
and U3353 (N_3353,In_326,N_1682);
or U3354 (N_3354,N_953,N_932);
nor U3355 (N_3355,N_1640,N_1706);
nand U3356 (N_3356,In_501,In_2344);
nor U3357 (N_3357,N_1051,In_632);
nor U3358 (N_3358,N_678,N_1479);
or U3359 (N_3359,N_1331,N_1748);
and U3360 (N_3360,N_580,In_762);
and U3361 (N_3361,In_4579,In_4477);
or U3362 (N_3362,In_4331,N_831);
or U3363 (N_3363,In_2657,In_1709);
nand U3364 (N_3364,In_3304,N_765);
or U3365 (N_3365,N_1495,In_377);
nor U3366 (N_3366,N_1566,N_1741);
or U3367 (N_3367,N_594,N_1596);
nor U3368 (N_3368,In_2577,In_494);
and U3369 (N_3369,In_4244,In_1588);
xor U3370 (N_3370,N_414,N_1276);
nand U3371 (N_3371,N_460,In_3915);
or U3372 (N_3372,In_768,N_1627);
and U3373 (N_3373,N_1211,N_1794);
and U3374 (N_3374,N_35,N_756);
and U3375 (N_3375,N_226,N_1515);
or U3376 (N_3376,N_787,N_499);
nand U3377 (N_3377,In_4710,In_2398);
and U3378 (N_3378,In_3568,N_966);
nor U3379 (N_3379,N_105,In_628);
nand U3380 (N_3380,N_599,N_615);
nor U3381 (N_3381,N_1647,In_991);
and U3382 (N_3382,N_535,In_1863);
nand U3383 (N_3383,N_884,In_2089);
nand U3384 (N_3384,In_1382,N_1182);
or U3385 (N_3385,N_54,N_1333);
xor U3386 (N_3386,N_1006,In_3144);
nand U3387 (N_3387,N_559,N_857);
and U3388 (N_3388,In_3133,N_627);
nor U3389 (N_3389,In_3507,N_1383);
or U3390 (N_3390,N_1556,N_892);
and U3391 (N_3391,In_936,N_554);
nand U3392 (N_3392,In_2897,In_2870);
and U3393 (N_3393,In_2174,N_1773);
nand U3394 (N_3394,N_13,In_79);
and U3395 (N_3395,N_1580,N_1531);
or U3396 (N_3396,N_910,In_3856);
xnor U3397 (N_3397,N_1920,N_1763);
nor U3398 (N_3398,N_1721,N_440);
nor U3399 (N_3399,N_1422,N_192);
or U3400 (N_3400,In_3955,In_977);
nor U3401 (N_3401,In_3973,In_3504);
or U3402 (N_3402,N_993,N_796);
or U3403 (N_3403,N_866,N_474);
nor U3404 (N_3404,N_1430,In_1168);
nand U3405 (N_3405,In_153,N_1234);
nor U3406 (N_3406,N_1411,In_141);
xor U3407 (N_3407,N_332,In_1270);
nor U3408 (N_3408,N_951,N_316);
or U3409 (N_3409,N_443,N_1305);
nand U3410 (N_3410,N_1453,N_920);
nor U3411 (N_3411,N_533,In_2779);
or U3412 (N_3412,N_1668,N_1742);
or U3413 (N_3413,N_1892,In_4117);
and U3414 (N_3414,In_744,N_727);
and U3415 (N_3415,In_2940,N_1382);
or U3416 (N_3416,N_802,In_2698);
nor U3417 (N_3417,N_811,In_4448);
nand U3418 (N_3418,In_3762,In_1639);
or U3419 (N_3419,N_1307,In_2674);
nand U3420 (N_3420,In_4738,In_4232);
nand U3421 (N_3421,N_911,N_655);
nor U3422 (N_3422,N_1780,In_2271);
and U3423 (N_3423,In_1955,In_2457);
or U3424 (N_3424,In_587,N_1511);
and U3425 (N_3425,N_1633,N_1148);
and U3426 (N_3426,N_1313,N_1508);
or U3427 (N_3427,In_2131,N_955);
nand U3428 (N_3428,In_3842,N_26);
and U3429 (N_3429,In_4093,N_358);
and U3430 (N_3430,N_913,N_384);
nor U3431 (N_3431,N_611,N_531);
and U3432 (N_3432,In_1481,N_986);
nor U3433 (N_3433,N_1684,N_1325);
nand U3434 (N_3434,In_2014,N_835);
nor U3435 (N_3435,N_1169,N_1594);
and U3436 (N_3436,N_1796,N_1944);
or U3437 (N_3437,N_1885,In_3700);
or U3438 (N_3438,N_992,In_4835);
and U3439 (N_3439,In_3136,N_181);
or U3440 (N_3440,N_1093,N_1557);
and U3441 (N_3441,N_949,N_1054);
or U3442 (N_3442,N_1734,In_4165);
and U3443 (N_3443,In_1617,N_189);
and U3444 (N_3444,N_528,N_1152);
nand U3445 (N_3445,In_569,N_1924);
nand U3446 (N_3446,In_4765,N_1337);
and U3447 (N_3447,In_1905,In_2033);
or U3448 (N_3448,N_788,N_1589);
and U3449 (N_3449,N_80,N_515);
and U3450 (N_3450,In_336,In_2204);
nor U3451 (N_3451,N_1328,N_333);
and U3452 (N_3452,In_4120,In_3607);
and U3453 (N_3453,N_997,In_3910);
nand U3454 (N_3454,N_1348,In_2668);
nor U3455 (N_3455,N_1905,In_4853);
and U3456 (N_3456,In_2273,N_1554);
nor U3457 (N_3457,N_853,N_180);
and U3458 (N_3458,N_184,N_939);
or U3459 (N_3459,N_704,In_3941);
nor U3460 (N_3460,In_4945,N_1529);
nand U3461 (N_3461,N_1285,In_1312);
nor U3462 (N_3462,N_707,In_486);
nor U3463 (N_3463,N_311,N_1486);
xor U3464 (N_3464,N_442,N_969);
or U3465 (N_3465,N_1544,N_56);
nor U3466 (N_3466,In_2363,In_2562);
nand U3467 (N_3467,N_1127,In_1182);
nor U3468 (N_3468,In_554,N_517);
nor U3469 (N_3469,N_1241,N_1899);
and U3470 (N_3470,N_621,N_1952);
or U3471 (N_3471,N_1282,N_1506);
nand U3472 (N_3472,N_61,N_1426);
or U3473 (N_3473,N_667,N_1050);
or U3474 (N_3474,N_1131,N_186);
and U3475 (N_3475,N_1754,In_639);
and U3476 (N_3476,N_1126,N_432);
or U3477 (N_3477,N_1053,In_4517);
or U3478 (N_3478,N_90,N_9);
and U3479 (N_3479,In_1048,N_1317);
and U3480 (N_3480,N_746,In_2165);
and U3481 (N_3481,N_347,N_349);
nor U3482 (N_3482,In_966,In_2778);
and U3483 (N_3483,N_1745,N_1605);
and U3484 (N_3484,N_1683,N_790);
or U3485 (N_3485,N_377,N_1179);
nand U3486 (N_3486,In_4162,N_1243);
nand U3487 (N_3487,N_980,In_3828);
or U3488 (N_3488,N_354,N_821);
nor U3489 (N_3489,In_1460,In_13);
and U3490 (N_3490,N_1853,N_373);
and U3491 (N_3491,In_2266,N_147);
or U3492 (N_3492,In_2862,In_1524);
and U3493 (N_3493,N_973,In_3727);
and U3494 (N_3494,N_926,N_1720);
nand U3495 (N_3495,N_101,In_3281);
nand U3496 (N_3496,N_1237,N_270);
or U3497 (N_3497,N_942,N_1517);
nand U3498 (N_3498,N_1825,In_1302);
and U3499 (N_3499,N_941,N_1790);
nor U3500 (N_3500,N_372,In_2685);
nor U3501 (N_3501,In_1099,N_153);
nor U3502 (N_3502,N_1107,In_191);
nand U3503 (N_3503,N_730,N_874);
or U3504 (N_3504,N_273,N_514);
nor U3505 (N_3505,In_3986,N_1424);
nand U3506 (N_3506,In_4028,In_4502);
and U3507 (N_3507,N_1700,N_1198);
nand U3508 (N_3508,In_4593,N_1869);
and U3509 (N_3509,N_1323,N_1122);
or U3510 (N_3510,N_1724,In_3464);
xor U3511 (N_3511,N_459,N_918);
and U3512 (N_3512,N_117,N_681);
nand U3513 (N_3513,N_1849,In_3835);
nor U3514 (N_3514,N_1211,N_270);
nor U3515 (N_3515,In_3064,N_445);
and U3516 (N_3516,N_189,In_3976);
nand U3517 (N_3517,N_695,In_3842);
and U3518 (N_3518,In_3018,In_2253);
and U3519 (N_3519,N_439,N_1603);
nand U3520 (N_3520,In_1622,N_504);
or U3521 (N_3521,N_1201,In_2285);
nand U3522 (N_3522,N_70,N_4);
xnor U3523 (N_3523,N_156,N_285);
nand U3524 (N_3524,In_3253,N_41);
or U3525 (N_3525,N_627,In_2654);
nor U3526 (N_3526,N_754,In_600);
or U3527 (N_3527,N_1627,N_1132);
or U3528 (N_3528,N_1822,N_475);
nor U3529 (N_3529,N_1379,In_4742);
or U3530 (N_3530,N_691,N_59);
and U3531 (N_3531,In_3955,N_1243);
nand U3532 (N_3532,N_1035,N_1360);
or U3533 (N_3533,In_212,N_397);
nand U3534 (N_3534,N_1470,N_548);
or U3535 (N_3535,N_269,In_3076);
and U3536 (N_3536,N_499,N_204);
nor U3537 (N_3537,In_3064,In_1275);
nor U3538 (N_3538,N_1024,In_1726);
nand U3539 (N_3539,N_388,In_589);
nand U3540 (N_3540,N_1948,N_688);
nor U3541 (N_3541,N_565,N_1125);
nor U3542 (N_3542,N_1618,N_5);
and U3543 (N_3543,In_3267,N_1282);
nand U3544 (N_3544,N_874,N_464);
nand U3545 (N_3545,N_134,N_1932);
nand U3546 (N_3546,N_66,In_4093);
nand U3547 (N_3547,N_785,In_4412);
or U3548 (N_3548,N_1809,In_4335);
or U3549 (N_3549,N_260,In_1851);
and U3550 (N_3550,N_1622,N_1722);
or U3551 (N_3551,N_1837,N_1038);
nand U3552 (N_3552,N_423,N_761);
nand U3553 (N_3553,N_184,N_1361);
and U3554 (N_3554,In_1896,In_3878);
and U3555 (N_3555,N_157,In_640);
nand U3556 (N_3556,In_169,In_4010);
nand U3557 (N_3557,N_1803,In_1731);
or U3558 (N_3558,In_3181,In_2685);
nand U3559 (N_3559,N_1939,N_1428);
nand U3560 (N_3560,In_1032,N_344);
or U3561 (N_3561,In_1622,N_1716);
or U3562 (N_3562,N_1984,In_4877);
xnor U3563 (N_3563,N_164,N_672);
nor U3564 (N_3564,In_2668,N_1769);
or U3565 (N_3565,N_575,N_1276);
nor U3566 (N_3566,In_679,In_1465);
nand U3567 (N_3567,In_4333,N_1574);
or U3568 (N_3568,N_1635,In_1355);
or U3569 (N_3569,In_3276,In_4335);
nor U3570 (N_3570,N_747,In_4020);
or U3571 (N_3571,N_1119,N_406);
or U3572 (N_3572,N_1996,In_4743);
or U3573 (N_3573,N_564,In_2734);
or U3574 (N_3574,N_277,In_2303);
nor U3575 (N_3575,N_1653,N_201);
nor U3576 (N_3576,N_1252,In_2742);
nand U3577 (N_3577,N_1467,N_1863);
nor U3578 (N_3578,In_1886,In_639);
and U3579 (N_3579,N_217,N_533);
nand U3580 (N_3580,In_3700,In_1474);
and U3581 (N_3581,N_250,In_3696);
nand U3582 (N_3582,N_1764,N_1406);
nand U3583 (N_3583,N_1263,N_451);
and U3584 (N_3584,In_1469,N_162);
nand U3585 (N_3585,N_273,In_1879);
and U3586 (N_3586,N_703,In_1402);
nor U3587 (N_3587,N_1535,N_1645);
and U3588 (N_3588,N_8,N_1066);
or U3589 (N_3589,N_579,N_1081);
nor U3590 (N_3590,N_897,In_3540);
nor U3591 (N_3591,In_2037,N_322);
nand U3592 (N_3592,N_355,In_4392);
or U3593 (N_3593,N_1843,N_252);
and U3594 (N_3594,N_1547,In_1278);
nand U3595 (N_3595,In_4358,In_4481);
or U3596 (N_3596,In_4771,N_360);
nor U3597 (N_3597,N_562,In_2668);
nor U3598 (N_3598,N_1227,In_1832);
nand U3599 (N_3599,In_2547,N_1187);
and U3600 (N_3600,N_541,In_2620);
and U3601 (N_3601,N_1520,In_366);
or U3602 (N_3602,N_246,In_55);
nor U3603 (N_3603,In_3330,In_825);
nand U3604 (N_3604,N_1465,In_4747);
or U3605 (N_3605,N_1249,In_342);
nor U3606 (N_3606,N_1468,N_967);
or U3607 (N_3607,N_629,In_4010);
or U3608 (N_3608,In_425,N_1002);
and U3609 (N_3609,N_902,In_1406);
or U3610 (N_3610,In_1632,N_1200);
or U3611 (N_3611,In_2199,N_897);
and U3612 (N_3612,N_319,In_1917);
nor U3613 (N_3613,In_587,N_347);
or U3614 (N_3614,In_1051,In_4587);
or U3615 (N_3615,In_2959,In_1465);
nand U3616 (N_3616,N_1157,In_978);
and U3617 (N_3617,In_1724,In_4130);
nor U3618 (N_3618,In_1824,N_1966);
and U3619 (N_3619,N_808,N_1263);
or U3620 (N_3620,N_1158,In_813);
nor U3621 (N_3621,N_1504,In_3093);
xnor U3622 (N_3622,In_3167,N_436);
and U3623 (N_3623,In_1119,In_1361);
or U3624 (N_3624,N_1602,In_483);
and U3625 (N_3625,N_1792,In_744);
nand U3626 (N_3626,N_1812,N_207);
xor U3627 (N_3627,In_3113,In_4765);
nor U3628 (N_3628,N_269,In_1465);
and U3629 (N_3629,N_1531,N_376);
and U3630 (N_3630,N_1251,N_98);
or U3631 (N_3631,In_3570,N_468);
and U3632 (N_3632,N_1673,N_1895);
or U3633 (N_3633,N_1403,N_149);
nand U3634 (N_3634,N_1861,N_578);
and U3635 (N_3635,In_4058,N_515);
xor U3636 (N_3636,N_141,In_330);
nand U3637 (N_3637,N_1692,N_192);
or U3638 (N_3638,In_3532,In_4358);
and U3639 (N_3639,N_1050,N_724);
or U3640 (N_3640,N_973,N_1910);
nand U3641 (N_3641,In_1639,N_376);
or U3642 (N_3642,N_1171,N_1197);
nand U3643 (N_3643,N_442,N_1723);
or U3644 (N_3644,N_959,N_779);
and U3645 (N_3645,N_1551,In_4347);
or U3646 (N_3646,In_592,In_2751);
nor U3647 (N_3647,N_806,N_1877);
nand U3648 (N_3648,N_968,In_1267);
xor U3649 (N_3649,N_68,N_1964);
and U3650 (N_3650,N_231,N_413);
nor U3651 (N_3651,N_1355,N_656);
nor U3652 (N_3652,N_535,N_1396);
nand U3653 (N_3653,In_3768,N_53);
and U3654 (N_3654,N_1110,N_731);
or U3655 (N_3655,N_726,N_1268);
or U3656 (N_3656,N_7,N_919);
or U3657 (N_3657,In_629,N_643);
or U3658 (N_3658,N_1626,In_4412);
nor U3659 (N_3659,In_4400,N_1562);
nor U3660 (N_3660,N_395,N_491);
and U3661 (N_3661,N_1266,N_531);
and U3662 (N_3662,N_695,N_714);
or U3663 (N_3663,In_483,N_1135);
nand U3664 (N_3664,N_316,N_717);
nand U3665 (N_3665,In_2938,N_1624);
and U3666 (N_3666,In_112,N_541);
nand U3667 (N_3667,N_310,In_3211);
or U3668 (N_3668,N_979,N_1980);
nor U3669 (N_3669,In_3267,N_974);
and U3670 (N_3670,N_1631,N_588);
nor U3671 (N_3671,N_889,In_1447);
and U3672 (N_3672,N_735,In_1924);
xnor U3673 (N_3673,N_1831,N_1851);
or U3674 (N_3674,In_4934,In_3050);
nor U3675 (N_3675,N_1577,N_1113);
nand U3676 (N_3676,N_665,N_44);
and U3677 (N_3677,N_1671,In_1406);
nand U3678 (N_3678,N_1075,N_1365);
nand U3679 (N_3679,In_202,N_318);
and U3680 (N_3680,N_1913,N_838);
nand U3681 (N_3681,N_1907,N_1973);
nor U3682 (N_3682,In_4448,N_799);
or U3683 (N_3683,N_1972,In_3905);
or U3684 (N_3684,In_494,N_1361);
nor U3685 (N_3685,N_1110,In_748);
nor U3686 (N_3686,N_1478,N_312);
and U3687 (N_3687,In_153,N_1569);
xnor U3688 (N_3688,N_843,In_1926);
nand U3689 (N_3689,In_3793,N_1698);
or U3690 (N_3690,N_329,N_1226);
and U3691 (N_3691,N_348,N_620);
or U3692 (N_3692,N_56,In_3281);
nand U3693 (N_3693,N_962,N_1288);
nor U3694 (N_3694,N_172,N_344);
and U3695 (N_3695,N_659,N_1507);
and U3696 (N_3696,In_337,N_842);
and U3697 (N_3697,N_1758,In_1739);
and U3698 (N_3698,In_4477,N_1905);
nor U3699 (N_3699,N_650,N_1772);
or U3700 (N_3700,In_4712,N_1692);
nand U3701 (N_3701,N_1241,N_1026);
nor U3702 (N_3702,N_1060,In_4358);
or U3703 (N_3703,N_1315,N_1512);
nand U3704 (N_3704,N_1491,N_1411);
nor U3705 (N_3705,In_2273,N_818);
nand U3706 (N_3706,N_428,N_1342);
nand U3707 (N_3707,N_1756,N_1286);
and U3708 (N_3708,N_1339,In_1124);
nand U3709 (N_3709,N_514,In_1465);
nand U3710 (N_3710,N_1181,N_1410);
xnor U3711 (N_3711,In_3195,N_500);
and U3712 (N_3712,In_2204,N_1908);
and U3713 (N_3713,N_1024,N_531);
or U3714 (N_3714,In_750,N_175);
nor U3715 (N_3715,N_342,N_252);
and U3716 (N_3716,In_1156,N_552);
nor U3717 (N_3717,In_1708,In_3637);
and U3718 (N_3718,N_1006,N_60);
or U3719 (N_3719,N_1717,In_3419);
nand U3720 (N_3720,In_880,N_1479);
nor U3721 (N_3721,N_709,In_1632);
nor U3722 (N_3722,N_1156,N_58);
nor U3723 (N_3723,In_3152,In_1148);
nand U3724 (N_3724,N_440,N_86);
nor U3725 (N_3725,N_1610,In_3478);
and U3726 (N_3726,N_961,In_3792);
and U3727 (N_3727,In_435,In_2366);
or U3728 (N_3728,N_1848,N_475);
and U3729 (N_3729,N_1954,N_26);
or U3730 (N_3730,N_1992,N_634);
or U3731 (N_3731,N_1016,N_1107);
nand U3732 (N_3732,N_111,N_277);
nand U3733 (N_3733,In_3654,N_307);
or U3734 (N_3734,N_1110,In_2276);
or U3735 (N_3735,In_2710,N_1565);
and U3736 (N_3736,In_3464,N_954);
nor U3737 (N_3737,N_1469,N_1982);
nor U3738 (N_3738,N_1691,In_899);
nor U3739 (N_3739,In_625,N_864);
or U3740 (N_3740,N_948,N_125);
and U3741 (N_3741,In_1616,N_1419);
and U3742 (N_3742,In_3580,In_4837);
and U3743 (N_3743,N_1044,In_2418);
and U3744 (N_3744,N_1671,N_1093);
nand U3745 (N_3745,In_2779,In_1608);
nor U3746 (N_3746,In_2762,In_309);
and U3747 (N_3747,N_1685,In_2328);
nand U3748 (N_3748,N_1854,In_782);
nor U3749 (N_3749,In_2864,N_448);
or U3750 (N_3750,N_333,N_1708);
or U3751 (N_3751,N_1579,N_1646);
nor U3752 (N_3752,N_66,In_68);
nand U3753 (N_3753,In_3507,In_1561);
nor U3754 (N_3754,N_1102,N_1976);
nand U3755 (N_3755,N_894,N_331);
or U3756 (N_3756,N_707,In_3050);
xor U3757 (N_3757,In_4810,In_1405);
and U3758 (N_3758,In_1032,N_1940);
nand U3759 (N_3759,In_3478,In_254);
xnor U3760 (N_3760,N_1545,N_31);
or U3761 (N_3761,In_4623,N_983);
or U3762 (N_3762,N_1648,N_1342);
and U3763 (N_3763,In_2988,N_295);
nor U3764 (N_3764,N_1050,N_546);
nor U3765 (N_3765,In_3707,N_1512);
nand U3766 (N_3766,N_521,In_3211);
nand U3767 (N_3767,N_1930,N_1083);
or U3768 (N_3768,In_3337,In_330);
nand U3769 (N_3769,N_978,N_1653);
and U3770 (N_3770,N_1443,In_3050);
or U3771 (N_3771,In_3303,In_2424);
nor U3772 (N_3772,In_4520,In_4502);
or U3773 (N_3773,N_502,N_62);
or U3774 (N_3774,N_839,N_391);
nand U3775 (N_3775,N_470,N_1279);
nor U3776 (N_3776,N_124,N_1854);
nand U3777 (N_3777,N_1997,N_1457);
nand U3778 (N_3778,In_860,In_1784);
and U3779 (N_3779,In_321,In_881);
nor U3780 (N_3780,In_222,In_1765);
and U3781 (N_3781,N_1025,N_386);
nand U3782 (N_3782,N_816,In_4390);
or U3783 (N_3783,In_1317,N_695);
and U3784 (N_3784,In_4977,N_1331);
or U3785 (N_3785,N_1932,In_477);
and U3786 (N_3786,N_80,N_1134);
nor U3787 (N_3787,In_4838,N_1123);
or U3788 (N_3788,N_1502,In_4478);
nand U3789 (N_3789,N_361,N_481);
or U3790 (N_3790,N_1248,N_1920);
nand U3791 (N_3791,N_639,N_580);
or U3792 (N_3792,N_308,In_1168);
nand U3793 (N_3793,In_1062,N_1139);
nand U3794 (N_3794,N_1364,N_1222);
nand U3795 (N_3795,N_1631,In_2161);
and U3796 (N_3796,In_1533,N_1911);
nand U3797 (N_3797,In_3986,N_1456);
or U3798 (N_3798,N_1427,In_4517);
and U3799 (N_3799,In_3862,N_1947);
nand U3800 (N_3800,N_1862,N_1315);
nor U3801 (N_3801,In_4630,N_944);
nand U3802 (N_3802,In_1642,In_1599);
nor U3803 (N_3803,N_1868,N_531);
or U3804 (N_3804,In_773,N_684);
or U3805 (N_3805,N_219,In_2842);
nor U3806 (N_3806,In_1708,In_1993);
and U3807 (N_3807,N_1105,N_110);
nand U3808 (N_3808,N_913,N_553);
and U3809 (N_3809,N_959,In_4879);
nor U3810 (N_3810,In_3064,In_2366);
or U3811 (N_3811,In_106,In_4977);
or U3812 (N_3812,N_736,In_4441);
or U3813 (N_3813,In_2297,N_1085);
or U3814 (N_3814,In_4585,In_800);
or U3815 (N_3815,N_170,N_18);
and U3816 (N_3816,In_3066,In_2307);
and U3817 (N_3817,N_182,N_1373);
nor U3818 (N_3818,N_375,N_1249);
or U3819 (N_3819,N_1986,N_442);
nand U3820 (N_3820,In_3358,N_1810);
nand U3821 (N_3821,N_514,N_399);
nand U3822 (N_3822,N_455,N_1400);
or U3823 (N_3823,N_1453,N_934);
and U3824 (N_3824,N_993,N_1818);
nand U3825 (N_3825,N_1125,N_1179);
nor U3826 (N_3826,In_889,In_3064);
and U3827 (N_3827,N_602,In_2763);
nand U3828 (N_3828,N_431,N_1075);
or U3829 (N_3829,In_4207,N_1938);
nor U3830 (N_3830,N_1774,In_3696);
or U3831 (N_3831,In_1522,In_39);
nand U3832 (N_3832,N_168,N_373);
nand U3833 (N_3833,N_1918,In_2787);
nor U3834 (N_3834,N_212,N_314);
and U3835 (N_3835,N_1148,In_953);
nand U3836 (N_3836,N_1895,N_1033);
and U3837 (N_3837,N_1660,N_1595);
or U3838 (N_3838,N_132,In_1137);
and U3839 (N_3839,N_664,In_3771);
nand U3840 (N_3840,In_1057,N_39);
nor U3841 (N_3841,In_4693,N_971);
nor U3842 (N_3842,N_1642,In_3870);
or U3843 (N_3843,N_288,N_1533);
nor U3844 (N_3844,N_355,N_251);
and U3845 (N_3845,N_774,N_1218);
and U3846 (N_3846,N_364,N_1210);
and U3847 (N_3847,In_496,N_1912);
and U3848 (N_3848,In_3809,N_605);
or U3849 (N_3849,N_1071,N_1390);
nor U3850 (N_3850,In_4565,N_930);
or U3851 (N_3851,N_594,In_1171);
and U3852 (N_3852,N_906,N_1570);
nor U3853 (N_3853,In_489,N_1860);
or U3854 (N_3854,N_573,N_1540);
or U3855 (N_3855,N_1229,N_1642);
or U3856 (N_3856,In_2037,N_364);
nand U3857 (N_3857,In_3423,N_1288);
nand U3858 (N_3858,N_198,N_1591);
nor U3859 (N_3859,N_153,In_2034);
nor U3860 (N_3860,N_105,N_732);
nand U3861 (N_3861,N_1078,In_2494);
nand U3862 (N_3862,N_1886,N_479);
nor U3863 (N_3863,In_3442,N_1116);
and U3864 (N_3864,N_1432,In_3986);
and U3865 (N_3865,In_4132,In_3020);
nor U3866 (N_3866,In_2847,N_805);
nand U3867 (N_3867,In_4634,N_524);
nand U3868 (N_3868,N_1992,In_1398);
nand U3869 (N_3869,N_705,In_2037);
or U3870 (N_3870,N_1832,N_1813);
or U3871 (N_3871,In_987,N_1382);
nand U3872 (N_3872,N_980,N_845);
and U3873 (N_3873,N_327,N_1497);
or U3874 (N_3874,In_3347,N_1369);
nand U3875 (N_3875,In_2119,In_1675);
and U3876 (N_3876,In_2505,N_499);
and U3877 (N_3877,N_1274,In_2976);
and U3878 (N_3878,In_2847,N_710);
or U3879 (N_3879,In_4360,In_2383);
nand U3880 (N_3880,N_149,In_3759);
nand U3881 (N_3881,N_679,N_1560);
and U3882 (N_3882,In_4147,N_1904);
nand U3883 (N_3883,N_1111,N_1224);
nor U3884 (N_3884,N_1066,N_1109);
or U3885 (N_3885,N_650,In_3615);
and U3886 (N_3886,N_508,N_484);
nor U3887 (N_3887,N_1834,In_1099);
nand U3888 (N_3888,In_2129,In_2917);
or U3889 (N_3889,In_715,In_2658);
and U3890 (N_3890,N_1419,In_3084);
nor U3891 (N_3891,N_609,N_364);
nor U3892 (N_3892,In_1198,N_519);
nor U3893 (N_3893,In_1572,N_101);
nor U3894 (N_3894,N_262,In_4613);
or U3895 (N_3895,N_685,In_1894);
and U3896 (N_3896,N_1830,N_1927);
or U3897 (N_3897,N_1490,N_1096);
or U3898 (N_3898,N_1391,N_1317);
or U3899 (N_3899,In_400,N_1943);
nand U3900 (N_3900,In_3856,N_1628);
nand U3901 (N_3901,In_1608,N_1246);
or U3902 (N_3902,In_234,In_825);
nand U3903 (N_3903,N_982,In_634);
nand U3904 (N_3904,N_512,N_1725);
nor U3905 (N_3905,N_1761,N_1852);
nand U3906 (N_3906,In_4167,N_596);
nor U3907 (N_3907,N_81,N_1915);
nand U3908 (N_3908,In_1382,In_1042);
and U3909 (N_3909,N_1606,N_1531);
nor U3910 (N_3910,N_1890,N_527);
and U3911 (N_3911,N_1990,N_493);
or U3912 (N_3912,In_1339,N_592);
and U3913 (N_3913,N_1562,In_3527);
or U3914 (N_3914,N_1161,N_1930);
nor U3915 (N_3915,N_1653,N_1304);
or U3916 (N_3916,N_250,N_1308);
nand U3917 (N_3917,N_1869,N_1333);
nand U3918 (N_3918,N_26,In_2288);
or U3919 (N_3919,N_1088,N_1985);
or U3920 (N_3920,N_200,N_1746);
nor U3921 (N_3921,N_1556,N_1411);
and U3922 (N_3922,N_808,N_27);
nand U3923 (N_3923,N_1394,In_1491);
or U3924 (N_3924,N_1352,N_1303);
and U3925 (N_3925,In_4838,N_822);
nor U3926 (N_3926,In_4626,N_1262);
and U3927 (N_3927,N_1476,N_913);
nand U3928 (N_3928,N_194,In_55);
and U3929 (N_3929,N_384,In_2646);
nor U3930 (N_3930,N_1736,In_868);
nor U3931 (N_3931,N_383,N_1152);
and U3932 (N_3932,In_4623,In_2765);
or U3933 (N_3933,N_1843,In_838);
nor U3934 (N_3934,In_1992,N_1434);
nor U3935 (N_3935,N_1213,N_598);
and U3936 (N_3936,N_145,N_1682);
and U3937 (N_3937,N_1082,In_2870);
nand U3938 (N_3938,N_1623,In_4997);
or U3939 (N_3939,N_433,N_931);
or U3940 (N_3940,In_2306,N_159);
nor U3941 (N_3941,In_2383,N_1556);
and U3942 (N_3942,N_826,N_1410);
xnor U3943 (N_3943,N_440,In_4108);
or U3944 (N_3944,N_829,N_170);
xor U3945 (N_3945,N_714,N_1879);
nor U3946 (N_3946,In_2771,N_189);
and U3947 (N_3947,N_268,N_160);
and U3948 (N_3948,N_1172,N_244);
nand U3949 (N_3949,In_1547,In_55);
and U3950 (N_3950,N_1191,In_496);
and U3951 (N_3951,N_911,In_2660);
or U3952 (N_3952,N_40,N_770);
and U3953 (N_3953,In_2328,N_1237);
and U3954 (N_3954,N_1615,In_825);
nand U3955 (N_3955,N_1280,N_543);
nand U3956 (N_3956,N_34,N_217);
and U3957 (N_3957,In_1522,N_1715);
or U3958 (N_3958,In_1747,N_1004);
and U3959 (N_3959,N_498,In_2037);
nor U3960 (N_3960,In_3068,N_185);
nand U3961 (N_3961,In_31,N_1652);
or U3962 (N_3962,N_781,N_73);
nand U3963 (N_3963,N_1507,N_1810);
nor U3964 (N_3964,In_3452,N_316);
nor U3965 (N_3965,In_2062,N_1229);
xor U3966 (N_3966,N_1853,N_1265);
and U3967 (N_3967,N_1299,N_1154);
nand U3968 (N_3968,N_249,N_1900);
nand U3969 (N_3969,N_172,N_1760);
and U3970 (N_3970,N_116,In_1724);
xnor U3971 (N_3971,N_216,N_404);
nand U3972 (N_3972,In_611,N_1505);
nand U3973 (N_3973,N_125,N_405);
nand U3974 (N_3974,In_1420,N_1029);
or U3975 (N_3975,N_957,N_1275);
or U3976 (N_3976,N_1484,N_282);
nor U3977 (N_3977,N_1255,In_2246);
or U3978 (N_3978,In_2246,N_1655);
nand U3979 (N_3979,N_1223,N_1207);
or U3980 (N_3980,N_1122,N_899);
nor U3981 (N_3981,N_477,N_1314);
nor U3982 (N_3982,In_4390,N_1306);
or U3983 (N_3983,N_1883,In_2288);
nor U3984 (N_3984,N_1101,N_641);
nor U3985 (N_3985,N_276,In_4540);
nand U3986 (N_3986,N_592,N_534);
or U3987 (N_3987,N_1372,N_202);
and U3988 (N_3988,N_746,N_1229);
xnor U3989 (N_3989,N_1574,N_1505);
or U3990 (N_3990,In_824,In_486);
and U3991 (N_3991,N_1397,N_1823);
and U3992 (N_3992,In_3925,N_786);
nand U3993 (N_3993,N_1936,In_4634);
nand U3994 (N_3994,N_679,N_411);
nand U3995 (N_3995,N_1502,N_858);
or U3996 (N_3996,N_1120,In_3862);
nand U3997 (N_3997,In_3870,N_1973);
nand U3998 (N_3998,In_2084,N_153);
and U3999 (N_3999,N_573,N_1036);
or U4000 (N_4000,N_2129,N_3871);
nand U4001 (N_4001,N_3238,N_3656);
nand U4002 (N_4002,N_2494,N_2477);
or U4003 (N_4003,N_2158,N_3802);
nor U4004 (N_4004,N_3374,N_2107);
nand U4005 (N_4005,N_3733,N_3738);
and U4006 (N_4006,N_3072,N_3890);
and U4007 (N_4007,N_3628,N_2985);
nand U4008 (N_4008,N_2416,N_2659);
and U4009 (N_4009,N_3322,N_2551);
or U4010 (N_4010,N_3271,N_3017);
nand U4011 (N_4011,N_2971,N_2160);
nor U4012 (N_4012,N_3346,N_2501);
nand U4013 (N_4013,N_3800,N_3601);
or U4014 (N_4014,N_2064,N_2113);
and U4015 (N_4015,N_3670,N_3371);
nand U4016 (N_4016,N_3023,N_3648);
nor U4017 (N_4017,N_2530,N_3986);
or U4018 (N_4018,N_2697,N_3555);
nand U4019 (N_4019,N_3360,N_2749);
and U4020 (N_4020,N_2110,N_3095);
nand U4021 (N_4021,N_2678,N_3012);
or U4022 (N_4022,N_3908,N_2790);
or U4023 (N_4023,N_2184,N_2376);
nor U4024 (N_4024,N_2937,N_2900);
or U4025 (N_4025,N_2926,N_2849);
xor U4026 (N_4026,N_2084,N_2941);
and U4027 (N_4027,N_2031,N_3968);
and U4028 (N_4028,N_2723,N_2743);
or U4029 (N_4029,N_2180,N_3508);
or U4030 (N_4030,N_3454,N_3070);
nor U4031 (N_4031,N_2325,N_3214);
and U4032 (N_4032,N_2015,N_3062);
and U4033 (N_4033,N_2652,N_3492);
nor U4034 (N_4034,N_3893,N_2375);
nand U4035 (N_4035,N_2228,N_3803);
or U4036 (N_4036,N_2498,N_2673);
nand U4037 (N_4037,N_3898,N_2062);
nand U4038 (N_4038,N_3328,N_3318);
xor U4039 (N_4039,N_3874,N_2271);
nand U4040 (N_4040,N_3566,N_2568);
nor U4041 (N_4041,N_3189,N_2818);
nor U4042 (N_4042,N_3806,N_3166);
nor U4043 (N_4043,N_2493,N_3600);
nand U4044 (N_4044,N_3515,N_2117);
and U4045 (N_4045,N_3570,N_2579);
nand U4046 (N_4046,N_3462,N_3080);
nand U4047 (N_4047,N_2753,N_3365);
nor U4048 (N_4048,N_2317,N_3042);
nand U4049 (N_4049,N_2936,N_2209);
xor U4050 (N_4050,N_3152,N_2897);
xor U4051 (N_4051,N_3305,N_3644);
and U4052 (N_4052,N_3688,N_2126);
or U4053 (N_4053,N_2448,N_3219);
or U4054 (N_4054,N_3827,N_2267);
or U4055 (N_4055,N_2982,N_2332);
nor U4056 (N_4056,N_3684,N_2385);
and U4057 (N_4057,N_3993,N_2420);
xor U4058 (N_4058,N_3003,N_3220);
nand U4059 (N_4059,N_2205,N_3263);
nand U4060 (N_4060,N_2224,N_2421);
or U4061 (N_4061,N_3426,N_2513);
nor U4062 (N_4062,N_2452,N_2475);
nor U4063 (N_4063,N_2237,N_2447);
or U4064 (N_4064,N_3541,N_3856);
nand U4065 (N_4065,N_2973,N_3063);
and U4066 (N_4066,N_2724,N_2812);
nor U4067 (N_4067,N_3341,N_2518);
nand U4068 (N_4068,N_3417,N_3580);
nand U4069 (N_4069,N_2217,N_2140);
or U4070 (N_4070,N_3414,N_2087);
nor U4071 (N_4071,N_3966,N_3604);
or U4072 (N_4072,N_3257,N_3234);
and U4073 (N_4073,N_2902,N_2100);
or U4074 (N_4074,N_2063,N_3217);
and U4075 (N_4075,N_2042,N_2044);
and U4076 (N_4076,N_2961,N_2757);
or U4077 (N_4077,N_3696,N_2457);
nand U4078 (N_4078,N_3721,N_3737);
or U4079 (N_4079,N_2067,N_2861);
nand U4080 (N_4080,N_3209,N_3973);
and U4081 (N_4081,N_3106,N_3598);
or U4082 (N_4082,N_3048,N_3101);
nand U4083 (N_4083,N_2685,N_2384);
and U4084 (N_4084,N_3490,N_2988);
or U4085 (N_4085,N_2574,N_3897);
nor U4086 (N_4086,N_2735,N_3694);
nand U4087 (N_4087,N_2965,N_3825);
nand U4088 (N_4088,N_3573,N_3997);
nor U4089 (N_4089,N_3211,N_2388);
and U4090 (N_4090,N_3819,N_3218);
nor U4091 (N_4091,N_3995,N_2169);
nor U4092 (N_4092,N_2689,N_3470);
nor U4093 (N_4093,N_3449,N_3677);
or U4094 (N_4094,N_2230,N_3581);
or U4095 (N_4095,N_3979,N_3693);
or U4096 (N_4096,N_2868,N_2709);
and U4097 (N_4097,N_2444,N_3407);
and U4098 (N_4098,N_3061,N_3536);
nor U4099 (N_4099,N_3611,N_3941);
or U4100 (N_4100,N_2045,N_2731);
nor U4101 (N_4101,N_2762,N_2281);
and U4102 (N_4102,N_3561,N_3041);
nand U4103 (N_4103,N_2650,N_3722);
or U4104 (N_4104,N_2144,N_3911);
and U4105 (N_4105,N_3148,N_3394);
and U4106 (N_4106,N_3633,N_3437);
and U4107 (N_4107,N_3781,N_2060);
and U4108 (N_4108,N_2086,N_3950);
or U4109 (N_4109,N_3790,N_2078);
and U4110 (N_4110,N_2472,N_3491);
or U4111 (N_4111,N_2360,N_3546);
and U4112 (N_4112,N_2565,N_2622);
nor U4113 (N_4113,N_2041,N_2030);
nor U4114 (N_4114,N_3196,N_3430);
and U4115 (N_4115,N_3554,N_2901);
or U4116 (N_4116,N_2567,N_3000);
nor U4117 (N_4117,N_3504,N_3547);
nand U4118 (N_4118,N_2666,N_2744);
and U4119 (N_4119,N_2223,N_3735);
nor U4120 (N_4120,N_3351,N_2729);
nand U4121 (N_4121,N_2034,N_3047);
or U4122 (N_4122,N_2279,N_2634);
and U4123 (N_4123,N_2337,N_3882);
and U4124 (N_4124,N_3009,N_3512);
or U4125 (N_4125,N_2584,N_2798);
nand U4126 (N_4126,N_2779,N_3232);
and U4127 (N_4127,N_3625,N_2502);
nor U4128 (N_4128,N_2688,N_3422);
nand U4129 (N_4129,N_3103,N_3946);
or U4130 (N_4130,N_2512,N_2197);
and U4131 (N_4131,N_3499,N_3181);
nand U4132 (N_4132,N_3732,N_2268);
nand U4133 (N_4133,N_3794,N_2202);
nand U4134 (N_4134,N_2250,N_3169);
nor U4135 (N_4135,N_2508,N_3076);
and U4136 (N_4136,N_3475,N_3496);
nor U4137 (N_4137,N_3237,N_3918);
nor U4138 (N_4138,N_2137,N_3355);
and U4139 (N_4139,N_3354,N_2733);
nor U4140 (N_4140,N_2708,N_3105);
nor U4141 (N_4141,N_2806,N_2663);
or U4142 (N_4142,N_3311,N_3087);
and U4143 (N_4143,N_3746,N_3309);
and U4144 (N_4144,N_3823,N_3117);
xor U4145 (N_4145,N_2528,N_3524);
nor U4146 (N_4146,N_3659,N_3368);
and U4147 (N_4147,N_2185,N_2639);
nor U4148 (N_4148,N_2213,N_3944);
nor U4149 (N_4149,N_2032,N_3165);
and U4150 (N_4150,N_2767,N_2782);
or U4151 (N_4151,N_2800,N_2231);
nand U4152 (N_4152,N_3246,N_3976);
nor U4153 (N_4153,N_2758,N_2934);
nand U4154 (N_4154,N_2641,N_3016);
nor U4155 (N_4155,N_3223,N_2296);
and U4156 (N_4156,N_3534,N_3099);
nor U4157 (N_4157,N_3847,N_3431);
xor U4158 (N_4158,N_2057,N_3613);
and U4159 (N_4159,N_3846,N_3637);
and U4160 (N_4160,N_2092,N_2823);
nor U4161 (N_4161,N_3353,N_2953);
nand U4162 (N_4162,N_2880,N_3467);
and U4163 (N_4163,N_3359,N_2661);
or U4164 (N_4164,N_2065,N_2895);
nor U4165 (N_4165,N_3844,N_2395);
nand U4166 (N_4166,N_3521,N_2349);
or U4167 (N_4167,N_3975,N_3939);
nand U4168 (N_4168,N_2235,N_3182);
nor U4169 (N_4169,N_2326,N_3765);
nand U4170 (N_4170,N_2949,N_2777);
nor U4171 (N_4171,N_3100,N_2108);
nand U4172 (N_4172,N_2370,N_3610);
nand U4173 (N_4173,N_3956,N_2910);
and U4174 (N_4174,N_2099,N_3129);
or U4175 (N_4175,N_2648,N_3502);
and U4176 (N_4176,N_3098,N_2970);
or U4177 (N_4177,N_3205,N_2525);
and U4178 (N_4178,N_3878,N_2262);
and U4179 (N_4179,N_3093,N_3964);
and U4180 (N_4180,N_2682,N_2431);
or U4181 (N_4181,N_3690,N_2357);
xor U4182 (N_4182,N_2399,N_2499);
nand U4183 (N_4183,N_2856,N_2581);
nand U4184 (N_4184,N_2911,N_3477);
or U4185 (N_4185,N_3378,N_3327);
nand U4186 (N_4186,N_3867,N_2667);
nand U4187 (N_4187,N_3402,N_3828);
nand U4188 (N_4188,N_2429,N_2162);
nor U4189 (N_4189,N_2462,N_3367);
nor U4190 (N_4190,N_3933,N_2321);
nor U4191 (N_4191,N_3658,N_2719);
nand U4192 (N_4192,N_3317,N_3830);
and U4193 (N_4193,N_3667,N_3319);
or U4194 (N_4194,N_2024,N_2869);
or U4195 (N_4195,N_2134,N_3291);
or U4196 (N_4196,N_2542,N_3817);
and U4197 (N_4197,N_2786,N_3591);
and U4198 (N_4198,N_3734,N_3358);
and U4199 (N_4199,N_3653,N_3789);
nor U4200 (N_4200,N_2964,N_3410);
nand U4201 (N_4201,N_2526,N_3938);
and U4202 (N_4202,N_2163,N_3382);
nand U4203 (N_4203,N_2585,N_3224);
nand U4204 (N_4204,N_2920,N_2559);
or U4205 (N_4205,N_3719,N_2538);
and U4206 (N_4206,N_2784,N_2925);
nor U4207 (N_4207,N_2956,N_2621);
nand U4208 (N_4208,N_3195,N_3969);
or U4209 (N_4209,N_2963,N_3880);
nand U4210 (N_4210,N_3162,N_3060);
nor U4211 (N_4211,N_2258,N_2437);
or U4212 (N_4212,N_3756,N_3935);
and U4213 (N_4213,N_2625,N_3068);
nor U4214 (N_4214,N_3481,N_3930);
or U4215 (N_4215,N_3122,N_2272);
or U4216 (N_4216,N_2788,N_3302);
or U4217 (N_4217,N_2742,N_2280);
nand U4218 (N_4218,N_2875,N_2571);
nor U4219 (N_4219,N_2587,N_3123);
nor U4220 (N_4220,N_2781,N_3339);
or U4221 (N_4221,N_3249,N_3574);
or U4222 (N_4222,N_2527,N_2051);
nor U4223 (N_4223,N_3198,N_2674);
and U4224 (N_4224,N_2717,N_2705);
nor U4225 (N_4225,N_3620,N_3888);
and U4226 (N_4226,N_3362,N_3836);
or U4227 (N_4227,N_2684,N_3233);
nand U4228 (N_4228,N_3344,N_2403);
xor U4229 (N_4229,N_2860,N_2830);
nand U4230 (N_4230,N_3260,N_2374);
and U4231 (N_4231,N_2341,N_3032);
and U4232 (N_4232,N_2642,N_3266);
and U4233 (N_4233,N_2362,N_3379);
nor U4234 (N_4234,N_3961,N_2241);
xnor U4235 (N_4235,N_2643,N_3283);
nand U4236 (N_4236,N_2871,N_2396);
nor U4237 (N_4237,N_3672,N_3511);
nand U4238 (N_4238,N_3370,N_2995);
and U4239 (N_4239,N_3928,N_3927);
nor U4240 (N_4240,N_2245,N_2836);
nand U4241 (N_4241,N_2566,N_3241);
nor U4242 (N_4242,N_3288,N_2750);
nor U4243 (N_4243,N_2894,N_3810);
and U4244 (N_4244,N_2293,N_3717);
or U4245 (N_4245,N_2948,N_3069);
nor U4246 (N_4246,N_3284,N_3043);
and U4247 (N_4247,N_3300,N_2549);
or U4248 (N_4248,N_3133,N_2632);
nand U4249 (N_4249,N_3204,N_3548);
or U4250 (N_4250,N_2408,N_2737);
xor U4251 (N_4251,N_3952,N_2738);
nand U4252 (N_4252,N_3024,N_3977);
or U4253 (N_4253,N_3139,N_2255);
and U4254 (N_4254,N_3974,N_3177);
nand U4255 (N_4255,N_3783,N_3669);
or U4256 (N_4256,N_2101,N_3796);
nor U4257 (N_4257,N_3290,N_2016);
and U4258 (N_4258,N_2294,N_2766);
nor U4259 (N_4259,N_3877,N_2819);
nor U4260 (N_4260,N_3683,N_2921);
nor U4261 (N_4261,N_2851,N_2390);
xnor U4262 (N_4262,N_2583,N_3759);
or U4263 (N_4263,N_2591,N_3630);
and U4264 (N_4264,N_3923,N_2019);
or U4265 (N_4265,N_3229,N_3978);
nand U4266 (N_4266,N_3662,N_2993);
or U4267 (N_4267,N_2404,N_3942);
nor U4268 (N_4268,N_3203,N_2852);
and U4269 (N_4269,N_3622,N_2001);
nor U4270 (N_4270,N_3797,N_3022);
nand U4271 (N_4271,N_3347,N_2138);
and U4272 (N_4272,N_3231,N_2473);
and U4273 (N_4273,N_3632,N_3001);
nor U4274 (N_4274,N_3804,N_3035);
and U4275 (N_4275,N_3583,N_2589);
nor U4276 (N_4276,N_3155,N_2487);
and U4277 (N_4277,N_3352,N_3831);
nand U4278 (N_4278,N_2668,N_3255);
or U4279 (N_4279,N_3616,N_2679);
nor U4280 (N_4280,N_2713,N_2198);
nand U4281 (N_4281,N_2468,N_2345);
nor U4282 (N_4282,N_3326,N_3143);
nor U4283 (N_4283,N_3623,N_3909);
nand U4284 (N_4284,N_2485,N_3543);
and U4285 (N_4285,N_2789,N_3277);
nor U4286 (N_4286,N_2515,N_3349);
nand U4287 (N_4287,N_3807,N_3599);
nand U4288 (N_4288,N_2827,N_3275);
or U4289 (N_4289,N_2547,N_2139);
nor U4290 (N_4290,N_3798,N_3709);
or U4291 (N_4291,N_2870,N_2662);
nand U4292 (N_4292,N_3842,N_3748);
nor U4293 (N_4293,N_2531,N_2211);
or U4294 (N_4294,N_3645,N_3618);
and U4295 (N_4295,N_2038,N_2402);
or U4296 (N_4296,N_2156,N_2930);
and U4297 (N_4297,N_2103,N_3274);
or U4298 (N_4298,N_3818,N_3313);
xor U4299 (N_4299,N_3592,N_2602);
nor U4300 (N_4300,N_3651,N_3350);
nand U4301 (N_4301,N_3212,N_3936);
nor U4302 (N_4302,N_2026,N_3739);
xnor U4303 (N_4303,N_2481,N_2633);
or U4304 (N_4304,N_3901,N_2972);
nor U4305 (N_4305,N_3951,N_2543);
nor U4306 (N_4306,N_3102,N_2843);
or U4307 (N_4307,N_3466,N_3862);
or U4308 (N_4308,N_2675,N_3227);
nor U4309 (N_4309,N_3532,N_3400);
or U4310 (N_4310,N_3285,N_2355);
or U4311 (N_4311,N_2425,N_2014);
nor U4312 (N_4312,N_3408,N_3985);
and U4313 (N_4313,N_2152,N_3920);
nand U4314 (N_4314,N_3784,N_2414);
or U4315 (N_4315,N_3235,N_3480);
and U4316 (N_4316,N_3999,N_2619);
or U4317 (N_4317,N_3766,N_2056);
and U4318 (N_4318,N_2569,N_3436);
nor U4319 (N_4319,N_2888,N_2389);
nor U4320 (N_4320,N_3404,N_3593);
nor U4321 (N_4321,N_3210,N_3779);
or U4322 (N_4322,N_3833,N_3465);
nor U4323 (N_4323,N_3805,N_3160);
nand U4324 (N_4324,N_2453,N_2336);
or U4325 (N_4325,N_2933,N_2826);
xor U4326 (N_4326,N_2623,N_2540);
or U4327 (N_4327,N_2315,N_3700);
nor U4328 (N_4328,N_2415,N_2669);
nand U4329 (N_4329,N_2149,N_2302);
or U4330 (N_4330,N_3770,N_2975);
nand U4331 (N_4331,N_2104,N_3471);
or U4332 (N_4332,N_2997,N_2610);
nand U4333 (N_4333,N_3419,N_3483);
nand U4334 (N_4334,N_2809,N_2210);
or U4335 (N_4335,N_2079,N_3896);
or U4336 (N_4336,N_3820,N_2102);
nand U4337 (N_4337,N_2381,N_3922);
nor U4338 (N_4338,N_3692,N_3340);
nor U4339 (N_4339,N_2655,N_2700);
nand U4340 (N_4340,N_2520,N_3086);
and U4341 (N_4341,N_3164,N_3046);
nand U4342 (N_4342,N_2096,N_3673);
nor U4343 (N_4343,N_2984,N_2489);
or U4344 (N_4344,N_2599,N_3058);
nand U4345 (N_4345,N_2470,N_3411);
and U4346 (N_4346,N_2859,N_3453);
or U4347 (N_4347,N_2146,N_2720);
and U4348 (N_4348,N_2514,N_3640);
nand U4349 (N_4349,N_3082,N_2855);
or U4350 (N_4350,N_2833,N_2906);
nand U4351 (N_4351,N_2368,N_3056);
xnor U4352 (N_4352,N_2524,N_2270);
and U4353 (N_4353,N_2168,N_3460);
nand U4354 (N_4354,N_3540,N_2838);
or U4355 (N_4355,N_3854,N_3256);
nor U4356 (N_4356,N_3868,N_3663);
and U4357 (N_4357,N_3903,N_2564);
nor U4358 (N_4358,N_3074,N_2776);
nor U4359 (N_4359,N_2919,N_2557);
nor U4360 (N_4360,N_2863,N_3170);
and U4361 (N_4361,N_2745,N_2842);
xor U4362 (N_4362,N_3708,N_3731);
nand U4363 (N_4363,N_3097,N_2333);
or U4364 (N_4364,N_2486,N_3110);
nand U4365 (N_4365,N_2507,N_3495);
and U4366 (N_4366,N_3121,N_3916);
or U4367 (N_4367,N_3059,N_2174);
xnor U4368 (N_4368,N_2885,N_3179);
and U4369 (N_4369,N_2068,N_2273);
or U4370 (N_4370,N_3364,N_2406);
nand U4371 (N_4371,N_3773,N_2968);
or U4372 (N_4372,N_3065,N_3085);
and U4373 (N_4373,N_2534,N_2841);
nor U4374 (N_4374,N_2710,N_2857);
or U4375 (N_4375,N_3201,N_3163);
nor U4376 (N_4376,N_2066,N_2318);
or U4377 (N_4377,N_2077,N_3438);
or U4378 (N_4378,N_3627,N_3306);
nand U4379 (N_4379,N_2006,N_3753);
and U4380 (N_4380,N_3641,N_2119);
or U4381 (N_4381,N_2133,N_2931);
and U4382 (N_4382,N_2094,N_3252);
nand U4383 (N_4383,N_3221,N_2831);
and U4384 (N_4384,N_3468,N_3811);
xnor U4385 (N_4385,N_3391,N_3006);
and U4386 (N_4386,N_3990,N_3487);
and U4387 (N_4387,N_3712,N_3760);
nor U4388 (N_4388,N_2876,N_3075);
or U4389 (N_4389,N_2221,N_3791);
and U4390 (N_4390,N_2131,N_2496);
nor U4391 (N_4391,N_2291,N_2282);
nand U4392 (N_4392,N_3751,N_2834);
or U4393 (N_4393,N_3792,N_2994);
and U4394 (N_4394,N_2482,N_2116);
nand U4395 (N_4395,N_2867,N_2264);
nor U4396 (N_4396,N_2035,N_3655);
nor U4397 (N_4397,N_2696,N_2234);
and U4398 (N_4398,N_3715,N_3387);
nand U4399 (N_4399,N_2986,N_2635);
and U4400 (N_4400,N_3366,N_2106);
nor U4401 (N_4401,N_2124,N_2627);
nor U4402 (N_4402,N_3176,N_3560);
nor U4403 (N_4403,N_3572,N_2218);
nor U4404 (N_4404,N_3900,N_3559);
and U4405 (N_4405,N_2275,N_2778);
nand U4406 (N_4406,N_2358,N_2554);
and U4407 (N_4407,N_3297,N_2216);
or U4408 (N_4408,N_3057,N_2979);
or U4409 (N_4409,N_2492,N_3192);
and U4410 (N_4410,N_3191,N_2027);
and U4411 (N_4411,N_2795,N_3259);
or U4412 (N_4412,N_3718,N_2850);
and U4413 (N_4413,N_3484,N_2153);
nand U4414 (N_4414,N_2483,N_2322);
or U4415 (N_4415,N_2186,N_3154);
nor U4416 (N_4416,N_3435,N_2017);
and U4417 (N_4417,N_2397,N_2242);
and U4418 (N_4418,N_2200,N_3158);
and U4419 (N_4419,N_3631,N_2394);
nor U4420 (N_4420,N_2418,N_3567);
nand U4421 (N_4421,N_2076,N_3464);
nor U4422 (N_4422,N_3373,N_2866);
nor U4423 (N_4423,N_2128,N_3914);
or U4424 (N_4424,N_3958,N_3845);
nor U4425 (N_4425,N_3747,N_2265);
nand U4426 (N_4426,N_2891,N_2509);
and U4427 (N_4427,N_3517,N_2334);
and U4428 (N_4428,N_3857,N_3873);
nor U4429 (N_4429,N_2922,N_2354);
nand U4430 (N_4430,N_2207,N_2284);
nor U4431 (N_4431,N_3758,N_2539);
nand U4432 (N_4432,N_3984,N_2261);
nor U4433 (N_4433,N_3409,N_3850);
or U4434 (N_4434,N_2154,N_2011);
or U4435 (N_4435,N_2792,N_3614);
and U4436 (N_4436,N_3582,N_3740);
nor U4437 (N_4437,N_2159,N_3859);
and U4438 (N_4438,N_3416,N_2810);
or U4439 (N_4439,N_2718,N_2908);
nor U4440 (N_4440,N_2594,N_2952);
nand U4441 (N_4441,N_3463,N_2835);
nand U4442 (N_4442,N_3126,N_3073);
nor U4443 (N_4443,N_2435,N_3034);
nor U4444 (N_4444,N_3421,N_3308);
nand U4445 (N_4445,N_3537,N_3183);
nand U4446 (N_4446,N_2939,N_3994);
or U4447 (N_4447,N_2433,N_3316);
nand U4448 (N_4448,N_2111,N_3486);
or U4449 (N_4449,N_2365,N_3094);
nor U4450 (N_4450,N_3138,N_3595);
nand U4451 (N_4451,N_3125,N_2423);
or U4452 (N_4452,N_3834,N_3795);
or U4453 (N_4453,N_2458,N_2148);
and U4454 (N_4454,N_2191,N_3187);
nand U4455 (N_4455,N_2563,N_3225);
nor U4456 (N_4456,N_2872,N_2614);
nand U4457 (N_4457,N_2353,N_3552);
and U4458 (N_4458,N_3334,N_3472);
or U4459 (N_4459,N_2058,N_2712);
nor U4460 (N_4460,N_3479,N_2794);
and U4461 (N_4461,N_3703,N_3931);
and U4462 (N_4462,N_3425,N_3096);
nand U4463 (N_4463,N_2658,N_2962);
and U4464 (N_4464,N_2575,N_3115);
nand U4465 (N_4465,N_3741,N_2081);
and U4466 (N_4466,N_3743,N_3242);
and U4467 (N_4467,N_2127,N_2383);
or U4468 (N_4468,N_2944,N_3962);
nand U4469 (N_4469,N_3886,N_2638);
nor U4470 (N_4470,N_2990,N_2410);
and U4471 (N_4471,N_3375,N_2611);
or U4472 (N_4472,N_3907,N_3423);
and U4473 (N_4473,N_2367,N_3039);
or U4474 (N_4474,N_2677,N_2441);
and U4475 (N_4475,N_2828,N_3925);
or U4476 (N_4476,N_3149,N_3014);
nor U4477 (N_4477,N_2259,N_3396);
and U4478 (N_4478,N_2455,N_3498);
or U4479 (N_4479,N_3119,N_2340);
and U4480 (N_4480,N_3937,N_2824);
nand U4481 (N_4481,N_3077,N_3533);
nand U4482 (N_4482,N_2747,N_3771);
nand U4483 (N_4483,N_2532,N_2883);
nand U4484 (N_4484,N_2351,N_2248);
nand U4485 (N_4485,N_3705,N_3587);
and U4486 (N_4486,N_3776,N_3565);
nand U4487 (N_4487,N_2225,N_2232);
and U4488 (N_4488,N_3714,N_2233);
or U4489 (N_4489,N_2491,N_2523);
and U4490 (N_4490,N_2844,N_2135);
and U4491 (N_4491,N_3775,N_3838);
or U4492 (N_4492,N_3755,N_3084);
and U4493 (N_4493,N_3276,N_3934);
nand U4494 (N_4494,N_3821,N_2061);
nor U4495 (N_4495,N_2671,N_2624);
or U4496 (N_4496,N_3294,N_2151);
or U4497 (N_4497,N_2243,N_2003);
and U4498 (N_4498,N_2327,N_3852);
nor U4499 (N_4499,N_3385,N_3839);
nand U4500 (N_4500,N_3654,N_2252);
nor U4501 (N_4501,N_3136,N_2172);
nand U4502 (N_4502,N_3178,N_3500);
and U4503 (N_4503,N_3206,N_3159);
nand U4504 (N_4504,N_2996,N_3542);
nor U4505 (N_4505,N_2466,N_3282);
nor U4506 (N_4506,N_2821,N_2846);
nand U4507 (N_4507,N_3505,N_3432);
or U4508 (N_4508,N_3701,N_3638);
or U4509 (N_4509,N_3109,N_2391);
and U4510 (N_4510,N_2346,N_3501);
or U4511 (N_4511,N_2500,N_2479);
nand U4512 (N_4512,N_3588,N_3891);
xnor U4513 (N_4513,N_2028,N_3647);
and U4514 (N_4514,N_3027,N_3298);
and U4515 (N_4515,N_2664,N_2167);
or U4516 (N_4516,N_3369,N_2945);
or U4517 (N_4517,N_3268,N_2175);
and U4518 (N_4518,N_3482,N_3895);
xnor U4519 (N_4519,N_2007,N_3280);
nand U4520 (N_4520,N_2319,N_3851);
and U4521 (N_4521,N_3348,N_2903);
and U4522 (N_4522,N_2913,N_3356);
nor U4523 (N_4523,N_2636,N_2864);
nor U4524 (N_4524,N_3131,N_3167);
nor U4525 (N_4525,N_2536,N_3389);
nand U4526 (N_4526,N_2657,N_3112);
nor U4527 (N_4527,N_2683,N_2085);
and U4528 (N_4528,N_2046,N_2484);
or U4529 (N_4529,N_3473,N_3853);
and U4530 (N_4530,N_2311,N_3456);
or U4531 (N_4531,N_2445,N_3026);
nor U4532 (N_4532,N_3513,N_2763);
nor U4533 (N_4533,N_3965,N_3585);
or U4534 (N_4534,N_3292,N_3768);
or U4535 (N_4535,N_2344,N_2115);
nor U4536 (N_4536,N_3571,N_3822);
nand U4537 (N_4537,N_3018,N_2693);
and U4538 (N_4538,N_3970,N_2439);
nand U4539 (N_4539,N_3392,N_2130);
or U4540 (N_4540,N_2048,N_2759);
and U4541 (N_4541,N_2887,N_3503);
or U4542 (N_4542,N_2430,N_2558);
nor U4543 (N_4543,N_3007,N_3689);
or U4544 (N_4544,N_2785,N_3824);
nand U4545 (N_4545,N_2050,N_2025);
or U4546 (N_4546,N_2097,N_3675);
and U4547 (N_4547,N_2460,N_2651);
xor U4548 (N_4548,N_2432,N_2393);
nand U4549 (N_4549,N_2804,N_2227);
nor U4550 (N_4550,N_2917,N_3253);
and U4551 (N_4551,N_2644,N_2817);
xor U4552 (N_4552,N_3960,N_2413);
and U4553 (N_4553,N_3955,N_2238);
nand U4554 (N_4554,N_2829,N_3881);
nand U4555 (N_4555,N_2194,N_2692);
and U4556 (N_4556,N_3067,N_2791);
or U4557 (N_4557,N_2967,N_3052);
nand U4558 (N_4558,N_3629,N_2283);
nand U4559 (N_4559,N_3296,N_3972);
and U4560 (N_4560,N_2862,N_2405);
and U4561 (N_4561,N_2721,N_3849);
and U4562 (N_4562,N_2630,N_3008);
nor U4563 (N_4563,N_3837,N_3321);
nand U4564 (N_4564,N_3202,N_2907);
nand U4565 (N_4565,N_3444,N_2417);
nor U4566 (N_4566,N_3707,N_3384);
nand U4567 (N_4567,N_2257,N_2298);
and U4568 (N_4568,N_2576,N_3772);
nand U4569 (N_4569,N_3295,N_3769);
or U4570 (N_4570,N_2957,N_2020);
nand U4571 (N_4571,N_3025,N_3750);
or U4572 (N_4572,N_2595,N_2896);
nand U4573 (N_4573,N_2879,N_3730);
nand U4574 (N_4574,N_2854,N_2927);
nor U4575 (N_4575,N_3066,N_3594);
xnor U4576 (N_4576,N_2313,N_2924);
or U4577 (N_4577,N_3528,N_2647);
nor U4578 (N_4578,N_2178,N_2400);
nand U4579 (N_4579,N_3681,N_2940);
and U4580 (N_4580,N_3390,N_3702);
nand U4581 (N_4581,N_3013,N_3089);
or U4582 (N_4582,N_3345,N_2022);
or U4583 (N_4583,N_2722,N_2299);
nor U4584 (N_4584,N_2161,N_2214);
or U4585 (N_4585,N_3679,N_3461);
or U4586 (N_4586,N_3064,N_3695);
or U4587 (N_4587,N_2157,N_2716);
and U4588 (N_4588,N_2506,N_3265);
nand U4589 (N_4589,N_2343,N_2331);
nor U4590 (N_4590,N_2519,N_3342);
nor U4591 (N_4591,N_2726,N_2805);
nor U4592 (N_4592,N_3383,N_3539);
nand U4593 (N_4593,N_2082,N_2454);
nor U4594 (N_4594,N_2411,N_3104);
nor U4595 (N_4595,N_3200,N_3147);
nor U4596 (N_4596,N_3040,N_2768);
nand U4597 (N_4597,N_2029,N_2164);
nor U4598 (N_4598,N_2604,N_2813);
nor U4599 (N_4599,N_2545,N_3697);
nand U4600 (N_4600,N_3002,N_3446);
nand U4601 (N_4601,N_3488,N_2053);
and U4602 (N_4602,N_3021,N_3826);
or U4603 (N_4603,N_3108,N_2338);
nand U4604 (N_4604,N_2438,N_3459);
and U4605 (N_4605,N_3980,N_3568);
nor U4606 (N_4606,N_2605,N_3742);
and U4607 (N_4607,N_2699,N_2649);
nand U4608 (N_4608,N_2301,N_3151);
and U4609 (N_4609,N_2199,N_3666);
and U4610 (N_4610,N_2488,N_3236);
nor U4611 (N_4611,N_3682,N_2873);
nor U4612 (N_4612,N_3030,N_2316);
nand U4613 (N_4613,N_3652,N_3835);
nand U4614 (N_4614,N_3902,N_2339);
nand U4615 (N_4615,N_2220,N_2573);
or U4616 (N_4616,N_3329,N_2533);
or U4617 (N_4617,N_2951,N_2276);
nand U4618 (N_4618,N_3286,N_3264);
and U4619 (N_4619,N_2613,N_3493);
nand U4620 (N_4620,N_2730,N_2803);
nor U4621 (N_4621,N_3180,N_2287);
nand U4622 (N_4622,N_3273,N_2935);
nand U4623 (N_4623,N_2461,N_3428);
xnor U4624 (N_4624,N_3301,N_3981);
nor U4625 (N_4625,N_2089,N_2274);
or U4626 (N_4626,N_3619,N_2608);
nor U4627 (N_4627,N_2597,N_3447);
and U4628 (N_4628,N_2371,N_2328);
xnor U4629 (N_4629,N_2471,N_3932);
or U4630 (N_4630,N_2858,N_2640);
nor U4631 (N_4631,N_2687,N_2387);
nor U4632 (N_4632,N_3720,N_2561);
nand U4633 (N_4633,N_2449,N_2929);
nand U4634 (N_4634,N_3194,N_3757);
nand U4635 (N_4635,N_2229,N_2797);
nand U4636 (N_4636,N_2165,N_3199);
and U4637 (N_4637,N_3244,N_3140);
or U4638 (N_4638,N_3439,N_3186);
nand U4639 (N_4639,N_3841,N_2978);
nand U4640 (N_4640,N_2681,N_2556);
nand U4641 (N_4641,N_3312,N_3153);
or U4642 (N_4642,N_2728,N_2711);
nor U4643 (N_4643,N_2814,N_2845);
xor U4644 (N_4644,N_3289,N_3293);
nor U4645 (N_4645,N_2977,N_3128);
nand U4646 (N_4646,N_2069,N_2769);
and U4647 (N_4647,N_3157,N_3727);
and U4648 (N_4648,N_3848,N_2018);
or U4649 (N_4649,N_2456,N_3917);
nor U4650 (N_4650,N_2989,N_2114);
nor U4651 (N_4651,N_2409,N_2451);
or U4652 (N_4652,N_2847,N_2356);
or U4653 (N_4653,N_3188,N_2330);
and U4654 (N_4654,N_3535,N_3530);
nand U4655 (N_4655,N_3892,N_2918);
nand U4656 (N_4656,N_2010,N_3250);
nand U4657 (N_4657,N_2761,N_3596);
and U4658 (N_4658,N_3357,N_3615);
and U4659 (N_4659,N_3281,N_3081);
and U4660 (N_4660,N_3905,N_2204);
nor U4661 (N_4661,N_2928,N_3398);
and U4662 (N_4662,N_3424,N_2266);
or U4663 (N_4663,N_2882,N_3782);
nor U4664 (N_4664,N_3563,N_3996);
or U4665 (N_4665,N_3745,N_3509);
nor U4666 (N_4666,N_3660,N_3228);
or U4667 (N_4667,N_3926,N_3808);
nor U4668 (N_4668,N_3729,N_3906);
xor U4669 (N_4669,N_2521,N_2039);
nand U4670 (N_4670,N_3992,N_2755);
nor U4671 (N_4671,N_2109,N_3184);
and U4672 (N_4672,N_2480,N_2323);
nand U4673 (N_4673,N_2645,N_3457);
xnor U4674 (N_4674,N_2631,N_3377);
nand U4675 (N_4675,N_3912,N_2646);
nand U4676 (N_4676,N_3603,N_3132);
or U4677 (N_4677,N_3325,N_2201);
or U4678 (N_4678,N_3450,N_3989);
and U4679 (N_4679,N_3545,N_3469);
nor U4680 (N_4680,N_2401,N_2382);
nor U4681 (N_4681,N_3406,N_2021);
or U4682 (N_4682,N_3576,N_3982);
nor U4683 (N_4683,N_2553,N_3921);
and U4684 (N_4684,N_2054,N_2307);
nand U4685 (N_4685,N_2748,N_2522);
xor U4686 (N_4686,N_2324,N_3736);
nor U4687 (N_4687,N_2916,N_3724);
nand U4688 (N_4688,N_3668,N_3333);
nand U4689 (N_4689,N_2497,N_2959);
or U4690 (N_4690,N_3005,N_2544);
nand U4691 (N_4691,N_3711,N_2770);
nor U4692 (N_4692,N_3142,N_3710);
or U4693 (N_4693,N_2653,N_2516);
nand U4694 (N_4694,N_2348,N_2459);
or U4695 (N_4695,N_3706,N_2898);
nand U4696 (N_4696,N_2598,N_3078);
nand U4697 (N_4697,N_2503,N_3948);
nor U4698 (N_4698,N_3763,N_3676);
or U4699 (N_4699,N_3332,N_3686);
nor U4700 (N_4700,N_2023,N_3448);
nand U4701 (N_4701,N_3324,N_2954);
and U4702 (N_4702,N_2407,N_3919);
and U4703 (N_4703,N_2080,N_3476);
and U4704 (N_4704,N_2125,N_2966);
nor U4705 (N_4705,N_3038,N_2120);
nor U4706 (N_4706,N_2088,N_3885);
or U4707 (N_4707,N_3767,N_2143);
nor U4708 (N_4708,N_2190,N_3114);
nand U4709 (N_4709,N_3650,N_3015);
nand U4710 (N_4710,N_3883,N_3840);
nor U4711 (N_4711,N_2603,N_2825);
nor U4712 (N_4712,N_2212,N_2305);
and U4713 (N_4713,N_2422,N_3331);
or U4714 (N_4714,N_2442,N_2091);
nand U4715 (N_4715,N_3780,N_2580);
or U4716 (N_4716,N_3088,N_2095);
and U4717 (N_4717,N_2297,N_2136);
nand U4718 (N_4718,N_3597,N_3403);
nor U4719 (N_4719,N_3141,N_3987);
or U4720 (N_4720,N_3636,N_2193);
nand U4721 (N_4721,N_2801,N_2208);
nand U4722 (N_4722,N_2796,N_3954);
xor U4723 (N_4723,N_3872,N_2739);
and U4724 (N_4724,N_2426,N_2070);
or U4725 (N_4725,N_2774,N_2177);
nor U4726 (N_4726,N_2617,N_2799);
and U4727 (N_4727,N_3744,N_2412);
nand U4728 (N_4728,N_3544,N_2173);
nor U4729 (N_4729,N_3943,N_2578);
nand U4730 (N_4730,N_3083,N_3399);
or U4731 (N_4731,N_2386,N_2040);
xnor U4732 (N_4732,N_3156,N_2446);
and U4733 (N_4733,N_3474,N_3704);
nor U4734 (N_4734,N_3788,N_3412);
nand U4735 (N_4735,N_2147,N_3314);
and U4736 (N_4736,N_2950,N_2246);
nand U4737 (N_4737,N_3320,N_2955);
or U4738 (N_4738,N_3361,N_2980);
or U4739 (N_4739,N_3278,N_3029);
nor U4740 (N_4740,N_2976,N_2474);
nand U4741 (N_4741,N_2450,N_3553);
or U4742 (N_4742,N_3251,N_3814);
nand U4743 (N_4743,N_3858,N_2601);
or U4744 (N_4744,N_2132,N_3578);
or U4745 (N_4745,N_3624,N_2765);
or U4746 (N_4746,N_3749,N_2600);
and U4747 (N_4747,N_2036,N_3516);
xor U4748 (N_4748,N_2822,N_2596);
nor U4749 (N_4749,N_3971,N_2347);
or U4750 (N_4750,N_3116,N_3634);
nand U4751 (N_4751,N_3381,N_2912);
and U4752 (N_4752,N_3118,N_3725);
nand U4753 (N_4753,N_2607,N_2877);
and U4754 (N_4754,N_3441,N_2808);
nand U4755 (N_4755,N_2701,N_3226);
nand U4756 (N_4756,N_3589,N_2884);
nor U4757 (N_4757,N_2771,N_2286);
or U4758 (N_4758,N_3413,N_3124);
and U4759 (N_4759,N_3879,N_3372);
nand U4760 (N_4760,N_2277,N_2467);
nor U4761 (N_4761,N_3036,N_2071);
nand U4762 (N_4762,N_2052,N_3643);
or U4763 (N_4763,N_2155,N_3609);
xor U4764 (N_4764,N_3304,N_2793);
nor U4765 (N_4765,N_3393,N_3161);
or U4766 (N_4766,N_3664,N_2419);
nor U4767 (N_4767,N_3612,N_2141);
nor U4768 (N_4768,N_3699,N_2572);
nand U4769 (N_4769,N_3728,N_3564);
xor U4770 (N_4770,N_3174,N_3816);
nand U4771 (N_4771,N_2329,N_2787);
nor U4772 (N_4772,N_3330,N_2183);
and U4773 (N_4773,N_3869,N_2440);
nand U4774 (N_4774,N_2308,N_2727);
nand U4775 (N_4775,N_2878,N_2181);
or U4776 (N_4776,N_3549,N_3983);
nand U4777 (N_4777,N_3929,N_3860);
and U4778 (N_4778,N_3272,N_3020);
nand U4779 (N_4779,N_2260,N_3894);
and U4780 (N_4780,N_3111,N_2263);
nor U4781 (N_4781,N_3605,N_3208);
and U4782 (N_4782,N_3173,N_2304);
nand U4783 (N_4783,N_3307,N_3809);
nand U4784 (N_4784,N_3861,N_2059);
nand U4785 (N_4785,N_2269,N_3497);
nor U4786 (N_4786,N_2893,N_3395);
or U4787 (N_4787,N_2150,N_2012);
nor U4788 (N_4788,N_3678,N_3107);
or U4789 (N_4789,N_2754,N_3988);
or U4790 (N_4790,N_3445,N_3113);
nand U4791 (N_4791,N_3338,N_2802);
or U4792 (N_4792,N_3323,N_3754);
nand U4793 (N_4793,N_2074,N_3522);
nand U4794 (N_4794,N_2535,N_2002);
nand U4795 (N_4795,N_3786,N_2892);
nor U4796 (N_4796,N_2075,N_2142);
nor U4797 (N_4797,N_2772,N_3091);
nor U4798 (N_4798,N_2550,N_3621);
nor U4799 (N_4799,N_2592,N_2314);
nor U4800 (N_4800,N_3506,N_2342);
and U4801 (N_4801,N_2947,N_2049);
nand U4802 (N_4802,N_2424,N_3586);
or U4803 (N_4803,N_2510,N_3054);
nand U4804 (N_4804,N_2033,N_2773);
nand U4805 (N_4805,N_2098,N_3092);
nand U4806 (N_4806,N_2434,N_2288);
xnor U4807 (N_4807,N_2005,N_3870);
nor U4808 (N_4808,N_3953,N_3518);
and U4809 (N_4809,N_3761,N_3050);
xnor U4810 (N_4810,N_2189,N_3420);
or U4811 (N_4811,N_3248,N_3579);
nand U4812 (N_4812,N_3130,N_2469);
or U4813 (N_4813,N_2987,N_2443);
or U4814 (N_4814,N_3033,N_2310);
or U4815 (N_4815,N_3380,N_2593);
and U4816 (N_4816,N_2932,N_2378);
nor U4817 (N_4817,N_3434,N_2226);
nor U4818 (N_4818,N_3945,N_2247);
nand U4819 (N_4819,N_3713,N_3055);
xnor U4820 (N_4820,N_2093,N_3947);
or U4821 (N_4821,N_2239,N_2974);
and U4822 (N_4822,N_2118,N_3863);
nand U4823 (N_4823,N_3267,N_3866);
or U4824 (N_4824,N_3053,N_3924);
xor U4825 (N_4825,N_2236,N_3049);
nor U4826 (N_4826,N_3031,N_2171);
nor U4827 (N_4827,N_2905,N_3144);
nand U4828 (N_4828,N_2582,N_3813);
nand U4829 (N_4829,N_2004,N_3243);
nand U4830 (N_4830,N_3254,N_2166);
or U4831 (N_4831,N_3671,N_3793);
or U4832 (N_4832,N_2490,N_2832);
nand U4833 (N_4833,N_3440,N_2560);
nand U4834 (N_4834,N_3335,N_2240);
or U4835 (N_4835,N_2192,N_2428);
nand U4836 (N_4836,N_2626,N_3137);
and U4837 (N_4837,N_2364,N_2629);
or U4838 (N_4838,N_3247,N_2292);
nand U4839 (N_4839,N_3649,N_3494);
nand U4840 (N_4840,N_2312,N_3299);
nand U4841 (N_4841,N_3019,N_3172);
or U4842 (N_4842,N_2256,N_2840);
nor U4843 (N_4843,N_2915,N_3010);
nand U4844 (N_4844,N_3998,N_3489);
and U4845 (N_4845,N_2182,N_3171);
nand U4846 (N_4846,N_2000,N_2616);
or U4847 (N_4847,N_2706,N_2960);
and U4848 (N_4848,N_2694,N_3239);
nand U4849 (N_4849,N_2734,N_3458);
or U4850 (N_4850,N_2073,N_2300);
nand U4851 (N_4851,N_3698,N_2463);
nand U4852 (N_4852,N_3270,N_3642);
or U4853 (N_4853,N_2686,N_3815);
nand U4854 (N_4854,N_2588,N_2698);
nand U4855 (N_4855,N_2546,N_2783);
nor U4856 (N_4856,N_2691,N_2751);
or U4857 (N_4857,N_2335,N_2904);
nor U4858 (N_4858,N_3556,N_3884);
nor U4859 (N_4859,N_2637,N_2811);
nor U4860 (N_4860,N_2848,N_3045);
or U4861 (N_4861,N_3940,N_2309);
or U4862 (N_4862,N_3764,N_3037);
nand U4863 (N_4863,N_3531,N_2704);
nand U4864 (N_4864,N_3261,N_3150);
nor U4865 (N_4865,N_3575,N_3887);
and U4866 (N_4866,N_2380,N_3674);
nor U4867 (N_4867,N_2740,N_3028);
nand U4868 (N_4868,N_3785,N_3691);
nor U4869 (N_4869,N_3608,N_3778);
and U4870 (N_4870,N_3452,N_2676);
nor U4871 (N_4871,N_3376,N_3523);
nor U4872 (N_4872,N_3957,N_2890);
xor U4873 (N_4873,N_2586,N_2570);
or U4874 (N_4874,N_2752,N_2505);
nor U4875 (N_4875,N_2881,N_3386);
nand U4876 (N_4876,N_2372,N_3433);
xor U4877 (N_4877,N_3635,N_3185);
or U4878 (N_4878,N_2807,N_2981);
nand U4879 (N_4879,N_2703,N_3397);
nor U4880 (N_4880,N_2620,N_3577);
or U4881 (N_4881,N_2760,N_3197);
nand U4882 (N_4882,N_2427,N_2816);
nand U4883 (N_4883,N_3716,N_2874);
nor U4884 (N_4884,N_2363,N_3418);
or U4885 (N_4885,N_2725,N_3336);
nor U4886 (N_4886,N_2373,N_2656);
or U4887 (N_4887,N_3538,N_3626);
nor U4888 (N_4888,N_2865,N_3963);
and U4889 (N_4889,N_2714,N_2290);
and U4890 (N_4890,N_3262,N_3602);
nand U4891 (N_4891,N_3843,N_2361);
nand U4892 (N_4892,N_3415,N_2008);
nand U4893 (N_4893,N_3562,N_2612);
nor U4894 (N_4894,N_2820,N_2215);
and U4895 (N_4895,N_2047,N_2665);
nand U4896 (N_4896,N_3915,N_2537);
and U4897 (N_4897,N_2853,N_2244);
or U4898 (N_4898,N_3240,N_3899);
and U4899 (N_4899,N_3507,N_3685);
nor U4900 (N_4900,N_2511,N_2958);
or U4901 (N_4901,N_3485,N_3617);
nor U4902 (N_4902,N_2909,N_2562);
and U4903 (N_4903,N_2715,N_2222);
or U4904 (N_4904,N_3752,N_2249);
or U4905 (N_4905,N_3723,N_2121);
and U4906 (N_4906,N_3193,N_2476);
nor U4907 (N_4907,N_3646,N_3120);
and U4908 (N_4908,N_2746,N_2775);
nand U4909 (N_4909,N_3510,N_2707);
and U4910 (N_4910,N_3550,N_3363);
and U4911 (N_4911,N_3527,N_2009);
or U4912 (N_4912,N_2839,N_2495);
or U4913 (N_4913,N_3801,N_2529);
nor U4914 (N_4914,N_2690,N_3525);
nand U4915 (N_4915,N_3429,N_3442);
and U4916 (N_4916,N_3913,N_3443);
nand U4917 (N_4917,N_2914,N_3812);
or U4918 (N_4918,N_3168,N_3215);
nand U4919 (N_4919,N_3388,N_2609);
or U4920 (N_4920,N_2889,N_2366);
nand U4921 (N_4921,N_2983,N_2303);
nand U4922 (N_4922,N_3071,N_3551);
nand U4923 (N_4923,N_3145,N_2123);
nand U4924 (N_4924,N_3216,N_2254);
and U4925 (N_4925,N_3146,N_3607);
nor U4926 (N_4926,N_2478,N_2122);
xnor U4927 (N_4927,N_2923,N_2203);
nand U4928 (N_4928,N_3557,N_3478);
or U4929 (N_4929,N_3657,N_2464);
nand U4930 (N_4930,N_2577,N_3090);
nand U4931 (N_4931,N_3337,N_2320);
and U4932 (N_4932,N_3590,N_3687);
nand U4933 (N_4933,N_3526,N_3310);
or U4934 (N_4934,N_3343,N_2253);
and U4935 (N_4935,N_2037,N_3230);
and U4936 (N_4936,N_3401,N_3726);
or U4937 (N_4937,N_2206,N_2289);
nor U4938 (N_4938,N_3315,N_3044);
and U4939 (N_4939,N_2815,N_2369);
nand U4940 (N_4940,N_2285,N_2083);
and U4941 (N_4941,N_3222,N_3832);
nand U4942 (N_4942,N_3606,N_2938);
nand U4943 (N_4943,N_3584,N_3051);
nor U4944 (N_4944,N_3258,N_3762);
nor U4945 (N_4945,N_2306,N_3799);
nand U4946 (N_4946,N_3529,N_2170);
and U4947 (N_4947,N_2590,N_3287);
or U4948 (N_4948,N_3967,N_2732);
or U4949 (N_4949,N_2195,N_2552);
nor U4950 (N_4950,N_3865,N_3519);
and U4951 (N_4951,N_2736,N_3569);
nand U4952 (N_4952,N_2998,N_2943);
or U4953 (N_4953,N_3269,N_2072);
nor U4954 (N_4954,N_2359,N_2899);
or U4955 (N_4955,N_3991,N_2398);
or U4956 (N_4956,N_2295,N_2660);
nor U4957 (N_4957,N_2377,N_2278);
or U4958 (N_4958,N_2196,N_2055);
or U4959 (N_4959,N_2999,N_3864);
nor U4960 (N_4960,N_2672,N_2702);
xor U4961 (N_4961,N_2628,N_2145);
or U4962 (N_4962,N_3875,N_3949);
and U4963 (N_4963,N_2946,N_3245);
nor U4964 (N_4964,N_2680,N_3876);
nand U4965 (N_4965,N_3661,N_3427);
and U4966 (N_4966,N_2251,N_3829);
or U4967 (N_4967,N_2392,N_2187);
or U4968 (N_4968,N_2043,N_3135);
or U4969 (N_4969,N_3405,N_2013);
xor U4970 (N_4970,N_2517,N_2352);
and U4971 (N_4971,N_2555,N_2436);
or U4972 (N_4972,N_2112,N_3127);
and U4973 (N_4973,N_3787,N_2105);
nand U4974 (N_4974,N_3455,N_3514);
nor U4975 (N_4975,N_2991,N_2837);
nand U4976 (N_4976,N_3680,N_2780);
and U4977 (N_4977,N_2541,N_3004);
nor U4978 (N_4978,N_3774,N_2969);
or U4979 (N_4979,N_3175,N_3910);
and U4980 (N_4980,N_3303,N_2756);
and U4981 (N_4981,N_3134,N_2618);
xor U4982 (N_4982,N_3889,N_3959);
nor U4983 (N_4983,N_2350,N_2379);
or U4984 (N_4984,N_3190,N_2942);
or U4985 (N_4985,N_2504,N_2886);
nor U4986 (N_4986,N_2188,N_2615);
nor U4987 (N_4987,N_2219,N_3079);
and U4988 (N_4988,N_3279,N_3777);
nor U4989 (N_4989,N_2764,N_2992);
nand U4990 (N_4990,N_2606,N_2090);
nand U4991 (N_4991,N_3665,N_3207);
and U4992 (N_4992,N_2465,N_3639);
or U4993 (N_4993,N_3011,N_3904);
nand U4994 (N_4994,N_2176,N_3558);
nor U4995 (N_4995,N_3451,N_3855);
nor U4996 (N_4996,N_2741,N_3213);
nand U4997 (N_4997,N_2179,N_2654);
and U4998 (N_4998,N_2670,N_2548);
nor U4999 (N_4999,N_2695,N_3520);
and U5000 (N_5000,N_3716,N_3427);
or U5001 (N_5001,N_2463,N_2453);
and U5002 (N_5002,N_3128,N_3325);
or U5003 (N_5003,N_3708,N_3472);
or U5004 (N_5004,N_3148,N_2028);
or U5005 (N_5005,N_2497,N_2473);
nor U5006 (N_5006,N_3081,N_2120);
nor U5007 (N_5007,N_3741,N_3757);
nor U5008 (N_5008,N_3554,N_2821);
and U5009 (N_5009,N_3025,N_2025);
or U5010 (N_5010,N_3709,N_2914);
nor U5011 (N_5011,N_2647,N_3818);
and U5012 (N_5012,N_2553,N_2260);
nor U5013 (N_5013,N_3908,N_2726);
nor U5014 (N_5014,N_3073,N_3111);
or U5015 (N_5015,N_2157,N_2239);
or U5016 (N_5016,N_2497,N_2195);
nor U5017 (N_5017,N_3620,N_2066);
nand U5018 (N_5018,N_2596,N_3096);
or U5019 (N_5019,N_2967,N_3187);
nand U5020 (N_5020,N_2456,N_3059);
or U5021 (N_5021,N_2469,N_3591);
and U5022 (N_5022,N_2473,N_2165);
nor U5023 (N_5023,N_2762,N_3195);
nor U5024 (N_5024,N_3992,N_2791);
nor U5025 (N_5025,N_2805,N_3295);
or U5026 (N_5026,N_2106,N_2180);
and U5027 (N_5027,N_3706,N_2127);
and U5028 (N_5028,N_3730,N_3740);
nand U5029 (N_5029,N_3544,N_2073);
and U5030 (N_5030,N_2277,N_3540);
and U5031 (N_5031,N_3368,N_3366);
and U5032 (N_5032,N_3496,N_2786);
and U5033 (N_5033,N_3365,N_3537);
or U5034 (N_5034,N_3885,N_3248);
nand U5035 (N_5035,N_3728,N_3890);
nand U5036 (N_5036,N_2561,N_2574);
nor U5037 (N_5037,N_3399,N_2855);
nor U5038 (N_5038,N_3141,N_3326);
nor U5039 (N_5039,N_2238,N_2010);
nand U5040 (N_5040,N_2294,N_3503);
or U5041 (N_5041,N_3843,N_3748);
nand U5042 (N_5042,N_3982,N_2188);
nor U5043 (N_5043,N_3987,N_2070);
nor U5044 (N_5044,N_2629,N_3350);
nand U5045 (N_5045,N_2163,N_3622);
and U5046 (N_5046,N_2754,N_3775);
nor U5047 (N_5047,N_2332,N_2400);
nor U5048 (N_5048,N_2272,N_2639);
or U5049 (N_5049,N_2060,N_3906);
nand U5050 (N_5050,N_3653,N_2677);
nor U5051 (N_5051,N_3802,N_3106);
and U5052 (N_5052,N_3754,N_3705);
or U5053 (N_5053,N_2377,N_2491);
or U5054 (N_5054,N_2055,N_3987);
and U5055 (N_5055,N_2121,N_2211);
nor U5056 (N_5056,N_2001,N_3812);
or U5057 (N_5057,N_3376,N_3831);
nor U5058 (N_5058,N_2085,N_3488);
or U5059 (N_5059,N_3588,N_2770);
nor U5060 (N_5060,N_3777,N_3482);
or U5061 (N_5061,N_3626,N_3078);
or U5062 (N_5062,N_3387,N_2403);
nand U5063 (N_5063,N_3626,N_3175);
nor U5064 (N_5064,N_3327,N_2571);
nand U5065 (N_5065,N_2827,N_3687);
and U5066 (N_5066,N_2103,N_3607);
and U5067 (N_5067,N_2219,N_3772);
or U5068 (N_5068,N_3466,N_2425);
nand U5069 (N_5069,N_2627,N_3444);
nor U5070 (N_5070,N_3493,N_2923);
xor U5071 (N_5071,N_2593,N_2144);
nand U5072 (N_5072,N_2254,N_3865);
or U5073 (N_5073,N_2144,N_2503);
and U5074 (N_5074,N_2077,N_3341);
or U5075 (N_5075,N_3733,N_3943);
and U5076 (N_5076,N_2107,N_2177);
or U5077 (N_5077,N_3948,N_2472);
nor U5078 (N_5078,N_3773,N_2625);
and U5079 (N_5079,N_2496,N_2291);
nand U5080 (N_5080,N_2958,N_3579);
or U5081 (N_5081,N_2759,N_3049);
and U5082 (N_5082,N_2379,N_2869);
and U5083 (N_5083,N_2691,N_2603);
nand U5084 (N_5084,N_2874,N_2307);
or U5085 (N_5085,N_2502,N_2782);
nand U5086 (N_5086,N_2118,N_3848);
nor U5087 (N_5087,N_3424,N_2003);
nor U5088 (N_5088,N_2825,N_2281);
and U5089 (N_5089,N_3118,N_3325);
or U5090 (N_5090,N_3457,N_2401);
or U5091 (N_5091,N_2994,N_2660);
or U5092 (N_5092,N_3709,N_3763);
nor U5093 (N_5093,N_3967,N_2742);
xor U5094 (N_5094,N_3693,N_2583);
nor U5095 (N_5095,N_3146,N_3855);
and U5096 (N_5096,N_2041,N_2079);
nand U5097 (N_5097,N_3695,N_2532);
or U5098 (N_5098,N_3806,N_2348);
or U5099 (N_5099,N_3669,N_3008);
nand U5100 (N_5100,N_3012,N_3274);
or U5101 (N_5101,N_2648,N_2661);
nor U5102 (N_5102,N_3220,N_2341);
or U5103 (N_5103,N_3981,N_3870);
or U5104 (N_5104,N_2334,N_2192);
or U5105 (N_5105,N_2212,N_3566);
nand U5106 (N_5106,N_3682,N_3356);
nor U5107 (N_5107,N_2905,N_2827);
and U5108 (N_5108,N_3889,N_2357);
nand U5109 (N_5109,N_3427,N_3068);
or U5110 (N_5110,N_3355,N_3987);
nor U5111 (N_5111,N_2302,N_3869);
or U5112 (N_5112,N_2714,N_2448);
or U5113 (N_5113,N_3543,N_2148);
or U5114 (N_5114,N_2851,N_3986);
and U5115 (N_5115,N_3856,N_2294);
and U5116 (N_5116,N_3424,N_3856);
or U5117 (N_5117,N_2903,N_3462);
nor U5118 (N_5118,N_3275,N_2272);
or U5119 (N_5119,N_2441,N_3023);
nor U5120 (N_5120,N_3217,N_2577);
and U5121 (N_5121,N_3180,N_2688);
and U5122 (N_5122,N_3378,N_2294);
or U5123 (N_5123,N_3819,N_3347);
nand U5124 (N_5124,N_2050,N_3367);
nor U5125 (N_5125,N_2419,N_3558);
or U5126 (N_5126,N_3986,N_2558);
and U5127 (N_5127,N_2927,N_2314);
and U5128 (N_5128,N_3847,N_3682);
nand U5129 (N_5129,N_3534,N_3704);
or U5130 (N_5130,N_2262,N_3190);
and U5131 (N_5131,N_3472,N_3762);
nand U5132 (N_5132,N_2342,N_2987);
nor U5133 (N_5133,N_3469,N_3870);
and U5134 (N_5134,N_2319,N_2440);
nand U5135 (N_5135,N_3346,N_3766);
and U5136 (N_5136,N_3714,N_2505);
or U5137 (N_5137,N_3036,N_2093);
nor U5138 (N_5138,N_3931,N_3542);
nor U5139 (N_5139,N_2161,N_3336);
nor U5140 (N_5140,N_3019,N_2265);
nor U5141 (N_5141,N_3517,N_2805);
and U5142 (N_5142,N_3879,N_3633);
or U5143 (N_5143,N_2355,N_3689);
xnor U5144 (N_5144,N_3476,N_2174);
or U5145 (N_5145,N_2523,N_2433);
nor U5146 (N_5146,N_2524,N_2964);
and U5147 (N_5147,N_2756,N_2590);
and U5148 (N_5148,N_3907,N_3253);
nor U5149 (N_5149,N_2349,N_3628);
xor U5150 (N_5150,N_3903,N_3549);
or U5151 (N_5151,N_3584,N_3809);
or U5152 (N_5152,N_2420,N_3726);
nor U5153 (N_5153,N_3109,N_2780);
nand U5154 (N_5154,N_3269,N_2759);
nor U5155 (N_5155,N_2494,N_3338);
or U5156 (N_5156,N_2399,N_3773);
nand U5157 (N_5157,N_3077,N_3865);
nand U5158 (N_5158,N_3211,N_2845);
or U5159 (N_5159,N_3913,N_2127);
nand U5160 (N_5160,N_2774,N_2415);
or U5161 (N_5161,N_3128,N_3307);
or U5162 (N_5162,N_2766,N_2040);
and U5163 (N_5163,N_2110,N_3745);
nor U5164 (N_5164,N_2895,N_3324);
and U5165 (N_5165,N_3642,N_2563);
and U5166 (N_5166,N_3331,N_2752);
and U5167 (N_5167,N_3471,N_2929);
or U5168 (N_5168,N_2880,N_2515);
and U5169 (N_5169,N_2457,N_3923);
nor U5170 (N_5170,N_3383,N_2213);
or U5171 (N_5171,N_2525,N_2534);
or U5172 (N_5172,N_2975,N_3668);
xor U5173 (N_5173,N_3630,N_2020);
or U5174 (N_5174,N_2231,N_3601);
nand U5175 (N_5175,N_2052,N_2849);
or U5176 (N_5176,N_2381,N_3973);
nand U5177 (N_5177,N_2017,N_3163);
nand U5178 (N_5178,N_3222,N_2892);
and U5179 (N_5179,N_3339,N_3964);
or U5180 (N_5180,N_2933,N_3766);
and U5181 (N_5181,N_3880,N_3241);
nand U5182 (N_5182,N_3056,N_2965);
nand U5183 (N_5183,N_3280,N_3822);
or U5184 (N_5184,N_3954,N_2983);
and U5185 (N_5185,N_3990,N_3179);
nand U5186 (N_5186,N_2938,N_2998);
and U5187 (N_5187,N_2540,N_2701);
or U5188 (N_5188,N_2719,N_2642);
or U5189 (N_5189,N_3339,N_3967);
nand U5190 (N_5190,N_3150,N_2395);
nand U5191 (N_5191,N_3013,N_2745);
or U5192 (N_5192,N_2761,N_2090);
nand U5193 (N_5193,N_2376,N_3746);
nand U5194 (N_5194,N_2361,N_2798);
and U5195 (N_5195,N_3716,N_2644);
and U5196 (N_5196,N_3320,N_3980);
or U5197 (N_5197,N_2028,N_3406);
and U5198 (N_5198,N_3308,N_3943);
and U5199 (N_5199,N_2155,N_2942);
and U5200 (N_5200,N_3575,N_2512);
nor U5201 (N_5201,N_3755,N_2794);
nand U5202 (N_5202,N_2775,N_3601);
nand U5203 (N_5203,N_3864,N_3049);
and U5204 (N_5204,N_2243,N_2873);
nand U5205 (N_5205,N_3990,N_3560);
nand U5206 (N_5206,N_2529,N_3479);
nor U5207 (N_5207,N_3753,N_2102);
nand U5208 (N_5208,N_3489,N_3342);
or U5209 (N_5209,N_3342,N_2183);
or U5210 (N_5210,N_2876,N_2753);
and U5211 (N_5211,N_2412,N_2098);
and U5212 (N_5212,N_2104,N_2846);
or U5213 (N_5213,N_2793,N_3884);
nand U5214 (N_5214,N_2206,N_3835);
or U5215 (N_5215,N_2670,N_2459);
and U5216 (N_5216,N_3223,N_3949);
nand U5217 (N_5217,N_3950,N_2272);
nand U5218 (N_5218,N_3061,N_2194);
nand U5219 (N_5219,N_2870,N_3640);
and U5220 (N_5220,N_2141,N_2893);
and U5221 (N_5221,N_3836,N_3964);
nor U5222 (N_5222,N_2834,N_2087);
nand U5223 (N_5223,N_2994,N_3908);
nand U5224 (N_5224,N_3390,N_3360);
or U5225 (N_5225,N_2025,N_3079);
or U5226 (N_5226,N_2101,N_3115);
nand U5227 (N_5227,N_2260,N_2093);
nor U5228 (N_5228,N_2995,N_3316);
or U5229 (N_5229,N_3931,N_2381);
or U5230 (N_5230,N_3027,N_2475);
or U5231 (N_5231,N_3020,N_3203);
and U5232 (N_5232,N_2277,N_3886);
nor U5233 (N_5233,N_2477,N_3181);
and U5234 (N_5234,N_2336,N_3999);
or U5235 (N_5235,N_3249,N_2445);
or U5236 (N_5236,N_3369,N_2996);
and U5237 (N_5237,N_2841,N_3744);
nand U5238 (N_5238,N_2047,N_3476);
or U5239 (N_5239,N_3201,N_2815);
and U5240 (N_5240,N_3376,N_2204);
nor U5241 (N_5241,N_2653,N_2590);
xnor U5242 (N_5242,N_2018,N_2517);
or U5243 (N_5243,N_2497,N_3719);
nand U5244 (N_5244,N_2842,N_2975);
and U5245 (N_5245,N_2712,N_3801);
nor U5246 (N_5246,N_3588,N_2214);
nor U5247 (N_5247,N_2803,N_3936);
or U5248 (N_5248,N_2064,N_2157);
nor U5249 (N_5249,N_3862,N_3827);
nor U5250 (N_5250,N_3889,N_2939);
and U5251 (N_5251,N_2086,N_2737);
and U5252 (N_5252,N_2832,N_2496);
nor U5253 (N_5253,N_2102,N_2636);
nand U5254 (N_5254,N_3089,N_3334);
nor U5255 (N_5255,N_3160,N_3300);
nand U5256 (N_5256,N_3089,N_2344);
and U5257 (N_5257,N_3389,N_3470);
nor U5258 (N_5258,N_2932,N_3334);
nor U5259 (N_5259,N_3010,N_3282);
nor U5260 (N_5260,N_3564,N_3848);
nand U5261 (N_5261,N_3599,N_2685);
xnor U5262 (N_5262,N_3849,N_2622);
and U5263 (N_5263,N_2750,N_2774);
or U5264 (N_5264,N_3412,N_3772);
nand U5265 (N_5265,N_2377,N_2368);
nand U5266 (N_5266,N_2186,N_2888);
xnor U5267 (N_5267,N_2330,N_2535);
nand U5268 (N_5268,N_2262,N_3650);
nor U5269 (N_5269,N_2772,N_3029);
nor U5270 (N_5270,N_2791,N_3646);
or U5271 (N_5271,N_3929,N_3146);
or U5272 (N_5272,N_2302,N_2764);
nor U5273 (N_5273,N_3100,N_3599);
and U5274 (N_5274,N_2356,N_3378);
and U5275 (N_5275,N_3630,N_2625);
and U5276 (N_5276,N_3272,N_3625);
or U5277 (N_5277,N_2078,N_2769);
or U5278 (N_5278,N_3644,N_3856);
xor U5279 (N_5279,N_2986,N_2267);
nor U5280 (N_5280,N_2597,N_3949);
nand U5281 (N_5281,N_2592,N_2983);
nand U5282 (N_5282,N_3737,N_3763);
xor U5283 (N_5283,N_2916,N_2661);
nor U5284 (N_5284,N_3355,N_3314);
xnor U5285 (N_5285,N_3691,N_2307);
and U5286 (N_5286,N_2083,N_3932);
or U5287 (N_5287,N_3936,N_3163);
xor U5288 (N_5288,N_3253,N_2668);
nor U5289 (N_5289,N_3836,N_2396);
and U5290 (N_5290,N_2247,N_2365);
nor U5291 (N_5291,N_2320,N_2736);
nand U5292 (N_5292,N_3985,N_3550);
and U5293 (N_5293,N_3037,N_2318);
nor U5294 (N_5294,N_2714,N_2338);
nor U5295 (N_5295,N_3983,N_2287);
nand U5296 (N_5296,N_3548,N_3677);
nor U5297 (N_5297,N_2156,N_3448);
or U5298 (N_5298,N_2779,N_2774);
or U5299 (N_5299,N_2069,N_3589);
nand U5300 (N_5300,N_3969,N_3206);
or U5301 (N_5301,N_2767,N_2377);
and U5302 (N_5302,N_2157,N_3932);
and U5303 (N_5303,N_3255,N_3151);
nand U5304 (N_5304,N_2738,N_2909);
nand U5305 (N_5305,N_3051,N_3019);
nand U5306 (N_5306,N_2683,N_2709);
nand U5307 (N_5307,N_3102,N_3174);
nor U5308 (N_5308,N_3440,N_3793);
nor U5309 (N_5309,N_2210,N_3527);
or U5310 (N_5310,N_2826,N_2338);
nand U5311 (N_5311,N_3525,N_2490);
and U5312 (N_5312,N_2974,N_2741);
or U5313 (N_5313,N_3030,N_2885);
and U5314 (N_5314,N_3140,N_3059);
or U5315 (N_5315,N_3629,N_3139);
xor U5316 (N_5316,N_3099,N_2615);
nand U5317 (N_5317,N_3709,N_2080);
nand U5318 (N_5318,N_3100,N_2369);
nand U5319 (N_5319,N_3032,N_3205);
or U5320 (N_5320,N_3761,N_2354);
nor U5321 (N_5321,N_2762,N_3216);
nand U5322 (N_5322,N_2043,N_3286);
nand U5323 (N_5323,N_3232,N_3719);
or U5324 (N_5324,N_2983,N_2115);
and U5325 (N_5325,N_2536,N_2063);
nand U5326 (N_5326,N_2059,N_3636);
nor U5327 (N_5327,N_3957,N_2128);
xor U5328 (N_5328,N_3084,N_3200);
nor U5329 (N_5329,N_3017,N_2345);
nand U5330 (N_5330,N_2919,N_3465);
nor U5331 (N_5331,N_3921,N_2736);
nand U5332 (N_5332,N_3301,N_2453);
nand U5333 (N_5333,N_2501,N_3001);
or U5334 (N_5334,N_3502,N_2616);
nand U5335 (N_5335,N_2736,N_2882);
xnor U5336 (N_5336,N_2824,N_3792);
or U5337 (N_5337,N_2742,N_2531);
or U5338 (N_5338,N_2827,N_2372);
or U5339 (N_5339,N_3668,N_3783);
or U5340 (N_5340,N_3995,N_3846);
nor U5341 (N_5341,N_2979,N_3044);
or U5342 (N_5342,N_3251,N_2312);
nor U5343 (N_5343,N_2222,N_2052);
nand U5344 (N_5344,N_2847,N_2276);
nor U5345 (N_5345,N_3922,N_3354);
nor U5346 (N_5346,N_2309,N_3729);
and U5347 (N_5347,N_3819,N_3006);
and U5348 (N_5348,N_3787,N_3124);
xor U5349 (N_5349,N_2311,N_2285);
and U5350 (N_5350,N_3410,N_3382);
nor U5351 (N_5351,N_3431,N_3728);
or U5352 (N_5352,N_3235,N_3384);
and U5353 (N_5353,N_3545,N_2940);
or U5354 (N_5354,N_2200,N_2027);
nor U5355 (N_5355,N_2882,N_3542);
or U5356 (N_5356,N_3114,N_3504);
nor U5357 (N_5357,N_2777,N_3848);
or U5358 (N_5358,N_2378,N_3798);
nor U5359 (N_5359,N_3168,N_3828);
and U5360 (N_5360,N_2985,N_2089);
nor U5361 (N_5361,N_3958,N_2884);
or U5362 (N_5362,N_3816,N_2309);
or U5363 (N_5363,N_2532,N_2261);
nor U5364 (N_5364,N_3057,N_3276);
or U5365 (N_5365,N_3679,N_3419);
or U5366 (N_5366,N_3239,N_2395);
or U5367 (N_5367,N_2263,N_3699);
or U5368 (N_5368,N_2780,N_2493);
nand U5369 (N_5369,N_2085,N_2160);
xnor U5370 (N_5370,N_2808,N_3134);
or U5371 (N_5371,N_2525,N_2887);
nand U5372 (N_5372,N_2241,N_2499);
and U5373 (N_5373,N_3346,N_2258);
nor U5374 (N_5374,N_2220,N_3989);
or U5375 (N_5375,N_2560,N_3662);
nand U5376 (N_5376,N_3550,N_2760);
and U5377 (N_5377,N_2375,N_3367);
or U5378 (N_5378,N_3831,N_2793);
nor U5379 (N_5379,N_2346,N_3299);
nand U5380 (N_5380,N_2855,N_2712);
or U5381 (N_5381,N_3743,N_3084);
nand U5382 (N_5382,N_3309,N_3228);
and U5383 (N_5383,N_3304,N_2257);
nor U5384 (N_5384,N_2242,N_3293);
or U5385 (N_5385,N_2048,N_3906);
and U5386 (N_5386,N_3344,N_3997);
nor U5387 (N_5387,N_2363,N_2497);
or U5388 (N_5388,N_2760,N_2950);
nor U5389 (N_5389,N_3067,N_3217);
or U5390 (N_5390,N_2744,N_2894);
or U5391 (N_5391,N_3842,N_2683);
nor U5392 (N_5392,N_3831,N_3250);
and U5393 (N_5393,N_2764,N_2554);
nor U5394 (N_5394,N_3671,N_2717);
nor U5395 (N_5395,N_3615,N_3424);
nor U5396 (N_5396,N_3737,N_3905);
nor U5397 (N_5397,N_3748,N_3682);
and U5398 (N_5398,N_3945,N_3109);
and U5399 (N_5399,N_3175,N_3918);
or U5400 (N_5400,N_2026,N_2935);
and U5401 (N_5401,N_3311,N_3090);
and U5402 (N_5402,N_2105,N_2605);
and U5403 (N_5403,N_3083,N_3275);
nor U5404 (N_5404,N_3828,N_3485);
or U5405 (N_5405,N_2723,N_3053);
or U5406 (N_5406,N_3545,N_3370);
or U5407 (N_5407,N_2199,N_2716);
or U5408 (N_5408,N_2779,N_2105);
or U5409 (N_5409,N_2207,N_2588);
nor U5410 (N_5410,N_3991,N_3589);
nand U5411 (N_5411,N_3573,N_2493);
nand U5412 (N_5412,N_3060,N_3947);
nor U5413 (N_5413,N_3942,N_2952);
and U5414 (N_5414,N_2050,N_2510);
and U5415 (N_5415,N_2925,N_3803);
nand U5416 (N_5416,N_3049,N_3836);
and U5417 (N_5417,N_3720,N_2504);
nand U5418 (N_5418,N_2172,N_2549);
or U5419 (N_5419,N_2015,N_3052);
nand U5420 (N_5420,N_3283,N_3511);
nor U5421 (N_5421,N_3401,N_3122);
and U5422 (N_5422,N_2339,N_2985);
nand U5423 (N_5423,N_3938,N_3406);
nand U5424 (N_5424,N_2166,N_3441);
nor U5425 (N_5425,N_3842,N_3332);
xor U5426 (N_5426,N_2824,N_3074);
nand U5427 (N_5427,N_3381,N_3980);
nand U5428 (N_5428,N_2787,N_3227);
or U5429 (N_5429,N_3044,N_3623);
and U5430 (N_5430,N_2001,N_2335);
nand U5431 (N_5431,N_3806,N_2672);
nor U5432 (N_5432,N_3040,N_2140);
nand U5433 (N_5433,N_3304,N_2989);
nor U5434 (N_5434,N_2080,N_3481);
and U5435 (N_5435,N_2211,N_3171);
nand U5436 (N_5436,N_3301,N_3594);
nor U5437 (N_5437,N_3264,N_2668);
or U5438 (N_5438,N_3992,N_2855);
nand U5439 (N_5439,N_3990,N_2419);
and U5440 (N_5440,N_3199,N_3850);
or U5441 (N_5441,N_3619,N_2436);
and U5442 (N_5442,N_3817,N_3520);
nand U5443 (N_5443,N_2390,N_2821);
or U5444 (N_5444,N_3752,N_2575);
nand U5445 (N_5445,N_2827,N_2343);
and U5446 (N_5446,N_2686,N_3997);
xor U5447 (N_5447,N_3794,N_3831);
or U5448 (N_5448,N_2956,N_2678);
and U5449 (N_5449,N_3775,N_3458);
nand U5450 (N_5450,N_3639,N_2536);
nor U5451 (N_5451,N_3311,N_2919);
nand U5452 (N_5452,N_2308,N_2969);
nand U5453 (N_5453,N_2373,N_2545);
or U5454 (N_5454,N_2976,N_3354);
or U5455 (N_5455,N_3544,N_3493);
nand U5456 (N_5456,N_2329,N_3168);
nand U5457 (N_5457,N_2708,N_3790);
nor U5458 (N_5458,N_3269,N_2422);
or U5459 (N_5459,N_2294,N_2255);
nand U5460 (N_5460,N_3705,N_3659);
and U5461 (N_5461,N_2068,N_3191);
nor U5462 (N_5462,N_3040,N_2139);
nand U5463 (N_5463,N_3873,N_3542);
or U5464 (N_5464,N_2908,N_2821);
nor U5465 (N_5465,N_2199,N_3405);
nand U5466 (N_5466,N_2585,N_3438);
and U5467 (N_5467,N_3255,N_3179);
or U5468 (N_5468,N_3141,N_2866);
and U5469 (N_5469,N_3087,N_2125);
nand U5470 (N_5470,N_2786,N_2861);
or U5471 (N_5471,N_2022,N_3561);
or U5472 (N_5472,N_3859,N_2249);
nand U5473 (N_5473,N_3110,N_2670);
nor U5474 (N_5474,N_3196,N_2192);
nor U5475 (N_5475,N_3313,N_2591);
and U5476 (N_5476,N_2043,N_2596);
and U5477 (N_5477,N_2754,N_3503);
and U5478 (N_5478,N_3804,N_3872);
or U5479 (N_5479,N_2750,N_2522);
nor U5480 (N_5480,N_3114,N_3971);
and U5481 (N_5481,N_3315,N_2040);
xor U5482 (N_5482,N_3248,N_2901);
nor U5483 (N_5483,N_2292,N_2649);
nor U5484 (N_5484,N_3674,N_3849);
nand U5485 (N_5485,N_2201,N_3953);
nor U5486 (N_5486,N_2648,N_3421);
or U5487 (N_5487,N_3860,N_3217);
nand U5488 (N_5488,N_2444,N_2845);
nor U5489 (N_5489,N_3573,N_2194);
nor U5490 (N_5490,N_3816,N_3586);
and U5491 (N_5491,N_2559,N_2509);
nand U5492 (N_5492,N_3327,N_2953);
and U5493 (N_5493,N_2598,N_2832);
nor U5494 (N_5494,N_2875,N_2688);
and U5495 (N_5495,N_2237,N_2438);
nor U5496 (N_5496,N_2268,N_2203);
nor U5497 (N_5497,N_2919,N_2321);
or U5498 (N_5498,N_2402,N_2787);
nor U5499 (N_5499,N_3372,N_3838);
or U5500 (N_5500,N_2241,N_2083);
or U5501 (N_5501,N_2092,N_3850);
nand U5502 (N_5502,N_3740,N_3211);
nand U5503 (N_5503,N_3324,N_3959);
or U5504 (N_5504,N_2935,N_3139);
nor U5505 (N_5505,N_2186,N_2796);
nor U5506 (N_5506,N_3258,N_2140);
nor U5507 (N_5507,N_3958,N_2668);
or U5508 (N_5508,N_3790,N_2955);
and U5509 (N_5509,N_2747,N_3243);
nand U5510 (N_5510,N_2803,N_2223);
and U5511 (N_5511,N_2884,N_3300);
nand U5512 (N_5512,N_3660,N_2302);
or U5513 (N_5513,N_3133,N_2504);
or U5514 (N_5514,N_2308,N_3482);
xnor U5515 (N_5515,N_2955,N_3645);
or U5516 (N_5516,N_2956,N_3623);
and U5517 (N_5517,N_2109,N_3751);
nor U5518 (N_5518,N_3883,N_2701);
nor U5519 (N_5519,N_3993,N_3381);
nand U5520 (N_5520,N_2073,N_2517);
or U5521 (N_5521,N_3348,N_3878);
and U5522 (N_5522,N_2037,N_2761);
and U5523 (N_5523,N_2972,N_3320);
nor U5524 (N_5524,N_3331,N_2070);
nor U5525 (N_5525,N_2782,N_3094);
nor U5526 (N_5526,N_2816,N_2868);
and U5527 (N_5527,N_3514,N_2905);
and U5528 (N_5528,N_2428,N_3257);
nand U5529 (N_5529,N_2278,N_2260);
nor U5530 (N_5530,N_2434,N_2829);
nor U5531 (N_5531,N_2264,N_2874);
nand U5532 (N_5532,N_2616,N_3702);
or U5533 (N_5533,N_2250,N_2144);
nand U5534 (N_5534,N_3306,N_2510);
and U5535 (N_5535,N_2376,N_3801);
and U5536 (N_5536,N_2943,N_3727);
and U5537 (N_5537,N_2384,N_2786);
and U5538 (N_5538,N_3017,N_2810);
nand U5539 (N_5539,N_3361,N_2889);
nor U5540 (N_5540,N_2491,N_2160);
nor U5541 (N_5541,N_2371,N_3830);
nand U5542 (N_5542,N_3322,N_3783);
and U5543 (N_5543,N_2629,N_2437);
nor U5544 (N_5544,N_3282,N_3629);
or U5545 (N_5545,N_3872,N_2170);
or U5546 (N_5546,N_3277,N_3746);
and U5547 (N_5547,N_3406,N_2989);
and U5548 (N_5548,N_3195,N_3009);
and U5549 (N_5549,N_3389,N_2151);
nor U5550 (N_5550,N_2024,N_3642);
nand U5551 (N_5551,N_3282,N_3265);
nor U5552 (N_5552,N_3733,N_2551);
and U5553 (N_5553,N_2189,N_3177);
nand U5554 (N_5554,N_3111,N_2680);
nor U5555 (N_5555,N_2131,N_2220);
and U5556 (N_5556,N_3650,N_3476);
nor U5557 (N_5557,N_3090,N_3937);
or U5558 (N_5558,N_2722,N_2984);
and U5559 (N_5559,N_2979,N_3419);
nor U5560 (N_5560,N_2877,N_3877);
and U5561 (N_5561,N_2665,N_2287);
or U5562 (N_5562,N_3835,N_3216);
and U5563 (N_5563,N_2969,N_2589);
nand U5564 (N_5564,N_3453,N_3575);
or U5565 (N_5565,N_3021,N_2509);
or U5566 (N_5566,N_2449,N_3757);
and U5567 (N_5567,N_2352,N_3426);
nand U5568 (N_5568,N_2629,N_3570);
or U5569 (N_5569,N_2156,N_2556);
or U5570 (N_5570,N_2700,N_3127);
xnor U5571 (N_5571,N_2023,N_2633);
and U5572 (N_5572,N_2049,N_2913);
nand U5573 (N_5573,N_3445,N_3897);
nor U5574 (N_5574,N_2977,N_2127);
nor U5575 (N_5575,N_2476,N_2369);
or U5576 (N_5576,N_3999,N_3793);
and U5577 (N_5577,N_2926,N_2648);
nor U5578 (N_5578,N_2478,N_2712);
nor U5579 (N_5579,N_2416,N_3226);
and U5580 (N_5580,N_3293,N_3002);
xnor U5581 (N_5581,N_2636,N_2913);
and U5582 (N_5582,N_2448,N_2680);
nand U5583 (N_5583,N_3043,N_3134);
nor U5584 (N_5584,N_2050,N_2513);
nand U5585 (N_5585,N_2883,N_2139);
nor U5586 (N_5586,N_3393,N_2184);
and U5587 (N_5587,N_2545,N_3677);
nand U5588 (N_5588,N_2358,N_3160);
or U5589 (N_5589,N_3476,N_3454);
nor U5590 (N_5590,N_2832,N_2756);
and U5591 (N_5591,N_3360,N_3863);
or U5592 (N_5592,N_2158,N_2676);
nand U5593 (N_5593,N_3328,N_2893);
nand U5594 (N_5594,N_3783,N_3498);
nand U5595 (N_5595,N_3953,N_3328);
or U5596 (N_5596,N_2776,N_3081);
nor U5597 (N_5597,N_3627,N_3046);
or U5598 (N_5598,N_2352,N_2738);
or U5599 (N_5599,N_3407,N_2683);
xor U5600 (N_5600,N_2980,N_3446);
nand U5601 (N_5601,N_2758,N_3349);
or U5602 (N_5602,N_2413,N_3364);
and U5603 (N_5603,N_2218,N_3847);
or U5604 (N_5604,N_2087,N_3773);
and U5605 (N_5605,N_2092,N_3606);
or U5606 (N_5606,N_2503,N_3034);
nand U5607 (N_5607,N_3936,N_3142);
nor U5608 (N_5608,N_2865,N_2839);
and U5609 (N_5609,N_3290,N_2947);
and U5610 (N_5610,N_3870,N_3645);
nor U5611 (N_5611,N_3235,N_3322);
nand U5612 (N_5612,N_2946,N_3127);
and U5613 (N_5613,N_2605,N_2338);
xnor U5614 (N_5614,N_2971,N_3225);
nor U5615 (N_5615,N_3357,N_2105);
and U5616 (N_5616,N_3232,N_3094);
nand U5617 (N_5617,N_2375,N_3873);
nor U5618 (N_5618,N_3974,N_2798);
or U5619 (N_5619,N_2673,N_3978);
nor U5620 (N_5620,N_2254,N_2388);
nand U5621 (N_5621,N_3816,N_3476);
nand U5622 (N_5622,N_2349,N_3649);
and U5623 (N_5623,N_3934,N_2998);
nor U5624 (N_5624,N_2221,N_2398);
or U5625 (N_5625,N_2045,N_3086);
nor U5626 (N_5626,N_3675,N_3680);
nor U5627 (N_5627,N_3164,N_2152);
or U5628 (N_5628,N_3693,N_2355);
and U5629 (N_5629,N_3252,N_2620);
and U5630 (N_5630,N_3886,N_3850);
nand U5631 (N_5631,N_2243,N_3283);
or U5632 (N_5632,N_3150,N_3171);
or U5633 (N_5633,N_3391,N_2244);
nand U5634 (N_5634,N_3589,N_2502);
and U5635 (N_5635,N_3865,N_3075);
nor U5636 (N_5636,N_2133,N_2888);
nor U5637 (N_5637,N_2417,N_3427);
and U5638 (N_5638,N_2869,N_2181);
and U5639 (N_5639,N_2734,N_2528);
and U5640 (N_5640,N_2006,N_3555);
or U5641 (N_5641,N_2130,N_2777);
and U5642 (N_5642,N_2003,N_2548);
and U5643 (N_5643,N_2711,N_3008);
and U5644 (N_5644,N_3993,N_3378);
or U5645 (N_5645,N_3043,N_3436);
nand U5646 (N_5646,N_3676,N_3243);
and U5647 (N_5647,N_2739,N_3820);
nor U5648 (N_5648,N_3263,N_2236);
nor U5649 (N_5649,N_2947,N_2217);
nand U5650 (N_5650,N_3905,N_2246);
nand U5651 (N_5651,N_2851,N_3666);
nor U5652 (N_5652,N_2724,N_3690);
nand U5653 (N_5653,N_3158,N_3123);
nor U5654 (N_5654,N_3312,N_3300);
nand U5655 (N_5655,N_2191,N_3842);
nor U5656 (N_5656,N_2070,N_3964);
or U5657 (N_5657,N_3443,N_3441);
nand U5658 (N_5658,N_2695,N_3579);
nand U5659 (N_5659,N_2994,N_2319);
nand U5660 (N_5660,N_3075,N_3931);
and U5661 (N_5661,N_2198,N_2521);
nand U5662 (N_5662,N_3613,N_2814);
nand U5663 (N_5663,N_3226,N_3473);
or U5664 (N_5664,N_2580,N_3767);
and U5665 (N_5665,N_2324,N_3701);
and U5666 (N_5666,N_3182,N_2784);
or U5667 (N_5667,N_2817,N_3975);
and U5668 (N_5668,N_3928,N_2551);
and U5669 (N_5669,N_3941,N_3736);
nor U5670 (N_5670,N_3083,N_3726);
nand U5671 (N_5671,N_2014,N_2301);
or U5672 (N_5672,N_2965,N_2412);
nor U5673 (N_5673,N_3785,N_3957);
and U5674 (N_5674,N_2866,N_2965);
nor U5675 (N_5675,N_3925,N_2495);
nand U5676 (N_5676,N_3911,N_3398);
nor U5677 (N_5677,N_3302,N_2176);
nand U5678 (N_5678,N_3190,N_3554);
nand U5679 (N_5679,N_3680,N_3172);
nor U5680 (N_5680,N_2386,N_3466);
nor U5681 (N_5681,N_2793,N_3149);
nand U5682 (N_5682,N_3890,N_3205);
and U5683 (N_5683,N_3928,N_3914);
and U5684 (N_5684,N_2915,N_2522);
nand U5685 (N_5685,N_3656,N_2367);
or U5686 (N_5686,N_2997,N_3492);
nor U5687 (N_5687,N_2671,N_2517);
and U5688 (N_5688,N_2963,N_2859);
nor U5689 (N_5689,N_2553,N_3694);
and U5690 (N_5690,N_3534,N_2979);
or U5691 (N_5691,N_3977,N_3655);
nand U5692 (N_5692,N_2659,N_2071);
or U5693 (N_5693,N_2385,N_2759);
nor U5694 (N_5694,N_3220,N_3548);
and U5695 (N_5695,N_3993,N_2837);
nor U5696 (N_5696,N_3265,N_3869);
xor U5697 (N_5697,N_3989,N_3315);
and U5698 (N_5698,N_2585,N_2402);
and U5699 (N_5699,N_2533,N_2048);
nor U5700 (N_5700,N_3920,N_2525);
or U5701 (N_5701,N_3742,N_3478);
nand U5702 (N_5702,N_2773,N_3553);
nand U5703 (N_5703,N_2662,N_3457);
or U5704 (N_5704,N_2532,N_2184);
or U5705 (N_5705,N_2208,N_2980);
and U5706 (N_5706,N_3904,N_2891);
and U5707 (N_5707,N_2447,N_2837);
nand U5708 (N_5708,N_3165,N_2168);
or U5709 (N_5709,N_3624,N_2034);
or U5710 (N_5710,N_3258,N_2308);
nor U5711 (N_5711,N_3304,N_2004);
nor U5712 (N_5712,N_3187,N_3100);
nand U5713 (N_5713,N_3621,N_3227);
nand U5714 (N_5714,N_3835,N_3799);
or U5715 (N_5715,N_3524,N_3447);
nor U5716 (N_5716,N_3540,N_2440);
nand U5717 (N_5717,N_2980,N_2806);
nand U5718 (N_5718,N_2959,N_2319);
and U5719 (N_5719,N_3158,N_3491);
and U5720 (N_5720,N_2873,N_3953);
nor U5721 (N_5721,N_2033,N_3717);
nand U5722 (N_5722,N_3975,N_2483);
nand U5723 (N_5723,N_3988,N_2217);
and U5724 (N_5724,N_3291,N_3703);
nand U5725 (N_5725,N_3678,N_2895);
and U5726 (N_5726,N_2218,N_2848);
or U5727 (N_5727,N_3688,N_2666);
and U5728 (N_5728,N_2045,N_3030);
nand U5729 (N_5729,N_2945,N_2013);
or U5730 (N_5730,N_3669,N_2815);
or U5731 (N_5731,N_3536,N_2605);
nor U5732 (N_5732,N_2284,N_2349);
or U5733 (N_5733,N_3739,N_3187);
or U5734 (N_5734,N_3970,N_3402);
nor U5735 (N_5735,N_3071,N_3492);
or U5736 (N_5736,N_3467,N_2499);
xor U5737 (N_5737,N_2357,N_2013);
nor U5738 (N_5738,N_2523,N_2624);
nand U5739 (N_5739,N_2782,N_3403);
nor U5740 (N_5740,N_3224,N_2998);
or U5741 (N_5741,N_3896,N_3552);
nor U5742 (N_5742,N_3682,N_2081);
or U5743 (N_5743,N_2300,N_2615);
nand U5744 (N_5744,N_3805,N_2161);
nor U5745 (N_5745,N_2822,N_3528);
or U5746 (N_5746,N_2969,N_3304);
nor U5747 (N_5747,N_3150,N_3396);
and U5748 (N_5748,N_2277,N_2946);
nand U5749 (N_5749,N_3573,N_3702);
and U5750 (N_5750,N_2315,N_2491);
xor U5751 (N_5751,N_3764,N_2653);
or U5752 (N_5752,N_3198,N_2649);
or U5753 (N_5753,N_3126,N_2779);
or U5754 (N_5754,N_3375,N_2861);
nand U5755 (N_5755,N_2715,N_3323);
nor U5756 (N_5756,N_3457,N_2686);
nand U5757 (N_5757,N_2427,N_2027);
or U5758 (N_5758,N_3318,N_3881);
or U5759 (N_5759,N_2410,N_2314);
nand U5760 (N_5760,N_2959,N_2680);
nand U5761 (N_5761,N_3546,N_3890);
xor U5762 (N_5762,N_2759,N_3581);
and U5763 (N_5763,N_2078,N_2140);
or U5764 (N_5764,N_3766,N_2303);
nor U5765 (N_5765,N_2038,N_3810);
or U5766 (N_5766,N_2853,N_2414);
or U5767 (N_5767,N_3937,N_3637);
nor U5768 (N_5768,N_3798,N_2901);
nor U5769 (N_5769,N_3928,N_2950);
or U5770 (N_5770,N_3022,N_3439);
nand U5771 (N_5771,N_2354,N_2800);
or U5772 (N_5772,N_2399,N_3908);
nor U5773 (N_5773,N_2160,N_3415);
xor U5774 (N_5774,N_3201,N_3540);
or U5775 (N_5775,N_3495,N_3305);
and U5776 (N_5776,N_3888,N_2422);
and U5777 (N_5777,N_2429,N_2837);
nand U5778 (N_5778,N_3000,N_2301);
nand U5779 (N_5779,N_3097,N_3957);
and U5780 (N_5780,N_2535,N_3775);
and U5781 (N_5781,N_3669,N_2679);
nor U5782 (N_5782,N_3374,N_2371);
nand U5783 (N_5783,N_3917,N_3263);
nand U5784 (N_5784,N_3681,N_3367);
and U5785 (N_5785,N_3665,N_2290);
nor U5786 (N_5786,N_3035,N_3596);
nand U5787 (N_5787,N_2294,N_3938);
nor U5788 (N_5788,N_3331,N_3911);
xor U5789 (N_5789,N_2160,N_3292);
nor U5790 (N_5790,N_2515,N_3418);
nand U5791 (N_5791,N_2275,N_3569);
and U5792 (N_5792,N_2945,N_2539);
and U5793 (N_5793,N_3563,N_3897);
nor U5794 (N_5794,N_2006,N_3292);
nor U5795 (N_5795,N_3559,N_3401);
and U5796 (N_5796,N_3453,N_3925);
nor U5797 (N_5797,N_2499,N_2885);
nor U5798 (N_5798,N_3814,N_3534);
nand U5799 (N_5799,N_3636,N_3960);
nand U5800 (N_5800,N_2283,N_3353);
and U5801 (N_5801,N_2724,N_3368);
or U5802 (N_5802,N_2406,N_2799);
or U5803 (N_5803,N_3193,N_3108);
nor U5804 (N_5804,N_2783,N_2138);
or U5805 (N_5805,N_3191,N_3263);
or U5806 (N_5806,N_3307,N_2801);
nor U5807 (N_5807,N_3899,N_3697);
or U5808 (N_5808,N_2011,N_3398);
and U5809 (N_5809,N_2149,N_3443);
nand U5810 (N_5810,N_2613,N_2488);
or U5811 (N_5811,N_3187,N_3411);
and U5812 (N_5812,N_3419,N_2558);
nand U5813 (N_5813,N_3470,N_2401);
nand U5814 (N_5814,N_3453,N_2790);
nand U5815 (N_5815,N_3945,N_2411);
nand U5816 (N_5816,N_3407,N_2574);
and U5817 (N_5817,N_2807,N_2835);
and U5818 (N_5818,N_3818,N_2112);
and U5819 (N_5819,N_3712,N_3060);
nor U5820 (N_5820,N_2418,N_2688);
nor U5821 (N_5821,N_3081,N_3319);
nand U5822 (N_5822,N_2945,N_2180);
nand U5823 (N_5823,N_3887,N_3172);
nor U5824 (N_5824,N_2660,N_3840);
and U5825 (N_5825,N_3357,N_3959);
xnor U5826 (N_5826,N_3806,N_3552);
nand U5827 (N_5827,N_2484,N_3302);
nand U5828 (N_5828,N_2778,N_3521);
and U5829 (N_5829,N_2285,N_3105);
nand U5830 (N_5830,N_3528,N_3171);
nor U5831 (N_5831,N_3936,N_2094);
or U5832 (N_5832,N_3308,N_3181);
or U5833 (N_5833,N_2421,N_2390);
nor U5834 (N_5834,N_2137,N_3745);
or U5835 (N_5835,N_3976,N_3756);
nor U5836 (N_5836,N_3147,N_3923);
nand U5837 (N_5837,N_2933,N_3867);
nor U5838 (N_5838,N_3281,N_3936);
and U5839 (N_5839,N_3751,N_2495);
xnor U5840 (N_5840,N_2070,N_2578);
nand U5841 (N_5841,N_3281,N_3398);
nand U5842 (N_5842,N_3920,N_2573);
nor U5843 (N_5843,N_2634,N_2153);
nand U5844 (N_5844,N_2225,N_3258);
and U5845 (N_5845,N_2855,N_2087);
nand U5846 (N_5846,N_2800,N_2011);
and U5847 (N_5847,N_2084,N_3767);
nor U5848 (N_5848,N_2157,N_2084);
and U5849 (N_5849,N_2928,N_2946);
or U5850 (N_5850,N_3972,N_2799);
or U5851 (N_5851,N_3694,N_2224);
and U5852 (N_5852,N_3396,N_3073);
nor U5853 (N_5853,N_3232,N_3526);
and U5854 (N_5854,N_2840,N_3185);
xor U5855 (N_5855,N_2179,N_3341);
and U5856 (N_5856,N_3832,N_2776);
or U5857 (N_5857,N_2236,N_3138);
nand U5858 (N_5858,N_2305,N_2263);
or U5859 (N_5859,N_3956,N_3240);
and U5860 (N_5860,N_3280,N_2866);
and U5861 (N_5861,N_3695,N_3128);
nor U5862 (N_5862,N_2221,N_3567);
or U5863 (N_5863,N_2522,N_2330);
and U5864 (N_5864,N_2778,N_3489);
or U5865 (N_5865,N_2674,N_3255);
or U5866 (N_5866,N_2773,N_2673);
and U5867 (N_5867,N_2451,N_2469);
or U5868 (N_5868,N_2224,N_2583);
nand U5869 (N_5869,N_3452,N_3749);
nand U5870 (N_5870,N_3554,N_3135);
or U5871 (N_5871,N_2453,N_2167);
nor U5872 (N_5872,N_3835,N_2748);
or U5873 (N_5873,N_3788,N_3136);
or U5874 (N_5874,N_2233,N_3992);
and U5875 (N_5875,N_3050,N_3953);
nand U5876 (N_5876,N_3520,N_2119);
nand U5877 (N_5877,N_3192,N_3693);
or U5878 (N_5878,N_2015,N_2319);
nor U5879 (N_5879,N_2864,N_3772);
nor U5880 (N_5880,N_2501,N_2977);
nor U5881 (N_5881,N_3638,N_3054);
nand U5882 (N_5882,N_2894,N_3652);
nand U5883 (N_5883,N_2106,N_3580);
nor U5884 (N_5884,N_2470,N_2565);
or U5885 (N_5885,N_2655,N_3464);
nand U5886 (N_5886,N_2529,N_3054);
nand U5887 (N_5887,N_2888,N_3873);
and U5888 (N_5888,N_2718,N_2575);
or U5889 (N_5889,N_3551,N_3576);
and U5890 (N_5890,N_2403,N_3601);
or U5891 (N_5891,N_3572,N_3227);
nand U5892 (N_5892,N_2359,N_3155);
or U5893 (N_5893,N_3137,N_3226);
or U5894 (N_5894,N_2469,N_2906);
nor U5895 (N_5895,N_3419,N_3293);
and U5896 (N_5896,N_2944,N_3518);
or U5897 (N_5897,N_3290,N_2786);
or U5898 (N_5898,N_2747,N_3902);
and U5899 (N_5899,N_3787,N_3739);
and U5900 (N_5900,N_2860,N_2245);
nor U5901 (N_5901,N_3176,N_3876);
and U5902 (N_5902,N_3595,N_3672);
or U5903 (N_5903,N_3037,N_2415);
or U5904 (N_5904,N_2892,N_3381);
or U5905 (N_5905,N_2612,N_2087);
xor U5906 (N_5906,N_2262,N_3397);
nor U5907 (N_5907,N_3338,N_2760);
nor U5908 (N_5908,N_2422,N_2279);
nor U5909 (N_5909,N_2213,N_3753);
nand U5910 (N_5910,N_3945,N_2339);
and U5911 (N_5911,N_3440,N_3565);
nor U5912 (N_5912,N_2834,N_3391);
xor U5913 (N_5913,N_2430,N_3923);
or U5914 (N_5914,N_3708,N_2029);
nor U5915 (N_5915,N_3819,N_3365);
or U5916 (N_5916,N_3636,N_2874);
nor U5917 (N_5917,N_2708,N_3796);
or U5918 (N_5918,N_3371,N_3598);
nor U5919 (N_5919,N_2495,N_2449);
nand U5920 (N_5920,N_2728,N_2031);
or U5921 (N_5921,N_3908,N_3602);
nor U5922 (N_5922,N_3087,N_3819);
nand U5923 (N_5923,N_2733,N_2216);
or U5924 (N_5924,N_2199,N_2241);
nor U5925 (N_5925,N_2868,N_3553);
and U5926 (N_5926,N_3636,N_2575);
and U5927 (N_5927,N_2691,N_2580);
and U5928 (N_5928,N_3280,N_2693);
nor U5929 (N_5929,N_3490,N_2700);
or U5930 (N_5930,N_3571,N_2502);
nand U5931 (N_5931,N_2220,N_3746);
nand U5932 (N_5932,N_2204,N_2594);
nor U5933 (N_5933,N_2292,N_3810);
xor U5934 (N_5934,N_3773,N_3758);
nor U5935 (N_5935,N_3485,N_3173);
nor U5936 (N_5936,N_2196,N_2601);
nor U5937 (N_5937,N_3106,N_3977);
nand U5938 (N_5938,N_3710,N_3727);
nor U5939 (N_5939,N_3960,N_2380);
nand U5940 (N_5940,N_3205,N_2104);
nor U5941 (N_5941,N_2904,N_3435);
nor U5942 (N_5942,N_3908,N_2483);
nor U5943 (N_5943,N_2713,N_2332);
and U5944 (N_5944,N_3736,N_2918);
or U5945 (N_5945,N_2049,N_3999);
and U5946 (N_5946,N_2162,N_2246);
nand U5947 (N_5947,N_3387,N_2922);
and U5948 (N_5948,N_3816,N_2304);
nand U5949 (N_5949,N_2874,N_3258);
and U5950 (N_5950,N_2919,N_2603);
nor U5951 (N_5951,N_3144,N_2786);
and U5952 (N_5952,N_3864,N_2800);
nand U5953 (N_5953,N_3389,N_3845);
and U5954 (N_5954,N_3875,N_3516);
and U5955 (N_5955,N_2821,N_3965);
and U5956 (N_5956,N_2782,N_3428);
nand U5957 (N_5957,N_2395,N_3932);
or U5958 (N_5958,N_2107,N_3778);
nand U5959 (N_5959,N_2251,N_3789);
or U5960 (N_5960,N_2341,N_3138);
or U5961 (N_5961,N_2879,N_3437);
nand U5962 (N_5962,N_2190,N_3560);
nor U5963 (N_5963,N_2208,N_2474);
nand U5964 (N_5964,N_2016,N_3257);
or U5965 (N_5965,N_3440,N_3399);
nor U5966 (N_5966,N_2925,N_2139);
nand U5967 (N_5967,N_2164,N_2311);
and U5968 (N_5968,N_2323,N_3111);
and U5969 (N_5969,N_3226,N_2622);
nor U5970 (N_5970,N_2356,N_2705);
and U5971 (N_5971,N_3589,N_3420);
and U5972 (N_5972,N_3713,N_2317);
and U5973 (N_5973,N_3763,N_3904);
or U5974 (N_5974,N_3312,N_2251);
or U5975 (N_5975,N_3945,N_3288);
nor U5976 (N_5976,N_3429,N_2760);
and U5977 (N_5977,N_3460,N_2906);
nor U5978 (N_5978,N_2521,N_2712);
or U5979 (N_5979,N_3986,N_2286);
nand U5980 (N_5980,N_2612,N_3751);
nor U5981 (N_5981,N_3622,N_2171);
or U5982 (N_5982,N_3948,N_3335);
nand U5983 (N_5983,N_2710,N_3982);
or U5984 (N_5984,N_3789,N_3262);
xnor U5985 (N_5985,N_2211,N_3971);
nand U5986 (N_5986,N_3302,N_3607);
and U5987 (N_5987,N_2821,N_2288);
nand U5988 (N_5988,N_2566,N_3083);
nand U5989 (N_5989,N_2416,N_3653);
and U5990 (N_5990,N_3511,N_2874);
and U5991 (N_5991,N_3785,N_3939);
nor U5992 (N_5992,N_3744,N_2525);
nor U5993 (N_5993,N_2429,N_3457);
nor U5994 (N_5994,N_2424,N_2344);
and U5995 (N_5995,N_2592,N_2383);
or U5996 (N_5996,N_2147,N_3050);
and U5997 (N_5997,N_2912,N_2239);
or U5998 (N_5998,N_3217,N_3253);
nand U5999 (N_5999,N_2741,N_2655);
and U6000 (N_6000,N_4528,N_4226);
and U6001 (N_6001,N_4564,N_4537);
nand U6002 (N_6002,N_4823,N_4035);
nor U6003 (N_6003,N_5908,N_5891);
nand U6004 (N_6004,N_4286,N_4670);
nor U6005 (N_6005,N_4623,N_4615);
nor U6006 (N_6006,N_5315,N_5460);
nand U6007 (N_6007,N_4117,N_4168);
or U6008 (N_6008,N_5308,N_4403);
or U6009 (N_6009,N_4915,N_4078);
or U6010 (N_6010,N_4264,N_4404);
and U6011 (N_6011,N_4980,N_5352);
and U6012 (N_6012,N_5989,N_5396);
and U6013 (N_6013,N_4785,N_5482);
or U6014 (N_6014,N_4585,N_5689);
nor U6015 (N_6015,N_4231,N_5394);
and U6016 (N_6016,N_4002,N_4702);
or U6017 (N_6017,N_4727,N_5544);
and U6018 (N_6018,N_4989,N_4981);
nand U6019 (N_6019,N_4737,N_4825);
and U6020 (N_6020,N_5918,N_4960);
nor U6021 (N_6021,N_4714,N_5378);
nor U6022 (N_6022,N_4485,N_5234);
nor U6023 (N_6023,N_4071,N_5114);
nor U6024 (N_6024,N_5109,N_4255);
nor U6025 (N_6025,N_4445,N_4937);
nand U6026 (N_6026,N_5215,N_5546);
nand U6027 (N_6027,N_5216,N_4158);
and U6028 (N_6028,N_4868,N_5873);
nand U6029 (N_6029,N_5156,N_5831);
nand U6030 (N_6030,N_5984,N_4227);
and U6031 (N_6031,N_4665,N_5956);
nor U6032 (N_6032,N_4303,N_5011);
nor U6033 (N_6033,N_4838,N_4409);
or U6034 (N_6034,N_4085,N_4323);
nor U6035 (N_6035,N_4879,N_4632);
nand U6036 (N_6036,N_4617,N_4745);
and U6037 (N_6037,N_5195,N_4070);
and U6038 (N_6038,N_5213,N_5402);
nand U6039 (N_6039,N_5755,N_5963);
or U6040 (N_6040,N_4143,N_4173);
xnor U6041 (N_6041,N_5595,N_5037);
or U6042 (N_6042,N_5495,N_5436);
nand U6043 (N_6043,N_5660,N_5379);
and U6044 (N_6044,N_4010,N_4912);
xor U6045 (N_6045,N_5877,N_4633);
and U6046 (N_6046,N_4928,N_5977);
xor U6047 (N_6047,N_5609,N_4810);
and U6048 (N_6048,N_5064,N_5063);
or U6049 (N_6049,N_4663,N_4244);
and U6050 (N_6050,N_4197,N_5257);
and U6051 (N_6051,N_4342,N_5768);
nand U6052 (N_6052,N_5836,N_4424);
and U6053 (N_6053,N_5252,N_5543);
and U6054 (N_6054,N_5312,N_4700);
nor U6055 (N_6055,N_4771,N_4610);
nor U6056 (N_6056,N_4518,N_5926);
or U6057 (N_6057,N_4510,N_5448);
nor U6058 (N_6058,N_4640,N_4012);
or U6059 (N_6059,N_5611,N_5897);
and U6060 (N_6060,N_4198,N_5733);
or U6061 (N_6061,N_4209,N_4148);
xor U6062 (N_6062,N_5590,N_4907);
or U6063 (N_6063,N_5438,N_5497);
nand U6064 (N_6064,N_4536,N_4516);
or U6065 (N_6065,N_5382,N_5676);
and U6066 (N_6066,N_5682,N_4936);
nand U6067 (N_6067,N_5925,N_5842);
nor U6068 (N_6068,N_4312,N_4199);
nor U6069 (N_6069,N_4237,N_4666);
or U6070 (N_6070,N_4119,N_5367);
and U6071 (N_6071,N_4345,N_4067);
or U6072 (N_6072,N_4321,N_5454);
and U6073 (N_6073,N_4284,N_5734);
nand U6074 (N_6074,N_5605,N_4847);
and U6075 (N_6075,N_5393,N_5010);
nand U6076 (N_6076,N_4938,N_5957);
nor U6077 (N_6077,N_5596,N_5728);
nor U6078 (N_6078,N_5948,N_4798);
nor U6079 (N_6079,N_4719,N_4037);
or U6080 (N_6080,N_4011,N_5319);
and U6081 (N_6081,N_4102,N_5720);
xnor U6082 (N_6082,N_5714,N_4425);
nand U6083 (N_6083,N_4254,N_5444);
nor U6084 (N_6084,N_5480,N_5968);
and U6085 (N_6085,N_5289,N_4359);
or U6086 (N_6086,N_4099,N_4166);
xor U6087 (N_6087,N_5071,N_4175);
and U6088 (N_6088,N_4437,N_5964);
or U6089 (N_6089,N_5809,N_4178);
xor U6090 (N_6090,N_5539,N_4234);
nand U6091 (N_6091,N_4943,N_4688);
or U6092 (N_6092,N_5101,N_5725);
or U6093 (N_6093,N_4030,N_4660);
or U6094 (N_6094,N_4180,N_4863);
nor U6095 (N_6095,N_4162,N_4744);
nand U6096 (N_6096,N_4703,N_5426);
and U6097 (N_6097,N_4228,N_5098);
nor U6098 (N_6098,N_4899,N_4008);
and U6099 (N_6099,N_4794,N_4109);
or U6100 (N_6100,N_5620,N_4651);
nand U6101 (N_6101,N_5191,N_4776);
and U6102 (N_6102,N_5330,N_4426);
and U6103 (N_6103,N_4858,N_5028);
xnor U6104 (N_6104,N_4783,N_5411);
xnor U6105 (N_6105,N_5062,N_5067);
or U6106 (N_6106,N_5023,N_5787);
and U6107 (N_6107,N_5299,N_5392);
xnor U6108 (N_6108,N_4083,N_4818);
nand U6109 (N_6109,N_4310,N_4796);
and U6110 (N_6110,N_4271,N_5653);
nand U6111 (N_6111,N_4599,N_4133);
and U6112 (N_6112,N_5752,N_4276);
nor U6113 (N_6113,N_5073,N_5339);
or U6114 (N_6114,N_5827,N_5056);
and U6115 (N_6115,N_5236,N_5515);
and U6116 (N_6116,N_5980,N_5747);
and U6117 (N_6117,N_4925,N_5971);
and U6118 (N_6118,N_5796,N_4397);
nand U6119 (N_6119,N_4374,N_5223);
nand U6120 (N_6120,N_4056,N_4370);
xnor U6121 (N_6121,N_4479,N_4627);
nand U6122 (N_6122,N_5832,N_4969);
and U6123 (N_6123,N_5131,N_4324);
nor U6124 (N_6124,N_4095,N_5932);
and U6125 (N_6125,N_5342,N_4261);
and U6126 (N_6126,N_4467,N_4979);
nor U6127 (N_6127,N_4207,N_5401);
nand U6128 (N_6128,N_5400,N_4557);
or U6129 (N_6129,N_5084,N_5814);
or U6130 (N_6130,N_4563,N_5890);
nor U6131 (N_6131,N_5462,N_4545);
nor U6132 (N_6132,N_4317,N_5302);
or U6133 (N_6133,N_5091,N_5437);
or U6134 (N_6134,N_5014,N_5916);
nand U6135 (N_6135,N_4318,N_4944);
and U6136 (N_6136,N_5222,N_5095);
xnor U6137 (N_6137,N_5039,N_4931);
nand U6138 (N_6138,N_4210,N_4618);
or U6139 (N_6139,N_4740,N_5273);
and U6140 (N_6140,N_4890,N_5913);
nand U6141 (N_6141,N_4570,N_4320);
and U6142 (N_6142,N_4786,N_4878);
nand U6143 (N_6143,N_4401,N_4279);
nor U6144 (N_6144,N_5316,N_4494);
or U6145 (N_6145,N_5681,N_4471);
and U6146 (N_6146,N_5617,N_5074);
xor U6147 (N_6147,N_5475,N_4932);
or U6148 (N_6148,N_5876,N_5863);
and U6149 (N_6149,N_4909,N_4182);
nor U6150 (N_6150,N_5524,N_5615);
or U6151 (N_6151,N_5186,N_5512);
and U6152 (N_6152,N_4551,N_4144);
nor U6153 (N_6153,N_5002,N_5113);
and U6154 (N_6154,N_5120,N_5962);
or U6155 (N_6155,N_5790,N_4521);
and U6156 (N_6156,N_5711,N_4391);
and U6157 (N_6157,N_5469,N_5846);
nor U6158 (N_6158,N_4720,N_5922);
and U6159 (N_6159,N_4676,N_4832);
nand U6160 (N_6160,N_4681,N_4233);
or U6161 (N_6161,N_4253,N_5107);
nor U6162 (N_6162,N_5384,N_5516);
nand U6163 (N_6163,N_4435,N_4459);
or U6164 (N_6164,N_5703,N_4747);
or U6165 (N_6165,N_4590,N_4772);
or U6166 (N_6166,N_4171,N_5266);
or U6167 (N_6167,N_5804,N_4384);
or U6168 (N_6168,N_4045,N_5134);
or U6169 (N_6169,N_4281,N_4476);
or U6170 (N_6170,N_5938,N_4807);
nor U6171 (N_6171,N_4929,N_5381);
or U6172 (N_6172,N_4216,N_5121);
xor U6173 (N_6173,N_5993,N_4760);
and U6174 (N_6174,N_4713,N_4413);
nor U6175 (N_6175,N_4867,N_4027);
nor U6176 (N_6176,N_5662,N_5003);
nor U6177 (N_6177,N_4550,N_4218);
nand U6178 (N_6178,N_4788,N_4272);
and U6179 (N_6179,N_4031,N_5288);
xnor U6180 (N_6180,N_5430,N_5347);
xor U6181 (N_6181,N_4508,N_5053);
nor U6182 (N_6182,N_4137,N_5604);
nor U6183 (N_6183,N_4525,N_4603);
nand U6184 (N_6184,N_4195,N_5840);
and U6185 (N_6185,N_4015,N_5616);
or U6186 (N_6186,N_4736,N_4058);
or U6187 (N_6187,N_4654,N_5303);
nand U6188 (N_6188,N_5025,N_4492);
or U6189 (N_6189,N_5828,N_5641);
nor U6190 (N_6190,N_5363,N_4290);
and U6191 (N_6191,N_5738,N_4668);
nor U6192 (N_6192,N_4582,N_5797);
nand U6193 (N_6193,N_5936,N_5072);
or U6194 (N_6194,N_4396,N_5265);
nor U6195 (N_6195,N_4774,N_5552);
nor U6196 (N_6196,N_5189,N_5470);
nand U6197 (N_6197,N_5820,N_5767);
nor U6198 (N_6198,N_5661,N_4506);
or U6199 (N_6199,N_4115,N_5354);
or U6200 (N_6200,N_4438,N_5626);
nand U6201 (N_6201,N_5332,N_4808);
or U6202 (N_6202,N_4025,N_4001);
nand U6203 (N_6203,N_4515,N_4866);
nor U6204 (N_6204,N_5974,N_5415);
or U6205 (N_6205,N_4793,N_5867);
nor U6206 (N_6206,N_5465,N_4329);
xnor U6207 (N_6207,N_5920,N_5835);
nor U6208 (N_6208,N_4880,N_5581);
nor U6209 (N_6209,N_4962,N_4251);
and U6210 (N_6210,N_5455,N_4597);
or U6211 (N_6211,N_5730,N_4822);
nand U6212 (N_6212,N_5449,N_4411);
or U6213 (N_6213,N_5882,N_4268);
or U6214 (N_6214,N_5638,N_5937);
nand U6215 (N_6215,N_4717,N_5854);
nor U6216 (N_6216,N_5081,N_4652);
or U6217 (N_6217,N_5439,N_5205);
nor U6218 (N_6218,N_5076,N_5124);
nand U6219 (N_6219,N_4129,N_5671);
nand U6220 (N_6220,N_5294,N_5712);
or U6221 (N_6221,N_4241,N_4689);
and U6222 (N_6222,N_5245,N_4174);
and U6223 (N_6223,N_4007,N_4131);
or U6224 (N_6224,N_4604,N_5841);
and U6225 (N_6225,N_4856,N_5706);
and U6226 (N_6226,N_5663,N_5298);
or U6227 (N_6227,N_4883,N_4690);
nor U6228 (N_6228,N_4683,N_4327);
nor U6229 (N_6229,N_4677,N_4724);
nand U6230 (N_6230,N_4821,N_4337);
nor U6231 (N_6231,N_4019,N_4183);
or U6232 (N_6232,N_4270,N_5173);
nand U6233 (N_6233,N_4331,N_5614);
and U6234 (N_6234,N_5656,N_5669);
and U6235 (N_6235,N_5565,N_4816);
or U6236 (N_6236,N_5397,N_5260);
or U6237 (N_6237,N_5577,N_5583);
nand U6238 (N_6238,N_5696,N_5976);
or U6239 (N_6239,N_4498,N_4190);
nor U6240 (N_6240,N_4330,N_4947);
nand U6241 (N_6241,N_4824,N_4970);
or U6242 (N_6242,N_4366,N_4835);
nand U6243 (N_6243,N_5329,N_5575);
or U6244 (N_6244,N_5770,N_4975);
and U6245 (N_6245,N_4021,N_4420);
or U6246 (N_6246,N_5946,N_4135);
nor U6247 (N_6247,N_5097,N_4649);
and U6248 (N_6248,N_4507,N_5272);
nor U6249 (N_6249,N_5602,N_5017);
and U6250 (N_6250,N_4718,N_4311);
and U6251 (N_6251,N_4038,N_4283);
nor U6252 (N_6252,N_4361,N_5780);
and U6253 (N_6253,N_4555,N_5038);
nor U6254 (N_6254,N_5423,N_5117);
or U6255 (N_6255,N_5386,N_4988);
nor U6256 (N_6256,N_5709,N_5634);
nand U6257 (N_6257,N_5279,N_4836);
or U6258 (N_6258,N_5724,N_4893);
nand U6259 (N_6259,N_4855,N_5630);
or U6260 (N_6260,N_4065,N_5498);
xnor U6261 (N_6261,N_5421,N_4495);
nand U6262 (N_6262,N_5417,N_4850);
nor U6263 (N_6263,N_4904,N_4278);
and U6264 (N_6264,N_5704,N_4130);
nand U6265 (N_6265,N_5988,N_5678);
nor U6266 (N_6266,N_5307,N_4741);
and U6267 (N_6267,N_4579,N_5160);
or U6268 (N_6268,N_5677,N_5200);
and U6269 (N_6269,N_5226,N_5328);
or U6270 (N_6270,N_4296,N_5931);
and U6271 (N_6271,N_4902,N_5566);
or U6272 (N_6272,N_4319,N_5293);
or U6273 (N_6273,N_4371,N_4481);
or U6274 (N_6274,N_4161,N_5744);
nand U6275 (N_6275,N_5702,N_4338);
nor U6276 (N_6276,N_4051,N_5254);
nand U6277 (N_6277,N_4383,N_4646);
nand U6278 (N_6278,N_5281,N_5545);
or U6279 (N_6279,N_4256,N_5007);
xor U6280 (N_6280,N_5707,N_4598);
nor U6281 (N_6281,N_5594,N_4189);
nand U6282 (N_6282,N_4223,N_5954);
nor U6283 (N_6283,N_5691,N_4167);
nand U6284 (N_6284,N_4295,N_5208);
and U6285 (N_6285,N_4841,N_4995);
or U6286 (N_6286,N_4973,N_4795);
and U6287 (N_6287,N_4940,N_4770);
and U6288 (N_6288,N_4126,N_5871);
or U6289 (N_6289,N_5390,N_5180);
nand U6290 (N_6290,N_4349,N_4450);
nand U6291 (N_6291,N_5631,N_4987);
and U6292 (N_6292,N_4926,N_4307);
or U6293 (N_6293,N_5297,N_4385);
nor U6294 (N_6294,N_4346,N_5992);
and U6295 (N_6295,N_5051,N_5889);
or U6296 (N_6296,N_5822,N_5238);
xnor U6297 (N_6297,N_4952,N_4430);
and U6298 (N_6298,N_5162,N_4600);
or U6299 (N_6299,N_4358,N_4414);
nor U6300 (N_6300,N_5228,N_4339);
nor U6301 (N_6301,N_4122,N_5001);
nor U6302 (N_6302,N_5510,N_5810);
and U6303 (N_6303,N_5754,N_4016);
or U6304 (N_6304,N_5710,N_5099);
and U6305 (N_6305,N_5535,N_4073);
nor U6306 (N_6306,N_5243,N_4188);
and U6307 (N_6307,N_5060,N_4398);
and U6308 (N_6308,N_5323,N_5826);
or U6309 (N_6309,N_4939,N_4048);
nor U6310 (N_6310,N_5061,N_5021);
or U6311 (N_6311,N_4581,N_4363);
or U6312 (N_6312,N_5326,N_4451);
nor U6313 (N_6313,N_4326,N_5144);
and U6314 (N_6314,N_5533,N_5485);
nor U6315 (N_6315,N_5847,N_4591);
nand U6316 (N_6316,N_4275,N_4628);
nand U6317 (N_6317,N_5753,N_5659);
and U6318 (N_6318,N_4387,N_5250);
or U6319 (N_6319,N_5579,N_4444);
nor U6320 (N_6320,N_5472,N_5757);
and U6321 (N_6321,N_5959,N_4072);
nor U6322 (N_6322,N_5697,N_4204);
nor U6323 (N_6323,N_5325,N_4005);
and U6324 (N_6324,N_5406,N_4325);
or U6325 (N_6325,N_5939,N_4176);
nand U6326 (N_6326,N_4723,N_5395);
nand U6327 (N_6327,N_4517,N_4675);
or U6328 (N_6328,N_4674,N_5155);
nand U6329 (N_6329,N_5489,N_5619);
nand U6330 (N_6330,N_5079,N_4830);
and U6331 (N_6331,N_4142,N_4889);
nand U6332 (N_6332,N_4567,N_5077);
nor U6333 (N_6333,N_4972,N_5779);
nand U6334 (N_6334,N_4365,N_5657);
and U6335 (N_6335,N_4888,N_5562);
nor U6336 (N_6336,N_5532,N_4864);
or U6337 (N_6337,N_4735,N_4376);
nor U6338 (N_6338,N_4919,N_4657);
and U6339 (N_6339,N_4141,N_4607);
or U6340 (N_6340,N_5808,N_4853);
or U6341 (N_6341,N_4357,N_4520);
nand U6342 (N_6342,N_5821,N_4576);
nand U6343 (N_6343,N_5219,N_5150);
or U6344 (N_6344,N_4820,N_4419);
nand U6345 (N_6345,N_4250,N_5955);
or U6346 (N_6346,N_5774,N_5530);
xnor U6347 (N_6347,N_4814,N_4658);
nor U6348 (N_6348,N_5549,N_4448);
nor U6349 (N_6349,N_5139,N_4245);
nor U6350 (N_6350,N_5991,N_5012);
and U6351 (N_6351,N_4558,N_5306);
and U6352 (N_6352,N_4291,N_5679);
nor U6353 (N_6353,N_5389,N_4427);
and U6354 (N_6354,N_5942,N_5020);
nor U6355 (N_6355,N_4090,N_4589);
nand U6356 (N_6356,N_4285,N_4573);
xor U6357 (N_6357,N_4764,N_5314);
nand U6358 (N_6358,N_4196,N_4375);
and U6359 (N_6359,N_4047,N_4861);
or U6360 (N_6360,N_4769,N_5811);
and U6361 (N_6361,N_5979,N_4041);
and U6362 (N_6362,N_5737,N_4111);
nand U6363 (N_6363,N_5527,N_4453);
nand U6364 (N_6364,N_4819,N_5078);
nand U6365 (N_6365,N_4140,N_4063);
or U6366 (N_6366,N_4968,N_5305);
and U6367 (N_6367,N_5096,N_5966);
or U6368 (N_6368,N_5275,N_4201);
nand U6369 (N_6369,N_5351,N_4758);
and U6370 (N_6370,N_5912,N_5645);
and U6371 (N_6371,N_5255,N_4433);
and U6372 (N_6372,N_4635,N_5794);
nor U6373 (N_6373,N_5235,N_4739);
and U6374 (N_6374,N_5082,N_5277);
nand U6375 (N_6375,N_4695,N_5901);
xnor U6376 (N_6376,N_5068,N_4913);
or U6377 (N_6377,N_4449,N_4860);
or U6378 (N_6378,N_5563,N_4608);
or U6379 (N_6379,N_5945,N_5715);
or U6380 (N_6380,N_5588,N_5129);
and U6381 (N_6381,N_4750,N_4766);
nor U6382 (N_6382,N_5874,N_5815);
and U6383 (N_6383,N_5399,N_4461);
nand U6384 (N_6384,N_4500,N_4884);
nor U6385 (N_6385,N_5269,N_5838);
nand U6386 (N_6386,N_5597,N_5185);
nor U6387 (N_6387,N_5478,N_5783);
and U6388 (N_6388,N_5164,N_5324);
or U6389 (N_6389,N_4460,N_4725);
or U6390 (N_6390,N_4229,N_5457);
or U6391 (N_6391,N_4659,N_5206);
nor U6392 (N_6392,N_5452,N_4542);
and U6393 (N_6393,N_5207,N_4875);
or U6394 (N_6394,N_4803,N_4985);
or U6395 (N_6395,N_5199,N_4679);
nor U6396 (N_6396,N_4815,N_5561);
or U6397 (N_6397,N_4629,N_4918);
or U6398 (N_6398,N_4742,N_4594);
nor U6399 (N_6399,N_4812,N_5667);
nand U6400 (N_6400,N_5054,N_4230);
nand U6401 (N_6401,N_4678,N_4215);
nand U6402 (N_6402,N_4191,N_4205);
nand U6403 (N_6403,N_4052,N_4225);
and U6404 (N_6404,N_4773,N_5343);
and U6405 (N_6405,N_4466,N_4593);
nor U6406 (N_6406,N_4149,N_4302);
and U6407 (N_6407,N_4854,N_4958);
or U6408 (N_6408,N_5176,N_5798);
and U6409 (N_6409,N_5593,N_5420);
or U6410 (N_6410,N_5765,N_5987);
and U6411 (N_6411,N_4150,N_5845);
nor U6412 (N_6412,N_4871,N_5547);
nor U6413 (N_6413,N_5159,N_4344);
nor U6414 (N_6414,N_5380,N_5743);
and U6415 (N_6415,N_5151,N_5311);
or U6416 (N_6416,N_4526,N_4273);
nand U6417 (N_6417,N_5785,N_5253);
nor U6418 (N_6418,N_5049,N_4948);
and U6419 (N_6419,N_5726,N_5259);
and U6420 (N_6420,N_5116,N_4123);
nor U6421 (N_6421,N_5895,N_5652);
or U6422 (N_6422,N_5899,N_4722);
and U6423 (N_6423,N_5598,N_4869);
and U6424 (N_6424,N_4601,N_5748);
nand U6425 (N_6425,N_5763,N_4924);
nor U6426 (N_6426,N_4566,N_5006);
or U6427 (N_6427,N_4499,N_4288);
nand U6428 (N_6428,N_4262,N_5239);
and U6429 (N_6429,N_4511,N_4152);
nand U6430 (N_6430,N_4066,N_4896);
xnor U6431 (N_6431,N_4643,N_4691);
xor U6432 (N_6432,N_4033,N_5230);
or U6433 (N_6433,N_5232,N_5204);
nor U6434 (N_6434,N_4258,N_4921);
nor U6435 (N_6435,N_4829,N_5824);
nand U6436 (N_6436,N_4957,N_4502);
nor U6437 (N_6437,N_5027,N_4049);
nor U6438 (N_6438,N_4616,N_5026);
nor U6439 (N_6439,N_4709,N_4145);
or U6440 (N_6440,N_4165,N_4606);
nand U6441 (N_6441,N_5746,N_5924);
nand U6442 (N_6442,N_5031,N_5088);
and U6443 (N_6443,N_5930,N_5910);
and U6444 (N_6444,N_4332,N_4040);
and U6445 (N_6445,N_5112,N_4761);
nand U6446 (N_6446,N_4993,N_4335);
or U6447 (N_6447,N_4266,N_5556);
or U6448 (N_6448,N_4484,N_5359);
nor U6449 (N_6449,N_5414,N_5092);
nand U6450 (N_6450,N_5672,N_5042);
nand U6451 (N_6451,N_4927,N_5699);
nand U6452 (N_6452,N_4263,N_5203);
and U6453 (N_6453,N_4755,N_5066);
nand U6454 (N_6454,N_4574,N_4187);
nor U6455 (N_6455,N_4686,N_5885);
or U6456 (N_6456,N_5247,N_5100);
and U6457 (N_6457,N_4638,N_5683);
nor U6458 (N_6458,N_5943,N_4434);
nand U6459 (N_6459,N_4428,N_4153);
or U6460 (N_6460,N_5418,N_4315);
and U6461 (N_6461,N_4417,N_4351);
or U6462 (N_6462,N_4472,N_4294);
nand U6463 (N_6463,N_5148,N_5461);
and U6464 (N_6464,N_5990,N_5643);
nor U6465 (N_6465,N_5424,N_5587);
nor U6466 (N_6466,N_5736,N_4368);
or U6467 (N_6467,N_5701,N_5103);
xor U6468 (N_6468,N_5262,N_4124);
nand U6469 (N_6469,N_4032,N_4792);
or U6470 (N_6470,N_5708,N_4509);
nor U6471 (N_6471,N_4749,N_5806);
nor U6472 (N_6472,N_4217,N_4895);
and U6473 (N_6473,N_4077,N_5300);
nand U6474 (N_6474,N_5521,N_5086);
nor U6475 (N_6475,N_5130,N_5434);
or U6476 (N_6476,N_4355,N_5280);
nand U6477 (N_6477,N_4706,N_4842);
nor U6478 (N_6478,N_5152,N_5220);
or U6479 (N_6479,N_5511,N_4219);
nand U6480 (N_6480,N_4743,N_5944);
or U6481 (N_6481,N_4159,N_4300);
and U6482 (N_6482,N_5358,N_5490);
or U6483 (N_6483,N_4029,N_4614);
and U6484 (N_6484,N_4081,N_5621);
nor U6485 (N_6485,N_5009,N_4694);
and U6486 (N_6486,N_5610,N_4293);
nand U6487 (N_6487,N_4112,N_4249);
or U6488 (N_6488,N_4194,N_4478);
nor U6489 (N_6489,N_5799,N_4650);
nor U6490 (N_6490,N_4456,N_5198);
and U6491 (N_6491,N_4076,N_5034);
and U6492 (N_6492,N_4084,N_5348);
nor U6493 (N_6493,N_4292,N_4372);
and U6494 (N_6494,N_5224,N_5403);
or U6495 (N_6495,N_4394,N_4922);
and U6496 (N_6496,N_4333,N_5338);
or U6497 (N_6497,N_4017,N_4524);
nor U6498 (N_6498,N_4621,N_5141);
or U6499 (N_6499,N_4408,N_5453);
nor U6500 (N_6500,N_4314,N_4777);
xor U6501 (N_6501,N_5214,N_5513);
and U6502 (N_6502,N_5267,N_5443);
xor U6503 (N_6503,N_5331,N_5951);
nor U6504 (N_6504,N_5477,N_4903);
nand U6505 (N_6505,N_5819,N_4546);
or U6506 (N_6506,N_5914,N_5286);
nor U6507 (N_6507,N_5903,N_4220);
and U6508 (N_6508,N_4556,N_4698);
nor U6509 (N_6509,N_5165,N_5104);
nand U6510 (N_6510,N_4734,N_5555);
or U6511 (N_6511,N_5655,N_4806);
and U6512 (N_6512,N_5169,N_4496);
and U6513 (N_6513,N_5887,N_4523);
nor U6514 (N_6514,N_5187,N_5875);
nor U6515 (N_6515,N_5468,N_5741);
or U6516 (N_6516,N_4093,N_5857);
or U6517 (N_6517,N_4848,N_4107);
nand U6518 (N_6518,N_5376,N_4831);
nand U6519 (N_6519,N_5409,N_4089);
nand U6520 (N_6520,N_5290,N_4613);
nand U6521 (N_6521,N_5869,N_5705);
or U6522 (N_6522,N_5902,N_5132);
nand U6523 (N_6523,N_5830,N_5529);
nand U6524 (N_6524,N_5432,N_5483);
nand U6525 (N_6525,N_5240,N_4971);
or U6526 (N_6526,N_5333,N_4986);
and U6527 (N_6527,N_4619,N_5571);
nand U6528 (N_6528,N_5739,N_4642);
or U6529 (N_6529,N_5138,N_4956);
xnor U6530 (N_6530,N_5047,N_5750);
or U6531 (N_6531,N_5135,N_4114);
or U6532 (N_6532,N_5337,N_5852);
nand U6533 (N_6533,N_4791,N_5801);
nand U6534 (N_6534,N_5356,N_4645);
or U6535 (N_6535,N_5713,N_5295);
and U6536 (N_6536,N_4715,N_5296);
or U6537 (N_6537,N_4583,N_5717);
nor U6538 (N_6538,N_4000,N_4876);
or U6539 (N_6539,N_4892,N_4055);
or U6540 (N_6540,N_5126,N_4094);
nand U6541 (N_6541,N_5334,N_5133);
nand U6542 (N_6542,N_5933,N_5157);
and U6543 (N_6543,N_4061,N_4105);
nand U6544 (N_6544,N_5906,N_5301);
xnor U6545 (N_6545,N_5451,N_4134);
or U6546 (N_6546,N_5196,N_5177);
and U6547 (N_6547,N_4697,N_4547);
nand U6548 (N_6548,N_4911,N_5837);
or U6549 (N_6549,N_4157,N_5559);
nor U6550 (N_6550,N_4243,N_5033);
nand U6551 (N_6551,N_5928,N_5435);
or U6552 (N_6552,N_4442,N_4132);
nor U6553 (N_6553,N_4313,N_5355);
or U6554 (N_6554,N_4381,N_5868);
nor U6555 (N_6555,N_4655,N_4458);
or U6556 (N_6556,N_4147,N_4648);
or U6557 (N_6557,N_4138,N_4763);
or U6558 (N_6558,N_4274,N_5090);
nor U6559 (N_6559,N_5282,N_5413);
nand U6560 (N_6560,N_5270,N_4587);
nand U6561 (N_6561,N_4910,N_4512);
or U6562 (N_6562,N_4407,N_5410);
and U6563 (N_6563,N_5839,N_5686);
nor U6564 (N_6564,N_4440,N_5981);
or U6565 (N_6565,N_4421,N_4738);
or U6566 (N_6566,N_5637,N_4768);
or U6567 (N_6567,N_4113,N_5540);
and U6568 (N_6568,N_5057,N_5446);
nand U6569 (N_6569,N_4881,N_4530);
or U6570 (N_6570,N_5357,N_4999);
nand U6571 (N_6571,N_5694,N_4631);
nand U6572 (N_6572,N_5592,N_5572);
nor U6573 (N_6573,N_5526,N_5246);
or U6574 (N_6574,N_4282,N_5456);
nand U6575 (N_6575,N_5878,N_4489);
and U6576 (N_6576,N_4347,N_5856);
and U6577 (N_6577,N_5464,N_4505);
nor U6578 (N_6578,N_5005,N_5018);
nor U6579 (N_6579,N_4996,N_4559);
and U6580 (N_6580,N_4992,N_5408);
and U6581 (N_6581,N_4699,N_5491);
nand U6582 (N_6582,N_5622,N_4522);
nand U6583 (N_6583,N_5570,N_5404);
nand U6584 (N_6584,N_4942,N_4905);
nand U6585 (N_6585,N_4400,N_4897);
and U6586 (N_6586,N_5344,N_5167);
and U6587 (N_6587,N_5865,N_5782);
nor U6588 (N_6588,N_4859,N_5674);
nor U6589 (N_6589,N_5953,N_4042);
and U6590 (N_6590,N_5927,N_5052);
or U6591 (N_6591,N_4701,N_5536);
xor U6592 (N_6592,N_5375,N_5346);
nand U6593 (N_6593,N_4534,N_4994);
and U6594 (N_6594,N_5843,N_5921);
nor U6595 (N_6595,N_4179,N_4309);
and U6596 (N_6596,N_5648,N_5416);
nor U6597 (N_6597,N_5970,N_5855);
and U6598 (N_6598,N_4074,N_4353);
nor U6599 (N_6599,N_4732,N_5321);
or U6600 (N_6600,N_4751,N_5795);
or U6601 (N_6601,N_5761,N_5789);
or U6602 (N_6602,N_4535,N_5862);
nor U6603 (N_6603,N_4588,N_5476);
or U6604 (N_6604,N_4865,N_4493);
nand U6605 (N_6605,N_4809,N_4193);
nor U6606 (N_6606,N_4014,N_5440);
nand U6607 (N_6607,N_5517,N_5249);
nor U6608 (N_6608,N_4541,N_4578);
nand U6609 (N_6609,N_5140,N_5760);
nand U6610 (N_6610,N_5844,N_4961);
or U6611 (N_6611,N_5996,N_5202);
nand U6612 (N_6612,N_5591,N_5118);
or U6613 (N_6613,N_4386,N_4804);
or U6614 (N_6614,N_4963,N_5364);
nor U6615 (N_6615,N_5531,N_5447);
and U6616 (N_6616,N_4833,N_4377);
or U6617 (N_6617,N_5041,N_5184);
nand U6618 (N_6618,N_5823,N_5884);
or U6619 (N_6619,N_5197,N_5178);
and U6620 (N_6620,N_5506,N_4043);
nor U6621 (N_6621,N_5881,N_4436);
nand U6622 (N_6622,N_5507,N_5762);
and U6623 (N_6623,N_5473,N_5428);
nor U6624 (N_6624,N_4392,N_4224);
nor U6625 (N_6625,N_5600,N_4572);
or U6626 (N_6626,N_5646,N_4208);
and U6627 (N_6627,N_5735,N_5606);
or U6628 (N_6628,N_4488,N_5111);
nand U6629 (N_6629,N_5442,N_5649);
or U6630 (N_6630,N_4259,N_5285);
nand U6631 (N_6631,N_5551,N_5479);
or U6632 (N_6632,N_5560,N_5158);
or U6633 (N_6633,N_5756,N_4464);
nor U6634 (N_6634,N_4609,N_4920);
or U6635 (N_6635,N_5668,N_4527);
and U6636 (N_6636,N_5650,N_5048);
nand U6637 (N_6637,N_5175,N_4834);
nand U6638 (N_6638,N_5494,N_5568);
nand U6639 (N_6639,N_5125,N_5019);
nand U6640 (N_6640,N_5192,N_4104);
nor U6641 (N_6641,N_5522,N_5370);
nand U6642 (N_6642,N_4540,N_4336);
nor U6643 (N_6643,N_5463,N_4068);
or U6644 (N_6644,N_4468,N_4656);
xnor U6645 (N_6645,N_5859,N_4277);
nand U6646 (N_6646,N_5635,N_4172);
and U6647 (N_6647,N_5849,N_5853);
xnor U6648 (N_6648,N_4023,N_4232);
and U6649 (N_6649,N_5923,N_5727);
nand U6650 (N_6650,N_5664,N_4672);
and U6651 (N_6651,N_5684,N_5313);
nor U6652 (N_6652,N_5773,N_5212);
and U6653 (N_6653,N_5817,N_5143);
and U6654 (N_6654,N_5030,N_4354);
and U6655 (N_6655,N_5573,N_5624);
or U6656 (N_6656,N_5909,N_4299);
nand U6657 (N_6657,N_5229,N_4412);
nand U6658 (N_6658,N_4990,N_5317);
and U6659 (N_6659,N_4543,N_4839);
and U6660 (N_6660,N_4639,N_5309);
nor U6661 (N_6661,N_5850,N_5749);
nor U6662 (N_6662,N_4716,N_5558);
xor U6663 (N_6663,N_4091,N_4787);
xnor U6664 (N_6664,N_5287,N_4671);
or U6665 (N_6665,N_5171,N_4647);
and U6666 (N_6666,N_4886,N_5256);
nand U6667 (N_6667,N_5122,N_4060);
xnor U6668 (N_6668,N_4901,N_4977);
or U6669 (N_6669,N_5501,N_5986);
nand U6670 (N_6670,N_5567,N_5242);
nor U6671 (N_6671,N_4762,N_4446);
nor U6672 (N_6672,N_4602,N_4753);
and U6673 (N_6673,N_4729,N_5805);
or U6674 (N_6674,N_5872,N_5193);
and U6675 (N_6675,N_4260,N_5569);
xnor U6676 (N_6676,N_4531,N_4422);
and U6677 (N_6677,N_4894,N_4827);
nand U6678 (N_6678,N_5194,N_5700);
or U6679 (N_6679,N_4637,N_5471);
or U6680 (N_6680,N_4103,N_5675);
or U6681 (N_6681,N_5586,N_4955);
or U6682 (N_6682,N_5024,N_4811);
nand U6683 (N_6683,N_5508,N_5368);
or U6684 (N_6684,N_5985,N_5792);
nand U6685 (N_6685,N_4388,N_4721);
nor U6686 (N_6686,N_4605,N_5163);
nor U6687 (N_6687,N_4872,N_4826);
nand U6688 (N_6688,N_5016,N_4006);
or U6689 (N_6689,N_5388,N_5777);
nand U6690 (N_6690,N_5231,N_4086);
nand U6691 (N_6691,N_4661,N_4684);
and U6692 (N_6692,N_4186,N_4898);
and U6693 (N_6693,N_5274,N_4118);
and U6694 (N_6694,N_5934,N_5803);
and U6695 (N_6695,N_4873,N_5665);
nor U6696 (N_6696,N_5174,N_4470);
nand U6697 (N_6697,N_5182,N_5983);
or U6698 (N_6698,N_4004,N_4790);
or U6699 (N_6699,N_4018,N_4441);
nand U6700 (N_6700,N_4731,N_4235);
or U6701 (N_6701,N_4289,N_4475);
and U6702 (N_6702,N_5578,N_5745);
nand U6703 (N_6703,N_4486,N_5237);
nor U6704 (N_6704,N_4390,N_5304);
or U6705 (N_6705,N_4746,N_5168);
or U6706 (N_6706,N_5800,N_5861);
or U6707 (N_6707,N_5361,N_4389);
or U6708 (N_6708,N_4402,N_5632);
xnor U6709 (N_6709,N_4759,N_4192);
nor U6710 (N_6710,N_5044,N_4062);
or U6711 (N_6711,N_5369,N_5405);
nor U6712 (N_6712,N_4252,N_4415);
nand U6713 (N_6713,N_5893,N_4687);
nand U6714 (N_6714,N_5261,N_5387);
nor U6715 (N_6715,N_4064,N_5612);
or U6716 (N_6716,N_5069,N_5751);
nand U6717 (N_6717,N_5466,N_5525);
nand U6718 (N_6718,N_5102,N_5486);
and U6719 (N_6719,N_4214,N_5601);
nor U6720 (N_6720,N_5629,N_4108);
nor U6721 (N_6721,N_4611,N_4967);
or U6722 (N_6722,N_5015,N_4538);
and U6723 (N_6723,N_4953,N_4101);
and U6724 (N_6724,N_5105,N_4305);
and U6725 (N_6725,N_4906,N_5919);
and U6726 (N_6726,N_4406,N_4584);
nand U6727 (N_6727,N_4951,N_4480);
and U6728 (N_6728,N_4730,N_5283);
and U6729 (N_6729,N_4726,N_5350);
nor U6730 (N_6730,N_4304,N_4222);
or U6731 (N_6731,N_4877,N_5154);
or U6732 (N_6732,N_5633,N_4151);
nand U6733 (N_6733,N_4340,N_4634);
nand U6734 (N_6734,N_5905,N_4039);
and U6735 (N_6735,N_4034,N_4022);
nor U6736 (N_6736,N_5520,N_4998);
nand U6737 (N_6737,N_4160,N_4057);
or U6738 (N_6738,N_4088,N_5335);
and U6739 (N_6739,N_4705,N_4287);
nand U6740 (N_6740,N_5721,N_4682);
or U6741 (N_6741,N_4959,N_5613);
nor U6742 (N_6742,N_5080,N_5880);
and U6743 (N_6743,N_5147,N_4852);
nand U6744 (N_6744,N_4782,N_5929);
nand U6745 (N_6745,N_4935,N_5731);
xnor U6746 (N_6746,N_4954,N_4369);
nand U6747 (N_6747,N_5059,N_5040);
or U6748 (N_6748,N_5670,N_5848);
nor U6749 (N_6749,N_5915,N_4301);
nor U6750 (N_6750,N_4462,N_4373);
nand U6751 (N_6751,N_5554,N_4242);
nand U6752 (N_6752,N_4817,N_4046);
nand U6753 (N_6753,N_5032,N_5778);
nor U6754 (N_6754,N_5947,N_4474);
nor U6755 (N_6755,N_4707,N_5965);
nor U6756 (N_6756,N_4552,N_4828);
nand U6757 (N_6757,N_5431,N_5487);
and U6758 (N_6758,N_5488,N_4733);
xor U6759 (N_6759,N_4028,N_4248);
nor U6760 (N_6760,N_4775,N_5917);
nor U6761 (N_6761,N_5818,N_4221);
or U6762 (N_6762,N_5900,N_5029);
and U6763 (N_6763,N_4711,N_5504);
nor U6764 (N_6764,N_4641,N_4322);
nor U6765 (N_6765,N_4801,N_5271);
nor U6766 (N_6766,N_5972,N_5627);
nor U6767 (N_6767,N_4463,N_5716);
nand U6768 (N_6768,N_5625,N_5509);
nor U6769 (N_6769,N_5327,N_5888);
and U6770 (N_6770,N_4079,N_5647);
nand U6771 (N_6771,N_5264,N_5599);
and U6772 (N_6772,N_5911,N_4797);
and U6773 (N_6773,N_4667,N_5045);
nand U6774 (N_6774,N_4813,N_4982);
or U6775 (N_6775,N_4393,N_5788);
and U6776 (N_6776,N_4851,N_5166);
nor U6777 (N_6777,N_4423,N_4036);
and U6778 (N_6778,N_4170,N_5636);
nand U6779 (N_6779,N_4395,N_5385);
and U6780 (N_6780,N_5108,N_4455);
and U6781 (N_6781,N_5083,N_4352);
nor U6782 (N_6782,N_4075,N_4849);
and U6783 (N_6783,N_5374,N_5999);
and U6784 (N_6784,N_5758,N_4504);
or U6785 (N_6785,N_4306,N_5146);
nor U6786 (N_6786,N_4379,N_5772);
nor U6787 (N_6787,N_4100,N_5340);
nor U6788 (N_6788,N_5894,N_4367);
and U6789 (N_6789,N_5975,N_4708);
nor U6790 (N_6790,N_4664,N_5864);
nor U6791 (N_6791,N_4754,N_5542);
or U6792 (N_6792,N_5967,N_4857);
nand U6793 (N_6793,N_4514,N_4009);
nand U6794 (N_6794,N_4704,N_5623);
nand U6795 (N_6795,N_5484,N_4662);
or U6796 (N_6796,N_4364,N_5994);
and U6797 (N_6797,N_4267,N_5769);
or U6798 (N_6798,N_4206,N_5127);
and U6799 (N_6799,N_4900,N_4050);
nor U6800 (N_6800,N_4439,N_5978);
nor U6801 (N_6801,N_5322,N_4549);
nand U6802 (N_6802,N_5528,N_4110);
and U6803 (N_6803,N_4846,N_5941);
nand U6804 (N_6804,N_4184,N_5398);
nand U6805 (N_6805,N_4780,N_5085);
nor U6806 (N_6806,N_4519,N_4974);
xnor U6807 (N_6807,N_5580,N_5492);
nor U6808 (N_6808,N_4308,N_5043);
nand U6809 (N_6809,N_5391,N_5995);
or U6810 (N_6810,N_5961,N_4767);
and U6811 (N_6811,N_5425,N_4155);
and U6812 (N_6812,N_5589,N_5500);
nand U6813 (N_6813,N_5149,N_5952);
or U6814 (N_6814,N_4513,N_5585);
nand U6815 (N_6815,N_4539,N_4116);
or U6816 (N_6816,N_4568,N_5698);
or U6817 (N_6817,N_5371,N_4298);
nor U6818 (N_6818,N_4024,N_4003);
nand U6819 (N_6819,N_5433,N_4862);
and U6820 (N_6820,N_4154,N_5858);
nor U6821 (N_6821,N_4966,N_5557);
and U6822 (N_6822,N_4236,N_5407);
or U6823 (N_6823,N_4908,N_4991);
nor U6824 (N_6824,N_4874,N_5958);
or U6825 (N_6825,N_5502,N_5441);
and U6826 (N_6826,N_4343,N_5688);
or U6827 (N_6827,N_4548,N_5050);
or U6828 (N_6828,N_4693,N_4748);
nand U6829 (N_6829,N_5576,N_5251);
or U6830 (N_6830,N_4156,N_5218);
and U6831 (N_6831,N_5816,N_4457);
or U6832 (N_6832,N_4013,N_5022);
nand U6833 (N_6833,N_5268,N_5644);
nand U6834 (N_6834,N_5654,N_5362);
nor U6835 (N_6835,N_4612,N_4405);
and U6836 (N_6836,N_5372,N_4169);
nor U6837 (N_6837,N_5241,N_4483);
or U6838 (N_6838,N_5365,N_4964);
and U6839 (N_6839,N_4571,N_4328);
or U6840 (N_6840,N_5519,N_4680);
or U6841 (N_6841,N_4473,N_4020);
nor U6842 (N_6842,N_5211,N_4431);
nand U6843 (N_6843,N_5291,N_4098);
nor U6844 (N_6844,N_5886,N_4348);
xnor U6845 (N_6845,N_5383,N_5642);
nor U6846 (N_6846,N_5065,N_5935);
and U6847 (N_6847,N_4121,N_4533);
nand U6848 (N_6848,N_4120,N_4128);
xnor U6849 (N_6849,N_5366,N_5036);
or U6850 (N_6850,N_4080,N_4044);
nand U6851 (N_6851,N_5982,N_5784);
or U6852 (N_6852,N_4845,N_4799);
nand U6853 (N_6853,N_5960,N_4482);
xnor U6854 (N_6854,N_5136,N_5459);
nor U6855 (N_6855,N_5603,N_4026);
nor U6856 (N_6856,N_5227,N_4580);
nand U6857 (N_6857,N_4341,N_5070);
or U6858 (N_6858,N_5892,N_4418);
xor U6859 (N_6859,N_5467,N_5427);
xnor U6860 (N_6860,N_5258,N_4562);
and U6861 (N_6861,N_5493,N_5651);
or U6862 (N_6862,N_5360,N_5775);
nand U6863 (N_6863,N_4887,N_5248);
nand U6864 (N_6864,N_4239,N_4362);
nor U6865 (N_6865,N_4380,N_5349);
and U6866 (N_6866,N_5786,N_5541);
nor U6867 (N_6867,N_5742,N_5538);
nand U6868 (N_6868,N_4586,N_4497);
and U6869 (N_6869,N_4789,N_4561);
and U6870 (N_6870,N_4082,N_4779);
xor U6871 (N_6871,N_4781,N_4212);
and U6872 (N_6872,N_4916,N_4620);
nand U6873 (N_6873,N_5766,N_5183);
and U6874 (N_6874,N_4891,N_4784);
nand U6875 (N_6875,N_5035,N_5550);
nand U6876 (N_6876,N_5949,N_5666);
and U6877 (N_6877,N_4636,N_5263);
nand U6878 (N_6878,N_4503,N_5221);
nor U6879 (N_6879,N_5658,N_4452);
nand U6880 (N_6880,N_4265,N_5004);
and U6881 (N_6881,N_5687,N_4653);
nand U6882 (N_6882,N_4447,N_4840);
nor U6883 (N_6883,N_5445,N_5123);
nand U6884 (N_6884,N_5523,N_5496);
or U6885 (N_6885,N_5732,N_5693);
nand U6886 (N_6886,N_5718,N_4945);
and U6887 (N_6887,N_5680,N_5093);
nor U6888 (N_6888,N_5310,N_4097);
nor U6889 (N_6889,N_5373,N_4712);
or U6890 (N_6890,N_4240,N_4805);
or U6891 (N_6891,N_5320,N_4202);
or U6892 (N_6892,N_5336,N_5628);
and U6893 (N_6893,N_4429,N_4139);
nor U6894 (N_6894,N_5582,N_5474);
nand U6895 (N_6895,N_5210,N_5618);
or U6896 (N_6896,N_5172,N_4622);
nand U6897 (N_6897,N_5834,N_4532);
and U6898 (N_6898,N_5574,N_4399);
or U6899 (N_6899,N_4177,N_5450);
and U6900 (N_6900,N_5087,N_5690);
or U6901 (N_6901,N_5851,N_4630);
or U6902 (N_6902,N_4257,N_5518);
nor U6903 (N_6903,N_5128,N_5422);
or U6904 (N_6904,N_5233,N_5640);
nor U6905 (N_6905,N_5825,N_4802);
nor U6906 (N_6906,N_5278,N_4710);
or U6907 (N_6907,N_5584,N_5866);
or U6908 (N_6908,N_4553,N_4965);
nor U6909 (N_6909,N_4477,N_4756);
and U6910 (N_6910,N_4203,N_5685);
and U6911 (N_6911,N_5008,N_5771);
or U6912 (N_6912,N_5089,N_4934);
nor U6913 (N_6913,N_4125,N_5802);
and U6914 (N_6914,N_4930,N_5377);
or U6915 (N_6915,N_4569,N_4069);
nand U6916 (N_6916,N_5209,N_4554);
or U6917 (N_6917,N_5723,N_4416);
nor U6918 (N_6918,N_4469,N_4316);
and U6919 (N_6919,N_5740,N_5153);
or U6920 (N_6920,N_5137,N_4053);
nand U6921 (N_6921,N_4949,N_5318);
and U6922 (N_6922,N_5217,N_5458);
nor U6923 (N_6923,N_5781,N_5695);
or U6924 (N_6924,N_4269,N_5115);
nor U6925 (N_6925,N_5860,N_4185);
and U6926 (N_6926,N_5907,N_4200);
nor U6927 (N_6927,N_5179,N_4092);
xnor U6928 (N_6928,N_5534,N_4624);
and U6929 (N_6929,N_4454,N_5244);
and U6930 (N_6930,N_4334,N_4765);
nand U6931 (N_6931,N_4096,N_4778);
and U6932 (N_6932,N_4560,N_4844);
nor U6933 (N_6933,N_4946,N_5345);
nor U6934 (N_6934,N_4544,N_5170);
or U6935 (N_6935,N_4644,N_5046);
and U6936 (N_6936,N_4356,N_5106);
nor U6937 (N_6937,N_4685,N_4410);
and U6938 (N_6938,N_5142,N_4360);
or U6939 (N_6939,N_4087,N_4280);
nand U6940 (N_6940,N_5499,N_5190);
or U6941 (N_6941,N_5639,N_4978);
nand U6942 (N_6942,N_4692,N_5759);
xor U6943 (N_6943,N_4669,N_4501);
nand U6944 (N_6944,N_4800,N_4164);
nor U6945 (N_6945,N_5829,N_4565);
nor U6946 (N_6946,N_4983,N_5973);
and U6947 (N_6947,N_4843,N_5058);
nor U6948 (N_6948,N_5898,N_5145);
and U6949 (N_6949,N_5094,N_4914);
or U6950 (N_6950,N_4757,N_4885);
or U6951 (N_6951,N_5341,N_5870);
nor U6952 (N_6952,N_5793,N_4213);
and U6953 (N_6953,N_5883,N_4350);
nor U6954 (N_6954,N_5879,N_4673);
nor U6955 (N_6955,N_5225,N_5503);
or U6956 (N_6956,N_5429,N_5537);
or U6957 (N_6957,N_4933,N_5722);
nor U6958 (N_6958,N_4181,N_4487);
or U6959 (N_6959,N_5692,N_5950);
nor U6960 (N_6960,N_4596,N_4941);
nand U6961 (N_6961,N_5904,N_5833);
or U6962 (N_6962,N_5201,N_5729);
nand U6963 (N_6963,N_5161,N_4432);
and U6964 (N_6964,N_5013,N_5548);
nor U6965 (N_6965,N_5791,N_4882);
or U6966 (N_6966,N_5998,N_4059);
nand U6967 (N_6967,N_4297,N_5055);
nand U6968 (N_6968,N_4976,N_5000);
and U6969 (N_6969,N_5997,N_4246);
nand U6970 (N_6970,N_4211,N_4054);
nor U6971 (N_6971,N_5896,N_4238);
nand U6972 (N_6972,N_4592,N_5607);
or U6973 (N_6973,N_5276,N_4247);
or U6974 (N_6974,N_4917,N_5764);
or U6975 (N_6975,N_5776,N_4490);
nor U6976 (N_6976,N_4752,N_4136);
and U6977 (N_6977,N_5188,N_4595);
and U6978 (N_6978,N_4106,N_4923);
nand U6979 (N_6979,N_5969,N_5608);
nor U6980 (N_6980,N_4443,N_4950);
nor U6981 (N_6981,N_4728,N_4465);
or U6982 (N_6982,N_4984,N_5553);
and U6983 (N_6983,N_5564,N_4127);
nand U6984 (N_6984,N_4625,N_5353);
and U6985 (N_6985,N_4378,N_5940);
nor U6986 (N_6986,N_4577,N_5812);
or U6987 (N_6987,N_4696,N_5075);
and U6988 (N_6988,N_4575,N_5412);
nor U6989 (N_6989,N_5673,N_5284);
nor U6990 (N_6990,N_5119,N_5514);
nand U6991 (N_6991,N_4529,N_4870);
nand U6992 (N_6992,N_5813,N_5110);
nor U6993 (N_6993,N_5419,N_4837);
nand U6994 (N_6994,N_5807,N_5505);
nand U6995 (N_6995,N_4146,N_4997);
and U6996 (N_6996,N_5719,N_4626);
or U6997 (N_6997,N_4491,N_5292);
nand U6998 (N_6998,N_4382,N_5481);
nand U6999 (N_6999,N_5181,N_4163);
nand U7000 (N_7000,N_4418,N_4842);
and U7001 (N_7001,N_4021,N_4939);
nand U7002 (N_7002,N_5485,N_4542);
nor U7003 (N_7003,N_5513,N_4741);
nor U7004 (N_7004,N_5404,N_5997);
or U7005 (N_7005,N_5643,N_5719);
and U7006 (N_7006,N_5796,N_4740);
and U7007 (N_7007,N_5195,N_4818);
or U7008 (N_7008,N_5742,N_5351);
and U7009 (N_7009,N_5914,N_4498);
or U7010 (N_7010,N_5535,N_4878);
or U7011 (N_7011,N_5539,N_4629);
nor U7012 (N_7012,N_5658,N_4862);
or U7013 (N_7013,N_5599,N_5867);
and U7014 (N_7014,N_4027,N_4472);
or U7015 (N_7015,N_5310,N_4349);
nor U7016 (N_7016,N_5294,N_5126);
nand U7017 (N_7017,N_4784,N_5521);
and U7018 (N_7018,N_5213,N_5115);
nor U7019 (N_7019,N_5686,N_5301);
and U7020 (N_7020,N_5370,N_5612);
nand U7021 (N_7021,N_5151,N_5967);
nor U7022 (N_7022,N_4550,N_5638);
or U7023 (N_7023,N_5378,N_4528);
and U7024 (N_7024,N_5795,N_4171);
nand U7025 (N_7025,N_5867,N_4023);
or U7026 (N_7026,N_4139,N_5227);
nor U7027 (N_7027,N_4832,N_5732);
and U7028 (N_7028,N_5981,N_4914);
nand U7029 (N_7029,N_4156,N_5647);
xor U7030 (N_7030,N_4520,N_4499);
nand U7031 (N_7031,N_5496,N_5329);
nand U7032 (N_7032,N_5532,N_5538);
and U7033 (N_7033,N_4364,N_4128);
nand U7034 (N_7034,N_5678,N_4160);
and U7035 (N_7035,N_4535,N_4383);
nor U7036 (N_7036,N_5828,N_5523);
or U7037 (N_7037,N_5579,N_5965);
nand U7038 (N_7038,N_4205,N_5376);
or U7039 (N_7039,N_5010,N_5854);
or U7040 (N_7040,N_4278,N_4015);
nand U7041 (N_7041,N_4794,N_4727);
and U7042 (N_7042,N_5604,N_4482);
and U7043 (N_7043,N_4764,N_4025);
or U7044 (N_7044,N_4463,N_5393);
or U7045 (N_7045,N_5246,N_5937);
nand U7046 (N_7046,N_4686,N_4073);
nand U7047 (N_7047,N_4696,N_5142);
nand U7048 (N_7048,N_5221,N_5335);
and U7049 (N_7049,N_4942,N_4794);
xor U7050 (N_7050,N_5281,N_4248);
and U7051 (N_7051,N_5008,N_5893);
or U7052 (N_7052,N_4236,N_4344);
nor U7053 (N_7053,N_5303,N_4863);
nand U7054 (N_7054,N_5115,N_4695);
nor U7055 (N_7055,N_4738,N_5119);
nand U7056 (N_7056,N_4050,N_4046);
nor U7057 (N_7057,N_4129,N_5861);
nand U7058 (N_7058,N_4081,N_5676);
nand U7059 (N_7059,N_4069,N_4176);
nor U7060 (N_7060,N_4765,N_5300);
nand U7061 (N_7061,N_4765,N_5241);
or U7062 (N_7062,N_4788,N_5205);
nor U7063 (N_7063,N_5287,N_4569);
nor U7064 (N_7064,N_4440,N_4742);
or U7065 (N_7065,N_4726,N_4096);
nor U7066 (N_7066,N_4939,N_5859);
and U7067 (N_7067,N_5899,N_4348);
nor U7068 (N_7068,N_4039,N_5791);
nor U7069 (N_7069,N_5981,N_5115);
nor U7070 (N_7070,N_4263,N_5892);
and U7071 (N_7071,N_5375,N_5791);
nand U7072 (N_7072,N_4566,N_4348);
nand U7073 (N_7073,N_5562,N_4258);
nand U7074 (N_7074,N_5380,N_5876);
or U7075 (N_7075,N_4314,N_5320);
nand U7076 (N_7076,N_5666,N_5876);
or U7077 (N_7077,N_4625,N_4878);
and U7078 (N_7078,N_4179,N_5605);
nand U7079 (N_7079,N_5122,N_5465);
nand U7080 (N_7080,N_4948,N_4271);
nor U7081 (N_7081,N_5653,N_5986);
or U7082 (N_7082,N_4497,N_4466);
or U7083 (N_7083,N_5892,N_4920);
and U7084 (N_7084,N_5900,N_5899);
nand U7085 (N_7085,N_5249,N_5023);
nor U7086 (N_7086,N_5258,N_4433);
and U7087 (N_7087,N_5731,N_5134);
nor U7088 (N_7088,N_5086,N_5826);
or U7089 (N_7089,N_5691,N_5934);
and U7090 (N_7090,N_5354,N_4490);
and U7091 (N_7091,N_4234,N_4312);
and U7092 (N_7092,N_5909,N_4298);
nand U7093 (N_7093,N_5088,N_4292);
or U7094 (N_7094,N_5034,N_5843);
or U7095 (N_7095,N_4976,N_4691);
or U7096 (N_7096,N_4435,N_4437);
and U7097 (N_7097,N_4874,N_5732);
nor U7098 (N_7098,N_5084,N_4465);
nand U7099 (N_7099,N_4026,N_5356);
or U7100 (N_7100,N_5845,N_5707);
nor U7101 (N_7101,N_4938,N_4461);
and U7102 (N_7102,N_4479,N_4473);
and U7103 (N_7103,N_4772,N_4719);
or U7104 (N_7104,N_4215,N_5193);
nand U7105 (N_7105,N_4411,N_5913);
nand U7106 (N_7106,N_5915,N_4823);
nor U7107 (N_7107,N_4818,N_5731);
and U7108 (N_7108,N_4711,N_5436);
or U7109 (N_7109,N_5876,N_5963);
nor U7110 (N_7110,N_4503,N_4924);
and U7111 (N_7111,N_4851,N_4229);
and U7112 (N_7112,N_4873,N_5388);
nand U7113 (N_7113,N_4136,N_4919);
or U7114 (N_7114,N_5501,N_5490);
and U7115 (N_7115,N_5293,N_4011);
and U7116 (N_7116,N_5078,N_5868);
xnor U7117 (N_7117,N_5521,N_4527);
nand U7118 (N_7118,N_5733,N_5561);
and U7119 (N_7119,N_5281,N_4243);
or U7120 (N_7120,N_4497,N_5439);
and U7121 (N_7121,N_5082,N_4734);
nand U7122 (N_7122,N_4936,N_5357);
or U7123 (N_7123,N_4821,N_5758);
and U7124 (N_7124,N_5646,N_5421);
or U7125 (N_7125,N_4748,N_5308);
and U7126 (N_7126,N_5874,N_5602);
nand U7127 (N_7127,N_4432,N_5708);
nand U7128 (N_7128,N_4403,N_5822);
nor U7129 (N_7129,N_5015,N_5851);
nand U7130 (N_7130,N_4140,N_5088);
and U7131 (N_7131,N_4543,N_4587);
and U7132 (N_7132,N_4545,N_5628);
and U7133 (N_7133,N_5258,N_4600);
nor U7134 (N_7134,N_4796,N_4171);
or U7135 (N_7135,N_5397,N_5599);
nand U7136 (N_7136,N_4917,N_5910);
or U7137 (N_7137,N_4137,N_4414);
nor U7138 (N_7138,N_4193,N_4196);
nand U7139 (N_7139,N_4230,N_4419);
nand U7140 (N_7140,N_5532,N_4172);
nand U7141 (N_7141,N_4142,N_5429);
nand U7142 (N_7142,N_5192,N_4026);
or U7143 (N_7143,N_5021,N_5875);
or U7144 (N_7144,N_5290,N_5249);
or U7145 (N_7145,N_5987,N_4898);
nand U7146 (N_7146,N_5334,N_4324);
or U7147 (N_7147,N_4065,N_4225);
or U7148 (N_7148,N_5591,N_4481);
nand U7149 (N_7149,N_5932,N_5523);
or U7150 (N_7150,N_4114,N_5819);
or U7151 (N_7151,N_5684,N_4533);
and U7152 (N_7152,N_4512,N_5147);
or U7153 (N_7153,N_4178,N_4291);
nand U7154 (N_7154,N_5995,N_5703);
and U7155 (N_7155,N_5606,N_4850);
or U7156 (N_7156,N_4417,N_4539);
and U7157 (N_7157,N_4369,N_4759);
and U7158 (N_7158,N_5712,N_5132);
nor U7159 (N_7159,N_4023,N_5335);
or U7160 (N_7160,N_5559,N_4039);
nand U7161 (N_7161,N_5162,N_5644);
and U7162 (N_7162,N_4760,N_5290);
or U7163 (N_7163,N_5590,N_5655);
nor U7164 (N_7164,N_5477,N_4142);
nor U7165 (N_7165,N_4949,N_4732);
and U7166 (N_7166,N_4432,N_5462);
nand U7167 (N_7167,N_5872,N_5125);
or U7168 (N_7168,N_4443,N_5096);
or U7169 (N_7169,N_5245,N_5773);
or U7170 (N_7170,N_5780,N_5578);
nor U7171 (N_7171,N_5933,N_4612);
and U7172 (N_7172,N_4732,N_5202);
and U7173 (N_7173,N_5345,N_4558);
or U7174 (N_7174,N_5393,N_5178);
nor U7175 (N_7175,N_5662,N_5527);
and U7176 (N_7176,N_5944,N_5565);
nand U7177 (N_7177,N_5522,N_4259);
nor U7178 (N_7178,N_5646,N_5765);
xor U7179 (N_7179,N_5940,N_5838);
nand U7180 (N_7180,N_5049,N_5267);
or U7181 (N_7181,N_4914,N_5101);
nand U7182 (N_7182,N_4462,N_4336);
nand U7183 (N_7183,N_4229,N_4941);
nand U7184 (N_7184,N_4217,N_5939);
or U7185 (N_7185,N_4806,N_4555);
nor U7186 (N_7186,N_5585,N_5721);
or U7187 (N_7187,N_4402,N_4700);
nand U7188 (N_7188,N_4269,N_5204);
nor U7189 (N_7189,N_5108,N_5345);
nor U7190 (N_7190,N_4144,N_5983);
and U7191 (N_7191,N_4103,N_4790);
nand U7192 (N_7192,N_5614,N_5706);
nand U7193 (N_7193,N_5930,N_4173);
nand U7194 (N_7194,N_5882,N_4008);
and U7195 (N_7195,N_4330,N_4128);
or U7196 (N_7196,N_5763,N_5249);
nor U7197 (N_7197,N_5462,N_4352);
nor U7198 (N_7198,N_5508,N_5869);
nor U7199 (N_7199,N_5244,N_4615);
and U7200 (N_7200,N_5011,N_4681);
or U7201 (N_7201,N_4375,N_4386);
and U7202 (N_7202,N_5614,N_4902);
nand U7203 (N_7203,N_5486,N_4386);
or U7204 (N_7204,N_5865,N_5162);
nand U7205 (N_7205,N_4258,N_4014);
nand U7206 (N_7206,N_5295,N_5302);
or U7207 (N_7207,N_5469,N_5500);
or U7208 (N_7208,N_4688,N_5005);
or U7209 (N_7209,N_5267,N_4553);
nand U7210 (N_7210,N_5142,N_5853);
nand U7211 (N_7211,N_5936,N_4682);
nor U7212 (N_7212,N_4387,N_4152);
and U7213 (N_7213,N_4828,N_5954);
nand U7214 (N_7214,N_5463,N_4470);
and U7215 (N_7215,N_4670,N_4449);
or U7216 (N_7216,N_5620,N_4979);
nand U7217 (N_7217,N_5916,N_4916);
xor U7218 (N_7218,N_4612,N_5178);
or U7219 (N_7219,N_5509,N_5418);
xor U7220 (N_7220,N_4740,N_4886);
or U7221 (N_7221,N_4568,N_4276);
and U7222 (N_7222,N_5279,N_4902);
or U7223 (N_7223,N_4561,N_5090);
or U7224 (N_7224,N_5545,N_4835);
and U7225 (N_7225,N_5662,N_4748);
or U7226 (N_7226,N_4784,N_5552);
nand U7227 (N_7227,N_5394,N_4169);
nor U7228 (N_7228,N_4103,N_4542);
or U7229 (N_7229,N_5621,N_5623);
nand U7230 (N_7230,N_5286,N_5750);
nand U7231 (N_7231,N_4287,N_5643);
nand U7232 (N_7232,N_4977,N_4883);
or U7233 (N_7233,N_4653,N_4510);
nand U7234 (N_7234,N_5947,N_4260);
or U7235 (N_7235,N_4079,N_4713);
and U7236 (N_7236,N_5260,N_4813);
nor U7237 (N_7237,N_4022,N_5295);
and U7238 (N_7238,N_4829,N_5171);
or U7239 (N_7239,N_5713,N_4652);
and U7240 (N_7240,N_4088,N_5868);
and U7241 (N_7241,N_4938,N_5050);
or U7242 (N_7242,N_5744,N_5734);
or U7243 (N_7243,N_5016,N_4023);
nand U7244 (N_7244,N_4577,N_4067);
or U7245 (N_7245,N_5285,N_4726);
nand U7246 (N_7246,N_4887,N_5600);
and U7247 (N_7247,N_5216,N_4939);
and U7248 (N_7248,N_5276,N_4515);
and U7249 (N_7249,N_4280,N_5001);
nand U7250 (N_7250,N_4647,N_4385);
nand U7251 (N_7251,N_5843,N_5817);
nor U7252 (N_7252,N_5938,N_5195);
nand U7253 (N_7253,N_4699,N_4517);
and U7254 (N_7254,N_5966,N_5106);
or U7255 (N_7255,N_5990,N_4948);
and U7256 (N_7256,N_5266,N_5500);
and U7257 (N_7257,N_4343,N_5471);
and U7258 (N_7258,N_4891,N_4209);
nand U7259 (N_7259,N_4266,N_4106);
nand U7260 (N_7260,N_4481,N_4376);
nand U7261 (N_7261,N_4280,N_5306);
nor U7262 (N_7262,N_4391,N_5260);
nor U7263 (N_7263,N_4598,N_5339);
and U7264 (N_7264,N_5341,N_4429);
and U7265 (N_7265,N_5034,N_5170);
or U7266 (N_7266,N_4200,N_4899);
or U7267 (N_7267,N_4800,N_5983);
or U7268 (N_7268,N_5490,N_4870);
nand U7269 (N_7269,N_5865,N_5549);
or U7270 (N_7270,N_5552,N_4309);
nor U7271 (N_7271,N_4460,N_4132);
and U7272 (N_7272,N_4037,N_5172);
nor U7273 (N_7273,N_5239,N_5293);
and U7274 (N_7274,N_5089,N_5104);
and U7275 (N_7275,N_5969,N_4039);
or U7276 (N_7276,N_4631,N_4121);
and U7277 (N_7277,N_5156,N_4637);
and U7278 (N_7278,N_5757,N_5548);
and U7279 (N_7279,N_4529,N_5526);
nand U7280 (N_7280,N_4499,N_4783);
xor U7281 (N_7281,N_4358,N_4852);
nor U7282 (N_7282,N_5262,N_5087);
or U7283 (N_7283,N_5015,N_4406);
nand U7284 (N_7284,N_5397,N_5766);
nand U7285 (N_7285,N_4660,N_4870);
nand U7286 (N_7286,N_5913,N_4390);
and U7287 (N_7287,N_5487,N_5078);
nor U7288 (N_7288,N_5144,N_4776);
nand U7289 (N_7289,N_4946,N_5114);
or U7290 (N_7290,N_5338,N_5974);
nor U7291 (N_7291,N_5256,N_4436);
or U7292 (N_7292,N_4345,N_5774);
xor U7293 (N_7293,N_5826,N_5141);
nor U7294 (N_7294,N_4125,N_5081);
and U7295 (N_7295,N_4736,N_4141);
nand U7296 (N_7296,N_5559,N_5948);
nand U7297 (N_7297,N_5636,N_5429);
and U7298 (N_7298,N_5842,N_4520);
nor U7299 (N_7299,N_4618,N_5437);
and U7300 (N_7300,N_5118,N_4336);
and U7301 (N_7301,N_4812,N_5956);
nor U7302 (N_7302,N_5795,N_5598);
xnor U7303 (N_7303,N_4941,N_4554);
and U7304 (N_7304,N_4486,N_5187);
nor U7305 (N_7305,N_5197,N_4164);
nor U7306 (N_7306,N_4804,N_4056);
or U7307 (N_7307,N_4000,N_5024);
and U7308 (N_7308,N_4868,N_5702);
or U7309 (N_7309,N_5032,N_4115);
or U7310 (N_7310,N_4478,N_4638);
and U7311 (N_7311,N_5742,N_4896);
or U7312 (N_7312,N_5105,N_5268);
or U7313 (N_7313,N_5355,N_5665);
nand U7314 (N_7314,N_4202,N_5622);
nand U7315 (N_7315,N_4431,N_4333);
nor U7316 (N_7316,N_4289,N_5922);
nand U7317 (N_7317,N_5150,N_5931);
or U7318 (N_7318,N_5884,N_5952);
nand U7319 (N_7319,N_4183,N_5072);
nor U7320 (N_7320,N_4504,N_5465);
nand U7321 (N_7321,N_4009,N_4595);
nor U7322 (N_7322,N_5301,N_5754);
or U7323 (N_7323,N_5057,N_5590);
nand U7324 (N_7324,N_5235,N_5058);
or U7325 (N_7325,N_5538,N_5202);
and U7326 (N_7326,N_4802,N_5357);
or U7327 (N_7327,N_4687,N_5587);
nand U7328 (N_7328,N_5218,N_4836);
nor U7329 (N_7329,N_4119,N_4236);
nand U7330 (N_7330,N_4586,N_4463);
nand U7331 (N_7331,N_5932,N_4648);
and U7332 (N_7332,N_4647,N_4891);
or U7333 (N_7333,N_5347,N_5318);
xnor U7334 (N_7334,N_5588,N_4747);
and U7335 (N_7335,N_4067,N_5976);
nor U7336 (N_7336,N_4487,N_4784);
and U7337 (N_7337,N_5635,N_4983);
nor U7338 (N_7338,N_5009,N_5380);
and U7339 (N_7339,N_5617,N_4359);
nand U7340 (N_7340,N_5271,N_4291);
and U7341 (N_7341,N_4174,N_5462);
or U7342 (N_7342,N_4647,N_4461);
and U7343 (N_7343,N_5490,N_5045);
nor U7344 (N_7344,N_4953,N_4829);
or U7345 (N_7345,N_5886,N_4733);
nor U7346 (N_7346,N_5285,N_5626);
or U7347 (N_7347,N_5409,N_5987);
nor U7348 (N_7348,N_5389,N_4852);
nand U7349 (N_7349,N_4066,N_4473);
nand U7350 (N_7350,N_4916,N_5416);
nor U7351 (N_7351,N_5922,N_4096);
nand U7352 (N_7352,N_5249,N_5200);
and U7353 (N_7353,N_4853,N_5166);
or U7354 (N_7354,N_4409,N_5777);
nor U7355 (N_7355,N_5208,N_4284);
or U7356 (N_7356,N_5792,N_5026);
nor U7357 (N_7357,N_5186,N_4631);
or U7358 (N_7358,N_5769,N_5367);
or U7359 (N_7359,N_4374,N_5804);
nor U7360 (N_7360,N_5024,N_5248);
nor U7361 (N_7361,N_5356,N_4881);
xor U7362 (N_7362,N_5037,N_4076);
and U7363 (N_7363,N_4021,N_5194);
nor U7364 (N_7364,N_5283,N_4477);
or U7365 (N_7365,N_4746,N_5950);
nor U7366 (N_7366,N_4623,N_5769);
or U7367 (N_7367,N_4927,N_5695);
nor U7368 (N_7368,N_5802,N_4052);
or U7369 (N_7369,N_5724,N_4732);
nor U7370 (N_7370,N_5610,N_5993);
and U7371 (N_7371,N_5008,N_5871);
nor U7372 (N_7372,N_5112,N_4352);
nor U7373 (N_7373,N_5836,N_5383);
nand U7374 (N_7374,N_5293,N_4246);
or U7375 (N_7375,N_5803,N_4300);
nand U7376 (N_7376,N_5490,N_5990);
nand U7377 (N_7377,N_5594,N_4247);
and U7378 (N_7378,N_5601,N_5497);
or U7379 (N_7379,N_4075,N_4644);
or U7380 (N_7380,N_4670,N_4437);
nor U7381 (N_7381,N_4522,N_5025);
or U7382 (N_7382,N_5982,N_4462);
nor U7383 (N_7383,N_4649,N_4094);
or U7384 (N_7384,N_5045,N_4442);
and U7385 (N_7385,N_4534,N_5297);
and U7386 (N_7386,N_5443,N_5389);
or U7387 (N_7387,N_5936,N_5093);
and U7388 (N_7388,N_5345,N_5153);
or U7389 (N_7389,N_4899,N_4276);
or U7390 (N_7390,N_4071,N_5229);
or U7391 (N_7391,N_5228,N_4018);
and U7392 (N_7392,N_5434,N_5613);
and U7393 (N_7393,N_4206,N_5898);
nor U7394 (N_7394,N_4367,N_5342);
xor U7395 (N_7395,N_5137,N_4476);
nor U7396 (N_7396,N_5200,N_4987);
nor U7397 (N_7397,N_4254,N_4096);
and U7398 (N_7398,N_4710,N_5500);
or U7399 (N_7399,N_4711,N_5275);
and U7400 (N_7400,N_5127,N_4359);
nand U7401 (N_7401,N_5574,N_4557);
nor U7402 (N_7402,N_5050,N_5414);
and U7403 (N_7403,N_4269,N_5656);
and U7404 (N_7404,N_4304,N_5148);
or U7405 (N_7405,N_5457,N_4278);
nand U7406 (N_7406,N_4626,N_5108);
nand U7407 (N_7407,N_4108,N_4201);
nor U7408 (N_7408,N_5756,N_5380);
nand U7409 (N_7409,N_5816,N_5290);
nand U7410 (N_7410,N_5001,N_5339);
nor U7411 (N_7411,N_5827,N_4321);
nand U7412 (N_7412,N_4150,N_4082);
or U7413 (N_7413,N_5721,N_5402);
nor U7414 (N_7414,N_4390,N_5441);
nor U7415 (N_7415,N_4400,N_4700);
and U7416 (N_7416,N_5857,N_5371);
nand U7417 (N_7417,N_4265,N_5204);
and U7418 (N_7418,N_4412,N_4674);
nor U7419 (N_7419,N_4285,N_5626);
or U7420 (N_7420,N_5034,N_4863);
or U7421 (N_7421,N_5303,N_4772);
or U7422 (N_7422,N_4875,N_5705);
nor U7423 (N_7423,N_5676,N_5023);
or U7424 (N_7424,N_4091,N_5616);
or U7425 (N_7425,N_5594,N_5211);
or U7426 (N_7426,N_5733,N_4767);
and U7427 (N_7427,N_5427,N_4252);
and U7428 (N_7428,N_5306,N_5032);
nand U7429 (N_7429,N_5233,N_5425);
or U7430 (N_7430,N_5467,N_5025);
nor U7431 (N_7431,N_5542,N_5583);
or U7432 (N_7432,N_5841,N_5105);
nor U7433 (N_7433,N_5255,N_5868);
nor U7434 (N_7434,N_5495,N_4952);
nand U7435 (N_7435,N_5965,N_4178);
nor U7436 (N_7436,N_5654,N_4021);
and U7437 (N_7437,N_4562,N_4214);
nand U7438 (N_7438,N_5644,N_4889);
or U7439 (N_7439,N_5862,N_4675);
and U7440 (N_7440,N_4762,N_5737);
or U7441 (N_7441,N_4934,N_4873);
nand U7442 (N_7442,N_4737,N_4064);
and U7443 (N_7443,N_4539,N_5629);
nand U7444 (N_7444,N_4952,N_4398);
or U7445 (N_7445,N_4960,N_5342);
and U7446 (N_7446,N_4445,N_4678);
nand U7447 (N_7447,N_5370,N_5475);
nand U7448 (N_7448,N_4329,N_4705);
and U7449 (N_7449,N_5656,N_4635);
and U7450 (N_7450,N_5153,N_5581);
or U7451 (N_7451,N_4390,N_4678);
or U7452 (N_7452,N_4470,N_4665);
and U7453 (N_7453,N_5826,N_4287);
nand U7454 (N_7454,N_4392,N_4825);
nor U7455 (N_7455,N_4997,N_5011);
xnor U7456 (N_7456,N_4478,N_5327);
nor U7457 (N_7457,N_5020,N_4857);
nor U7458 (N_7458,N_5179,N_4169);
nand U7459 (N_7459,N_4921,N_4294);
or U7460 (N_7460,N_5295,N_4320);
or U7461 (N_7461,N_4673,N_5470);
or U7462 (N_7462,N_4076,N_5038);
nand U7463 (N_7463,N_4934,N_5364);
nor U7464 (N_7464,N_5649,N_5115);
nand U7465 (N_7465,N_4922,N_4728);
nor U7466 (N_7466,N_4406,N_4008);
or U7467 (N_7467,N_4969,N_4291);
nand U7468 (N_7468,N_4221,N_4171);
or U7469 (N_7469,N_4591,N_5372);
nand U7470 (N_7470,N_4114,N_4187);
or U7471 (N_7471,N_5410,N_4450);
or U7472 (N_7472,N_5214,N_5537);
nand U7473 (N_7473,N_4493,N_5962);
or U7474 (N_7474,N_5883,N_5098);
nand U7475 (N_7475,N_5112,N_5858);
nor U7476 (N_7476,N_4972,N_5370);
nand U7477 (N_7477,N_5732,N_5119);
nor U7478 (N_7478,N_5457,N_5235);
and U7479 (N_7479,N_4096,N_4377);
and U7480 (N_7480,N_5889,N_4303);
nand U7481 (N_7481,N_5596,N_5631);
or U7482 (N_7482,N_4111,N_5549);
nor U7483 (N_7483,N_4387,N_5839);
nand U7484 (N_7484,N_4585,N_4086);
xor U7485 (N_7485,N_4366,N_5902);
nor U7486 (N_7486,N_5626,N_5477);
or U7487 (N_7487,N_5607,N_4019);
and U7488 (N_7488,N_5201,N_5233);
nand U7489 (N_7489,N_4341,N_5401);
nor U7490 (N_7490,N_5889,N_5648);
nand U7491 (N_7491,N_4199,N_5043);
nand U7492 (N_7492,N_5496,N_5044);
nor U7493 (N_7493,N_5124,N_4961);
nor U7494 (N_7494,N_5286,N_4137);
nand U7495 (N_7495,N_4229,N_4881);
nand U7496 (N_7496,N_4203,N_5272);
nor U7497 (N_7497,N_5762,N_4369);
and U7498 (N_7498,N_5405,N_5980);
and U7499 (N_7499,N_5651,N_5585);
nor U7500 (N_7500,N_4187,N_5567);
or U7501 (N_7501,N_4529,N_4117);
or U7502 (N_7502,N_5649,N_5534);
nand U7503 (N_7503,N_5083,N_4294);
nand U7504 (N_7504,N_4395,N_4117);
and U7505 (N_7505,N_5783,N_5507);
or U7506 (N_7506,N_5039,N_5885);
nor U7507 (N_7507,N_5253,N_5519);
or U7508 (N_7508,N_5324,N_5594);
nor U7509 (N_7509,N_5140,N_5862);
or U7510 (N_7510,N_4832,N_4502);
nand U7511 (N_7511,N_4155,N_4855);
nor U7512 (N_7512,N_5341,N_4969);
nand U7513 (N_7513,N_5514,N_4298);
or U7514 (N_7514,N_4342,N_5022);
nand U7515 (N_7515,N_5416,N_5403);
nand U7516 (N_7516,N_4580,N_5488);
or U7517 (N_7517,N_5372,N_5090);
nor U7518 (N_7518,N_5406,N_5597);
nor U7519 (N_7519,N_5190,N_5168);
and U7520 (N_7520,N_4955,N_5280);
nor U7521 (N_7521,N_4377,N_5735);
nand U7522 (N_7522,N_5546,N_5423);
nand U7523 (N_7523,N_5619,N_5467);
or U7524 (N_7524,N_4206,N_5741);
and U7525 (N_7525,N_5107,N_5611);
nor U7526 (N_7526,N_4591,N_4029);
and U7527 (N_7527,N_4636,N_4557);
xor U7528 (N_7528,N_5933,N_5565);
nand U7529 (N_7529,N_4244,N_5556);
nor U7530 (N_7530,N_5295,N_5660);
nand U7531 (N_7531,N_5740,N_4743);
nand U7532 (N_7532,N_4300,N_5383);
nand U7533 (N_7533,N_4429,N_5773);
nor U7534 (N_7534,N_5308,N_4308);
and U7535 (N_7535,N_5917,N_4373);
or U7536 (N_7536,N_4799,N_5401);
or U7537 (N_7537,N_4567,N_4118);
or U7538 (N_7538,N_5961,N_5068);
or U7539 (N_7539,N_4964,N_5303);
nor U7540 (N_7540,N_4216,N_5982);
nand U7541 (N_7541,N_4666,N_4474);
nand U7542 (N_7542,N_4100,N_4150);
or U7543 (N_7543,N_4196,N_4632);
nand U7544 (N_7544,N_4941,N_4715);
or U7545 (N_7545,N_4816,N_4748);
or U7546 (N_7546,N_4057,N_5572);
nor U7547 (N_7547,N_5318,N_4660);
nor U7548 (N_7548,N_4739,N_4636);
and U7549 (N_7549,N_4374,N_4555);
and U7550 (N_7550,N_4148,N_4931);
and U7551 (N_7551,N_4861,N_5344);
or U7552 (N_7552,N_4320,N_4486);
and U7553 (N_7553,N_5471,N_5949);
nor U7554 (N_7554,N_4970,N_5491);
nand U7555 (N_7555,N_5781,N_5250);
nor U7556 (N_7556,N_4823,N_5877);
and U7557 (N_7557,N_4603,N_5421);
nand U7558 (N_7558,N_4109,N_5284);
nand U7559 (N_7559,N_5813,N_5075);
and U7560 (N_7560,N_5887,N_4144);
and U7561 (N_7561,N_4354,N_5516);
nand U7562 (N_7562,N_4262,N_5040);
nand U7563 (N_7563,N_4100,N_4992);
or U7564 (N_7564,N_4055,N_4814);
nor U7565 (N_7565,N_4509,N_4350);
or U7566 (N_7566,N_5117,N_4687);
and U7567 (N_7567,N_4841,N_5472);
or U7568 (N_7568,N_5896,N_5212);
nor U7569 (N_7569,N_4806,N_5404);
nand U7570 (N_7570,N_4967,N_5649);
nand U7571 (N_7571,N_5041,N_4995);
nor U7572 (N_7572,N_4734,N_5345);
xor U7573 (N_7573,N_5141,N_5522);
nor U7574 (N_7574,N_5728,N_4172);
nand U7575 (N_7575,N_5322,N_4290);
nand U7576 (N_7576,N_5163,N_5612);
nand U7577 (N_7577,N_5289,N_4120);
xor U7578 (N_7578,N_5124,N_5343);
nor U7579 (N_7579,N_5455,N_4768);
or U7580 (N_7580,N_4297,N_4893);
and U7581 (N_7581,N_4674,N_4772);
nand U7582 (N_7582,N_5110,N_5643);
and U7583 (N_7583,N_4427,N_5460);
nor U7584 (N_7584,N_4916,N_5810);
and U7585 (N_7585,N_5341,N_5896);
and U7586 (N_7586,N_5244,N_5282);
nor U7587 (N_7587,N_4770,N_4580);
nor U7588 (N_7588,N_5802,N_5101);
or U7589 (N_7589,N_5585,N_5130);
or U7590 (N_7590,N_4840,N_5582);
nor U7591 (N_7591,N_5453,N_4450);
nor U7592 (N_7592,N_4736,N_4914);
or U7593 (N_7593,N_5467,N_4696);
nor U7594 (N_7594,N_4315,N_5659);
or U7595 (N_7595,N_5399,N_4160);
nor U7596 (N_7596,N_5382,N_4976);
xnor U7597 (N_7597,N_5954,N_4271);
xor U7598 (N_7598,N_5004,N_5203);
and U7599 (N_7599,N_4376,N_5836);
and U7600 (N_7600,N_4246,N_4228);
or U7601 (N_7601,N_4386,N_4842);
and U7602 (N_7602,N_4366,N_5561);
and U7603 (N_7603,N_5421,N_4706);
nand U7604 (N_7604,N_4886,N_4507);
nor U7605 (N_7605,N_5793,N_4602);
or U7606 (N_7606,N_5387,N_4142);
or U7607 (N_7607,N_5085,N_4856);
nor U7608 (N_7608,N_4885,N_5631);
nor U7609 (N_7609,N_5390,N_5006);
nand U7610 (N_7610,N_5464,N_5734);
or U7611 (N_7611,N_4859,N_5652);
nor U7612 (N_7612,N_5051,N_4817);
or U7613 (N_7613,N_4454,N_5070);
and U7614 (N_7614,N_4620,N_4901);
nor U7615 (N_7615,N_5818,N_5089);
and U7616 (N_7616,N_5396,N_5072);
xnor U7617 (N_7617,N_4227,N_4689);
nor U7618 (N_7618,N_5491,N_5867);
nor U7619 (N_7619,N_4907,N_5342);
and U7620 (N_7620,N_5130,N_4594);
nor U7621 (N_7621,N_5167,N_4651);
or U7622 (N_7622,N_4768,N_4041);
or U7623 (N_7623,N_5991,N_4206);
and U7624 (N_7624,N_5784,N_4800);
or U7625 (N_7625,N_4315,N_5129);
and U7626 (N_7626,N_4699,N_4512);
or U7627 (N_7627,N_4352,N_4912);
and U7628 (N_7628,N_5544,N_4959);
nor U7629 (N_7629,N_4865,N_5599);
or U7630 (N_7630,N_4942,N_5550);
nor U7631 (N_7631,N_5180,N_5245);
nand U7632 (N_7632,N_4098,N_4730);
xor U7633 (N_7633,N_4203,N_4453);
and U7634 (N_7634,N_5693,N_4065);
nand U7635 (N_7635,N_5419,N_4063);
nor U7636 (N_7636,N_4013,N_5400);
xnor U7637 (N_7637,N_5571,N_5457);
and U7638 (N_7638,N_4240,N_4550);
and U7639 (N_7639,N_4162,N_5008);
nor U7640 (N_7640,N_5626,N_4365);
and U7641 (N_7641,N_5494,N_4483);
nand U7642 (N_7642,N_5944,N_4467);
nor U7643 (N_7643,N_5583,N_4560);
xnor U7644 (N_7644,N_4833,N_4248);
or U7645 (N_7645,N_4543,N_4178);
nand U7646 (N_7646,N_5487,N_5872);
and U7647 (N_7647,N_5050,N_4141);
xor U7648 (N_7648,N_5274,N_4506);
xor U7649 (N_7649,N_5252,N_4896);
or U7650 (N_7650,N_4173,N_4791);
xor U7651 (N_7651,N_5390,N_5861);
and U7652 (N_7652,N_5870,N_5716);
nand U7653 (N_7653,N_5910,N_4466);
nor U7654 (N_7654,N_4281,N_5747);
nor U7655 (N_7655,N_5734,N_4039);
nand U7656 (N_7656,N_4062,N_4844);
nor U7657 (N_7657,N_4994,N_4249);
xor U7658 (N_7658,N_5552,N_5258);
nand U7659 (N_7659,N_5796,N_5545);
or U7660 (N_7660,N_5633,N_5251);
nand U7661 (N_7661,N_5869,N_5152);
or U7662 (N_7662,N_5277,N_5946);
nand U7663 (N_7663,N_4133,N_4495);
nor U7664 (N_7664,N_5667,N_5058);
nand U7665 (N_7665,N_4464,N_5227);
nand U7666 (N_7666,N_4502,N_4669);
nand U7667 (N_7667,N_4224,N_5446);
nor U7668 (N_7668,N_5188,N_4484);
and U7669 (N_7669,N_5656,N_5692);
xnor U7670 (N_7670,N_4137,N_5085);
or U7671 (N_7671,N_5879,N_4158);
nand U7672 (N_7672,N_4486,N_4289);
nor U7673 (N_7673,N_5084,N_4108);
and U7674 (N_7674,N_4246,N_4127);
nor U7675 (N_7675,N_4230,N_5936);
nand U7676 (N_7676,N_5247,N_5681);
nor U7677 (N_7677,N_5121,N_5152);
nand U7678 (N_7678,N_5321,N_5802);
and U7679 (N_7679,N_5592,N_5336);
nand U7680 (N_7680,N_5997,N_5334);
and U7681 (N_7681,N_4419,N_5483);
nor U7682 (N_7682,N_5000,N_4647);
nand U7683 (N_7683,N_5516,N_4242);
nor U7684 (N_7684,N_4228,N_5450);
nor U7685 (N_7685,N_5412,N_4830);
and U7686 (N_7686,N_4023,N_4540);
or U7687 (N_7687,N_4516,N_5598);
nand U7688 (N_7688,N_5151,N_4143);
or U7689 (N_7689,N_4015,N_5470);
nand U7690 (N_7690,N_5922,N_4211);
or U7691 (N_7691,N_4134,N_4969);
and U7692 (N_7692,N_4531,N_5367);
or U7693 (N_7693,N_4971,N_5789);
or U7694 (N_7694,N_5608,N_4116);
nand U7695 (N_7695,N_5039,N_4880);
or U7696 (N_7696,N_4132,N_5158);
xnor U7697 (N_7697,N_5613,N_5924);
and U7698 (N_7698,N_5309,N_5324);
and U7699 (N_7699,N_4729,N_4943);
or U7700 (N_7700,N_5916,N_5627);
and U7701 (N_7701,N_4869,N_4180);
and U7702 (N_7702,N_5909,N_5159);
and U7703 (N_7703,N_5505,N_5208);
or U7704 (N_7704,N_4283,N_5514);
and U7705 (N_7705,N_5929,N_5012);
nor U7706 (N_7706,N_5379,N_4937);
or U7707 (N_7707,N_4434,N_4849);
nor U7708 (N_7708,N_4204,N_5299);
nand U7709 (N_7709,N_5828,N_5315);
nor U7710 (N_7710,N_4060,N_4322);
or U7711 (N_7711,N_5261,N_4807);
and U7712 (N_7712,N_5940,N_4864);
or U7713 (N_7713,N_5264,N_5159);
or U7714 (N_7714,N_5938,N_4186);
nand U7715 (N_7715,N_5832,N_5861);
nor U7716 (N_7716,N_4033,N_5161);
nor U7717 (N_7717,N_5945,N_5311);
or U7718 (N_7718,N_4725,N_5851);
nor U7719 (N_7719,N_4237,N_5691);
nand U7720 (N_7720,N_4205,N_5124);
and U7721 (N_7721,N_4520,N_5619);
and U7722 (N_7722,N_4574,N_4764);
nor U7723 (N_7723,N_5658,N_5805);
nor U7724 (N_7724,N_5974,N_5267);
nor U7725 (N_7725,N_5080,N_5169);
nand U7726 (N_7726,N_4354,N_4682);
and U7727 (N_7727,N_5390,N_5258);
or U7728 (N_7728,N_4804,N_4290);
nor U7729 (N_7729,N_5851,N_5650);
nor U7730 (N_7730,N_4036,N_4718);
nor U7731 (N_7731,N_5413,N_4907);
nor U7732 (N_7732,N_4414,N_4791);
or U7733 (N_7733,N_4234,N_4104);
nor U7734 (N_7734,N_5633,N_5481);
nor U7735 (N_7735,N_4400,N_5315);
nor U7736 (N_7736,N_5560,N_5344);
or U7737 (N_7737,N_5097,N_4820);
or U7738 (N_7738,N_4180,N_4724);
and U7739 (N_7739,N_5226,N_4138);
or U7740 (N_7740,N_5548,N_5736);
or U7741 (N_7741,N_5813,N_5323);
or U7742 (N_7742,N_5174,N_5235);
or U7743 (N_7743,N_4056,N_5586);
nand U7744 (N_7744,N_5984,N_5250);
and U7745 (N_7745,N_5789,N_4443);
nor U7746 (N_7746,N_5332,N_4747);
xor U7747 (N_7747,N_4263,N_5604);
and U7748 (N_7748,N_4646,N_4411);
nand U7749 (N_7749,N_4233,N_4237);
and U7750 (N_7750,N_4168,N_4629);
or U7751 (N_7751,N_4705,N_4935);
nor U7752 (N_7752,N_4946,N_5765);
nor U7753 (N_7753,N_5263,N_4265);
or U7754 (N_7754,N_4989,N_5631);
or U7755 (N_7755,N_5445,N_4972);
or U7756 (N_7756,N_5325,N_4646);
nor U7757 (N_7757,N_5858,N_4641);
or U7758 (N_7758,N_4490,N_5963);
nor U7759 (N_7759,N_4460,N_5237);
or U7760 (N_7760,N_4676,N_4882);
and U7761 (N_7761,N_5574,N_5716);
nand U7762 (N_7762,N_4389,N_5280);
or U7763 (N_7763,N_5164,N_4988);
xnor U7764 (N_7764,N_4244,N_4081);
and U7765 (N_7765,N_5778,N_5895);
and U7766 (N_7766,N_4922,N_4650);
and U7767 (N_7767,N_5364,N_5380);
and U7768 (N_7768,N_5419,N_4023);
nor U7769 (N_7769,N_4920,N_5114);
and U7770 (N_7770,N_4801,N_4368);
and U7771 (N_7771,N_4682,N_5175);
nand U7772 (N_7772,N_5540,N_5936);
or U7773 (N_7773,N_4811,N_5249);
nor U7774 (N_7774,N_4092,N_5950);
nand U7775 (N_7775,N_4112,N_4889);
nor U7776 (N_7776,N_4494,N_4945);
nor U7777 (N_7777,N_4163,N_5455);
nand U7778 (N_7778,N_5444,N_4952);
or U7779 (N_7779,N_4686,N_4027);
nor U7780 (N_7780,N_4099,N_5031);
or U7781 (N_7781,N_4074,N_5926);
nand U7782 (N_7782,N_4698,N_4147);
nand U7783 (N_7783,N_5414,N_4045);
nand U7784 (N_7784,N_4889,N_4354);
xor U7785 (N_7785,N_5064,N_4008);
nor U7786 (N_7786,N_5310,N_4440);
nand U7787 (N_7787,N_5164,N_5760);
nand U7788 (N_7788,N_4517,N_4044);
or U7789 (N_7789,N_5200,N_5435);
nand U7790 (N_7790,N_4206,N_4915);
xor U7791 (N_7791,N_5534,N_4654);
nand U7792 (N_7792,N_4732,N_5264);
or U7793 (N_7793,N_5287,N_4858);
or U7794 (N_7794,N_5842,N_5040);
or U7795 (N_7795,N_4751,N_5610);
nand U7796 (N_7796,N_5499,N_5039);
nor U7797 (N_7797,N_4445,N_5164);
nor U7798 (N_7798,N_4535,N_4360);
or U7799 (N_7799,N_5275,N_4067);
or U7800 (N_7800,N_4431,N_5356);
nand U7801 (N_7801,N_4927,N_4394);
xor U7802 (N_7802,N_4217,N_5958);
or U7803 (N_7803,N_5413,N_5430);
or U7804 (N_7804,N_5787,N_4240);
and U7805 (N_7805,N_4310,N_5906);
or U7806 (N_7806,N_4132,N_5011);
or U7807 (N_7807,N_5393,N_5547);
or U7808 (N_7808,N_4834,N_5605);
or U7809 (N_7809,N_4628,N_5486);
nor U7810 (N_7810,N_5513,N_5805);
nor U7811 (N_7811,N_4369,N_5993);
and U7812 (N_7812,N_5340,N_4934);
nand U7813 (N_7813,N_5447,N_5304);
and U7814 (N_7814,N_4623,N_4539);
nor U7815 (N_7815,N_5260,N_4328);
nand U7816 (N_7816,N_5827,N_5368);
and U7817 (N_7817,N_5622,N_5120);
or U7818 (N_7818,N_4275,N_5197);
or U7819 (N_7819,N_5050,N_4747);
and U7820 (N_7820,N_5695,N_4819);
nand U7821 (N_7821,N_4020,N_5216);
xnor U7822 (N_7822,N_4532,N_4479);
nor U7823 (N_7823,N_5870,N_4159);
nand U7824 (N_7824,N_4717,N_4763);
nor U7825 (N_7825,N_5021,N_4132);
nor U7826 (N_7826,N_4491,N_4668);
nand U7827 (N_7827,N_4978,N_5717);
or U7828 (N_7828,N_5704,N_5992);
and U7829 (N_7829,N_5635,N_4211);
nor U7830 (N_7830,N_5074,N_4728);
and U7831 (N_7831,N_4813,N_5038);
nand U7832 (N_7832,N_4077,N_5669);
and U7833 (N_7833,N_5885,N_4034);
nor U7834 (N_7834,N_5753,N_4184);
and U7835 (N_7835,N_4108,N_4492);
and U7836 (N_7836,N_5943,N_5919);
and U7837 (N_7837,N_4793,N_5087);
or U7838 (N_7838,N_5445,N_4885);
nor U7839 (N_7839,N_4902,N_5828);
nand U7840 (N_7840,N_5509,N_5229);
and U7841 (N_7841,N_5663,N_4622);
or U7842 (N_7842,N_4058,N_5652);
or U7843 (N_7843,N_4071,N_4637);
nor U7844 (N_7844,N_4564,N_4887);
or U7845 (N_7845,N_4098,N_4524);
and U7846 (N_7846,N_4783,N_4468);
and U7847 (N_7847,N_4837,N_4365);
nand U7848 (N_7848,N_4299,N_5090);
nand U7849 (N_7849,N_5924,N_4649);
nor U7850 (N_7850,N_4119,N_5155);
nand U7851 (N_7851,N_5714,N_5408);
or U7852 (N_7852,N_4259,N_5997);
or U7853 (N_7853,N_5286,N_4325);
and U7854 (N_7854,N_4872,N_4620);
nor U7855 (N_7855,N_4497,N_4116);
or U7856 (N_7856,N_4039,N_5293);
or U7857 (N_7857,N_5994,N_4879);
and U7858 (N_7858,N_4810,N_5121);
nand U7859 (N_7859,N_5248,N_4747);
nand U7860 (N_7860,N_5486,N_5058);
and U7861 (N_7861,N_4605,N_4383);
or U7862 (N_7862,N_4669,N_5761);
and U7863 (N_7863,N_5111,N_5848);
nand U7864 (N_7864,N_4082,N_5190);
or U7865 (N_7865,N_4577,N_5916);
and U7866 (N_7866,N_5704,N_4555);
nand U7867 (N_7867,N_5224,N_5699);
or U7868 (N_7868,N_5592,N_4748);
and U7869 (N_7869,N_5432,N_4157);
and U7870 (N_7870,N_5276,N_5344);
or U7871 (N_7871,N_5766,N_4050);
or U7872 (N_7872,N_4825,N_4945);
nand U7873 (N_7873,N_4043,N_5628);
nand U7874 (N_7874,N_4600,N_4417);
and U7875 (N_7875,N_5770,N_5746);
or U7876 (N_7876,N_5521,N_5302);
or U7877 (N_7877,N_5888,N_5732);
nor U7878 (N_7878,N_5493,N_5597);
nor U7879 (N_7879,N_4636,N_5285);
nand U7880 (N_7880,N_5341,N_4015);
or U7881 (N_7881,N_5943,N_5792);
nor U7882 (N_7882,N_5441,N_4196);
or U7883 (N_7883,N_5108,N_5708);
nand U7884 (N_7884,N_4976,N_5052);
and U7885 (N_7885,N_5051,N_4794);
and U7886 (N_7886,N_4872,N_4670);
or U7887 (N_7887,N_5405,N_5579);
nor U7888 (N_7888,N_4740,N_5710);
and U7889 (N_7889,N_4681,N_5630);
nor U7890 (N_7890,N_4287,N_5257);
nor U7891 (N_7891,N_5739,N_5700);
nand U7892 (N_7892,N_4914,N_5229);
nand U7893 (N_7893,N_5947,N_4039);
nand U7894 (N_7894,N_5412,N_5351);
xor U7895 (N_7895,N_4535,N_5449);
or U7896 (N_7896,N_5220,N_4204);
or U7897 (N_7897,N_4221,N_5372);
or U7898 (N_7898,N_4094,N_5709);
nand U7899 (N_7899,N_5073,N_5193);
xor U7900 (N_7900,N_4487,N_4486);
and U7901 (N_7901,N_4004,N_4121);
and U7902 (N_7902,N_4380,N_4264);
and U7903 (N_7903,N_5855,N_5907);
nand U7904 (N_7904,N_5422,N_4764);
and U7905 (N_7905,N_4797,N_4113);
or U7906 (N_7906,N_4211,N_4359);
nand U7907 (N_7907,N_5509,N_5544);
xnor U7908 (N_7908,N_5385,N_4025);
nand U7909 (N_7909,N_4765,N_5470);
nor U7910 (N_7910,N_5007,N_5670);
or U7911 (N_7911,N_5852,N_5400);
and U7912 (N_7912,N_4731,N_5175);
and U7913 (N_7913,N_5785,N_5689);
or U7914 (N_7914,N_4943,N_4872);
and U7915 (N_7915,N_4810,N_4331);
nand U7916 (N_7916,N_5585,N_5653);
nor U7917 (N_7917,N_5363,N_5467);
xor U7918 (N_7918,N_4324,N_5592);
xnor U7919 (N_7919,N_5996,N_5715);
and U7920 (N_7920,N_5483,N_4812);
or U7921 (N_7921,N_4247,N_5749);
and U7922 (N_7922,N_4839,N_5380);
or U7923 (N_7923,N_5361,N_4443);
nor U7924 (N_7924,N_5027,N_5270);
nor U7925 (N_7925,N_4005,N_5422);
and U7926 (N_7926,N_5570,N_4198);
nor U7927 (N_7927,N_4394,N_4982);
and U7928 (N_7928,N_4877,N_4044);
and U7929 (N_7929,N_5613,N_4641);
nand U7930 (N_7930,N_5103,N_5718);
nor U7931 (N_7931,N_4066,N_4598);
nand U7932 (N_7932,N_4491,N_5462);
or U7933 (N_7933,N_4926,N_5909);
nor U7934 (N_7934,N_4598,N_5112);
and U7935 (N_7935,N_4025,N_4986);
or U7936 (N_7936,N_5794,N_5589);
and U7937 (N_7937,N_5444,N_4953);
nand U7938 (N_7938,N_4562,N_5900);
and U7939 (N_7939,N_4808,N_4802);
nand U7940 (N_7940,N_5111,N_4747);
and U7941 (N_7941,N_5544,N_5892);
nor U7942 (N_7942,N_4334,N_5332);
or U7943 (N_7943,N_5240,N_5151);
nor U7944 (N_7944,N_4708,N_4671);
or U7945 (N_7945,N_5939,N_5097);
nor U7946 (N_7946,N_4607,N_4895);
nor U7947 (N_7947,N_5134,N_5945);
nand U7948 (N_7948,N_5529,N_5304);
nand U7949 (N_7949,N_4201,N_5151);
nor U7950 (N_7950,N_4782,N_5538);
nor U7951 (N_7951,N_4042,N_5065);
nor U7952 (N_7952,N_5888,N_4650);
nand U7953 (N_7953,N_4325,N_5399);
or U7954 (N_7954,N_5561,N_5641);
nor U7955 (N_7955,N_4525,N_4497);
and U7956 (N_7956,N_5210,N_4768);
and U7957 (N_7957,N_4133,N_5876);
nand U7958 (N_7958,N_5341,N_5322);
and U7959 (N_7959,N_5846,N_4606);
nor U7960 (N_7960,N_4546,N_4698);
and U7961 (N_7961,N_5304,N_5523);
nand U7962 (N_7962,N_4783,N_5857);
nand U7963 (N_7963,N_5976,N_4815);
nor U7964 (N_7964,N_5668,N_5742);
or U7965 (N_7965,N_5603,N_5905);
and U7966 (N_7966,N_4421,N_4162);
and U7967 (N_7967,N_4555,N_5635);
nor U7968 (N_7968,N_4181,N_5363);
or U7969 (N_7969,N_4622,N_5900);
or U7970 (N_7970,N_5759,N_5227);
nand U7971 (N_7971,N_4717,N_4789);
nand U7972 (N_7972,N_4177,N_5772);
or U7973 (N_7973,N_4776,N_4007);
nor U7974 (N_7974,N_4659,N_4067);
and U7975 (N_7975,N_4115,N_5815);
nor U7976 (N_7976,N_4636,N_4721);
and U7977 (N_7977,N_4323,N_4759);
nor U7978 (N_7978,N_4151,N_4995);
nand U7979 (N_7979,N_4715,N_5962);
nor U7980 (N_7980,N_5718,N_4219);
or U7981 (N_7981,N_5722,N_4411);
nor U7982 (N_7982,N_4386,N_4549);
nand U7983 (N_7983,N_4838,N_5118);
nor U7984 (N_7984,N_5912,N_5474);
nor U7985 (N_7985,N_4385,N_4904);
nor U7986 (N_7986,N_5371,N_5042);
or U7987 (N_7987,N_4457,N_5824);
and U7988 (N_7988,N_4660,N_4958);
nor U7989 (N_7989,N_5345,N_5113);
nand U7990 (N_7990,N_5328,N_4506);
and U7991 (N_7991,N_5196,N_4949);
nor U7992 (N_7992,N_5083,N_5557);
or U7993 (N_7993,N_5801,N_4722);
nor U7994 (N_7994,N_5385,N_4386);
or U7995 (N_7995,N_4729,N_5838);
or U7996 (N_7996,N_5048,N_5451);
or U7997 (N_7997,N_4854,N_4512);
or U7998 (N_7998,N_5886,N_4493);
nand U7999 (N_7999,N_4033,N_4840);
nor U8000 (N_8000,N_6387,N_6459);
nor U8001 (N_8001,N_6015,N_7244);
and U8002 (N_8002,N_6100,N_7205);
and U8003 (N_8003,N_6507,N_7324);
and U8004 (N_8004,N_7301,N_6179);
or U8005 (N_8005,N_7201,N_7991);
and U8006 (N_8006,N_6174,N_6045);
or U8007 (N_8007,N_6866,N_6151);
or U8008 (N_8008,N_6340,N_6125);
nor U8009 (N_8009,N_7926,N_7628);
and U8010 (N_8010,N_6709,N_6912);
nand U8011 (N_8011,N_6162,N_6733);
nor U8012 (N_8012,N_7231,N_6799);
nor U8013 (N_8013,N_7100,N_6403);
and U8014 (N_8014,N_7128,N_7455);
and U8015 (N_8015,N_7573,N_7714);
nor U8016 (N_8016,N_6558,N_7618);
and U8017 (N_8017,N_7196,N_6604);
nor U8018 (N_8018,N_6822,N_7059);
and U8019 (N_8019,N_6482,N_7509);
nor U8020 (N_8020,N_6770,N_7843);
and U8021 (N_8021,N_7235,N_6897);
nor U8022 (N_8022,N_7846,N_6580);
nand U8023 (N_8023,N_7898,N_7526);
or U8024 (N_8024,N_7853,N_6810);
nand U8025 (N_8025,N_6239,N_7890);
and U8026 (N_8026,N_6644,N_6855);
or U8027 (N_8027,N_6910,N_7871);
and U8028 (N_8028,N_6964,N_6540);
or U8029 (N_8029,N_6296,N_6607);
or U8030 (N_8030,N_6003,N_6868);
nor U8031 (N_8031,N_7099,N_6590);
nor U8032 (N_8032,N_7503,N_7213);
nor U8033 (N_8033,N_6758,N_7824);
or U8034 (N_8034,N_7191,N_7688);
nor U8035 (N_8035,N_6889,N_7807);
or U8036 (N_8036,N_7287,N_6640);
or U8037 (N_8037,N_7036,N_6450);
nand U8038 (N_8038,N_6428,N_7698);
and U8039 (N_8039,N_7261,N_7922);
and U8040 (N_8040,N_7047,N_6588);
nor U8041 (N_8041,N_6158,N_7692);
and U8042 (N_8042,N_7916,N_7366);
or U8043 (N_8043,N_6738,N_7765);
or U8044 (N_8044,N_7470,N_7415);
nand U8045 (N_8045,N_7716,N_7315);
nand U8046 (N_8046,N_7617,N_7646);
nor U8047 (N_8047,N_7314,N_6355);
and U8048 (N_8048,N_6857,N_7747);
nor U8049 (N_8049,N_6114,N_7773);
nand U8050 (N_8050,N_6562,N_6009);
and U8051 (N_8051,N_7331,N_7375);
nor U8052 (N_8052,N_7740,N_6985);
nor U8053 (N_8053,N_7606,N_7277);
nand U8054 (N_8054,N_6299,N_6731);
nand U8055 (N_8055,N_7552,N_6210);
and U8056 (N_8056,N_6375,N_6197);
nand U8057 (N_8057,N_6776,N_7670);
nor U8058 (N_8058,N_6863,N_6165);
nand U8059 (N_8059,N_6156,N_6067);
and U8060 (N_8060,N_7891,N_7385);
nand U8061 (N_8061,N_6809,N_7312);
and U8062 (N_8062,N_6423,N_7997);
nor U8063 (N_8063,N_6603,N_7654);
and U8064 (N_8064,N_7419,N_6662);
and U8065 (N_8065,N_6225,N_6219);
nand U8066 (N_8066,N_6885,N_6668);
and U8067 (N_8067,N_7177,N_6675);
nor U8068 (N_8068,N_6460,N_6339);
or U8069 (N_8069,N_6846,N_7995);
and U8070 (N_8070,N_7474,N_6907);
nand U8071 (N_8071,N_7251,N_6443);
and U8072 (N_8072,N_7323,N_6650);
nor U8073 (N_8073,N_7561,N_7071);
and U8074 (N_8074,N_6998,N_7781);
and U8075 (N_8075,N_7004,N_7220);
nand U8076 (N_8076,N_6622,N_6494);
or U8077 (N_8077,N_7808,N_7631);
or U8078 (N_8078,N_7106,N_6745);
nand U8079 (N_8079,N_6040,N_7844);
nor U8080 (N_8080,N_7369,N_7318);
and U8081 (N_8081,N_6752,N_6262);
and U8082 (N_8082,N_6913,N_6116);
nor U8083 (N_8083,N_6038,N_7248);
nor U8084 (N_8084,N_7992,N_7786);
nor U8085 (N_8085,N_6353,N_6363);
nor U8086 (N_8086,N_6395,N_6371);
nor U8087 (N_8087,N_7156,N_6892);
nand U8088 (N_8088,N_6688,N_6726);
or U8089 (N_8089,N_7704,N_6856);
nor U8090 (N_8090,N_7407,N_7738);
nand U8091 (N_8091,N_6596,N_6908);
nor U8092 (N_8092,N_6970,N_7398);
or U8093 (N_8093,N_6663,N_6259);
nand U8094 (N_8094,N_6397,N_7712);
or U8095 (N_8095,N_7865,N_6333);
or U8096 (N_8096,N_6775,N_6656);
and U8097 (N_8097,N_6585,N_7157);
nand U8098 (N_8098,N_6851,N_7791);
or U8099 (N_8099,N_6323,N_6773);
and U8100 (N_8100,N_7972,N_6876);
nand U8101 (N_8101,N_7687,N_6666);
and U8102 (N_8102,N_7061,N_7505);
nor U8103 (N_8103,N_7246,N_6651);
and U8104 (N_8104,N_7999,N_6115);
nor U8105 (N_8105,N_7651,N_6360);
nor U8106 (N_8106,N_7496,N_6101);
nor U8107 (N_8107,N_7906,N_6105);
nand U8108 (N_8108,N_7311,N_7001);
xnor U8109 (N_8109,N_7927,N_6514);
nand U8110 (N_8110,N_7471,N_6138);
nor U8111 (N_8111,N_7335,N_7804);
or U8112 (N_8112,N_7284,N_7150);
or U8113 (N_8113,N_6700,N_7896);
nor U8114 (N_8114,N_7152,N_7852);
and U8115 (N_8115,N_6248,N_7727);
or U8116 (N_8116,N_6418,N_6078);
nor U8117 (N_8117,N_7459,N_6634);
nand U8118 (N_8118,N_6571,N_7836);
and U8119 (N_8119,N_7500,N_7695);
nor U8120 (N_8120,N_6432,N_6281);
or U8121 (N_8121,N_7523,N_6229);
nand U8122 (N_8122,N_6919,N_7214);
nor U8123 (N_8123,N_7831,N_7599);
or U8124 (N_8124,N_6419,N_7476);
and U8125 (N_8125,N_7632,N_6936);
nor U8126 (N_8126,N_6699,N_7153);
nand U8127 (N_8127,N_7298,N_6811);
or U8128 (N_8128,N_6121,N_7166);
and U8129 (N_8129,N_6721,N_6109);
nand U8130 (N_8130,N_6316,N_7519);
nor U8131 (N_8131,N_6245,N_7203);
nand U8132 (N_8132,N_6161,N_6090);
nand U8133 (N_8133,N_6918,N_6513);
nand U8134 (N_8134,N_7862,N_7942);
nor U8135 (N_8135,N_7325,N_6737);
xnor U8136 (N_8136,N_7326,N_7608);
nor U8137 (N_8137,N_7619,N_7445);
or U8138 (N_8138,N_7031,N_7147);
nor U8139 (N_8139,N_6952,N_7368);
nand U8140 (N_8140,N_6043,N_7431);
or U8141 (N_8141,N_7188,N_7572);
or U8142 (N_8142,N_7780,N_6785);
nor U8143 (N_8143,N_7557,N_6004);
and U8144 (N_8144,N_7696,N_7902);
and U8145 (N_8145,N_7208,N_6808);
nor U8146 (N_8146,N_6670,N_6960);
nor U8147 (N_8147,N_7330,N_6530);
and U8148 (N_8148,N_6012,N_6236);
nor U8149 (N_8149,N_6969,N_7593);
nor U8150 (N_8150,N_6388,N_6155);
and U8151 (N_8151,N_6768,N_7034);
xor U8152 (N_8152,N_7946,N_6764);
nand U8153 (N_8153,N_7160,N_7771);
nand U8154 (N_8154,N_7603,N_6169);
or U8155 (N_8155,N_6519,N_7443);
nand U8156 (N_8156,N_6232,N_6391);
and U8157 (N_8157,N_6914,N_7777);
xor U8158 (N_8158,N_7452,N_7488);
nand U8159 (N_8159,N_6329,N_6303);
and U8160 (N_8160,N_7276,N_6937);
and U8161 (N_8161,N_7532,N_7810);
nor U8162 (N_8162,N_7017,N_7650);
nand U8163 (N_8163,N_7332,N_7805);
nand U8164 (N_8164,N_6006,N_7477);
nand U8165 (N_8165,N_7511,N_7333);
or U8166 (N_8166,N_7855,N_7327);
nor U8167 (N_8167,N_6087,N_6801);
or U8168 (N_8168,N_6124,N_7190);
and U8169 (N_8169,N_7905,N_6746);
nor U8170 (N_8170,N_7897,N_7577);
or U8171 (N_8171,N_6869,N_6933);
nor U8172 (N_8172,N_7581,N_7685);
or U8173 (N_8173,N_6658,N_7764);
or U8174 (N_8174,N_7535,N_7155);
or U8175 (N_8175,N_6207,N_7874);
xnor U8176 (N_8176,N_6199,N_6744);
nor U8177 (N_8177,N_7390,N_6832);
nor U8178 (N_8178,N_6615,N_7612);
or U8179 (N_8179,N_7982,N_6535);
or U8180 (N_8180,N_6212,N_7506);
nand U8181 (N_8181,N_6905,N_7198);
and U8182 (N_8182,N_6356,N_7342);
nand U8183 (N_8183,N_6163,N_7337);
nor U8184 (N_8184,N_6137,N_7064);
nor U8185 (N_8185,N_7711,N_7648);
or U8186 (N_8186,N_7232,N_6023);
nand U8187 (N_8187,N_6583,N_6057);
or U8188 (N_8188,N_7879,N_6267);
and U8189 (N_8189,N_7847,N_6258);
or U8190 (N_8190,N_6018,N_7627);
nand U8191 (N_8191,N_7515,N_7253);
or U8192 (N_8192,N_7349,N_6170);
or U8193 (N_8193,N_7045,N_6926);
nor U8194 (N_8194,N_6471,N_7021);
or U8195 (N_8195,N_7374,N_6820);
nand U8196 (N_8196,N_7564,N_7126);
nor U8197 (N_8197,N_6036,N_7384);
nor U8198 (N_8198,N_7204,N_6176);
or U8199 (N_8199,N_6415,N_6787);
and U8200 (N_8200,N_6383,N_6728);
nor U8201 (N_8201,N_7175,N_7923);
nor U8202 (N_8202,N_6623,N_7768);
and U8203 (N_8203,N_7555,N_7566);
and U8204 (N_8204,N_7334,N_6445);
nand U8205 (N_8205,N_6024,N_7217);
and U8206 (N_8206,N_7142,N_7255);
nand U8207 (N_8207,N_6243,N_7812);
nand U8208 (N_8208,N_7114,N_6903);
nand U8209 (N_8209,N_7222,N_6453);
nor U8210 (N_8210,N_6382,N_7453);
and U8211 (N_8211,N_7209,N_7393);
nand U8212 (N_8212,N_6050,N_6895);
or U8213 (N_8213,N_6093,N_6702);
and U8214 (N_8214,N_6493,N_7362);
nor U8215 (N_8215,N_7241,N_6111);
and U8216 (N_8216,N_6107,N_7661);
nor U8217 (N_8217,N_7259,N_6888);
nand U8218 (N_8218,N_7534,N_6426);
nor U8219 (N_8219,N_6135,N_6049);
nand U8220 (N_8220,N_6160,N_6478);
nor U8221 (N_8221,N_6435,N_6496);
nor U8222 (N_8222,N_6975,N_7483);
xor U8223 (N_8223,N_6468,N_7850);
or U8224 (N_8224,N_6748,N_6630);
nor U8225 (N_8225,N_7469,N_7060);
or U8226 (N_8226,N_6191,N_6991);
and U8227 (N_8227,N_6480,N_7310);
or U8228 (N_8228,N_7624,N_7767);
or U8229 (N_8229,N_6216,N_7551);
nor U8230 (N_8230,N_7909,N_7359);
and U8231 (N_8231,N_7880,N_7914);
and U8232 (N_8232,N_7075,N_7200);
and U8233 (N_8233,N_7528,N_7401);
nand U8234 (N_8234,N_6440,N_7814);
or U8235 (N_8235,N_7547,N_6805);
or U8236 (N_8236,N_7371,N_7788);
nor U8237 (N_8237,N_6774,N_7585);
and U8238 (N_8238,N_7095,N_6102);
nand U8239 (N_8239,N_7270,N_6446);
xnor U8240 (N_8240,N_6777,N_6891);
nand U8241 (N_8241,N_6365,N_7647);
nor U8242 (N_8242,N_6437,N_7077);
or U8243 (N_8243,N_6048,N_7245);
and U8244 (N_8244,N_7266,N_7122);
nand U8245 (N_8245,N_7389,N_7102);
or U8246 (N_8246,N_7838,N_6421);
or U8247 (N_8247,N_7728,N_7822);
nor U8248 (N_8248,N_7729,N_7404);
nand U8249 (N_8249,N_6920,N_6999);
nor U8250 (N_8250,N_6182,N_7257);
or U8251 (N_8251,N_6927,N_7662);
nor U8252 (N_8252,N_6899,N_6767);
nand U8253 (N_8253,N_7187,N_6639);
nand U8254 (N_8254,N_6020,N_6416);
nand U8255 (N_8255,N_6501,N_7939);
nor U8256 (N_8256,N_7722,N_7974);
or U8257 (N_8257,N_7278,N_7546);
or U8258 (N_8258,N_6698,N_7953);
or U8259 (N_8259,N_7306,N_7464);
nand U8260 (N_8260,N_6136,N_7886);
and U8261 (N_8261,N_6942,N_7533);
xnor U8262 (N_8262,N_7833,N_6217);
and U8263 (N_8263,N_7985,N_6322);
nor U8264 (N_8264,N_6171,N_7604);
or U8265 (N_8265,N_6921,N_6987);
nand U8266 (N_8266,N_7888,N_7652);
nand U8267 (N_8267,N_6842,N_7826);
and U8268 (N_8268,N_7872,N_7499);
and U8269 (N_8269,N_6747,N_7525);
nor U8270 (N_8270,N_7146,N_6119);
or U8271 (N_8271,N_7116,N_6466);
and U8272 (N_8272,N_6481,N_7405);
nand U8273 (N_8273,N_7737,N_6625);
and U8274 (N_8274,N_6643,N_7172);
nand U8275 (N_8275,N_7319,N_7396);
and U8276 (N_8276,N_7364,N_6112);
or U8277 (N_8277,N_6330,N_6257);
nor U8278 (N_8278,N_6237,N_6000);
and U8279 (N_8279,N_6696,N_6598);
or U8280 (N_8280,N_6828,N_6962);
xnor U8281 (N_8281,N_7613,N_6277);
nand U8282 (N_8282,N_6543,N_6310);
nor U8283 (N_8283,N_7983,N_7524);
and U8284 (N_8284,N_7089,N_7731);
or U8285 (N_8285,N_6807,N_7913);
nor U8286 (N_8286,N_6380,N_7908);
nor U8287 (N_8287,N_6410,N_7543);
nor U8288 (N_8288,N_6994,N_7352);
or U8289 (N_8289,N_6081,N_6691);
nor U8290 (N_8290,N_6974,N_6701);
nor U8291 (N_8291,N_7361,N_7799);
nand U8292 (N_8292,N_7262,N_6997);
nand U8293 (N_8293,N_7039,N_6384);
or U8294 (N_8294,N_6821,N_6189);
nand U8295 (N_8295,N_7752,N_6061);
nor U8296 (N_8296,N_6106,N_6282);
nand U8297 (N_8297,N_6404,N_7171);
nor U8298 (N_8298,N_7430,N_6177);
nand U8299 (N_8299,N_7305,N_7479);
and U8300 (N_8300,N_6373,N_6358);
or U8301 (N_8301,N_6693,N_7821);
or U8302 (N_8302,N_6250,N_7081);
nand U8303 (N_8303,N_7783,N_7286);
nand U8304 (N_8304,N_6569,N_6291);
or U8305 (N_8305,N_7328,N_6594);
nand U8306 (N_8306,N_6327,N_6678);
or U8307 (N_8307,N_6979,N_7290);
or U8308 (N_8308,N_6390,N_6185);
or U8309 (N_8309,N_7529,N_7709);
nand U8310 (N_8310,N_7736,N_7707);
nand U8311 (N_8311,N_6328,N_6204);
or U8312 (N_8312,N_7565,N_6032);
xnor U8313 (N_8313,N_6576,N_7616);
nor U8314 (N_8314,N_7829,N_7406);
or U8315 (N_8315,N_7597,N_7094);
nor U8316 (N_8316,N_6680,N_7123);
or U8317 (N_8317,N_6720,N_6088);
nor U8318 (N_8318,N_6213,N_7986);
and U8319 (N_8319,N_6676,N_7050);
nor U8320 (N_8320,N_6686,N_7795);
nand U8321 (N_8321,N_6948,N_6035);
nand U8322 (N_8322,N_7441,N_7436);
and U8323 (N_8323,N_6130,N_7302);
and U8324 (N_8324,N_6859,N_7980);
nor U8325 (N_8325,N_6195,N_7966);
and U8326 (N_8326,N_6218,N_6029);
nor U8327 (N_8327,N_6167,N_6347);
and U8328 (N_8328,N_7733,N_7485);
and U8329 (N_8329,N_7184,N_7678);
or U8330 (N_8330,N_7580,N_7074);
nand U8331 (N_8331,N_7239,N_6346);
or U8332 (N_8332,N_6186,N_7068);
and U8333 (N_8333,N_6642,N_6261);
nand U8334 (N_8334,N_6126,N_7033);
and U8335 (N_8335,N_6089,N_6749);
or U8336 (N_8336,N_7932,N_7046);
nor U8337 (N_8337,N_6683,N_7801);
nor U8338 (N_8338,N_6472,N_6528);
nor U8339 (N_8339,N_7756,N_6713);
nor U8340 (N_8340,N_7975,N_6986);
nor U8341 (N_8341,N_7092,N_7868);
or U8342 (N_8342,N_7296,N_7358);
or U8343 (N_8343,N_6886,N_6022);
and U8344 (N_8344,N_7981,N_6315);
or U8345 (N_8345,N_7484,N_6694);
or U8346 (N_8346,N_7426,N_6249);
nand U8347 (N_8347,N_6474,N_6794);
or U8348 (N_8348,N_6076,N_6063);
and U8349 (N_8349,N_7757,N_6251);
nand U8350 (N_8350,N_6645,N_6394);
and U8351 (N_8351,N_6127,N_7224);
nand U8352 (N_8352,N_7947,N_6619);
nand U8353 (N_8353,N_7462,N_7588);
and U8354 (N_8354,N_6646,N_6305);
nor U8355 (N_8355,N_7811,N_6414);
or U8356 (N_8356,N_6504,N_6843);
nand U8357 (N_8357,N_6484,N_7892);
and U8358 (N_8358,N_6348,N_6362);
and U8359 (N_8359,N_7223,N_7141);
nand U8360 (N_8360,N_7762,N_6795);
and U8361 (N_8361,N_7904,N_7165);
or U8362 (N_8362,N_6238,N_6564);
nor U8363 (N_8363,N_7351,N_7027);
or U8364 (N_8364,N_6629,N_7069);
nor U8365 (N_8365,N_7867,N_6944);
or U8366 (N_8366,N_6546,N_6168);
nor U8367 (N_8367,N_7634,N_6424);
nand U8368 (N_8368,N_6848,N_7813);
nand U8369 (N_8369,N_6376,N_7877);
or U8370 (N_8370,N_7410,N_7776);
nand U8371 (N_8371,N_6108,N_7024);
nand U8372 (N_8372,N_7548,N_7589);
nand U8373 (N_8373,N_7281,N_6684);
or U8374 (N_8374,N_7096,N_7316);
xnor U8375 (N_8375,N_7660,N_7878);
xnor U8376 (N_8376,N_7668,N_6943);
nor U8377 (N_8377,N_7549,N_6381);
and U8378 (N_8378,N_6104,N_7989);
and U8379 (N_8379,N_6231,N_7193);
nor U8380 (N_8380,N_7113,N_7249);
nand U8381 (N_8381,N_7693,N_6046);
xor U8382 (N_8382,N_6878,N_6741);
or U8383 (N_8383,N_6429,N_7067);
nor U8384 (N_8384,N_7520,N_7120);
and U8385 (N_8385,N_6730,N_6797);
nand U8386 (N_8386,N_6627,N_6862);
or U8387 (N_8387,N_7512,N_6761);
or U8388 (N_8388,N_7595,N_7713);
nand U8389 (N_8389,N_6617,N_6722);
and U8390 (N_8390,N_6705,N_6368);
nor U8391 (N_8391,N_6624,N_6313);
or U8392 (N_8392,N_7769,N_7420);
nand U8393 (N_8393,N_7683,N_6957);
or U8394 (N_8394,N_6792,N_7424);
and U8395 (N_8395,N_7115,N_6091);
nor U8396 (N_8396,N_6042,N_7542);
nor U8397 (N_8397,N_7667,N_7273);
nand U8398 (N_8398,N_6537,N_6477);
or U8399 (N_8399,N_7107,N_7093);
or U8400 (N_8400,N_6253,N_6657);
or U8401 (N_8401,N_6021,N_7216);
nand U8402 (N_8402,N_7635,N_6893);
or U8403 (N_8403,N_6240,N_6601);
nand U8404 (N_8404,N_6479,N_6274);
nand U8405 (N_8405,N_6953,N_6354);
nor U8406 (N_8406,N_6463,N_7994);
and U8407 (N_8407,N_6951,N_6495);
nor U8408 (N_8408,N_6110,N_6019);
nor U8409 (N_8409,N_6704,N_6485);
nor U8410 (N_8410,N_6659,N_7447);
nor U8411 (N_8411,N_6781,N_6379);
nand U8412 (N_8412,N_6915,N_7288);
and U8413 (N_8413,N_7457,N_7583);
nand U8414 (N_8414,N_6727,N_7108);
or U8415 (N_8415,N_7517,N_7976);
and U8416 (N_8416,N_7041,N_6900);
or U8417 (N_8417,N_6870,N_6144);
or U8418 (N_8418,N_7044,N_7303);
or U8419 (N_8419,N_7003,N_6469);
or U8420 (N_8420,N_6802,N_6592);
nor U8421 (N_8421,N_6149,N_6187);
nor U8422 (N_8422,N_6616,N_6669);
nand U8423 (N_8423,N_6196,N_6928);
nand U8424 (N_8424,N_7959,N_6014);
and U8425 (N_8425,N_6060,N_6307);
nor U8426 (N_8426,N_6286,N_7438);
nand U8427 (N_8427,N_6304,N_7292);
nand U8428 (N_8428,N_7051,N_7117);
nor U8429 (N_8429,N_7367,N_7630);
or U8430 (N_8430,N_7507,N_7990);
xor U8431 (N_8431,N_7414,N_7154);
nor U8432 (N_8432,N_7354,N_7856);
nand U8433 (N_8433,N_6007,N_7356);
and U8434 (N_8434,N_6448,N_7759);
or U8435 (N_8435,N_7965,N_7828);
or U8436 (N_8436,N_6252,N_7416);
or U8437 (N_8437,N_6534,N_7121);
and U8438 (N_8438,N_7864,N_6692);
nor U8439 (N_8439,N_7225,N_7633);
and U8440 (N_8440,N_6605,N_6561);
or U8441 (N_8441,N_6652,N_6420);
or U8442 (N_8442,N_6436,N_6406);
nand U8443 (N_8443,N_6509,N_6923);
and U8444 (N_8444,N_6385,N_6541);
and U8445 (N_8445,N_6298,N_6852);
and U8446 (N_8446,N_6393,N_7465);
nor U8447 (N_8447,N_7189,N_7238);
nand U8448 (N_8448,N_7080,N_7882);
nor U8449 (N_8449,N_7504,N_7148);
nand U8450 (N_8450,N_6877,N_6826);
nor U8451 (N_8451,N_7900,N_6386);
nand U8452 (N_8452,N_7967,N_6739);
nor U8453 (N_8453,N_7937,N_6524);
nand U8454 (N_8454,N_6192,N_7014);
and U8455 (N_8455,N_7596,N_7194);
nor U8456 (N_8456,N_6208,N_7012);
nor U8457 (N_8457,N_6896,N_7659);
and U8458 (N_8458,N_6636,N_6835);
or U8459 (N_8459,N_7007,N_7212);
xnor U8460 (N_8460,N_6140,N_7387);
xnor U8461 (N_8461,N_7579,N_7112);
or U8462 (N_8462,N_7026,N_6289);
nand U8463 (N_8463,N_6378,N_6766);
or U8464 (N_8464,N_6278,N_7848);
and U8465 (N_8465,N_6844,N_6413);
or U8466 (N_8466,N_7468,N_6188);
or U8467 (N_8467,N_7894,N_6934);
nor U8468 (N_8468,N_7948,N_7817);
nor U8469 (N_8469,N_7682,N_6756);
and U8470 (N_8470,N_6041,N_7700);
nor U8471 (N_8471,N_6201,N_6577);
and U8472 (N_8472,N_7065,N_6335);
and U8473 (N_8473,N_7735,N_6925);
nor U8474 (N_8474,N_7574,N_6655);
or U8475 (N_8475,N_7860,N_7778);
nor U8476 (N_8476,N_6300,N_7675);
nor U8477 (N_8477,N_6719,N_7009);
nand U8478 (N_8478,N_6013,N_6244);
nor U8479 (N_8479,N_6297,N_7043);
or U8480 (N_8480,N_6465,N_6945);
nand U8481 (N_8481,N_7625,N_6568);
nor U8482 (N_8482,N_6031,N_6319);
or U8483 (N_8483,N_6827,N_6366);
nor U8484 (N_8484,N_6591,N_7011);
or U8485 (N_8485,N_6336,N_7028);
nor U8486 (N_8486,N_7875,N_6980);
or U8487 (N_8487,N_7708,N_7677);
nor U8488 (N_8488,N_7293,N_7744);
or U8489 (N_8489,N_6983,N_7793);
or U8490 (N_8490,N_7040,N_6825);
and U8491 (N_8491,N_6492,N_7516);
nor U8492 (N_8492,N_6784,N_7761);
nand U8493 (N_8493,N_6173,N_7917);
nor U8494 (N_8494,N_6553,N_6671);
and U8495 (N_8495,N_6612,N_7563);
nand U8496 (N_8496,N_7823,N_6226);
or U8497 (N_8497,N_7919,N_6181);
or U8498 (N_8498,N_7492,N_6778);
and U8499 (N_8499,N_7285,N_7726);
nor U8500 (N_8500,N_6295,N_6120);
or U8501 (N_8501,N_6294,N_7019);
nand U8502 (N_8502,N_6971,N_6814);
nand U8503 (N_8503,N_6573,N_6990);
nand U8504 (N_8504,N_7941,N_6412);
and U8505 (N_8505,N_6593,N_7181);
or U8506 (N_8506,N_6337,N_7815);
nand U8507 (N_8507,N_6648,N_6451);
nor U8508 (N_8508,N_7857,N_6940);
nand U8509 (N_8509,N_7639,N_7427);
nand U8510 (N_8510,N_6981,N_7598);
or U8511 (N_8511,N_6054,N_7931);
nand U8512 (N_8512,N_7883,N_7086);
and U8513 (N_8513,N_7806,N_7163);
or U8514 (N_8514,N_7956,N_6707);
or U8515 (N_8515,N_7104,N_7139);
nand U8516 (N_8516,N_6517,N_6672);
nor U8517 (N_8517,N_7308,N_6887);
or U8518 (N_8518,N_7421,N_6628);
nand U8519 (N_8519,N_7615,N_6052);
and U8520 (N_8520,N_7395,N_6708);
nand U8521 (N_8521,N_7949,N_6467);
or U8522 (N_8522,N_6224,N_6989);
nand U8523 (N_8523,N_6861,N_6309);
or U8524 (N_8524,N_7267,N_6341);
xor U8525 (N_8525,N_6079,N_6142);
and U8526 (N_8526,N_7481,N_7841);
and U8527 (N_8527,N_7412,N_7934);
nand U8528 (N_8528,N_7397,N_6118);
nor U8529 (N_8529,N_7984,N_7048);
nor U8530 (N_8530,N_7621,N_7785);
or U8531 (N_8531,N_7513,N_6010);
or U8532 (N_8532,N_6051,N_7386);
and U8533 (N_8533,N_6153,N_6500);
or U8534 (N_8534,N_7680,N_7056);
or U8535 (N_8535,N_6521,N_7432);
or U8536 (N_8536,N_6071,N_7940);
nor U8537 (N_8537,N_6717,N_7763);
nand U8538 (N_8538,N_7030,N_7789);
or U8539 (N_8539,N_6830,N_6026);
or U8540 (N_8540,N_7706,N_6560);
nor U8541 (N_8541,N_6364,N_7610);
nand U8542 (N_8542,N_6392,N_7347);
nor U8543 (N_8543,N_6681,N_7015);
and U8544 (N_8544,N_7629,N_6408);
and U8545 (N_8545,N_6270,N_6551);
or U8546 (N_8546,N_7674,N_6600);
nand U8547 (N_8547,N_6922,N_7211);
nand U8548 (N_8548,N_7062,N_6139);
or U8549 (N_8549,N_7458,N_7025);
and U8550 (N_8550,N_7037,N_6028);
or U8551 (N_8551,N_6898,N_6200);
or U8552 (N_8552,N_7049,N_6417);
nand U8553 (N_8553,N_7388,N_6190);
and U8554 (N_8554,N_6241,N_6864);
or U8555 (N_8555,N_7690,N_6407);
nand U8556 (N_8556,N_6935,N_6084);
nor U8557 (N_8557,N_7605,N_7537);
and U8558 (N_8558,N_7380,N_6867);
and U8559 (N_8559,N_6609,N_6575);
nand U8560 (N_8560,N_7070,N_7642);
xnor U8561 (N_8561,N_7002,N_6334);
and U8562 (N_8562,N_7839,N_7291);
nand U8563 (N_8563,N_7226,N_7353);
and U8564 (N_8564,N_6377,N_7666);
and U8565 (N_8565,N_6972,N_6449);
nor U8566 (N_8566,N_7620,N_7467);
nor U8567 (N_8567,N_7697,N_7979);
and U8568 (N_8568,N_6847,N_7178);
nand U8569 (N_8569,N_7460,N_6595);
or U8570 (N_8570,N_7772,N_6875);
or U8571 (N_8571,N_7313,N_7144);
xnor U8572 (N_8572,N_6796,N_7103);
and U8573 (N_8573,N_6523,N_6512);
nor U8574 (N_8574,N_6725,N_7394);
nand U8575 (N_8575,N_6002,N_7592);
nand U8576 (N_8576,N_7863,N_6882);
nand U8577 (N_8577,N_6790,N_7428);
nand U8578 (N_8578,N_7701,N_6924);
or U8579 (N_8579,N_7988,N_6344);
or U8580 (N_8580,N_7299,N_7343);
nand U8581 (N_8581,N_6077,N_6613);
nand U8582 (N_8582,N_7372,N_7186);
or U8583 (N_8583,N_6320,N_6475);
and U8584 (N_8584,N_6771,N_7218);
nand U8585 (N_8585,N_7422,N_6273);
or U8586 (N_8586,N_6098,N_7575);
nand U8587 (N_8587,N_6703,N_7766);
and U8588 (N_8588,N_6357,N_7307);
and U8589 (N_8589,N_7724,N_6456);
or U8590 (N_8590,N_6312,N_7254);
or U8591 (N_8591,N_6890,N_6194);
and U8592 (N_8592,N_6917,N_7229);
nand U8593 (N_8593,N_6505,N_7755);
xor U8594 (N_8594,N_6996,N_7669);
nor U8595 (N_8595,N_6198,N_7247);
nand U8596 (N_8596,N_6401,N_7915);
and U8597 (N_8597,N_6222,N_7567);
nand U8598 (N_8598,N_6881,N_6715);
and U8599 (N_8599,N_7725,N_6058);
nor U8600 (N_8600,N_7022,N_7796);
nor U8601 (N_8601,N_7559,N_6017);
or U8602 (N_8602,N_6075,N_6586);
and U8603 (N_8603,N_7206,N_6027);
or U8604 (N_8604,N_6538,N_7952);
nand U8605 (N_8605,N_7962,N_7322);
or U8606 (N_8606,N_6016,N_7748);
nor U8607 (N_8607,N_7739,N_7448);
or U8608 (N_8608,N_7066,N_6959);
and U8609 (N_8609,N_7199,N_7444);
nor U8610 (N_8610,N_7672,N_7578);
nor U8611 (N_8611,N_6039,N_7545);
or U8612 (N_8612,N_7429,N_7720);
nand U8613 (N_8613,N_7373,N_7568);
and U8614 (N_8614,N_6180,N_6047);
and U8615 (N_8615,N_7461,N_6288);
nor U8616 (N_8616,N_6255,N_6982);
and U8617 (N_8617,N_7151,N_7032);
or U8618 (N_8618,N_6488,N_7694);
nand U8619 (N_8619,N_6499,N_7357);
nor U8620 (N_8620,N_7784,N_6117);
or U8621 (N_8621,N_7055,N_7754);
xor U8622 (N_8622,N_7363,N_6183);
and U8623 (N_8623,N_7973,N_6508);
or U8624 (N_8624,N_6400,N_7275);
or U8625 (N_8625,N_7381,N_7161);
nand U8626 (N_8626,N_7522,N_6860);
nand U8627 (N_8627,N_6425,N_7859);
and U8628 (N_8628,N_7501,N_7434);
nor U8629 (N_8629,N_7718,N_6487);
nor U8630 (N_8630,N_7887,N_6444);
and U8631 (N_8631,N_6823,N_6732);
or U8632 (N_8632,N_7182,N_7173);
or U8633 (N_8633,N_7237,N_6589);
nor U8634 (N_8634,N_6718,N_6818);
nand U8635 (N_8635,N_6559,N_7215);
and U8636 (N_8636,N_6929,N_7136);
and U8637 (N_8637,N_7623,N_6324);
nor U8638 (N_8638,N_7138,N_7899);
nor U8639 (N_8639,N_7091,N_7491);
nor U8640 (N_8640,N_7072,N_7876);
and U8641 (N_8641,N_7076,N_6497);
nand U8642 (N_8642,N_6542,N_6399);
or U8643 (N_8643,N_7480,N_6438);
and U8644 (N_8644,N_6470,N_6911);
nand U8645 (N_8645,N_6306,N_6332);
nor U8646 (N_8646,N_7145,N_6164);
or U8647 (N_8647,N_6260,N_7782);
nor U8648 (N_8648,N_6995,N_6581);
nor U8649 (N_8649,N_7297,N_6783);
nand U8650 (N_8650,N_6742,N_6325);
nand U8651 (N_8651,N_7958,N_7192);
and U8652 (N_8652,N_7282,N_7673);
or U8653 (N_8653,N_7038,N_7174);
or U8654 (N_8654,N_6234,N_7518);
and U8655 (N_8655,N_7935,N_6146);
nand U8656 (N_8656,N_6833,N_7383);
xnor U8657 (N_8657,N_7008,N_6280);
and U8658 (N_8658,N_6723,N_6263);
nand U8659 (N_8659,N_7912,N_7300);
and U8660 (N_8660,N_7236,N_6131);
nor U8661 (N_8661,N_7870,N_7435);
nor U8662 (N_8662,N_6374,N_6800);
nor U8663 (N_8663,N_7149,N_7329);
nor U8664 (N_8664,N_6473,N_6086);
and U8665 (N_8665,N_6434,N_7977);
and U8666 (N_8666,N_7382,N_6476);
nor U8667 (N_8667,N_7195,N_7197);
or U8668 (N_8668,N_7576,N_7391);
nor U8669 (N_8669,N_6452,N_6734);
or U8670 (N_8670,N_7889,N_7553);
nor U8671 (N_8671,N_6272,N_7819);
nand U8672 (N_8672,N_6103,N_6954);
or U8673 (N_8673,N_6254,N_7230);
or U8674 (N_8674,N_7794,N_7221);
and U8675 (N_8675,N_7269,N_6527);
or U8676 (N_8676,N_6791,N_6070);
and U8677 (N_8677,N_7514,N_7399);
or U8678 (N_8678,N_7978,N_7449);
nand U8679 (N_8679,N_6008,N_6901);
or U8680 (N_8680,N_6963,N_7964);
and U8681 (N_8681,N_6753,N_6956);
and U8682 (N_8682,N_7179,N_7042);
nand U8683 (N_8683,N_7943,N_7234);
nor U8684 (N_8684,N_7350,N_7760);
nor U8685 (N_8685,N_6283,N_7294);
and U8686 (N_8686,N_7751,N_6884);
or U8687 (N_8687,N_7536,N_7925);
or U8688 (N_8688,N_6660,N_6638);
xor U8689 (N_8689,N_7510,N_7242);
nand U8690 (N_8690,N_6788,N_6606);
nand U8691 (N_8691,N_6955,N_6967);
or U8692 (N_8692,N_6361,N_6269);
nor U8693 (N_8693,N_7998,N_7732);
or U8694 (N_8694,N_6949,N_7280);
and U8695 (N_8695,N_6025,N_6290);
nand U8696 (N_8696,N_7265,N_6958);
or U8697 (N_8697,N_7111,N_6930);
xor U8698 (N_8698,N_7866,N_7918);
xnor U8699 (N_8699,N_6193,N_7582);
and U8700 (N_8700,N_6839,N_6351);
nor U8701 (N_8701,N_6398,N_7130);
nand U8702 (N_8702,N_6547,N_6779);
and U8703 (N_8703,N_7392,N_7167);
nand U8704 (N_8704,N_6129,N_6872);
and U8705 (N_8705,N_6275,N_6946);
nand U8706 (N_8706,N_7960,N_7903);
or U8707 (N_8707,N_6205,N_7938);
or U8708 (N_8708,N_7827,N_6690);
or U8709 (N_8709,N_6916,N_7893);
nand U8710 (N_8710,N_7869,N_7425);
nor U8711 (N_8711,N_7473,N_7450);
and U8712 (N_8712,N_7168,N_7442);
or U8713 (N_8713,N_6080,N_7183);
or U8714 (N_8714,N_6667,N_6813);
nor U8715 (N_8715,N_6633,N_6533);
nor U8716 (N_8716,N_7750,N_6735);
nand U8717 (N_8717,N_7745,N_7554);
and U8718 (N_8718,N_7360,N_6854);
nor U8719 (N_8719,N_7018,N_6128);
nor U8720 (N_8720,N_6242,N_7684);
and U8721 (N_8721,N_7971,N_7016);
nand U8722 (N_8722,N_6372,N_7417);
or U8723 (N_8723,N_6871,N_6211);
nor U8724 (N_8724,N_6318,N_6712);
or U8725 (N_8725,N_7185,N_6510);
nor U8726 (N_8726,N_7207,N_6442);
xnor U8727 (N_8727,N_7109,N_6653);
nor U8728 (N_8728,N_6141,N_6276);
or U8729 (N_8729,N_6743,N_6812);
or U8730 (N_8730,N_7774,N_6834);
nor U8731 (N_8731,N_7798,N_7858);
nor U8732 (N_8732,N_6369,N_7643);
and U8733 (N_8733,N_6582,N_6976);
and U8734 (N_8734,N_7134,N_6166);
nand U8735 (N_8735,N_6359,N_6763);
nand U8736 (N_8736,N_7344,N_7105);
nor U8737 (N_8737,N_6062,N_7283);
and U8738 (N_8738,N_7475,N_7345);
xnor U8739 (N_8739,N_7950,N_6570);
or U8740 (N_8740,N_7271,N_7851);
nor U8741 (N_8741,N_7258,N_6610);
nand U8742 (N_8742,N_7490,N_6789);
and U8743 (N_8743,N_7256,N_6687);
nand U8744 (N_8744,N_6545,N_7968);
and U8745 (N_8745,N_6486,N_7527);
and U8746 (N_8746,N_7901,N_7264);
and U8747 (N_8747,N_6447,N_7498);
nor U8748 (N_8748,N_6556,N_6961);
or U8749 (N_8749,N_7955,N_6706);
or U8750 (N_8750,N_7140,N_6483);
nand U8751 (N_8751,N_6256,N_7494);
nor U8752 (N_8752,N_7820,N_7054);
nand U8753 (N_8753,N_7854,N_7341);
or U8754 (N_8754,N_6695,N_6431);
nor U8755 (N_8755,N_6206,N_6614);
or U8756 (N_8756,N_7159,N_6544);
and U8757 (N_8757,N_7721,N_7723);
and U8758 (N_8758,N_6620,N_6059);
nand U8759 (N_8759,N_6711,N_7378);
nor U8760 (N_8760,N_6133,N_6247);
and U8761 (N_8761,N_6458,N_6579);
or U8762 (N_8762,N_6661,N_6906);
nor U8763 (N_8763,N_6554,N_7691);
and U8764 (N_8764,N_6082,N_6824);
and U8765 (N_8765,N_6525,N_7119);
and U8766 (N_8766,N_7180,N_7320);
and U8767 (N_8767,N_6502,N_6411);
or U8768 (N_8768,N_7656,N_6178);
and U8769 (N_8769,N_7930,N_7558);
and U8770 (N_8770,N_6685,N_6909);
and U8771 (N_8771,N_7309,N_6550);
or U8772 (N_8772,N_6873,N_7370);
nand U8773 (N_8773,N_6154,N_7570);
or U8774 (N_8774,N_6266,N_6430);
and U8775 (N_8775,N_7907,N_7073);
nand U8776 (N_8776,N_7835,N_6172);
and U8777 (N_8777,N_6113,N_7655);
and U8778 (N_8778,N_7645,N_7000);
nand U8779 (N_8779,N_7742,N_7679);
or U8780 (N_8780,N_7703,N_6836);
nor U8781 (N_8781,N_6441,N_7158);
and U8782 (N_8782,N_6635,N_7289);
nand U8783 (N_8783,N_7569,N_7243);
or U8784 (N_8784,N_7837,N_7987);
nand U8785 (N_8785,N_6287,N_6815);
or U8786 (N_8786,N_6068,N_6314);
xnor U8787 (N_8787,N_6066,N_7591);
nor U8788 (N_8788,N_6433,N_6665);
and U8789 (N_8789,N_6457,N_6175);
or U8790 (N_8790,N_6491,N_7818);
and U8791 (N_8791,N_7079,N_6850);
or U8792 (N_8792,N_7274,N_7715);
or U8793 (N_8793,N_6880,N_7614);
or U8794 (N_8794,N_7944,N_7689);
nor U8795 (N_8795,N_7641,N_6932);
nand U8796 (N_8796,N_7873,N_6677);
xor U8797 (N_8797,N_6755,N_6221);
or U8798 (N_8798,N_6396,N_6902);
and U8799 (N_8799,N_7210,N_7408);
and U8800 (N_8800,N_7466,N_6710);
nand U8801 (N_8801,N_6342,N_6555);
and U8802 (N_8802,N_7304,N_6637);
nand U8803 (N_8803,N_6782,N_7749);
nand U8804 (N_8804,N_6030,N_7590);
nor U8805 (N_8805,N_6515,N_7454);
and U8806 (N_8806,N_6083,N_6134);
or U8807 (N_8807,N_6841,N_7885);
xnor U8808 (N_8808,N_6308,N_7063);
and U8809 (N_8809,N_7169,N_6150);
nand U8810 (N_8810,N_7338,N_6697);
nor U8811 (N_8811,N_7743,N_6065);
and U8812 (N_8812,N_7802,N_6874);
or U8813 (N_8813,N_6367,N_6674);
nand U8814 (N_8814,N_6268,N_6608);
and U8815 (N_8815,N_7133,N_6724);
and U8816 (N_8816,N_7402,N_7078);
or U8817 (N_8817,N_6806,N_6034);
nor U8818 (N_8818,N_6740,N_7636);
or U8819 (N_8819,N_6064,N_6786);
and U8820 (N_8820,N_6302,N_7502);
nor U8821 (N_8821,N_7686,N_6641);
nand U8822 (N_8822,N_6529,N_6409);
nor U8823 (N_8823,N_6152,N_7101);
and U8824 (N_8824,N_7088,N_6829);
nand U8825 (N_8825,N_6817,N_7933);
nor U8826 (N_8826,N_6602,N_7993);
nor U8827 (N_8827,N_7832,N_7508);
and U8828 (N_8828,N_7493,N_6845);
nand U8829 (N_8829,N_7521,N_7176);
nand U8830 (N_8830,N_7849,N_6055);
nor U8831 (N_8831,N_6271,N_7770);
nor U8832 (N_8832,N_7594,N_7637);
or U8833 (N_8833,N_6439,N_6572);
nor U8834 (N_8834,N_7600,N_7911);
nand U8835 (N_8835,N_7340,N_7082);
xnor U8836 (N_8836,N_6148,N_7472);
nor U8837 (N_8837,N_6389,N_6563);
or U8838 (N_8838,N_6780,N_6798);
or U8839 (N_8839,N_7809,N_6837);
nand U8840 (N_8840,N_7790,N_6235);
nor U8841 (N_8841,N_7321,N_7057);
and U8842 (N_8842,N_7840,N_6301);
nand U8843 (N_8843,N_6649,N_6757);
or U8844 (N_8844,N_7090,N_6264);
nand U8845 (N_8845,N_6285,N_6729);
nand U8846 (N_8846,N_7834,N_6565);
nor U8847 (N_8847,N_6293,N_6498);
or U8848 (N_8848,N_7663,N_7098);
or U8849 (N_8849,N_6405,N_6455);
and U8850 (N_8850,N_7143,N_6931);
nand U8851 (N_8851,N_6402,N_6552);
or U8852 (N_8852,N_6978,N_6220);
nor U8853 (N_8853,N_6716,N_6621);
nor U8854 (N_8854,N_7135,N_7951);
nor U8855 (N_8855,N_7945,N_7336);
or U8856 (N_8856,N_7446,N_6350);
or U8857 (N_8857,N_6831,N_6793);
and U8858 (N_8858,N_7681,N_7058);
nor U8859 (N_8859,N_7705,N_7348);
or U8860 (N_8860,N_7550,N_6338);
or U8861 (N_8861,N_6992,N_7263);
and U8862 (N_8862,N_7418,N_6074);
nor U8863 (N_8863,N_6760,N_6011);
and U8864 (N_8864,N_6518,N_6037);
nand U8865 (N_8865,N_6326,N_7936);
nand U8866 (N_8866,N_7317,N_6227);
xor U8867 (N_8867,N_7638,N_7830);
xor U8868 (N_8868,N_7845,N_7957);
or U8869 (N_8869,N_7538,N_6085);
nand U8870 (N_8870,N_6143,N_6849);
or U8871 (N_8871,N_7029,N_6977);
or U8872 (N_8872,N_6759,N_6526);
and U8873 (N_8873,N_6215,N_7734);
or U8874 (N_8874,N_6894,N_7928);
or U8875 (N_8875,N_6865,N_6228);
or U8876 (N_8876,N_6966,N_7006);
nor U8877 (N_8877,N_7792,N_6069);
nand U8878 (N_8878,N_7702,N_7929);
nand U8879 (N_8879,N_7970,N_7437);
nand U8880 (N_8880,N_6984,N_7601);
and U8881 (N_8881,N_7376,N_6246);
nor U8882 (N_8882,N_7996,N_6765);
or U8883 (N_8883,N_6223,N_7346);
or U8884 (N_8884,N_6097,N_7825);
and U8885 (N_8885,N_7676,N_6096);
or U8886 (N_8886,N_6073,N_6147);
nand U8887 (N_8887,N_7252,N_6549);
or U8888 (N_8888,N_7451,N_6950);
nor U8889 (N_8889,N_7556,N_6673);
and U8890 (N_8890,N_7653,N_7954);
or U8891 (N_8891,N_6567,N_7433);
nand U8892 (N_8892,N_7560,N_6202);
nor U8893 (N_8893,N_7087,N_7440);
nand U8894 (N_8894,N_7083,N_6853);
and U8895 (N_8895,N_6879,N_7295);
and U8896 (N_8896,N_6566,N_6345);
nand U8897 (N_8897,N_6033,N_6574);
nor U8898 (N_8898,N_6427,N_7881);
or U8899 (N_8899,N_6044,N_6284);
nor U8900 (N_8900,N_7228,N_6611);
nor U8901 (N_8901,N_6005,N_7413);
or U8902 (N_8902,N_6343,N_7400);
nand U8903 (N_8903,N_6548,N_7456);
or U8904 (N_8904,N_6132,N_6938);
nand U8905 (N_8905,N_7775,N_6536);
nor U8906 (N_8906,N_7531,N_6631);
nand U8907 (N_8907,N_6506,N_7010);
nor U8908 (N_8908,N_6762,N_7562);
nand U8909 (N_8909,N_7699,N_7411);
nor U8910 (N_8910,N_6203,N_6754);
and U8911 (N_8911,N_6532,N_7125);
or U8912 (N_8912,N_6265,N_7495);
nor U8913 (N_8913,N_6001,N_7961);
nor U8914 (N_8914,N_7649,N_6230);
nand U8915 (N_8915,N_6099,N_6292);
nand U8916 (N_8916,N_7377,N_7611);
nor U8917 (N_8917,N_6233,N_7409);
nand U8918 (N_8918,N_7586,N_6819);
nor U8919 (N_8919,N_7482,N_6647);
nand U8920 (N_8920,N_6599,N_7921);
nand U8921 (N_8921,N_6531,N_6157);
and U8922 (N_8922,N_6654,N_7365);
xnor U8923 (N_8923,N_6965,N_7717);
or U8924 (N_8924,N_7497,N_7463);
nor U8925 (N_8925,N_7787,N_7170);
nand U8926 (N_8926,N_7884,N_6352);
and U8927 (N_8927,N_6750,N_7797);
nor U8928 (N_8928,N_6664,N_7439);
and U8929 (N_8929,N_7544,N_6993);
or U8930 (N_8930,N_6516,N_7719);
nor U8931 (N_8931,N_7423,N_6279);
or U8932 (N_8932,N_7219,N_6370);
or U8933 (N_8933,N_7602,N_6464);
nand U8934 (N_8934,N_6679,N_6092);
and U8935 (N_8935,N_7640,N_7530);
and U8936 (N_8936,N_7118,N_6557);
nand U8937 (N_8937,N_6184,N_6321);
and U8938 (N_8938,N_7053,N_6522);
and U8939 (N_8939,N_6947,N_7035);
nor U8940 (N_8940,N_7671,N_6682);
and U8941 (N_8941,N_6736,N_7842);
or U8942 (N_8942,N_7861,N_6095);
or U8943 (N_8943,N_7478,N_6939);
nand U8944 (N_8944,N_7969,N_7910);
nor U8945 (N_8945,N_7052,N_6973);
and U8946 (N_8946,N_7753,N_6883);
nand U8947 (N_8947,N_6587,N_6988);
or U8948 (N_8948,N_6632,N_7540);
and U8949 (N_8949,N_7403,N_7085);
nor U8950 (N_8950,N_7730,N_7963);
and U8951 (N_8951,N_7110,N_6816);
nand U8952 (N_8952,N_6422,N_6072);
or U8953 (N_8953,N_7268,N_6803);
and U8954 (N_8954,N_7227,N_7005);
nor U8955 (N_8955,N_7233,N_6626);
nor U8956 (N_8956,N_6539,N_7584);
nand U8957 (N_8957,N_6858,N_7124);
nor U8958 (N_8958,N_6094,N_6503);
nand U8959 (N_8959,N_7202,N_7587);
and U8960 (N_8960,N_7250,N_6461);
or U8961 (N_8961,N_6597,N_7137);
or U8962 (N_8962,N_7664,N_6159);
or U8963 (N_8963,N_7539,N_7609);
or U8964 (N_8964,N_7097,N_7023);
or U8965 (N_8965,N_7084,N_6122);
and U8966 (N_8966,N_6056,N_7279);
and U8967 (N_8967,N_7127,N_7129);
nor U8968 (N_8968,N_6053,N_6489);
nor U8969 (N_8969,N_6209,N_7355);
nor U8970 (N_8970,N_7131,N_6490);
nor U8971 (N_8971,N_6840,N_6511);
and U8972 (N_8972,N_7644,N_7741);
or U8973 (N_8973,N_7710,N_6123);
or U8974 (N_8974,N_6349,N_6689);
nor U8975 (N_8975,N_7816,N_6145);
or U8976 (N_8976,N_6331,N_6772);
nor U8977 (N_8977,N_7803,N_6578);
or U8978 (N_8978,N_7895,N_7162);
nor U8979 (N_8979,N_6311,N_7489);
and U8980 (N_8980,N_7487,N_6714);
nor U8981 (N_8981,N_7260,N_7622);
nor U8982 (N_8982,N_7924,N_7240);
nor U8983 (N_8983,N_7657,N_6454);
and U8984 (N_8984,N_6838,N_7920);
and U8985 (N_8985,N_6214,N_7379);
nand U8986 (N_8986,N_7626,N_7665);
and U8987 (N_8987,N_7746,N_7339);
nand U8988 (N_8988,N_6317,N_7541);
nor U8989 (N_8989,N_7164,N_6520);
nand U8990 (N_8990,N_7800,N_6584);
nor U8991 (N_8991,N_7272,N_6904);
nor U8992 (N_8992,N_6462,N_6804);
nor U8993 (N_8993,N_7779,N_6968);
nand U8994 (N_8994,N_6941,N_7758);
nor U8995 (N_8995,N_6618,N_7020);
and U8996 (N_8996,N_7571,N_6769);
nand U8997 (N_8997,N_7486,N_7658);
or U8998 (N_8998,N_7607,N_7132);
nand U8999 (N_8999,N_7013,N_6751);
nor U9000 (N_9000,N_6109,N_6577);
and U9001 (N_9001,N_7741,N_6494);
and U9002 (N_9002,N_6673,N_7394);
nor U9003 (N_9003,N_6575,N_6207);
nand U9004 (N_9004,N_7293,N_7020);
or U9005 (N_9005,N_6615,N_7616);
nand U9006 (N_9006,N_6495,N_7941);
nand U9007 (N_9007,N_6548,N_6339);
nor U9008 (N_9008,N_6757,N_6226);
and U9009 (N_9009,N_6884,N_7261);
or U9010 (N_9010,N_7548,N_7957);
or U9011 (N_9011,N_7270,N_7180);
or U9012 (N_9012,N_7823,N_7913);
or U9013 (N_9013,N_6333,N_7101);
or U9014 (N_9014,N_6052,N_6447);
nor U9015 (N_9015,N_7749,N_7461);
and U9016 (N_9016,N_7547,N_6713);
nand U9017 (N_9017,N_7156,N_6628);
nand U9018 (N_9018,N_6557,N_7763);
and U9019 (N_9019,N_6348,N_6698);
and U9020 (N_9020,N_7557,N_7423);
or U9021 (N_9021,N_6278,N_6812);
and U9022 (N_9022,N_6956,N_6542);
or U9023 (N_9023,N_6355,N_7252);
or U9024 (N_9024,N_7860,N_6983);
and U9025 (N_9025,N_6274,N_7600);
nand U9026 (N_9026,N_6055,N_6611);
and U9027 (N_9027,N_7951,N_6414);
xor U9028 (N_9028,N_7685,N_6760);
or U9029 (N_9029,N_7219,N_7493);
nand U9030 (N_9030,N_6024,N_7630);
and U9031 (N_9031,N_7626,N_7004);
nand U9032 (N_9032,N_7312,N_7868);
or U9033 (N_9033,N_7758,N_6074);
and U9034 (N_9034,N_7436,N_7080);
or U9035 (N_9035,N_6285,N_6465);
and U9036 (N_9036,N_7703,N_7547);
or U9037 (N_9037,N_6595,N_7063);
xnor U9038 (N_9038,N_7362,N_6448);
nand U9039 (N_9039,N_6443,N_6007);
xor U9040 (N_9040,N_6313,N_7925);
or U9041 (N_9041,N_7576,N_6589);
nand U9042 (N_9042,N_7478,N_7615);
nand U9043 (N_9043,N_7873,N_7388);
nand U9044 (N_9044,N_6037,N_7966);
nor U9045 (N_9045,N_7329,N_6784);
nand U9046 (N_9046,N_7119,N_7577);
and U9047 (N_9047,N_7621,N_6655);
nand U9048 (N_9048,N_7029,N_6178);
or U9049 (N_9049,N_7523,N_6139);
and U9050 (N_9050,N_7697,N_7276);
nor U9051 (N_9051,N_6336,N_6034);
or U9052 (N_9052,N_7257,N_6053);
nand U9053 (N_9053,N_6697,N_7109);
nor U9054 (N_9054,N_6266,N_6020);
nor U9055 (N_9055,N_6587,N_6539);
nand U9056 (N_9056,N_7793,N_6698);
and U9057 (N_9057,N_6768,N_7617);
or U9058 (N_9058,N_6983,N_7344);
and U9059 (N_9059,N_6893,N_7887);
and U9060 (N_9060,N_7093,N_7765);
nand U9061 (N_9061,N_6604,N_7739);
nand U9062 (N_9062,N_7750,N_6339);
nor U9063 (N_9063,N_6888,N_6400);
nand U9064 (N_9064,N_6189,N_6864);
nor U9065 (N_9065,N_6787,N_7919);
or U9066 (N_9066,N_6890,N_6125);
nand U9067 (N_9067,N_7547,N_6681);
nor U9068 (N_9068,N_6336,N_6629);
nor U9069 (N_9069,N_7779,N_6855);
or U9070 (N_9070,N_6597,N_7190);
and U9071 (N_9071,N_7987,N_6211);
and U9072 (N_9072,N_6963,N_6842);
nand U9073 (N_9073,N_7413,N_6405);
and U9074 (N_9074,N_6687,N_6212);
and U9075 (N_9075,N_6344,N_7785);
nand U9076 (N_9076,N_6072,N_6662);
nand U9077 (N_9077,N_6177,N_6585);
nand U9078 (N_9078,N_7864,N_6158);
and U9079 (N_9079,N_7789,N_6566);
nand U9080 (N_9080,N_6267,N_7962);
nand U9081 (N_9081,N_7549,N_7774);
and U9082 (N_9082,N_6415,N_7659);
or U9083 (N_9083,N_6657,N_7093);
nand U9084 (N_9084,N_6928,N_7611);
or U9085 (N_9085,N_6961,N_6073);
and U9086 (N_9086,N_6297,N_7888);
nand U9087 (N_9087,N_6962,N_7698);
or U9088 (N_9088,N_7440,N_6517);
nor U9089 (N_9089,N_7509,N_7049);
or U9090 (N_9090,N_7508,N_7619);
or U9091 (N_9091,N_7379,N_6154);
nor U9092 (N_9092,N_6210,N_6615);
and U9093 (N_9093,N_7239,N_6657);
or U9094 (N_9094,N_7980,N_7506);
or U9095 (N_9095,N_6965,N_7942);
and U9096 (N_9096,N_6863,N_7358);
nand U9097 (N_9097,N_7543,N_7557);
nor U9098 (N_9098,N_6059,N_6034);
nor U9099 (N_9099,N_6413,N_7415);
nand U9100 (N_9100,N_6816,N_7106);
and U9101 (N_9101,N_6112,N_7616);
or U9102 (N_9102,N_7172,N_7675);
or U9103 (N_9103,N_6344,N_7146);
and U9104 (N_9104,N_6426,N_6449);
or U9105 (N_9105,N_7543,N_6322);
nand U9106 (N_9106,N_7807,N_7812);
nand U9107 (N_9107,N_6413,N_6225);
and U9108 (N_9108,N_7410,N_6591);
nand U9109 (N_9109,N_6094,N_7079);
or U9110 (N_9110,N_7559,N_6515);
or U9111 (N_9111,N_6936,N_6704);
nand U9112 (N_9112,N_6569,N_7046);
nor U9113 (N_9113,N_7471,N_7693);
nand U9114 (N_9114,N_7863,N_7225);
or U9115 (N_9115,N_7546,N_7410);
or U9116 (N_9116,N_7283,N_7535);
or U9117 (N_9117,N_6327,N_7740);
and U9118 (N_9118,N_6927,N_7689);
nand U9119 (N_9119,N_7538,N_7281);
nor U9120 (N_9120,N_7367,N_7241);
nor U9121 (N_9121,N_7791,N_7807);
or U9122 (N_9122,N_7197,N_6418);
nand U9123 (N_9123,N_6832,N_6582);
xnor U9124 (N_9124,N_7074,N_7107);
nand U9125 (N_9125,N_6135,N_7777);
and U9126 (N_9126,N_6887,N_7807);
nor U9127 (N_9127,N_7048,N_7751);
or U9128 (N_9128,N_6227,N_6704);
and U9129 (N_9129,N_7277,N_7386);
or U9130 (N_9130,N_7619,N_6054);
and U9131 (N_9131,N_6305,N_7759);
nand U9132 (N_9132,N_6243,N_7910);
or U9133 (N_9133,N_6154,N_7701);
nand U9134 (N_9134,N_6970,N_6805);
nor U9135 (N_9135,N_7641,N_7534);
nor U9136 (N_9136,N_7390,N_7575);
nor U9137 (N_9137,N_6402,N_6631);
and U9138 (N_9138,N_6959,N_6833);
and U9139 (N_9139,N_7282,N_6074);
nor U9140 (N_9140,N_6983,N_7147);
nor U9141 (N_9141,N_7103,N_6118);
nand U9142 (N_9142,N_6145,N_7482);
or U9143 (N_9143,N_7886,N_6765);
nand U9144 (N_9144,N_7990,N_7308);
and U9145 (N_9145,N_7582,N_7726);
nand U9146 (N_9146,N_7948,N_6626);
nor U9147 (N_9147,N_6874,N_6023);
nor U9148 (N_9148,N_7074,N_6151);
nor U9149 (N_9149,N_6085,N_6789);
xnor U9150 (N_9150,N_6591,N_7607);
nor U9151 (N_9151,N_7762,N_6330);
nand U9152 (N_9152,N_6318,N_6216);
and U9153 (N_9153,N_7393,N_6679);
nor U9154 (N_9154,N_7416,N_6457);
nand U9155 (N_9155,N_6800,N_7962);
or U9156 (N_9156,N_7960,N_6690);
nor U9157 (N_9157,N_7988,N_6276);
or U9158 (N_9158,N_7808,N_6572);
nor U9159 (N_9159,N_6654,N_6993);
or U9160 (N_9160,N_7431,N_6073);
nand U9161 (N_9161,N_6361,N_7406);
or U9162 (N_9162,N_6230,N_7062);
nand U9163 (N_9163,N_6507,N_6865);
nor U9164 (N_9164,N_7144,N_7729);
or U9165 (N_9165,N_7862,N_6619);
and U9166 (N_9166,N_6711,N_6279);
nand U9167 (N_9167,N_6100,N_7773);
nand U9168 (N_9168,N_7334,N_7452);
nand U9169 (N_9169,N_6814,N_6836);
nor U9170 (N_9170,N_6666,N_7141);
and U9171 (N_9171,N_7309,N_7032);
nor U9172 (N_9172,N_6877,N_6782);
nor U9173 (N_9173,N_6661,N_6938);
nor U9174 (N_9174,N_7327,N_6572);
nor U9175 (N_9175,N_6526,N_6566);
nand U9176 (N_9176,N_7810,N_6442);
or U9177 (N_9177,N_6632,N_6584);
or U9178 (N_9178,N_7960,N_7091);
nand U9179 (N_9179,N_6114,N_7942);
or U9180 (N_9180,N_7140,N_7978);
nor U9181 (N_9181,N_7085,N_7188);
nor U9182 (N_9182,N_7027,N_7796);
nand U9183 (N_9183,N_6846,N_7695);
or U9184 (N_9184,N_6781,N_7524);
or U9185 (N_9185,N_6504,N_6791);
nand U9186 (N_9186,N_6560,N_6255);
nand U9187 (N_9187,N_6221,N_7135);
nor U9188 (N_9188,N_6316,N_6605);
nor U9189 (N_9189,N_6259,N_7268);
or U9190 (N_9190,N_6960,N_6295);
or U9191 (N_9191,N_7229,N_7466);
nand U9192 (N_9192,N_7206,N_6190);
or U9193 (N_9193,N_7626,N_7297);
xnor U9194 (N_9194,N_6654,N_6589);
nor U9195 (N_9195,N_7855,N_6270);
nor U9196 (N_9196,N_7133,N_6243);
nand U9197 (N_9197,N_7182,N_7273);
or U9198 (N_9198,N_6409,N_7957);
or U9199 (N_9199,N_7361,N_6198);
or U9200 (N_9200,N_7550,N_6557);
nor U9201 (N_9201,N_6547,N_7689);
or U9202 (N_9202,N_7978,N_6587);
and U9203 (N_9203,N_6031,N_7210);
or U9204 (N_9204,N_6369,N_6911);
and U9205 (N_9205,N_7439,N_7359);
xor U9206 (N_9206,N_7618,N_7728);
nor U9207 (N_9207,N_6093,N_7616);
and U9208 (N_9208,N_6092,N_7999);
and U9209 (N_9209,N_7554,N_7278);
nor U9210 (N_9210,N_7838,N_7365);
or U9211 (N_9211,N_7100,N_7719);
or U9212 (N_9212,N_7734,N_6345);
and U9213 (N_9213,N_7885,N_7614);
and U9214 (N_9214,N_7038,N_6543);
and U9215 (N_9215,N_7142,N_7627);
nor U9216 (N_9216,N_7219,N_6621);
nand U9217 (N_9217,N_7553,N_6278);
nor U9218 (N_9218,N_6459,N_7257);
or U9219 (N_9219,N_6933,N_6420);
or U9220 (N_9220,N_7953,N_7673);
or U9221 (N_9221,N_6040,N_6597);
or U9222 (N_9222,N_6934,N_6980);
nor U9223 (N_9223,N_6664,N_6168);
nor U9224 (N_9224,N_6771,N_6907);
nor U9225 (N_9225,N_6194,N_6515);
nand U9226 (N_9226,N_6493,N_7450);
nor U9227 (N_9227,N_6133,N_6323);
or U9228 (N_9228,N_7225,N_7136);
nor U9229 (N_9229,N_6532,N_6206);
xnor U9230 (N_9230,N_7570,N_7179);
nor U9231 (N_9231,N_7276,N_7719);
nand U9232 (N_9232,N_6937,N_6919);
nor U9233 (N_9233,N_7075,N_6939);
or U9234 (N_9234,N_6234,N_6652);
or U9235 (N_9235,N_6679,N_7672);
nor U9236 (N_9236,N_6801,N_6830);
and U9237 (N_9237,N_6486,N_7764);
nor U9238 (N_9238,N_6359,N_7488);
and U9239 (N_9239,N_6282,N_6443);
nand U9240 (N_9240,N_7702,N_7564);
and U9241 (N_9241,N_7833,N_7853);
and U9242 (N_9242,N_6071,N_7055);
and U9243 (N_9243,N_7183,N_6668);
nand U9244 (N_9244,N_6139,N_6044);
nor U9245 (N_9245,N_6830,N_6857);
nand U9246 (N_9246,N_6778,N_6245);
nor U9247 (N_9247,N_7612,N_6245);
and U9248 (N_9248,N_7081,N_6141);
nand U9249 (N_9249,N_6705,N_6844);
or U9250 (N_9250,N_6928,N_7803);
and U9251 (N_9251,N_7389,N_7605);
and U9252 (N_9252,N_7917,N_6842);
and U9253 (N_9253,N_6489,N_7695);
nor U9254 (N_9254,N_7526,N_6547);
or U9255 (N_9255,N_6459,N_6453);
or U9256 (N_9256,N_7025,N_6663);
or U9257 (N_9257,N_6360,N_7584);
or U9258 (N_9258,N_7184,N_7200);
nand U9259 (N_9259,N_7942,N_7330);
or U9260 (N_9260,N_6032,N_7749);
nand U9261 (N_9261,N_7960,N_6586);
nand U9262 (N_9262,N_6317,N_7783);
nor U9263 (N_9263,N_7577,N_7985);
or U9264 (N_9264,N_6779,N_7521);
nand U9265 (N_9265,N_7887,N_6615);
xnor U9266 (N_9266,N_6116,N_6088);
nand U9267 (N_9267,N_6643,N_7195);
nor U9268 (N_9268,N_7345,N_7829);
nand U9269 (N_9269,N_7090,N_7948);
and U9270 (N_9270,N_6333,N_7242);
nand U9271 (N_9271,N_7978,N_7156);
nor U9272 (N_9272,N_7573,N_7086);
nor U9273 (N_9273,N_6647,N_7299);
nor U9274 (N_9274,N_6584,N_7276);
nand U9275 (N_9275,N_7133,N_6028);
nand U9276 (N_9276,N_7770,N_7478);
or U9277 (N_9277,N_6465,N_6149);
nor U9278 (N_9278,N_6414,N_6598);
nand U9279 (N_9279,N_7944,N_6430);
or U9280 (N_9280,N_6667,N_6193);
nand U9281 (N_9281,N_6511,N_6932);
or U9282 (N_9282,N_7680,N_6127);
or U9283 (N_9283,N_7663,N_6014);
nor U9284 (N_9284,N_7244,N_6864);
or U9285 (N_9285,N_7683,N_6241);
or U9286 (N_9286,N_7632,N_6508);
nand U9287 (N_9287,N_6290,N_7398);
and U9288 (N_9288,N_7897,N_7319);
nand U9289 (N_9289,N_7681,N_6015);
or U9290 (N_9290,N_6940,N_6393);
or U9291 (N_9291,N_7545,N_7391);
or U9292 (N_9292,N_6480,N_6532);
nand U9293 (N_9293,N_6082,N_7459);
nand U9294 (N_9294,N_7096,N_7991);
or U9295 (N_9295,N_6687,N_7889);
or U9296 (N_9296,N_7613,N_7132);
nor U9297 (N_9297,N_7529,N_7735);
and U9298 (N_9298,N_6535,N_7309);
nand U9299 (N_9299,N_6471,N_6257);
nor U9300 (N_9300,N_6616,N_7043);
and U9301 (N_9301,N_7775,N_7466);
nand U9302 (N_9302,N_7385,N_7039);
nand U9303 (N_9303,N_7697,N_6818);
or U9304 (N_9304,N_7871,N_6504);
nand U9305 (N_9305,N_7594,N_7512);
and U9306 (N_9306,N_6378,N_7666);
nor U9307 (N_9307,N_7749,N_7451);
and U9308 (N_9308,N_7500,N_7156);
nand U9309 (N_9309,N_6712,N_7517);
or U9310 (N_9310,N_6691,N_6247);
and U9311 (N_9311,N_7123,N_7110);
nand U9312 (N_9312,N_6979,N_7429);
and U9313 (N_9313,N_7504,N_6557);
or U9314 (N_9314,N_6099,N_6576);
nor U9315 (N_9315,N_7672,N_6177);
or U9316 (N_9316,N_7394,N_6572);
nand U9317 (N_9317,N_6067,N_7960);
and U9318 (N_9318,N_6857,N_6681);
and U9319 (N_9319,N_6341,N_7846);
or U9320 (N_9320,N_6966,N_6061);
nor U9321 (N_9321,N_7587,N_7539);
nand U9322 (N_9322,N_6962,N_6591);
nor U9323 (N_9323,N_6915,N_6788);
xnor U9324 (N_9324,N_6019,N_7898);
nand U9325 (N_9325,N_6652,N_6705);
and U9326 (N_9326,N_6399,N_6662);
and U9327 (N_9327,N_6161,N_6737);
nor U9328 (N_9328,N_6805,N_6469);
and U9329 (N_9329,N_7700,N_7706);
nand U9330 (N_9330,N_6279,N_6218);
or U9331 (N_9331,N_7029,N_6030);
nor U9332 (N_9332,N_7764,N_6328);
nand U9333 (N_9333,N_6149,N_7583);
or U9334 (N_9334,N_6427,N_6138);
nor U9335 (N_9335,N_7806,N_6628);
nand U9336 (N_9336,N_7578,N_7806);
or U9337 (N_9337,N_7370,N_6635);
and U9338 (N_9338,N_6657,N_6474);
nor U9339 (N_9339,N_7919,N_6763);
nor U9340 (N_9340,N_7655,N_7270);
nand U9341 (N_9341,N_7059,N_7420);
nand U9342 (N_9342,N_6939,N_6646);
or U9343 (N_9343,N_7301,N_6575);
nand U9344 (N_9344,N_6501,N_7126);
xnor U9345 (N_9345,N_7521,N_7916);
nor U9346 (N_9346,N_7834,N_7882);
or U9347 (N_9347,N_6329,N_6356);
nor U9348 (N_9348,N_7871,N_6747);
nor U9349 (N_9349,N_7718,N_6710);
nor U9350 (N_9350,N_7339,N_7708);
and U9351 (N_9351,N_6858,N_7785);
and U9352 (N_9352,N_6892,N_7895);
nor U9353 (N_9353,N_7647,N_7134);
nand U9354 (N_9354,N_6196,N_6892);
nor U9355 (N_9355,N_7430,N_6006);
xnor U9356 (N_9356,N_7762,N_6924);
and U9357 (N_9357,N_7227,N_6315);
or U9358 (N_9358,N_6595,N_7228);
or U9359 (N_9359,N_7113,N_6725);
and U9360 (N_9360,N_7178,N_6166);
and U9361 (N_9361,N_7589,N_7050);
or U9362 (N_9362,N_7763,N_7490);
or U9363 (N_9363,N_7144,N_7658);
nand U9364 (N_9364,N_6492,N_6073);
or U9365 (N_9365,N_6750,N_6720);
nor U9366 (N_9366,N_7915,N_6309);
xor U9367 (N_9367,N_7243,N_6957);
and U9368 (N_9368,N_6777,N_7947);
and U9369 (N_9369,N_6382,N_7909);
and U9370 (N_9370,N_7953,N_7282);
nor U9371 (N_9371,N_7189,N_7115);
xor U9372 (N_9372,N_7050,N_7375);
nor U9373 (N_9373,N_7710,N_6368);
nor U9374 (N_9374,N_7356,N_7382);
nand U9375 (N_9375,N_6973,N_7507);
and U9376 (N_9376,N_6769,N_6500);
nand U9377 (N_9377,N_6202,N_7305);
or U9378 (N_9378,N_7482,N_7536);
or U9379 (N_9379,N_6295,N_7744);
or U9380 (N_9380,N_6319,N_6602);
or U9381 (N_9381,N_6865,N_6860);
nand U9382 (N_9382,N_6097,N_6001);
or U9383 (N_9383,N_7706,N_7741);
nor U9384 (N_9384,N_6630,N_6668);
nand U9385 (N_9385,N_7281,N_7991);
or U9386 (N_9386,N_7216,N_6345);
and U9387 (N_9387,N_7904,N_6610);
and U9388 (N_9388,N_7348,N_6413);
or U9389 (N_9389,N_6098,N_6825);
or U9390 (N_9390,N_7912,N_7863);
nor U9391 (N_9391,N_7696,N_6982);
nor U9392 (N_9392,N_6676,N_7053);
or U9393 (N_9393,N_6689,N_7760);
nor U9394 (N_9394,N_6473,N_7095);
nand U9395 (N_9395,N_6203,N_6224);
nand U9396 (N_9396,N_7725,N_6777);
and U9397 (N_9397,N_6075,N_7027);
xor U9398 (N_9398,N_6880,N_7058);
nor U9399 (N_9399,N_7599,N_7237);
and U9400 (N_9400,N_6538,N_7917);
or U9401 (N_9401,N_7617,N_6687);
or U9402 (N_9402,N_6795,N_6480);
and U9403 (N_9403,N_6286,N_7558);
and U9404 (N_9404,N_7543,N_7042);
or U9405 (N_9405,N_6041,N_6264);
and U9406 (N_9406,N_6632,N_6989);
and U9407 (N_9407,N_6896,N_7232);
and U9408 (N_9408,N_7682,N_6918);
or U9409 (N_9409,N_6994,N_6542);
or U9410 (N_9410,N_7260,N_7480);
nor U9411 (N_9411,N_6224,N_7354);
and U9412 (N_9412,N_7318,N_6945);
and U9413 (N_9413,N_6167,N_7722);
nor U9414 (N_9414,N_7878,N_6059);
and U9415 (N_9415,N_6857,N_6115);
or U9416 (N_9416,N_6177,N_7500);
or U9417 (N_9417,N_6890,N_6291);
nand U9418 (N_9418,N_7418,N_6912);
nand U9419 (N_9419,N_6874,N_6672);
or U9420 (N_9420,N_7691,N_7197);
or U9421 (N_9421,N_6496,N_7472);
nand U9422 (N_9422,N_6964,N_6081);
nand U9423 (N_9423,N_6614,N_7922);
nor U9424 (N_9424,N_7068,N_7126);
nor U9425 (N_9425,N_6169,N_6983);
or U9426 (N_9426,N_6116,N_7986);
nor U9427 (N_9427,N_6135,N_6764);
and U9428 (N_9428,N_6577,N_7349);
or U9429 (N_9429,N_6489,N_6573);
or U9430 (N_9430,N_7688,N_7120);
and U9431 (N_9431,N_6072,N_6815);
or U9432 (N_9432,N_7072,N_7340);
and U9433 (N_9433,N_6105,N_7817);
nand U9434 (N_9434,N_6170,N_7819);
nor U9435 (N_9435,N_6521,N_7075);
nor U9436 (N_9436,N_6458,N_7908);
and U9437 (N_9437,N_7060,N_6303);
nand U9438 (N_9438,N_7709,N_6233);
nand U9439 (N_9439,N_7707,N_6263);
and U9440 (N_9440,N_7434,N_6029);
nor U9441 (N_9441,N_6939,N_6748);
or U9442 (N_9442,N_6060,N_7652);
and U9443 (N_9443,N_7072,N_6123);
and U9444 (N_9444,N_7893,N_6197);
nor U9445 (N_9445,N_6616,N_7888);
nand U9446 (N_9446,N_6087,N_7338);
nor U9447 (N_9447,N_6202,N_6362);
nor U9448 (N_9448,N_6734,N_6796);
or U9449 (N_9449,N_6477,N_7109);
nand U9450 (N_9450,N_7782,N_7161);
nor U9451 (N_9451,N_6493,N_7923);
xor U9452 (N_9452,N_6078,N_6357);
nor U9453 (N_9453,N_7326,N_6699);
or U9454 (N_9454,N_6960,N_7368);
nor U9455 (N_9455,N_7916,N_7495);
nand U9456 (N_9456,N_6288,N_6810);
and U9457 (N_9457,N_7790,N_7078);
nand U9458 (N_9458,N_7228,N_6427);
and U9459 (N_9459,N_6002,N_7580);
nand U9460 (N_9460,N_7471,N_7202);
nand U9461 (N_9461,N_7538,N_7772);
or U9462 (N_9462,N_7286,N_7255);
xor U9463 (N_9463,N_7300,N_7351);
and U9464 (N_9464,N_7333,N_6186);
nand U9465 (N_9465,N_6888,N_7494);
or U9466 (N_9466,N_6137,N_7174);
nand U9467 (N_9467,N_7916,N_7663);
and U9468 (N_9468,N_7804,N_6645);
nor U9469 (N_9469,N_7724,N_6670);
nand U9470 (N_9470,N_6079,N_6089);
nand U9471 (N_9471,N_6541,N_7059);
nand U9472 (N_9472,N_7516,N_6127);
nor U9473 (N_9473,N_6215,N_7180);
and U9474 (N_9474,N_6303,N_7640);
or U9475 (N_9475,N_6794,N_7967);
and U9476 (N_9476,N_6385,N_6727);
and U9477 (N_9477,N_6705,N_7052);
or U9478 (N_9478,N_7795,N_7995);
nor U9479 (N_9479,N_6784,N_7270);
nor U9480 (N_9480,N_6795,N_6587);
and U9481 (N_9481,N_7947,N_7656);
or U9482 (N_9482,N_7473,N_6412);
nand U9483 (N_9483,N_6033,N_6812);
nand U9484 (N_9484,N_6435,N_6531);
or U9485 (N_9485,N_7153,N_6939);
nor U9486 (N_9486,N_6177,N_6031);
or U9487 (N_9487,N_6403,N_7177);
and U9488 (N_9488,N_6288,N_7175);
and U9489 (N_9489,N_7813,N_7131);
and U9490 (N_9490,N_6746,N_7319);
nand U9491 (N_9491,N_6285,N_7167);
and U9492 (N_9492,N_6536,N_6145);
or U9493 (N_9493,N_7405,N_6687);
nand U9494 (N_9494,N_6419,N_7468);
nor U9495 (N_9495,N_7621,N_7838);
nand U9496 (N_9496,N_7633,N_6477);
or U9497 (N_9497,N_6576,N_7978);
and U9498 (N_9498,N_7384,N_7278);
nor U9499 (N_9499,N_6849,N_7004);
nor U9500 (N_9500,N_7263,N_7149);
or U9501 (N_9501,N_7347,N_6094);
nand U9502 (N_9502,N_7959,N_7624);
and U9503 (N_9503,N_6128,N_6415);
and U9504 (N_9504,N_7144,N_7026);
nand U9505 (N_9505,N_7812,N_7003);
and U9506 (N_9506,N_7831,N_7397);
or U9507 (N_9507,N_6963,N_7549);
nand U9508 (N_9508,N_7259,N_7166);
nand U9509 (N_9509,N_6523,N_7087);
nand U9510 (N_9510,N_7892,N_7014);
and U9511 (N_9511,N_6049,N_7145);
or U9512 (N_9512,N_6715,N_6157);
nand U9513 (N_9513,N_7154,N_7268);
or U9514 (N_9514,N_6240,N_6979);
xnor U9515 (N_9515,N_6905,N_7963);
or U9516 (N_9516,N_7057,N_7645);
nor U9517 (N_9517,N_7614,N_7503);
and U9518 (N_9518,N_7892,N_7367);
nor U9519 (N_9519,N_7168,N_6491);
or U9520 (N_9520,N_6854,N_6311);
and U9521 (N_9521,N_6920,N_6244);
and U9522 (N_9522,N_6326,N_7302);
nor U9523 (N_9523,N_6744,N_7989);
nor U9524 (N_9524,N_6348,N_6392);
nor U9525 (N_9525,N_6844,N_6030);
and U9526 (N_9526,N_7861,N_6399);
nor U9527 (N_9527,N_6626,N_6366);
nand U9528 (N_9528,N_7182,N_7157);
nand U9529 (N_9529,N_6126,N_6665);
and U9530 (N_9530,N_6659,N_6055);
or U9531 (N_9531,N_7104,N_7164);
nor U9532 (N_9532,N_6170,N_6527);
or U9533 (N_9533,N_6128,N_7878);
or U9534 (N_9534,N_6060,N_6642);
nor U9535 (N_9535,N_6226,N_6980);
or U9536 (N_9536,N_7071,N_7986);
or U9537 (N_9537,N_6820,N_7563);
nand U9538 (N_9538,N_7892,N_7521);
or U9539 (N_9539,N_6572,N_6333);
and U9540 (N_9540,N_7783,N_6407);
and U9541 (N_9541,N_6298,N_7543);
and U9542 (N_9542,N_7583,N_6443);
and U9543 (N_9543,N_7842,N_7848);
and U9544 (N_9544,N_6187,N_6501);
nor U9545 (N_9545,N_7245,N_7991);
and U9546 (N_9546,N_6372,N_7414);
nand U9547 (N_9547,N_7154,N_7251);
or U9548 (N_9548,N_7016,N_6348);
or U9549 (N_9549,N_6604,N_7222);
nand U9550 (N_9550,N_6368,N_7301);
nor U9551 (N_9551,N_7785,N_6292);
or U9552 (N_9552,N_6684,N_7892);
or U9553 (N_9553,N_6898,N_6148);
nor U9554 (N_9554,N_7446,N_6677);
and U9555 (N_9555,N_6241,N_7860);
or U9556 (N_9556,N_7045,N_7888);
and U9557 (N_9557,N_6653,N_7296);
nor U9558 (N_9558,N_6566,N_6891);
nor U9559 (N_9559,N_7436,N_6748);
or U9560 (N_9560,N_6818,N_7877);
nor U9561 (N_9561,N_6250,N_6696);
nand U9562 (N_9562,N_7019,N_6316);
or U9563 (N_9563,N_6183,N_6633);
nor U9564 (N_9564,N_6339,N_7452);
or U9565 (N_9565,N_7486,N_7061);
or U9566 (N_9566,N_7301,N_6217);
or U9567 (N_9567,N_7438,N_7676);
nor U9568 (N_9568,N_7506,N_7868);
nand U9569 (N_9569,N_6735,N_7549);
nand U9570 (N_9570,N_6014,N_7934);
or U9571 (N_9571,N_6460,N_7919);
and U9572 (N_9572,N_7195,N_7211);
or U9573 (N_9573,N_7290,N_6997);
or U9574 (N_9574,N_7753,N_7584);
nand U9575 (N_9575,N_6052,N_7286);
nor U9576 (N_9576,N_6590,N_6553);
nand U9577 (N_9577,N_6771,N_7543);
or U9578 (N_9578,N_7804,N_7809);
and U9579 (N_9579,N_6114,N_6438);
nor U9580 (N_9580,N_7682,N_6549);
nor U9581 (N_9581,N_7128,N_6102);
nand U9582 (N_9582,N_6665,N_6107);
or U9583 (N_9583,N_7495,N_7057);
nand U9584 (N_9584,N_6402,N_7481);
nor U9585 (N_9585,N_6482,N_7963);
and U9586 (N_9586,N_7376,N_7310);
nand U9587 (N_9587,N_7167,N_7138);
or U9588 (N_9588,N_6368,N_7086);
or U9589 (N_9589,N_6630,N_6891);
and U9590 (N_9590,N_7425,N_6438);
or U9591 (N_9591,N_7647,N_7880);
nor U9592 (N_9592,N_7981,N_6219);
and U9593 (N_9593,N_7016,N_6641);
nor U9594 (N_9594,N_6640,N_6091);
or U9595 (N_9595,N_7579,N_7788);
nor U9596 (N_9596,N_7505,N_7464);
nor U9597 (N_9597,N_6910,N_7216);
nand U9598 (N_9598,N_6075,N_7597);
and U9599 (N_9599,N_7811,N_7963);
nor U9600 (N_9600,N_7587,N_7030);
or U9601 (N_9601,N_7743,N_7672);
nand U9602 (N_9602,N_7503,N_6233);
nand U9603 (N_9603,N_7450,N_6608);
nor U9604 (N_9604,N_6423,N_6264);
nor U9605 (N_9605,N_7289,N_7986);
and U9606 (N_9606,N_7126,N_7141);
nor U9607 (N_9607,N_7669,N_6704);
nor U9608 (N_9608,N_7952,N_6954);
nand U9609 (N_9609,N_6874,N_6614);
and U9610 (N_9610,N_6573,N_7632);
nand U9611 (N_9611,N_6789,N_6917);
or U9612 (N_9612,N_6994,N_7642);
nand U9613 (N_9613,N_6914,N_7534);
nor U9614 (N_9614,N_7822,N_7332);
or U9615 (N_9615,N_6178,N_6427);
nor U9616 (N_9616,N_7604,N_7370);
and U9617 (N_9617,N_7702,N_6649);
nor U9618 (N_9618,N_7025,N_6031);
nand U9619 (N_9619,N_6021,N_6398);
nand U9620 (N_9620,N_7705,N_6156);
nor U9621 (N_9621,N_6204,N_6114);
nand U9622 (N_9622,N_7937,N_7548);
nor U9623 (N_9623,N_7493,N_6932);
nor U9624 (N_9624,N_6274,N_7122);
or U9625 (N_9625,N_7338,N_7754);
nor U9626 (N_9626,N_7851,N_6137);
and U9627 (N_9627,N_6459,N_7283);
nand U9628 (N_9628,N_7713,N_6637);
nor U9629 (N_9629,N_6382,N_7265);
nor U9630 (N_9630,N_6695,N_6905);
nand U9631 (N_9631,N_6368,N_7702);
nand U9632 (N_9632,N_7128,N_7212);
nor U9633 (N_9633,N_6383,N_7965);
or U9634 (N_9634,N_7314,N_6497);
and U9635 (N_9635,N_6258,N_6263);
nor U9636 (N_9636,N_7688,N_7296);
nand U9637 (N_9637,N_7495,N_7869);
nand U9638 (N_9638,N_6741,N_6954);
nor U9639 (N_9639,N_7915,N_7857);
nand U9640 (N_9640,N_6211,N_6720);
or U9641 (N_9641,N_7963,N_7361);
xnor U9642 (N_9642,N_6827,N_6958);
nor U9643 (N_9643,N_7939,N_6792);
and U9644 (N_9644,N_6572,N_6042);
nor U9645 (N_9645,N_6413,N_6001);
and U9646 (N_9646,N_6280,N_6015);
nand U9647 (N_9647,N_7197,N_6667);
and U9648 (N_9648,N_6637,N_6052);
nor U9649 (N_9649,N_7216,N_6804);
or U9650 (N_9650,N_7947,N_6009);
nor U9651 (N_9651,N_7988,N_6729);
or U9652 (N_9652,N_7730,N_6522);
and U9653 (N_9653,N_7179,N_7364);
nor U9654 (N_9654,N_7405,N_7784);
and U9655 (N_9655,N_6846,N_7125);
or U9656 (N_9656,N_7543,N_6813);
and U9657 (N_9657,N_6411,N_7338);
nor U9658 (N_9658,N_7296,N_7106);
and U9659 (N_9659,N_7618,N_7311);
xor U9660 (N_9660,N_7026,N_7792);
or U9661 (N_9661,N_6429,N_6746);
or U9662 (N_9662,N_7305,N_7238);
nor U9663 (N_9663,N_7785,N_7889);
and U9664 (N_9664,N_7055,N_6148);
or U9665 (N_9665,N_6751,N_7678);
nor U9666 (N_9666,N_6695,N_7385);
nand U9667 (N_9667,N_6615,N_7290);
and U9668 (N_9668,N_6572,N_6699);
or U9669 (N_9669,N_7591,N_6664);
nand U9670 (N_9670,N_6943,N_7904);
and U9671 (N_9671,N_7198,N_7076);
nand U9672 (N_9672,N_6538,N_6754);
nand U9673 (N_9673,N_7576,N_7684);
nor U9674 (N_9674,N_7404,N_6521);
and U9675 (N_9675,N_6820,N_6459);
xor U9676 (N_9676,N_6587,N_6699);
xnor U9677 (N_9677,N_6340,N_7247);
xor U9678 (N_9678,N_7296,N_6477);
or U9679 (N_9679,N_7221,N_7442);
nor U9680 (N_9680,N_7225,N_7651);
nor U9681 (N_9681,N_6124,N_6188);
or U9682 (N_9682,N_7913,N_7056);
and U9683 (N_9683,N_6735,N_7496);
and U9684 (N_9684,N_7772,N_6877);
and U9685 (N_9685,N_6809,N_7519);
nand U9686 (N_9686,N_7045,N_7808);
nand U9687 (N_9687,N_6727,N_6047);
or U9688 (N_9688,N_6930,N_6671);
or U9689 (N_9689,N_7488,N_7283);
nor U9690 (N_9690,N_6266,N_6658);
and U9691 (N_9691,N_7797,N_7153);
nor U9692 (N_9692,N_6801,N_6977);
and U9693 (N_9693,N_7427,N_6359);
and U9694 (N_9694,N_7368,N_7623);
nand U9695 (N_9695,N_7193,N_7072);
nand U9696 (N_9696,N_7821,N_6378);
or U9697 (N_9697,N_6054,N_6297);
nor U9698 (N_9698,N_7772,N_6911);
or U9699 (N_9699,N_7829,N_6923);
nand U9700 (N_9700,N_7479,N_7802);
nand U9701 (N_9701,N_6397,N_6121);
nand U9702 (N_9702,N_6479,N_6280);
or U9703 (N_9703,N_6287,N_6181);
nor U9704 (N_9704,N_6390,N_6848);
nor U9705 (N_9705,N_7554,N_7124);
and U9706 (N_9706,N_7019,N_6983);
nand U9707 (N_9707,N_7314,N_6948);
nor U9708 (N_9708,N_6888,N_6530);
nand U9709 (N_9709,N_6729,N_7415);
nand U9710 (N_9710,N_7704,N_7247);
and U9711 (N_9711,N_7289,N_6365);
nor U9712 (N_9712,N_6066,N_6754);
or U9713 (N_9713,N_7622,N_6475);
nand U9714 (N_9714,N_7460,N_6530);
nor U9715 (N_9715,N_7421,N_7383);
nand U9716 (N_9716,N_7993,N_6370);
and U9717 (N_9717,N_6984,N_7538);
and U9718 (N_9718,N_7259,N_7870);
nand U9719 (N_9719,N_6155,N_7035);
nor U9720 (N_9720,N_6940,N_6133);
and U9721 (N_9721,N_6769,N_7943);
nor U9722 (N_9722,N_6945,N_7806);
or U9723 (N_9723,N_7095,N_7164);
nand U9724 (N_9724,N_7184,N_6971);
nor U9725 (N_9725,N_6611,N_7262);
nor U9726 (N_9726,N_6777,N_7824);
nand U9727 (N_9727,N_7749,N_7936);
nor U9728 (N_9728,N_7552,N_6816);
nor U9729 (N_9729,N_6956,N_6545);
nand U9730 (N_9730,N_6718,N_6419);
nand U9731 (N_9731,N_6312,N_7654);
nor U9732 (N_9732,N_7567,N_6658);
or U9733 (N_9733,N_7055,N_7094);
nand U9734 (N_9734,N_6223,N_6960);
or U9735 (N_9735,N_7973,N_7429);
nor U9736 (N_9736,N_7532,N_7720);
nor U9737 (N_9737,N_6415,N_7730);
and U9738 (N_9738,N_6547,N_6316);
nand U9739 (N_9739,N_6303,N_6465);
and U9740 (N_9740,N_7649,N_6916);
or U9741 (N_9741,N_6279,N_7063);
nor U9742 (N_9742,N_6056,N_7254);
and U9743 (N_9743,N_7839,N_6065);
and U9744 (N_9744,N_6096,N_7232);
and U9745 (N_9745,N_7884,N_6048);
and U9746 (N_9746,N_6510,N_6948);
or U9747 (N_9747,N_6826,N_6169);
nand U9748 (N_9748,N_7315,N_7308);
or U9749 (N_9749,N_6800,N_6717);
and U9750 (N_9750,N_7254,N_6900);
nand U9751 (N_9751,N_7630,N_7122);
nor U9752 (N_9752,N_6981,N_7757);
and U9753 (N_9753,N_7740,N_6266);
nand U9754 (N_9754,N_7009,N_6372);
nand U9755 (N_9755,N_7701,N_7231);
or U9756 (N_9756,N_7338,N_6574);
or U9757 (N_9757,N_7419,N_7620);
nand U9758 (N_9758,N_7021,N_6057);
nand U9759 (N_9759,N_7651,N_7491);
or U9760 (N_9760,N_7167,N_7973);
nor U9761 (N_9761,N_6795,N_7854);
and U9762 (N_9762,N_7022,N_6864);
nand U9763 (N_9763,N_7714,N_6180);
nand U9764 (N_9764,N_7901,N_7438);
or U9765 (N_9765,N_6284,N_6448);
nor U9766 (N_9766,N_6916,N_6533);
nand U9767 (N_9767,N_7757,N_6764);
nor U9768 (N_9768,N_6512,N_6279);
and U9769 (N_9769,N_6781,N_7749);
nor U9770 (N_9770,N_7787,N_7357);
and U9771 (N_9771,N_6159,N_7654);
and U9772 (N_9772,N_6448,N_6972);
nand U9773 (N_9773,N_6496,N_6288);
nor U9774 (N_9774,N_7011,N_7232);
nor U9775 (N_9775,N_6914,N_6107);
nor U9776 (N_9776,N_7755,N_7570);
or U9777 (N_9777,N_6885,N_6481);
nand U9778 (N_9778,N_7044,N_7218);
and U9779 (N_9779,N_7408,N_6211);
nand U9780 (N_9780,N_6006,N_7230);
or U9781 (N_9781,N_7100,N_6775);
nand U9782 (N_9782,N_7841,N_7067);
or U9783 (N_9783,N_6538,N_7766);
and U9784 (N_9784,N_7670,N_7604);
or U9785 (N_9785,N_6580,N_6673);
nor U9786 (N_9786,N_7961,N_7891);
and U9787 (N_9787,N_6548,N_7217);
and U9788 (N_9788,N_7044,N_7774);
xor U9789 (N_9789,N_7522,N_7189);
nand U9790 (N_9790,N_6499,N_7812);
or U9791 (N_9791,N_6519,N_7189);
nor U9792 (N_9792,N_6060,N_7715);
or U9793 (N_9793,N_7902,N_6613);
nand U9794 (N_9794,N_6211,N_7278);
and U9795 (N_9795,N_6282,N_7165);
nor U9796 (N_9796,N_7262,N_7139);
or U9797 (N_9797,N_6711,N_7270);
nor U9798 (N_9798,N_6275,N_6303);
and U9799 (N_9799,N_7170,N_7454);
and U9800 (N_9800,N_7867,N_7283);
and U9801 (N_9801,N_7157,N_7551);
and U9802 (N_9802,N_6319,N_6338);
or U9803 (N_9803,N_6785,N_7490);
nand U9804 (N_9804,N_6862,N_7073);
nand U9805 (N_9805,N_7797,N_6023);
and U9806 (N_9806,N_6833,N_6899);
nand U9807 (N_9807,N_7557,N_7996);
nand U9808 (N_9808,N_7319,N_7489);
and U9809 (N_9809,N_7505,N_7850);
and U9810 (N_9810,N_7656,N_6363);
or U9811 (N_9811,N_6861,N_7305);
or U9812 (N_9812,N_6834,N_6258);
or U9813 (N_9813,N_6519,N_6986);
or U9814 (N_9814,N_7074,N_6210);
and U9815 (N_9815,N_7520,N_7592);
nand U9816 (N_9816,N_6334,N_6764);
nand U9817 (N_9817,N_7874,N_6867);
or U9818 (N_9818,N_6895,N_7085);
and U9819 (N_9819,N_6113,N_6148);
and U9820 (N_9820,N_7040,N_6454);
and U9821 (N_9821,N_6281,N_6416);
or U9822 (N_9822,N_6690,N_7078);
or U9823 (N_9823,N_6342,N_7506);
nor U9824 (N_9824,N_6384,N_6044);
nand U9825 (N_9825,N_7177,N_7325);
or U9826 (N_9826,N_6837,N_7001);
nand U9827 (N_9827,N_7081,N_7424);
nand U9828 (N_9828,N_7516,N_7607);
and U9829 (N_9829,N_6146,N_6589);
and U9830 (N_9830,N_6645,N_7125);
or U9831 (N_9831,N_7125,N_7245);
nand U9832 (N_9832,N_6084,N_6346);
nand U9833 (N_9833,N_7413,N_7076);
nand U9834 (N_9834,N_7070,N_6725);
or U9835 (N_9835,N_7770,N_6516);
or U9836 (N_9836,N_6641,N_7934);
nor U9837 (N_9837,N_6045,N_7050);
nand U9838 (N_9838,N_7505,N_6896);
and U9839 (N_9839,N_6622,N_6550);
and U9840 (N_9840,N_6488,N_7278);
or U9841 (N_9841,N_7073,N_6260);
or U9842 (N_9842,N_7256,N_7896);
and U9843 (N_9843,N_6158,N_6291);
nor U9844 (N_9844,N_6626,N_6538);
nor U9845 (N_9845,N_7479,N_6793);
or U9846 (N_9846,N_6579,N_6315);
nor U9847 (N_9847,N_6911,N_7496);
or U9848 (N_9848,N_7196,N_6990);
and U9849 (N_9849,N_6988,N_7236);
and U9850 (N_9850,N_6041,N_7414);
xor U9851 (N_9851,N_7275,N_7672);
or U9852 (N_9852,N_7631,N_7463);
nand U9853 (N_9853,N_6150,N_7193);
nand U9854 (N_9854,N_7023,N_7856);
nor U9855 (N_9855,N_6110,N_6307);
or U9856 (N_9856,N_6824,N_7382);
or U9857 (N_9857,N_7142,N_7567);
nor U9858 (N_9858,N_7054,N_6642);
and U9859 (N_9859,N_6721,N_7347);
nand U9860 (N_9860,N_6960,N_7382);
nand U9861 (N_9861,N_6228,N_7350);
and U9862 (N_9862,N_6238,N_6823);
and U9863 (N_9863,N_7198,N_7233);
and U9864 (N_9864,N_7832,N_7497);
and U9865 (N_9865,N_7974,N_7257);
nor U9866 (N_9866,N_6832,N_6254);
or U9867 (N_9867,N_7324,N_6254);
nor U9868 (N_9868,N_6596,N_6678);
and U9869 (N_9869,N_6505,N_7148);
and U9870 (N_9870,N_6185,N_7493);
nand U9871 (N_9871,N_6096,N_7564);
or U9872 (N_9872,N_7934,N_6855);
nor U9873 (N_9873,N_6057,N_7012);
or U9874 (N_9874,N_7866,N_6849);
nor U9875 (N_9875,N_6173,N_7893);
and U9876 (N_9876,N_7367,N_7719);
or U9877 (N_9877,N_7803,N_6316);
nand U9878 (N_9878,N_6571,N_6144);
xnor U9879 (N_9879,N_6144,N_6841);
nor U9880 (N_9880,N_7066,N_7251);
or U9881 (N_9881,N_6551,N_6037);
nand U9882 (N_9882,N_7311,N_6542);
nor U9883 (N_9883,N_7623,N_7058);
nand U9884 (N_9884,N_7622,N_6547);
nand U9885 (N_9885,N_7925,N_6263);
nand U9886 (N_9886,N_7201,N_7754);
and U9887 (N_9887,N_7975,N_7203);
or U9888 (N_9888,N_7463,N_6383);
nand U9889 (N_9889,N_7940,N_7274);
nor U9890 (N_9890,N_6974,N_6588);
or U9891 (N_9891,N_7542,N_7154);
nor U9892 (N_9892,N_7520,N_7453);
nand U9893 (N_9893,N_6996,N_7874);
and U9894 (N_9894,N_7831,N_7245);
or U9895 (N_9895,N_6293,N_7756);
or U9896 (N_9896,N_7073,N_6717);
nor U9897 (N_9897,N_6803,N_6330);
and U9898 (N_9898,N_7603,N_6381);
nor U9899 (N_9899,N_6976,N_6963);
nand U9900 (N_9900,N_7078,N_6033);
and U9901 (N_9901,N_7796,N_7368);
nand U9902 (N_9902,N_6333,N_6902);
or U9903 (N_9903,N_6355,N_6520);
nand U9904 (N_9904,N_7344,N_7747);
and U9905 (N_9905,N_7141,N_6452);
nand U9906 (N_9906,N_7605,N_6959);
nand U9907 (N_9907,N_7502,N_6619);
nor U9908 (N_9908,N_6915,N_7966);
nor U9909 (N_9909,N_6998,N_6443);
or U9910 (N_9910,N_7806,N_7004);
nor U9911 (N_9911,N_7358,N_7623);
or U9912 (N_9912,N_7322,N_6044);
or U9913 (N_9913,N_7183,N_6739);
nand U9914 (N_9914,N_6692,N_7110);
and U9915 (N_9915,N_7814,N_6307);
nor U9916 (N_9916,N_6315,N_7432);
nand U9917 (N_9917,N_6555,N_7551);
and U9918 (N_9918,N_7260,N_6627);
and U9919 (N_9919,N_6479,N_7901);
and U9920 (N_9920,N_6247,N_7883);
and U9921 (N_9921,N_6877,N_7078);
nand U9922 (N_9922,N_6631,N_7574);
xor U9923 (N_9923,N_6279,N_6131);
nand U9924 (N_9924,N_6647,N_6709);
nand U9925 (N_9925,N_7971,N_6093);
or U9926 (N_9926,N_6261,N_7470);
nand U9927 (N_9927,N_7754,N_7932);
nand U9928 (N_9928,N_7918,N_6208);
nand U9929 (N_9929,N_7873,N_7074);
nor U9930 (N_9930,N_7531,N_7379);
nand U9931 (N_9931,N_6838,N_7916);
xor U9932 (N_9932,N_7091,N_7352);
nand U9933 (N_9933,N_7632,N_7809);
nor U9934 (N_9934,N_6088,N_7545);
nand U9935 (N_9935,N_6075,N_7031);
xnor U9936 (N_9936,N_6188,N_7355);
nor U9937 (N_9937,N_7514,N_6303);
nand U9938 (N_9938,N_7605,N_7340);
and U9939 (N_9939,N_6727,N_6514);
or U9940 (N_9940,N_6181,N_7683);
or U9941 (N_9941,N_6331,N_6284);
or U9942 (N_9942,N_6986,N_7510);
nand U9943 (N_9943,N_7527,N_6992);
and U9944 (N_9944,N_7677,N_7320);
and U9945 (N_9945,N_6711,N_7576);
xnor U9946 (N_9946,N_7396,N_7966);
or U9947 (N_9947,N_6383,N_7271);
nand U9948 (N_9948,N_7316,N_6281);
or U9949 (N_9949,N_7494,N_7096);
nor U9950 (N_9950,N_6644,N_7551);
and U9951 (N_9951,N_6729,N_6332);
or U9952 (N_9952,N_7915,N_6727);
nor U9953 (N_9953,N_6489,N_7011);
or U9954 (N_9954,N_7570,N_6108);
nor U9955 (N_9955,N_7567,N_6464);
or U9956 (N_9956,N_7505,N_7206);
and U9957 (N_9957,N_6046,N_6833);
nand U9958 (N_9958,N_7023,N_7462);
or U9959 (N_9959,N_7836,N_6190);
or U9960 (N_9960,N_7154,N_6662);
nand U9961 (N_9961,N_7821,N_7610);
and U9962 (N_9962,N_6501,N_6167);
nand U9963 (N_9963,N_7293,N_7392);
nand U9964 (N_9964,N_7739,N_7711);
nand U9965 (N_9965,N_7168,N_7832);
nand U9966 (N_9966,N_7280,N_6207);
nor U9967 (N_9967,N_6750,N_6968);
and U9968 (N_9968,N_6001,N_6503);
nor U9969 (N_9969,N_6354,N_7813);
nand U9970 (N_9970,N_6183,N_6877);
nor U9971 (N_9971,N_6531,N_7459);
nor U9972 (N_9972,N_6004,N_6409);
xnor U9973 (N_9973,N_6659,N_7980);
nand U9974 (N_9974,N_6196,N_7452);
nor U9975 (N_9975,N_7147,N_7647);
or U9976 (N_9976,N_7668,N_7516);
nor U9977 (N_9977,N_6617,N_7184);
nor U9978 (N_9978,N_6454,N_6071);
nand U9979 (N_9979,N_6508,N_6984);
and U9980 (N_9980,N_6669,N_7617);
and U9981 (N_9981,N_6957,N_6548);
nand U9982 (N_9982,N_6502,N_6110);
or U9983 (N_9983,N_6716,N_7667);
and U9984 (N_9984,N_6159,N_6628);
and U9985 (N_9985,N_6010,N_6972);
or U9986 (N_9986,N_6105,N_7995);
and U9987 (N_9987,N_6865,N_6319);
or U9988 (N_9988,N_6513,N_6620);
or U9989 (N_9989,N_6040,N_6794);
nor U9990 (N_9990,N_6335,N_6041);
or U9991 (N_9991,N_7279,N_7702);
and U9992 (N_9992,N_6529,N_7288);
and U9993 (N_9993,N_6994,N_6746);
nand U9994 (N_9994,N_7249,N_6096);
and U9995 (N_9995,N_6496,N_6531);
nor U9996 (N_9996,N_6008,N_7248);
nor U9997 (N_9997,N_6327,N_7264);
and U9998 (N_9998,N_6296,N_6078);
and U9999 (N_9999,N_6627,N_6643);
nand U10000 (N_10000,N_9441,N_9345);
nand U10001 (N_10001,N_9991,N_9837);
or U10002 (N_10002,N_9839,N_9537);
xnor U10003 (N_10003,N_9903,N_9484);
and U10004 (N_10004,N_9107,N_9931);
xor U10005 (N_10005,N_9965,N_8917);
or U10006 (N_10006,N_8809,N_8580);
nand U10007 (N_10007,N_9809,N_8683);
nand U10008 (N_10008,N_8091,N_8819);
nand U10009 (N_10009,N_9076,N_8174);
and U10010 (N_10010,N_8878,N_9246);
nor U10011 (N_10011,N_8473,N_8121);
nand U10012 (N_10012,N_9170,N_8745);
or U10013 (N_10013,N_9379,N_9130);
nand U10014 (N_10014,N_8669,N_9320);
or U10015 (N_10015,N_8957,N_8805);
and U10016 (N_10016,N_9531,N_8789);
nor U10017 (N_10017,N_8800,N_8196);
or U10018 (N_10018,N_8513,N_8936);
or U10019 (N_10019,N_8245,N_9672);
or U10020 (N_10020,N_9536,N_9619);
nand U10021 (N_10021,N_8737,N_8301);
and U10022 (N_10022,N_8511,N_9288);
and U10023 (N_10023,N_8066,N_8356);
nand U10024 (N_10024,N_9756,N_9408);
or U10025 (N_10025,N_9138,N_8489);
and U10026 (N_10026,N_8642,N_9272);
or U10027 (N_10027,N_9396,N_9593);
or U10028 (N_10028,N_9274,N_8775);
or U10029 (N_10029,N_8495,N_8432);
nand U10030 (N_10030,N_9277,N_8656);
and U10031 (N_10031,N_9407,N_9491);
nor U10032 (N_10032,N_8949,N_9662);
nand U10033 (N_10033,N_8488,N_9735);
nor U10034 (N_10034,N_9920,N_8524);
nand U10035 (N_10035,N_8793,N_9674);
nor U10036 (N_10036,N_9624,N_9861);
nor U10037 (N_10037,N_9368,N_9198);
and U10038 (N_10038,N_8001,N_9502);
and U10039 (N_10039,N_8869,N_8983);
nand U10040 (N_10040,N_8463,N_8294);
and U10041 (N_10041,N_8598,N_9853);
xor U10042 (N_10042,N_9646,N_8998);
nand U10043 (N_10043,N_9577,N_9060);
nand U10044 (N_10044,N_8994,N_9697);
or U10045 (N_10045,N_9715,N_9286);
nor U10046 (N_10046,N_8823,N_9582);
nor U10047 (N_10047,N_8373,N_9018);
nand U10048 (N_10048,N_8930,N_9367);
nand U10049 (N_10049,N_8280,N_9400);
and U10050 (N_10050,N_9605,N_8686);
nand U10051 (N_10051,N_9014,N_9559);
or U10052 (N_10052,N_8728,N_9771);
xor U10053 (N_10053,N_8098,N_9097);
nor U10054 (N_10054,N_8332,N_9857);
nand U10055 (N_10055,N_9164,N_9812);
nand U10056 (N_10056,N_8670,N_8904);
or U10057 (N_10057,N_9052,N_9166);
and U10058 (N_10058,N_9704,N_8677);
xor U10059 (N_10059,N_8216,N_9999);
and U10060 (N_10060,N_9355,N_9507);
and U10061 (N_10061,N_9448,N_9158);
nand U10062 (N_10062,N_9687,N_9008);
and U10063 (N_10063,N_8249,N_8239);
nand U10064 (N_10064,N_9244,N_8040);
nand U10065 (N_10065,N_9959,N_8036);
and U10066 (N_10066,N_9783,N_9343);
or U10067 (N_10067,N_8867,N_8662);
nor U10068 (N_10068,N_8747,N_9731);
nor U10069 (N_10069,N_8194,N_8515);
or U10070 (N_10070,N_8942,N_9952);
nand U10071 (N_10071,N_9137,N_8554);
or U10072 (N_10072,N_8237,N_9557);
and U10073 (N_10073,N_8629,N_9472);
and U10074 (N_10074,N_8619,N_9677);
or U10075 (N_10075,N_9808,N_9547);
and U10076 (N_10076,N_8141,N_9456);
nor U10077 (N_10077,N_9386,N_8816);
or U10078 (N_10078,N_9645,N_8400);
nand U10079 (N_10079,N_8312,N_8228);
nand U10080 (N_10080,N_9235,N_9720);
or U10081 (N_10081,N_8282,N_9990);
nand U10082 (N_10082,N_8401,N_9772);
or U10083 (N_10083,N_8022,N_9374);
nor U10084 (N_10084,N_8729,N_8416);
or U10085 (N_10085,N_9106,N_8296);
and U10086 (N_10086,N_8876,N_8344);
or U10087 (N_10087,N_8700,N_8922);
and U10088 (N_10088,N_8882,N_9887);
nor U10089 (N_10089,N_9785,N_9561);
and U10090 (N_10090,N_9128,N_9256);
nor U10091 (N_10091,N_8852,N_9849);
xnor U10092 (N_10092,N_8081,N_9404);
and U10093 (N_10093,N_8420,N_8811);
nor U10094 (N_10094,N_8364,N_9125);
and U10095 (N_10095,N_8292,N_9370);
nand U10096 (N_10096,N_9928,N_8360);
nand U10097 (N_10097,N_9746,N_9236);
nor U10098 (N_10098,N_8353,N_9180);
and U10099 (N_10099,N_8828,N_9243);
or U10100 (N_10100,N_9459,N_9840);
or U10101 (N_10101,N_8187,N_9978);
and U10102 (N_10102,N_8633,N_9475);
and U10103 (N_10103,N_8502,N_8647);
xor U10104 (N_10104,N_8252,N_8873);
and U10105 (N_10105,N_9961,N_9776);
nor U10106 (N_10106,N_9775,N_9831);
and U10107 (N_10107,N_8185,N_9035);
nor U10108 (N_10108,N_8972,N_9834);
or U10109 (N_10109,N_8701,N_9171);
or U10110 (N_10110,N_8863,N_8366);
and U10111 (N_10111,N_9197,N_8556);
nor U10112 (N_10112,N_8361,N_9628);
nor U10113 (N_10113,N_8143,N_9129);
or U10114 (N_10114,N_8050,N_8504);
nand U10115 (N_10115,N_8798,N_9784);
and U10116 (N_10116,N_9373,N_9023);
or U10117 (N_10117,N_8134,N_8525);
nand U10118 (N_10118,N_8964,N_8256);
xor U10119 (N_10119,N_8562,N_8838);
and U10120 (N_10120,N_9460,N_8948);
nor U10121 (N_10121,N_8711,N_8663);
and U10122 (N_10122,N_9564,N_8126);
and U10123 (N_10123,N_8906,N_9929);
nor U10124 (N_10124,N_9533,N_9290);
or U10125 (N_10125,N_8130,N_8343);
and U10126 (N_10126,N_8507,N_9705);
or U10127 (N_10127,N_9017,N_9165);
nand U10128 (N_10128,N_9868,N_8981);
xor U10129 (N_10129,N_8678,N_8450);
nor U10130 (N_10130,N_8573,N_9737);
and U10131 (N_10131,N_8183,N_9316);
nor U10132 (N_10132,N_9755,N_8116);
and U10133 (N_10133,N_9609,N_8626);
nor U10134 (N_10134,N_9254,N_8648);
nor U10135 (N_10135,N_9093,N_9412);
nor U10136 (N_10136,N_8202,N_8697);
or U10137 (N_10137,N_9769,N_8231);
and U10138 (N_10138,N_8108,N_9401);
nand U10139 (N_10139,N_8024,N_8063);
nor U10140 (N_10140,N_8466,N_8902);
nand U10141 (N_10141,N_9021,N_9631);
xnor U10142 (N_10142,N_9736,N_9930);
and U10143 (N_10143,N_9132,N_8821);
and U10144 (N_10144,N_8530,N_9001);
and U10145 (N_10145,N_9923,N_9711);
nand U10146 (N_10146,N_9391,N_9214);
nor U10147 (N_10147,N_8579,N_8424);
nor U10148 (N_10148,N_8848,N_8542);
nand U10149 (N_10149,N_8275,N_8272);
and U10150 (N_10150,N_9151,N_8792);
nand U10151 (N_10151,N_9947,N_8164);
xnor U10152 (N_10152,N_8897,N_9160);
nor U10153 (N_10153,N_9529,N_9543);
and U10154 (N_10154,N_9268,N_9416);
nand U10155 (N_10155,N_8068,N_9875);
nand U10156 (N_10156,N_9219,N_8969);
or U10157 (N_10157,N_8498,N_8399);
and U10158 (N_10158,N_8988,N_9780);
or U10159 (N_10159,N_9242,N_9377);
and U10160 (N_10160,N_8430,N_8672);
nor U10161 (N_10161,N_9925,N_9420);
nor U10162 (N_10162,N_8406,N_8449);
nand U10163 (N_10163,N_9234,N_9292);
or U10164 (N_10164,N_9602,N_9758);
nor U10165 (N_10165,N_9104,N_9415);
and U10166 (N_10166,N_8710,N_9541);
and U10167 (N_10167,N_8529,N_8370);
nand U10168 (N_10168,N_9912,N_9402);
or U10169 (N_10169,N_9464,N_9588);
nor U10170 (N_10170,N_8889,N_8995);
nand U10171 (N_10171,N_9392,N_9349);
or U10172 (N_10172,N_9346,N_8713);
xnor U10173 (N_10173,N_9492,N_9647);
nand U10174 (N_10174,N_9095,N_8467);
nor U10175 (N_10175,N_8115,N_9212);
nor U10176 (N_10176,N_8924,N_8225);
or U10177 (N_10177,N_9802,N_8382);
nand U10178 (N_10178,N_9625,N_9987);
nand U10179 (N_10179,N_8625,N_8864);
nor U10180 (N_10180,N_8060,N_9520);
and U10181 (N_10181,N_9438,N_9080);
nand U10182 (N_10182,N_8699,N_8552);
or U10183 (N_10183,N_8393,N_9157);
and U10184 (N_10184,N_9059,N_8991);
and U10185 (N_10185,N_8993,N_9922);
nor U10186 (N_10186,N_8703,N_8085);
nor U10187 (N_10187,N_8099,N_9584);
nor U10188 (N_10188,N_9297,N_9632);
nand U10189 (N_10189,N_8576,N_8680);
nor U10190 (N_10190,N_9227,N_8451);
nor U10191 (N_10191,N_8348,N_8434);
nand U10192 (N_10192,N_8764,N_9682);
or U10193 (N_10193,N_8762,N_9729);
and U10194 (N_10194,N_9908,N_8574);
nor U10195 (N_10195,N_8203,N_9535);
nand U10196 (N_10196,N_8169,N_9919);
or U10197 (N_10197,N_8522,N_9381);
nor U10198 (N_10198,N_8155,N_9838);
nand U10199 (N_10199,N_9960,N_9237);
nor U10200 (N_10200,N_8860,N_8455);
and U10201 (N_10201,N_9911,N_9989);
and U10202 (N_10202,N_8646,N_9067);
nand U10203 (N_10203,N_9465,N_9867);
or U10204 (N_10204,N_9707,N_8217);
and U10205 (N_10205,N_8073,N_8137);
or U10206 (N_10206,N_9612,N_9686);
nand U10207 (N_10207,N_9578,N_8814);
nand U10208 (N_10208,N_9556,N_8738);
nand U10209 (N_10209,N_9114,N_8956);
nand U10210 (N_10210,N_8242,N_8170);
or U10211 (N_10211,N_8271,N_8679);
nor U10212 (N_10212,N_8114,N_9889);
or U10213 (N_10213,N_9532,N_9082);
nor U10214 (N_10214,N_9016,N_8059);
and U10215 (N_10215,N_9692,N_9664);
nand U10216 (N_10216,N_8962,N_8362);
xnor U10217 (N_10217,N_9430,N_8311);
or U10218 (N_10218,N_8874,N_8381);
or U10219 (N_10219,N_8966,N_9096);
and U10220 (N_10220,N_8011,N_9045);
nor U10221 (N_10221,N_8611,N_8335);
or U10222 (N_10222,N_9659,N_8853);
or U10223 (N_10223,N_9604,N_8499);
nor U10224 (N_10224,N_9192,N_8349);
nand U10225 (N_10225,N_9905,N_9115);
or U10226 (N_10226,N_8568,N_9225);
or U10227 (N_10227,N_9006,N_9074);
nor U10228 (N_10228,N_8308,N_8384);
nor U10229 (N_10229,N_8019,N_8148);
and U10230 (N_10230,N_8501,N_8145);
nand U10231 (N_10231,N_9029,N_9918);
or U10232 (N_10232,N_9065,N_8965);
and U10233 (N_10233,N_8342,N_8591);
nor U10234 (N_10234,N_8487,N_8482);
or U10235 (N_10235,N_8291,N_8281);
nor U10236 (N_10236,N_9068,N_9708);
or U10237 (N_10237,N_8039,N_9757);
nor U10238 (N_10238,N_8152,N_8365);
nor U10239 (N_10239,N_8743,N_8305);
nand U10240 (N_10240,N_8290,N_8627);
nor U10241 (N_10241,N_8772,N_8493);
nand U10242 (N_10242,N_9866,N_9331);
nor U10243 (N_10243,N_8605,N_8946);
and U10244 (N_10244,N_9871,N_9289);
or U10245 (N_10245,N_9336,N_9305);
xor U10246 (N_10246,N_8199,N_8383);
nor U10247 (N_10247,N_8508,N_8074);
or U10248 (N_10248,N_9426,N_8794);
and U10249 (N_10249,N_8724,N_8535);
nor U10250 (N_10250,N_8620,N_8894);
or U10251 (N_10251,N_9550,N_8636);
nand U10252 (N_10252,N_8947,N_8248);
and U10253 (N_10253,N_8016,N_9260);
nor U10254 (N_10254,N_9716,N_9449);
and U10255 (N_10255,N_9741,N_8125);
nor U10256 (N_10256,N_9501,N_8954);
nor U10257 (N_10257,N_8140,N_9015);
or U10258 (N_10258,N_9497,N_8389);
and U10259 (N_10259,N_9865,N_9850);
or U10260 (N_10260,N_8767,N_9806);
nand U10261 (N_10261,N_8209,N_9820);
or U10262 (N_10262,N_9253,N_9897);
and U10263 (N_10263,N_9347,N_8425);
nand U10264 (N_10264,N_9187,N_9754);
nand U10265 (N_10265,N_9226,N_8223);
nand U10266 (N_10266,N_9496,N_8634);
and U10267 (N_10267,N_8566,N_9725);
and U10268 (N_10268,N_9051,N_9098);
nand U10269 (N_10269,N_9215,N_8083);
or U10270 (N_10270,N_8232,N_9603);
and U10271 (N_10271,N_8410,N_9092);
or U10272 (N_10272,N_8111,N_8048);
nand U10273 (N_10273,N_9993,N_9724);
nor U10274 (N_10274,N_8787,N_9299);
or U10275 (N_10275,N_9648,N_8950);
nor U10276 (N_10276,N_8505,N_9087);
xnor U10277 (N_10277,N_9940,N_8774);
or U10278 (N_10278,N_8053,N_9486);
nor U10279 (N_10279,N_9750,N_9474);
or U10280 (N_10280,N_9935,N_8684);
and U10281 (N_10281,N_9406,N_8409);
or U10282 (N_10282,N_8269,N_8624);
or U10283 (N_10283,N_8241,N_9701);
and U10284 (N_10284,N_8959,N_8915);
nand U10285 (N_10285,N_8491,N_8328);
or U10286 (N_10286,N_8741,N_8892);
nor U10287 (N_10287,N_9123,N_8698);
nand U10288 (N_10288,N_9970,N_9789);
or U10289 (N_10289,N_9342,N_8696);
xor U10290 (N_10290,N_9778,N_9764);
and U10291 (N_10291,N_9027,N_9567);
and U10292 (N_10292,N_9135,N_9079);
or U10293 (N_10293,N_9530,N_8303);
nor U10294 (N_10294,N_9283,N_9207);
or U10295 (N_10295,N_8154,N_8888);
or U10296 (N_10296,N_9505,N_8928);
nor U10297 (N_10297,N_8157,N_9032);
and U10298 (N_10298,N_9512,N_8551);
or U10299 (N_10299,N_8431,N_8105);
nor U10300 (N_10300,N_9781,N_9419);
nand U10301 (N_10301,N_8037,N_9688);
nand U10302 (N_10302,N_9360,N_8803);
or U10303 (N_10303,N_9804,N_9022);
or U10304 (N_10304,N_8144,N_8188);
nand U10305 (N_10305,N_8555,N_8771);
or U10306 (N_10306,N_9914,N_9836);
and U10307 (N_10307,N_8990,N_8388);
xor U10308 (N_10308,N_8931,N_8132);
nand U10309 (N_10309,N_9937,N_9179);
and U10310 (N_10310,N_9955,N_8458);
and U10311 (N_10311,N_9440,N_8604);
and U10312 (N_10312,N_8926,N_8259);
or U10313 (N_10313,N_8309,N_8200);
or U10314 (N_10314,N_8492,N_9359);
nor U10315 (N_10315,N_8795,N_8716);
nand U10316 (N_10316,N_8034,N_8087);
or U10317 (N_10317,N_8590,N_9152);
and U10318 (N_10318,N_8363,N_8230);
or U10319 (N_10319,N_9830,N_9493);
nand U10320 (N_10320,N_8751,N_8086);
nor U10321 (N_10321,N_8748,N_9884);
nor U10322 (N_10322,N_8671,N_9159);
or U10323 (N_10323,N_9186,N_8320);
or U10324 (N_10324,N_8843,N_9852);
or U10325 (N_10325,N_9037,N_8667);
nand U10326 (N_10326,N_8856,N_9994);
and U10327 (N_10327,N_8921,N_8235);
or U10328 (N_10328,N_9761,N_8005);
or U10329 (N_10329,N_9118,N_9172);
nor U10330 (N_10330,N_9432,N_9250);
and U10331 (N_10331,N_9281,N_9364);
and U10332 (N_10332,N_9767,N_9835);
nor U10333 (N_10333,N_8023,N_9458);
nor U10334 (N_10334,N_8456,N_9821);
nand U10335 (N_10335,N_8740,N_8031);
or U10336 (N_10336,N_9976,N_8189);
xnor U10337 (N_10337,N_8621,N_9385);
nor U10338 (N_10338,N_8462,N_9534);
nand U10339 (N_10339,N_8323,N_9307);
nor U10340 (N_10340,N_9615,N_8445);
nand U10341 (N_10341,N_9596,N_9770);
or U10342 (N_10342,N_8355,N_8368);
xor U10343 (N_10343,N_9061,N_9817);
and U10344 (N_10344,N_9069,N_9539);
or U10345 (N_10345,N_9702,N_9142);
and U10346 (N_10346,N_9880,N_9468);
nor U10347 (N_10347,N_9977,N_8347);
nand U10348 (N_10348,N_9969,N_9521);
or U10349 (N_10349,N_9362,N_8175);
nand U10350 (N_10350,N_8635,N_8734);
nor U10351 (N_10351,N_9954,N_8092);
nand U10352 (N_10352,N_9201,N_8687);
nand U10353 (N_10353,N_8958,N_8129);
xnor U10354 (N_10354,N_8661,N_8267);
xor U10355 (N_10355,N_9278,N_9803);
nand U10356 (N_10356,N_8655,N_8206);
or U10357 (N_10357,N_8637,N_9427);
nand U10358 (N_10358,N_8061,N_9902);
nand U10359 (N_10359,N_8405,N_9066);
nand U10360 (N_10360,N_8056,N_9109);
nand U10361 (N_10361,N_8118,N_8996);
nor U10362 (N_10362,N_8939,N_8791);
and U10363 (N_10363,N_8396,N_9816);
or U10364 (N_10364,N_9848,N_8136);
nor U10365 (N_10365,N_8788,N_9141);
nor U10366 (N_10366,N_9369,N_9100);
nor U10367 (N_10367,N_8089,N_8978);
and U10368 (N_10368,N_8166,N_8221);
nor U10369 (N_10369,N_8868,N_9700);
and U10370 (N_10370,N_9085,N_9621);
or U10371 (N_10371,N_9222,N_8520);
xor U10372 (N_10372,N_9590,N_9218);
nand U10373 (N_10373,N_9103,N_9088);
nand U10374 (N_10374,N_9311,N_9463);
nand U10375 (N_10375,N_9575,N_8193);
nor U10376 (N_10376,N_8330,N_8407);
and U10377 (N_10377,N_8763,N_8984);
or U10378 (N_10378,N_9284,N_9062);
nand U10379 (N_10379,N_8883,N_9586);
and U10380 (N_10380,N_9428,N_8142);
or U10381 (N_10381,N_8057,N_8801);
nand U10382 (N_10382,N_8338,N_9058);
or U10383 (N_10383,N_9689,N_9293);
xor U10384 (N_10384,N_8553,N_8881);
or U10385 (N_10385,N_9513,N_8970);
nand U10386 (N_10386,N_9594,N_9665);
and U10387 (N_10387,N_9760,N_8506);
nor U10388 (N_10388,N_9444,N_8916);
and U10389 (N_10389,N_9148,N_8614);
nand U10390 (N_10390,N_8538,N_9344);
and U10391 (N_10391,N_8742,N_9352);
nand U10392 (N_10392,N_9655,N_9693);
nand U10393 (N_10393,N_8238,N_9607);
nor U10394 (N_10394,N_9053,N_9083);
or U10395 (N_10395,N_8618,N_9042);
nand U10396 (N_10396,N_8264,N_9147);
nand U10397 (N_10397,N_8616,N_9791);
and U10398 (N_10398,N_8293,N_8133);
nand U10399 (N_10399,N_9601,N_8923);
nor U10400 (N_10400,N_8444,N_9699);
and U10401 (N_10401,N_9894,N_8885);
nor U10402 (N_10402,N_8101,N_9685);
nand U10403 (N_10403,N_8219,N_9562);
or U10404 (N_10404,N_9348,N_8460);
or U10405 (N_10405,N_9819,N_9451);
xor U10406 (N_10406,N_9231,N_8952);
or U10407 (N_10407,N_8503,N_8375);
nand U10408 (N_10408,N_8844,N_9202);
nor U10409 (N_10409,N_8029,N_8051);
nor U10410 (N_10410,N_8197,N_9863);
nor U10411 (N_10411,N_8736,N_8841);
nor U10412 (N_10412,N_8987,N_9879);
nand U10413 (N_10413,N_8107,N_8879);
nand U10414 (N_10414,N_9025,N_9309);
nand U10415 (N_10415,N_8766,N_8727);
or U10416 (N_10416,N_9571,N_8198);
nand U10417 (N_10417,N_8875,N_9728);
nor U10418 (N_10418,N_9313,N_8975);
and U10419 (N_10419,N_8599,N_8397);
or U10420 (N_10420,N_8543,N_9120);
xnor U10421 (N_10421,N_8173,N_8484);
and U10422 (N_10422,N_8770,N_9043);
nor U10423 (N_10423,N_8784,N_9548);
nand U10424 (N_10424,N_8827,N_9744);
or U10425 (N_10425,N_9936,N_8761);
or U10426 (N_10426,N_9657,N_8279);
and U10427 (N_10427,N_8999,N_8893);
nor U10428 (N_10428,N_8289,N_9613);
and U10429 (N_10429,N_9900,N_8643);
nand U10430 (N_10430,N_8427,N_8807);
nor U10431 (N_10431,N_9633,N_9992);
and U10432 (N_10432,N_8124,N_9136);
nor U10433 (N_10433,N_9240,N_9962);
or U10434 (N_10434,N_9579,N_9924);
nand U10435 (N_10435,N_8372,N_8842);
or U10436 (N_10436,N_9298,N_8376);
nand U10437 (N_10437,N_8707,N_8944);
nor U10438 (N_10438,N_8333,N_8009);
nor U10439 (N_10439,N_9050,N_9393);
or U10440 (N_10440,N_8865,N_8768);
xor U10441 (N_10441,N_8443,N_9494);
or U10442 (N_10442,N_9262,N_8652);
nor U10443 (N_10443,N_8536,N_8013);
or U10444 (N_10444,N_8840,N_8390);
or U10445 (N_10445,N_9623,N_8480);
and U10446 (N_10446,N_8709,N_9113);
nand U10447 (N_10447,N_9047,N_8000);
and U10448 (N_10448,N_9443,N_9239);
or U10449 (N_10449,N_8395,N_8908);
xor U10450 (N_10450,N_8069,N_8226);
or U10451 (N_10451,N_9445,N_8288);
and U10452 (N_10452,N_8120,N_9569);
and U10453 (N_10453,N_9126,N_8064);
or U10454 (N_10454,N_9241,N_8644);
nand U10455 (N_10455,N_8300,N_8117);
or U10456 (N_10456,N_8090,N_8632);
or U10457 (N_10457,N_9753,N_9358);
or U10458 (N_10458,N_9739,N_9985);
nand U10459 (N_10459,N_9980,N_9714);
and U10460 (N_10460,N_8464,N_9300);
nor U10461 (N_10461,N_9335,N_8184);
nand U10462 (N_10462,N_9599,N_9078);
or U10463 (N_10463,N_9673,N_8918);
and U10464 (N_10464,N_9200,N_9542);
nand U10465 (N_10465,N_8112,N_8314);
or U10466 (N_10466,N_8474,N_8191);
nand U10467 (N_10467,N_9382,N_8822);
or U10468 (N_10468,N_9629,N_8527);
nor U10469 (N_10469,N_8640,N_8457);
nand U10470 (N_10470,N_9503,N_8007);
or U10471 (N_10471,N_9933,N_8150);
nand U10472 (N_10472,N_9943,N_9127);
or U10473 (N_10473,N_9824,N_8419);
and U10474 (N_10474,N_8705,N_9473);
xnor U10475 (N_10475,N_9916,N_8018);
nand U10476 (N_10476,N_8909,N_9856);
or U10477 (N_10477,N_9324,N_9794);
nor U10478 (N_10478,N_9941,N_9630);
nand U10479 (N_10479,N_9002,N_9896);
and U10480 (N_10480,N_9323,N_8567);
nor U10481 (N_10481,N_9228,N_8891);
and U10482 (N_10482,N_9433,N_9030);
and U10483 (N_10483,N_8413,N_8517);
nor U10484 (N_10484,N_9696,N_8895);
and U10485 (N_10485,N_8673,N_8945);
and U10486 (N_10486,N_8593,N_9636);
xnor U10487 (N_10487,N_9094,N_8452);
or U10488 (N_10488,N_8247,N_8977);
nor U10489 (N_10489,N_9651,N_9585);
or U10490 (N_10490,N_9013,N_8479);
nand U10491 (N_10491,N_9188,N_8378);
nor U10492 (N_10492,N_8391,N_9191);
and U10493 (N_10493,N_8418,N_8104);
nand U10494 (N_10494,N_8569,N_8829);
and U10495 (N_10495,N_9679,N_9796);
nor U10496 (N_10496,N_8675,N_9447);
and U10497 (N_10497,N_9545,N_8210);
nand U10498 (N_10498,N_8799,N_9055);
or U10499 (N_10499,N_8352,N_9885);
or U10500 (N_10500,N_9927,N_8417);
nor U10501 (N_10501,N_9275,N_9026);
nand U10502 (N_10502,N_9611,N_8319);
nand U10503 (N_10503,N_8236,N_9351);
nor U10504 (N_10504,N_8354,N_8337);
nor U10505 (N_10505,N_9435,N_9627);
or U10506 (N_10506,N_8890,N_8317);
nor U10507 (N_10507,N_9518,N_8973);
nor U10508 (N_10508,N_8564,N_9938);
and U10509 (N_10509,N_9175,N_8777);
nor U10510 (N_10510,N_8730,N_9071);
and U10511 (N_10511,N_9617,N_9409);
or U10512 (N_10512,N_8980,N_9675);
nor U10513 (N_10513,N_9301,N_8030);
or U10514 (N_10514,N_8244,N_9827);
or U10515 (N_10515,N_8429,N_8327);
nand U10516 (N_10516,N_9797,N_9765);
nand U10517 (N_10517,N_8428,N_8100);
or U10518 (N_10518,N_8693,N_9442);
nor U10519 (N_10519,N_9048,N_8476);
nand U10520 (N_10520,N_8358,N_8521);
and U10521 (N_10521,N_9818,N_8298);
and U10522 (N_10522,N_8180,N_8558);
nand U10523 (N_10523,N_9888,N_9964);
nor U10524 (N_10524,N_8528,N_8859);
and U10525 (N_10525,N_9455,N_8717);
or U10526 (N_10526,N_9517,N_8113);
nor U10527 (N_10527,N_8442,N_8218);
nand U10528 (N_10528,N_8128,N_9102);
and U10529 (N_10529,N_8559,N_9552);
nand U10530 (N_10530,N_9295,N_9873);
nand U10531 (N_10531,N_9410,N_8369);
and U10532 (N_10532,N_8072,N_8321);
nor U10533 (N_10533,N_8855,N_9495);
and U10534 (N_10534,N_8695,N_8654);
or U10535 (N_10535,N_8886,N_8544);
nand U10536 (N_10536,N_9271,N_9898);
or U10537 (N_10537,N_9882,N_9121);
xor U10538 (N_10538,N_8570,N_9005);
or U10539 (N_10539,N_8276,N_8179);
nand U10540 (N_10540,N_9595,N_8547);
nand U10541 (N_10541,N_8645,N_8387);
nor U10542 (N_10542,N_8454,N_8028);
nor U10543 (N_10543,N_9671,N_9858);
nor U10544 (N_10544,N_8986,N_9205);
nand U10545 (N_10545,N_8953,N_9967);
or U10546 (N_10546,N_8940,N_8817);
nor U10547 (N_10547,N_9163,N_9658);
nand U10548 (N_10548,N_9553,N_8537);
nor U10549 (N_10549,N_9668,N_8602);
nor U10550 (N_10550,N_8694,N_9049);
nor U10551 (N_10551,N_8653,N_9425);
nor U10552 (N_10552,N_9527,N_8182);
or U10553 (N_10553,N_8765,N_8082);
nand U10554 (N_10554,N_8613,N_8531);
nand U10555 (N_10555,N_8224,N_9656);
or U10556 (N_10556,N_9653,N_8796);
and U10557 (N_10557,N_8834,N_8273);
nand U10558 (N_10558,N_8664,N_8651);
nand U10559 (N_10559,N_8212,N_9161);
xor U10560 (N_10560,N_9810,N_8749);
nor U10561 (N_10561,N_8565,N_9498);
and U10562 (N_10562,N_8516,N_8932);
nor U10563 (N_10563,N_8837,N_9551);
nand U10564 (N_10564,N_8512,N_8339);
nand U10565 (N_10565,N_8380,N_8167);
nor U10566 (N_10566,N_9457,N_9538);
xnor U10567 (N_10567,N_8609,N_9471);
nor U10568 (N_10568,N_8872,N_9904);
nor U10569 (N_10569,N_8571,N_8211);
nand U10570 (N_10570,N_9768,N_9398);
or U10571 (N_10571,N_8386,N_9860);
nor U10572 (N_10572,N_9745,N_8093);
or U10573 (N_10573,N_8340,N_9046);
and U10574 (N_10574,N_8781,N_9968);
xnor U10575 (N_10575,N_9608,N_8047);
and U10576 (N_10576,N_9318,N_8465);
and U10577 (N_10577,N_9007,N_8638);
nor U10578 (N_10578,N_8982,N_9216);
nor U10579 (N_10579,N_8153,N_9269);
or U10580 (N_10580,N_8403,N_8744);
nor U10581 (N_10581,N_8017,N_9146);
and U10582 (N_10582,N_9294,N_9851);
or U10583 (N_10583,N_9469,N_9470);
and U10584 (N_10584,N_9031,N_8316);
or U10585 (N_10585,N_8159,N_8268);
nor U10586 (N_10586,N_8733,N_8681);
nor U10587 (N_10587,N_9334,N_9365);
nor U10588 (N_10588,N_9876,N_9110);
nand U10589 (N_10589,N_9957,N_8753);
or U10590 (N_10590,N_9384,N_9354);
nand U10591 (N_10591,N_8639,N_8049);
or U10592 (N_10592,N_8746,N_9638);
and U10593 (N_10593,N_8446,N_8610);
nor U10594 (N_10594,N_8192,N_8607);
nand U10595 (N_10595,N_9826,N_8877);
or U10596 (N_10596,N_8127,N_8162);
nor U10597 (N_10597,N_9777,N_8577);
nand U10598 (N_10598,N_9972,N_8597);
or U10599 (N_10599,N_9718,N_9572);
nor U10600 (N_10600,N_9461,N_8315);
and U10601 (N_10601,N_9454,N_8204);
nor U10602 (N_10602,N_9650,N_9610);
nand U10603 (N_10603,N_8665,N_9555);
nand U10604 (N_10604,N_9759,N_8437);
nand U10605 (N_10605,N_8884,N_9546);
nand U10606 (N_10606,N_9945,N_9963);
and U10607 (N_10607,N_8481,N_9883);
nand U10608 (N_10608,N_9874,N_8010);
or U10609 (N_10609,N_9913,N_8336);
nor U10610 (N_10610,N_9644,N_9549);
or U10611 (N_10611,N_8588,N_9149);
nand U10612 (N_10612,N_8250,N_8812);
nand U10613 (N_10613,N_8139,N_8097);
nand U10614 (N_10614,N_8176,N_8096);
nor U10615 (N_10615,N_8968,N_8158);
or U10616 (N_10616,N_9832,N_9296);
or U10617 (N_10617,N_9798,N_8666);
and U10618 (N_10618,N_8900,N_9841);
nor U10619 (N_10619,N_8755,N_9847);
nor U10620 (N_10620,N_8657,N_9439);
nor U10621 (N_10621,N_9907,N_8682);
and U10622 (N_10622,N_9703,N_9249);
or U10623 (N_10623,N_8600,N_8606);
nand U10624 (N_10624,N_9452,N_8265);
nor U10625 (N_10625,N_9380,N_8234);
nor U10626 (N_10626,N_9910,N_9133);
nor U10627 (N_10627,N_8163,N_8270);
and U10628 (N_10628,N_8808,N_8692);
nand U10629 (N_10629,N_8195,N_8447);
nor U10630 (N_10630,N_9733,N_8612);
or U10631 (N_10631,N_9116,N_9956);
and U10632 (N_10632,N_8523,N_9075);
nor U10633 (N_10633,N_9862,N_8177);
nand U10634 (N_10634,N_9482,N_9054);
and U10635 (N_10635,N_9009,N_8002);
or U10636 (N_10636,N_8122,N_9680);
nand U10637 (N_10637,N_8341,N_9583);
nand U10638 (N_10638,N_8732,N_8519);
and U10639 (N_10639,N_8832,N_8898);
or U10640 (N_10640,N_8899,N_9799);
nand U10641 (N_10641,N_9932,N_8584);
or U10642 (N_10642,N_9811,N_8110);
nand U10643 (N_10643,N_9844,N_9403);
or U10644 (N_10644,N_9337,N_9070);
nand U10645 (N_10645,N_8769,N_9667);
nor U10646 (N_10646,N_8750,N_8790);
nand U10647 (N_10647,N_8423,N_8258);
and U10648 (N_10648,N_9773,N_8783);
nand U10649 (N_10649,N_9183,N_9353);
nor U10650 (N_10650,N_8813,N_9580);
nand U10651 (N_10651,N_8802,N_9516);
nor U10652 (N_10652,N_9229,N_9322);
nand U10653 (N_10653,N_9266,N_8820);
nand U10654 (N_10654,N_9641,N_9308);
nor U10655 (N_10655,N_9795,N_9248);
xnor U10656 (N_10656,N_9245,N_8026);
nand U10657 (N_10657,N_9762,N_9467);
and U10658 (N_10658,N_9376,N_9722);
nor U10659 (N_10659,N_9039,N_8261);
nor U10660 (N_10660,N_9314,N_8147);
nor U10661 (N_10661,N_9814,N_8421);
nand U10662 (N_10662,N_8911,N_9522);
and U10663 (N_10663,N_9639,N_9328);
nand U10664 (N_10664,N_8622,N_9652);
and U10665 (N_10665,N_8534,N_8367);
and U10666 (N_10666,N_8985,N_9828);
and U10667 (N_10667,N_8961,N_8545);
nor U10668 (N_10668,N_8160,N_8469);
nand U10669 (N_10669,N_8285,N_9174);
nand U10670 (N_10670,N_8779,N_9330);
and U10671 (N_10671,N_8941,N_8151);
and U10672 (N_10672,N_9338,N_9787);
nor U10673 (N_10673,N_8785,N_9131);
xnor U10674 (N_10674,N_8394,N_9105);
and U10675 (N_10675,N_8402,N_8913);
and U10676 (N_10676,N_8887,N_8773);
and U10677 (N_10677,N_9063,N_8937);
nor U10678 (N_10678,N_8222,N_8581);
or U10679 (N_10679,N_9740,N_8255);
or U10680 (N_10680,N_8065,N_8326);
nor U10681 (N_10681,N_9726,N_8229);
or U10682 (N_10682,N_9181,N_9949);
or U10683 (N_10683,N_9279,N_8871);
or U10684 (N_10684,N_9221,N_8572);
and U10685 (N_10685,N_8850,N_9944);
or U10686 (N_10686,N_8436,N_8412);
and U10687 (N_10687,N_8857,N_9825);
nor U10688 (N_10688,N_8470,N_8156);
and U10689 (N_10689,N_8052,N_8483);
or U10690 (N_10690,N_9434,N_9592);
nand U10691 (N_10691,N_8123,N_9917);
or U10692 (N_10692,N_8782,N_8833);
or U10693 (N_10693,N_9723,N_9626);
or U10694 (N_10694,N_9361,N_9984);
nor U10695 (N_10695,N_8201,N_9683);
nor U10696 (N_10696,N_9012,N_9500);
or U10697 (N_10697,N_9040,N_9350);
nand U10698 (N_10698,N_9939,N_8933);
nand U10699 (N_10699,N_8215,N_8062);
or U10700 (N_10700,N_9620,N_8518);
and U10701 (N_10701,N_8561,N_8408);
nor U10702 (N_10702,N_9122,N_9204);
nor U10703 (N_10703,N_8712,N_9000);
nand U10704 (N_10704,N_8778,N_9134);
nor U10705 (N_10705,N_8485,N_8735);
or U10706 (N_10706,N_9356,N_9663);
or U10707 (N_10707,N_8205,N_8976);
and U10708 (N_10708,N_9203,N_8533);
and U10709 (N_10709,N_8955,N_9606);
and U10710 (N_10710,N_8815,N_9366);
or U10711 (N_10711,N_9089,N_9233);
nor U10712 (N_10712,N_9388,N_8758);
nor U10713 (N_10713,N_8731,N_8278);
and U10714 (N_10714,N_8989,N_9975);
nand U10715 (N_10715,N_8960,N_9966);
nand U10716 (N_10716,N_9156,N_8274);
nor U10717 (N_10717,N_9394,N_9786);
and U10718 (N_10718,N_9666,N_9558);
and U10719 (N_10719,N_9508,N_9144);
nor U10720 (N_10720,N_9568,N_9525);
or U10721 (N_10721,N_8477,N_8441);
nand U10722 (N_10722,N_9267,N_9411);
nand U10723 (N_10723,N_9073,N_8071);
and U10724 (N_10724,N_8557,N_8027);
nand U10725 (N_10725,N_8539,N_9996);
and U10726 (N_10726,N_8084,N_9223);
and U10727 (N_10727,N_9719,N_9375);
and U10728 (N_10728,N_9807,N_8379);
nand U10729 (N_10729,N_8033,N_9423);
and U10730 (N_10730,N_8331,N_8161);
nand U10731 (N_10731,N_9036,N_9934);
and U10732 (N_10732,N_8689,N_9640);
and U10733 (N_10733,N_8582,N_9064);
or U10734 (N_10734,N_9024,N_8896);
or U10735 (N_10735,N_9263,N_9397);
nor U10736 (N_10736,N_9357,N_8297);
nor U10737 (N_10737,N_9217,N_9090);
nor U10738 (N_10738,N_8439,N_8251);
nor U10739 (N_10739,N_9869,N_9843);
nand U10740 (N_10740,N_8045,N_9511);
nor U10741 (N_10741,N_9694,N_8020);
and U10742 (N_10742,N_9143,N_9833);
or U10743 (N_10743,N_8078,N_8307);
nor U10744 (N_10744,N_8284,N_9635);
or U10745 (N_10745,N_8720,N_8854);
nor U10746 (N_10746,N_8905,N_8603);
xnor U10747 (N_10747,N_9589,N_8934);
nor U10748 (N_10748,N_8220,N_9890);
nor U10749 (N_10749,N_8979,N_9209);
nand U10750 (N_10750,N_9111,N_9418);
nand U10751 (N_10751,N_8912,N_8608);
and U10752 (N_10752,N_9119,N_8471);
or U10753 (N_10753,N_8514,N_8690);
or U10754 (N_10754,N_8149,N_9878);
nor U10755 (N_10755,N_8650,N_9854);
nand U10756 (N_10756,N_9921,N_8146);
or U10757 (N_10757,N_9782,N_8943);
nand U10758 (N_10758,N_9280,N_9565);
nor U10759 (N_10759,N_9845,N_9846);
or U10760 (N_10760,N_9951,N_8723);
or U10761 (N_10761,N_8254,N_8350);
nand U10762 (N_10762,N_9195,N_9056);
or U10763 (N_10763,N_8415,N_9734);
and U10764 (N_10764,N_8486,N_9091);
or U10765 (N_10765,N_9983,N_9598);
nor U10766 (N_10766,N_9084,N_9805);
or U10767 (N_10767,N_8546,N_9891);
and U10768 (N_10768,N_8243,N_8810);
nand U10769 (N_10769,N_9252,N_9020);
and U10770 (N_10770,N_9554,N_8266);
nand U10771 (N_10771,N_8722,N_8468);
nand U10772 (N_10772,N_8004,N_9751);
nor U10773 (N_10773,N_8702,N_9340);
nand U10774 (N_10774,N_8595,N_8575);
or U10775 (N_10775,N_8714,N_8997);
and U10776 (N_10776,N_8540,N_9870);
or U10777 (N_10777,N_9706,N_8668);
and U10778 (N_10778,N_8718,N_9238);
nand U10779 (N_10779,N_8497,N_8715);
and U10780 (N_10780,N_8076,N_9877);
nor U10781 (N_10781,N_8325,N_9193);
and U10782 (N_10782,N_9270,N_8398);
nand U10783 (N_10783,N_9117,N_9421);
or U10784 (N_10784,N_9872,N_9752);
nor U10785 (N_10785,N_8165,N_9788);
or U10786 (N_10786,N_9979,N_8870);
and U10787 (N_10787,N_9414,N_8257);
nor U10788 (N_10788,N_8726,N_9698);
and U10789 (N_10789,N_9339,N_9600);
or U10790 (N_10790,N_8752,N_9199);
nor U10791 (N_10791,N_9748,N_9864);
nand U10792 (N_10792,N_9540,N_9971);
and U10793 (N_10793,N_9466,N_9177);
and U10794 (N_10794,N_9713,N_8706);
nand U10795 (N_10795,N_8172,N_8131);
and U10796 (N_10796,N_9072,N_9948);
nand U10797 (N_10797,N_8262,N_9057);
and U10798 (N_10798,N_8207,N_8008);
nand U10799 (N_10799,N_9478,N_8038);
or U10800 (N_10800,N_9823,N_8587);
nand U10801 (N_10801,N_8845,N_8938);
and U10802 (N_10802,N_8910,N_9642);
or U10803 (N_10803,N_8641,N_9643);
nand U10804 (N_10804,N_9998,N_9429);
or U10805 (N_10805,N_9901,N_9779);
nand U10806 (N_10806,N_8756,N_8171);
and U10807 (N_10807,N_9622,N_8704);
xor U10808 (N_10808,N_8310,N_8095);
and U10809 (N_10809,N_9184,N_8659);
and U10810 (N_10810,N_9315,N_9034);
xnor U10811 (N_10811,N_9325,N_8601);
nand U10812 (N_10812,N_8260,N_9946);
nor U10813 (N_10813,N_9437,N_9506);
and U10814 (N_10814,N_9649,N_9413);
and U10815 (N_10815,N_9892,N_9259);
nor U10816 (N_10816,N_8676,N_8835);
and U10817 (N_10817,N_8371,N_9173);
xor U10818 (N_10818,N_9661,N_9637);
nand U10819 (N_10819,N_8776,N_9154);
nor U10820 (N_10820,N_9678,N_8914);
and U10821 (N_10821,N_8334,N_9855);
nor U10822 (N_10822,N_9101,N_9581);
xor U10823 (N_10823,N_8780,N_9742);
nand U10824 (N_10824,N_9004,N_8472);
and U10825 (N_10825,N_8119,N_9790);
and U10826 (N_10826,N_9801,N_9974);
and U10827 (N_10827,N_8578,N_9378);
and U10828 (N_10828,N_8549,N_8674);
nand U10829 (N_10829,N_9973,N_8649);
nor U10830 (N_10830,N_8974,N_8277);
nor U10831 (N_10831,N_8496,N_9395);
nor U10832 (N_10832,N_9185,N_9614);
or U10833 (N_10833,N_8560,N_9206);
nor U10834 (N_10834,N_8903,N_9302);
or U10835 (N_10835,N_8935,N_8426);
and U10836 (N_10836,N_8846,N_9766);
or U10837 (N_10837,N_9654,N_9926);
or U10838 (N_10838,N_9189,N_9519);
xor U10839 (N_10839,N_9446,N_9387);
or U10840 (N_10840,N_8630,N_9514);
or U10841 (N_10841,N_9196,N_9792);
nand U10842 (N_10842,N_9390,N_8615);
nand U10843 (N_10843,N_8302,N_8032);
nor U10844 (N_10844,N_9566,N_9893);
nor U10845 (N_10845,N_9405,N_8596);
nand U10846 (N_10846,N_8628,N_8847);
and U10847 (N_10847,N_8377,N_8929);
xnor U10848 (N_10848,N_8858,N_8826);
or U10849 (N_10849,N_8708,N_9363);
or U10850 (N_10850,N_8849,N_8586);
or U10851 (N_10851,N_9265,N_8862);
nor U10852 (N_10852,N_8433,N_8951);
nand U10853 (N_10853,N_8067,N_8088);
and U10854 (N_10854,N_8227,N_8208);
nor U10855 (N_10855,N_8006,N_8135);
nand U10856 (N_10856,N_9431,N_8851);
nor U10857 (N_10857,N_8880,N_9727);
xor U10858 (N_10858,N_9462,N_9660);
or U10859 (N_10859,N_9372,N_9261);
nor U10860 (N_10860,N_8825,N_8459);
nor U10861 (N_10861,N_8014,N_8329);
xnor U10862 (N_10862,N_8346,N_8583);
nand U10863 (N_10863,N_9182,N_8374);
nor U10864 (N_10864,N_9669,N_8757);
and U10865 (N_10865,N_9099,N_9162);
and U10866 (N_10866,N_9997,N_9774);
or U10867 (N_10867,N_9691,N_9489);
and U10868 (N_10868,N_9670,N_8526);
and U10869 (N_10869,N_9321,N_8920);
and U10870 (N_10870,N_9319,N_9436);
nor U10871 (N_10871,N_8404,N_9515);
or U10872 (N_10872,N_8631,N_9915);
or U10873 (N_10873,N_8589,N_8754);
nor U10874 (N_10874,N_8925,N_9304);
nor U10875 (N_10875,N_9895,N_9881);
nand U10876 (N_10876,N_8992,N_9327);
nand U10877 (N_10877,N_8836,N_9526);
or U10878 (N_10878,N_9587,N_8253);
nand U10879 (N_10879,N_9273,N_8438);
nor U10880 (N_10880,N_8861,N_9743);
nor U10881 (N_10881,N_9155,N_9450);
or U10882 (N_10882,N_9108,N_9618);
nand U10883 (N_10883,N_8240,N_9453);
and U10884 (N_10884,N_9086,N_9291);
or U10885 (N_10885,N_8015,N_9749);
xor U10886 (N_10886,N_8070,N_8971);
nor U10887 (N_10887,N_8214,N_8440);
nand U10888 (N_10888,N_9190,N_9528);
or U10889 (N_10889,N_8760,N_9942);
and U10890 (N_10890,N_8453,N_9829);
or U10891 (N_10891,N_9481,N_8797);
and U10892 (N_10892,N_8233,N_9317);
xor U10893 (N_10893,N_9224,N_9563);
nor U10894 (N_10894,N_8318,N_8824);
and U10895 (N_10895,N_8359,N_8688);
or U10896 (N_10896,N_9019,N_9033);
or U10897 (N_10897,N_9488,N_9690);
and U10898 (N_10898,N_8475,N_8306);
nand U10899 (N_10899,N_9485,N_9738);
and U10900 (N_10900,N_9676,N_8818);
nand U10901 (N_10901,N_8080,N_9333);
xor U10902 (N_10902,N_8287,N_8594);
nand U10903 (N_10903,N_9251,N_8003);
nand U10904 (N_10904,N_8500,N_9230);
or U10905 (N_10905,N_8963,N_9982);
nand U10906 (N_10906,N_8510,N_8759);
or U10907 (N_10907,N_9194,N_9312);
nand U10908 (N_10908,N_8411,N_9476);
or U10909 (N_10909,N_9483,N_9800);
xnor U10910 (N_10910,N_9813,N_8283);
nand U10911 (N_10911,N_8021,N_9168);
or U10912 (N_10912,N_9479,N_9721);
and U10913 (N_10913,N_9169,N_8357);
nor U10914 (N_10914,N_9287,N_9210);
xnor U10915 (N_10915,N_9524,N_9981);
and U10916 (N_10916,N_9211,N_8435);
or U10917 (N_10917,N_8286,N_9167);
or U10918 (N_10918,N_9842,N_8739);
nor U10919 (N_10919,N_8541,N_8044);
and U10920 (N_10920,N_9616,N_9124);
or U10921 (N_10921,N_8786,N_9995);
xnor U10922 (N_10922,N_9634,N_9258);
nor U10923 (N_10923,N_8025,N_9570);
or U10924 (N_10924,N_9003,N_9712);
nor U10925 (N_10925,N_8299,N_8721);
and U10926 (N_10926,N_8054,N_9953);
or U10927 (N_10927,N_9038,N_8103);
and U10928 (N_10928,N_9326,N_9988);
nand U10929 (N_10929,N_9504,N_8563);
nand U10930 (N_10930,N_9909,N_9329);
nor U10931 (N_10931,N_9341,N_8168);
and U10932 (N_10932,N_9332,N_9028);
or U10933 (N_10933,N_8102,N_8725);
and U10934 (N_10934,N_8509,N_9310);
nand U10935 (N_10935,N_8585,N_9424);
or U10936 (N_10936,N_9544,N_8181);
and U10937 (N_10937,N_8041,N_8106);
nor U10938 (N_10938,N_9011,N_8548);
nand U10939 (N_10939,N_9213,N_8345);
nor U10940 (N_10940,N_9178,N_8392);
or U10941 (N_10941,N_8295,N_9264);
and U10942 (N_10942,N_8213,N_9747);
nand U10943 (N_10943,N_9480,N_9986);
and U10944 (N_10944,N_9399,N_8901);
nand U10945 (N_10945,N_8046,N_9684);
nor U10946 (N_10946,N_9695,N_8691);
nor U10947 (N_10947,N_9732,N_9041);
nor U10948 (N_10948,N_8324,N_9730);
or U10949 (N_10949,N_9681,N_9710);
or U10950 (N_10950,N_9282,N_9208);
and U10951 (N_10951,N_9285,N_8478);
nor U10952 (N_10952,N_9717,N_9044);
and U10953 (N_10953,N_9077,N_8422);
nor U10954 (N_10954,N_9081,N_8190);
nor U10955 (N_10955,N_8058,N_9303);
nor U10956 (N_10956,N_8830,N_8055);
xnor U10957 (N_10957,N_9150,N_8804);
or U10958 (N_10958,N_8186,N_8660);
xor U10959 (N_10959,N_9815,N_8351);
and U10960 (N_10960,N_9490,N_9560);
nor U10961 (N_10961,N_8919,N_9822);
or U10962 (N_10962,N_9371,N_8138);
nand U10963 (N_10963,N_9139,N_9257);
nor U10964 (N_10964,N_9477,N_9276);
or U10965 (N_10965,N_9709,N_8685);
nor U10966 (N_10966,N_9499,N_9906);
nand U10967 (N_10967,N_9389,N_8494);
and U10968 (N_10968,N_9306,N_8178);
and U10969 (N_10969,N_9950,N_9958);
or U10970 (N_10970,N_8839,N_9763);
or U10971 (N_10971,N_8094,N_8322);
xor U10972 (N_10972,N_9574,N_9793);
and U10973 (N_10973,N_8075,N_9422);
and U10974 (N_10974,N_9576,N_8448);
nor U10975 (N_10975,N_8077,N_8831);
nor U10976 (N_10976,N_8532,N_8414);
and U10977 (N_10977,N_9247,N_8079);
or U10978 (N_10978,N_8658,N_9176);
and U10979 (N_10979,N_9487,N_8313);
nor U10980 (N_10980,N_9591,N_8866);
or U10981 (N_10981,N_9140,N_9255);
and U10982 (N_10982,N_8263,N_8304);
or U10983 (N_10983,N_9232,N_8385);
nand U10984 (N_10984,N_8461,N_9145);
nor U10985 (N_10985,N_8617,N_9112);
nor U10986 (N_10986,N_8623,N_8490);
nand U10987 (N_10987,N_8109,N_8927);
xnor U10988 (N_10988,N_9417,N_8246);
and U10989 (N_10989,N_9899,N_9573);
or U10990 (N_10990,N_8967,N_9220);
nor U10991 (N_10991,N_8550,N_9010);
and U10992 (N_10992,N_8907,N_8035);
nand U10993 (N_10993,N_9886,N_8042);
or U10994 (N_10994,N_9859,N_8719);
and U10995 (N_10995,N_8592,N_8043);
and U10996 (N_10996,N_9523,N_8012);
and U10997 (N_10997,N_9509,N_8806);
or U10998 (N_10998,N_9153,N_9383);
and U10999 (N_10999,N_9597,N_9510);
nor U11000 (N_11000,N_8812,N_8558);
and U11001 (N_11001,N_8274,N_8483);
nand U11002 (N_11002,N_9433,N_8087);
or U11003 (N_11003,N_9669,N_8812);
and U11004 (N_11004,N_9597,N_8309);
nand U11005 (N_11005,N_8816,N_9237);
or U11006 (N_11006,N_9578,N_9924);
nand U11007 (N_11007,N_8651,N_9665);
nand U11008 (N_11008,N_8648,N_9736);
and U11009 (N_11009,N_8850,N_8011);
nor U11010 (N_11010,N_8243,N_9251);
nor U11011 (N_11011,N_8723,N_8333);
nand U11012 (N_11012,N_9822,N_8876);
nor U11013 (N_11013,N_9429,N_8408);
or U11014 (N_11014,N_8615,N_8221);
nor U11015 (N_11015,N_9893,N_9617);
nor U11016 (N_11016,N_9882,N_9393);
nor U11017 (N_11017,N_8161,N_8799);
nand U11018 (N_11018,N_8919,N_8598);
or U11019 (N_11019,N_8901,N_9089);
nor U11020 (N_11020,N_9706,N_8734);
and U11021 (N_11021,N_8915,N_9855);
nand U11022 (N_11022,N_8357,N_9610);
and U11023 (N_11023,N_8338,N_9508);
and U11024 (N_11024,N_8435,N_9587);
nor U11025 (N_11025,N_9188,N_9224);
nand U11026 (N_11026,N_9014,N_9499);
nand U11027 (N_11027,N_9897,N_9642);
or U11028 (N_11028,N_9401,N_8548);
and U11029 (N_11029,N_9330,N_8665);
or U11030 (N_11030,N_9131,N_9499);
or U11031 (N_11031,N_8939,N_9535);
xnor U11032 (N_11032,N_8518,N_9217);
nand U11033 (N_11033,N_8440,N_8528);
or U11034 (N_11034,N_8906,N_9788);
and U11035 (N_11035,N_8049,N_9839);
nand U11036 (N_11036,N_8043,N_8980);
nand U11037 (N_11037,N_8936,N_9545);
nor U11038 (N_11038,N_9681,N_9850);
nand U11039 (N_11039,N_9631,N_9767);
nor U11040 (N_11040,N_9846,N_8320);
and U11041 (N_11041,N_8937,N_8278);
and U11042 (N_11042,N_8124,N_8087);
and U11043 (N_11043,N_8745,N_8066);
xnor U11044 (N_11044,N_8339,N_9365);
or U11045 (N_11045,N_9118,N_9007);
nor U11046 (N_11046,N_8281,N_9858);
or U11047 (N_11047,N_8555,N_8779);
nand U11048 (N_11048,N_8107,N_9863);
nand U11049 (N_11049,N_9019,N_9973);
nor U11050 (N_11050,N_8713,N_8464);
or U11051 (N_11051,N_8832,N_9226);
and U11052 (N_11052,N_8414,N_8989);
or U11053 (N_11053,N_8453,N_8242);
nand U11054 (N_11054,N_8935,N_9477);
or U11055 (N_11055,N_8170,N_8992);
and U11056 (N_11056,N_9600,N_9570);
and U11057 (N_11057,N_9066,N_8967);
and U11058 (N_11058,N_8381,N_9585);
nor U11059 (N_11059,N_8454,N_8468);
or U11060 (N_11060,N_9824,N_9152);
nor U11061 (N_11061,N_9873,N_8308);
nand U11062 (N_11062,N_9132,N_8684);
or U11063 (N_11063,N_8762,N_9758);
nand U11064 (N_11064,N_8478,N_9129);
nand U11065 (N_11065,N_8635,N_8524);
and U11066 (N_11066,N_8118,N_8252);
or U11067 (N_11067,N_8460,N_8630);
nand U11068 (N_11068,N_9692,N_8195);
nand U11069 (N_11069,N_8358,N_9341);
nand U11070 (N_11070,N_9677,N_8599);
nor U11071 (N_11071,N_8142,N_8112);
and U11072 (N_11072,N_8060,N_8235);
or U11073 (N_11073,N_9350,N_8898);
or U11074 (N_11074,N_8852,N_9726);
and U11075 (N_11075,N_9146,N_9592);
nor U11076 (N_11076,N_9568,N_9470);
and U11077 (N_11077,N_8390,N_9682);
nor U11078 (N_11078,N_8339,N_9812);
or U11079 (N_11079,N_9909,N_9171);
or U11080 (N_11080,N_8694,N_9183);
nand U11081 (N_11081,N_9094,N_9332);
nor U11082 (N_11082,N_9393,N_8568);
and U11083 (N_11083,N_9587,N_9903);
and U11084 (N_11084,N_8843,N_9044);
and U11085 (N_11085,N_8001,N_9485);
nor U11086 (N_11086,N_8516,N_8631);
nand U11087 (N_11087,N_8201,N_8100);
nor U11088 (N_11088,N_8987,N_8784);
nand U11089 (N_11089,N_8036,N_8175);
nor U11090 (N_11090,N_8958,N_9703);
nor U11091 (N_11091,N_8219,N_9917);
nor U11092 (N_11092,N_8972,N_9202);
and U11093 (N_11093,N_9395,N_9964);
and U11094 (N_11094,N_8598,N_9989);
nand U11095 (N_11095,N_9349,N_9292);
nand U11096 (N_11096,N_8795,N_9320);
and U11097 (N_11097,N_9798,N_8775);
nand U11098 (N_11098,N_8556,N_8007);
nor U11099 (N_11099,N_8480,N_9533);
or U11100 (N_11100,N_8256,N_8582);
and U11101 (N_11101,N_8764,N_9209);
or U11102 (N_11102,N_9336,N_8599);
and U11103 (N_11103,N_8404,N_8043);
or U11104 (N_11104,N_9282,N_8686);
nor U11105 (N_11105,N_9107,N_8540);
or U11106 (N_11106,N_8902,N_8923);
nand U11107 (N_11107,N_9752,N_8057);
nor U11108 (N_11108,N_9682,N_8813);
nor U11109 (N_11109,N_9026,N_8769);
nor U11110 (N_11110,N_9712,N_9617);
and U11111 (N_11111,N_9401,N_9544);
nand U11112 (N_11112,N_8682,N_9877);
or U11113 (N_11113,N_9417,N_8613);
or U11114 (N_11114,N_9454,N_8666);
and U11115 (N_11115,N_9374,N_8459);
and U11116 (N_11116,N_9042,N_9755);
nor U11117 (N_11117,N_9292,N_8191);
and U11118 (N_11118,N_8836,N_9967);
xnor U11119 (N_11119,N_8200,N_8475);
or U11120 (N_11120,N_9467,N_8447);
nor U11121 (N_11121,N_8899,N_8911);
and U11122 (N_11122,N_9188,N_9964);
and U11123 (N_11123,N_8582,N_9459);
nor U11124 (N_11124,N_8212,N_8335);
and U11125 (N_11125,N_9914,N_8877);
or U11126 (N_11126,N_9755,N_9116);
or U11127 (N_11127,N_8251,N_8913);
or U11128 (N_11128,N_9000,N_8693);
or U11129 (N_11129,N_9149,N_8372);
nor U11130 (N_11130,N_9971,N_8976);
nor U11131 (N_11131,N_9226,N_9806);
nand U11132 (N_11132,N_8179,N_8200);
nand U11133 (N_11133,N_8129,N_8903);
or U11134 (N_11134,N_9864,N_8848);
and U11135 (N_11135,N_9459,N_9254);
nor U11136 (N_11136,N_9947,N_8824);
nor U11137 (N_11137,N_9976,N_9007);
or U11138 (N_11138,N_8410,N_8944);
nor U11139 (N_11139,N_9454,N_8704);
nor U11140 (N_11140,N_9373,N_8315);
or U11141 (N_11141,N_9893,N_8145);
nand U11142 (N_11142,N_8299,N_8684);
and U11143 (N_11143,N_8562,N_9365);
nor U11144 (N_11144,N_9736,N_9168);
and U11145 (N_11145,N_9885,N_9827);
nand U11146 (N_11146,N_8766,N_9037);
or U11147 (N_11147,N_9721,N_8068);
and U11148 (N_11148,N_9617,N_9887);
nand U11149 (N_11149,N_8551,N_8905);
nand U11150 (N_11150,N_9455,N_9852);
and U11151 (N_11151,N_8831,N_8763);
or U11152 (N_11152,N_8619,N_9608);
nand U11153 (N_11153,N_9593,N_8079);
nor U11154 (N_11154,N_8947,N_8655);
or U11155 (N_11155,N_8464,N_8954);
xnor U11156 (N_11156,N_8941,N_9694);
xnor U11157 (N_11157,N_8522,N_8271);
or U11158 (N_11158,N_9620,N_8147);
or U11159 (N_11159,N_8806,N_9922);
nor U11160 (N_11160,N_9792,N_8700);
and U11161 (N_11161,N_8097,N_9053);
or U11162 (N_11162,N_9494,N_9493);
and U11163 (N_11163,N_9510,N_9323);
and U11164 (N_11164,N_8158,N_9446);
and U11165 (N_11165,N_8631,N_9265);
nand U11166 (N_11166,N_8448,N_8116);
or U11167 (N_11167,N_8967,N_8088);
nor U11168 (N_11168,N_8337,N_8544);
or U11169 (N_11169,N_9906,N_9289);
nor U11170 (N_11170,N_8288,N_9181);
and U11171 (N_11171,N_8409,N_8622);
or U11172 (N_11172,N_8570,N_9221);
and U11173 (N_11173,N_9024,N_8904);
or U11174 (N_11174,N_9672,N_9851);
and U11175 (N_11175,N_8760,N_8119);
nand U11176 (N_11176,N_9320,N_8203);
nor U11177 (N_11177,N_9071,N_8902);
nand U11178 (N_11178,N_8858,N_9967);
or U11179 (N_11179,N_8819,N_9329);
and U11180 (N_11180,N_8462,N_8959);
or U11181 (N_11181,N_8897,N_9619);
or U11182 (N_11182,N_8815,N_9206);
nand U11183 (N_11183,N_9287,N_9104);
or U11184 (N_11184,N_9321,N_9983);
and U11185 (N_11185,N_9467,N_9730);
or U11186 (N_11186,N_9072,N_9223);
nand U11187 (N_11187,N_9350,N_8860);
and U11188 (N_11188,N_9137,N_9474);
nor U11189 (N_11189,N_9528,N_9091);
nor U11190 (N_11190,N_8072,N_8766);
nor U11191 (N_11191,N_8399,N_8467);
and U11192 (N_11192,N_9414,N_8556);
or U11193 (N_11193,N_9663,N_9031);
or U11194 (N_11194,N_8331,N_8520);
nor U11195 (N_11195,N_8257,N_9080);
nand U11196 (N_11196,N_9197,N_8570);
and U11197 (N_11197,N_9089,N_8569);
and U11198 (N_11198,N_8159,N_9591);
and U11199 (N_11199,N_9782,N_8375);
nand U11200 (N_11200,N_8456,N_8567);
and U11201 (N_11201,N_8939,N_9040);
and U11202 (N_11202,N_9085,N_8148);
nor U11203 (N_11203,N_8673,N_8526);
or U11204 (N_11204,N_8359,N_8379);
or U11205 (N_11205,N_8990,N_9457);
or U11206 (N_11206,N_9148,N_8806);
nor U11207 (N_11207,N_9617,N_8063);
nand U11208 (N_11208,N_8580,N_8248);
or U11209 (N_11209,N_8743,N_9970);
nor U11210 (N_11210,N_9296,N_9712);
nand U11211 (N_11211,N_8131,N_8235);
nand U11212 (N_11212,N_9686,N_9598);
nand U11213 (N_11213,N_9450,N_8191);
xnor U11214 (N_11214,N_8207,N_8739);
nor U11215 (N_11215,N_9415,N_9755);
and U11216 (N_11216,N_8336,N_8083);
and U11217 (N_11217,N_8931,N_9068);
nand U11218 (N_11218,N_9965,N_9231);
nor U11219 (N_11219,N_9116,N_8388);
and U11220 (N_11220,N_8535,N_8878);
nor U11221 (N_11221,N_9262,N_9870);
nand U11222 (N_11222,N_8794,N_8208);
xnor U11223 (N_11223,N_8634,N_8180);
and U11224 (N_11224,N_9258,N_9281);
nor U11225 (N_11225,N_8217,N_9002);
or U11226 (N_11226,N_9622,N_8750);
or U11227 (N_11227,N_8721,N_9247);
and U11228 (N_11228,N_8846,N_9269);
nor U11229 (N_11229,N_8745,N_9973);
nand U11230 (N_11230,N_9546,N_8195);
nand U11231 (N_11231,N_9025,N_9996);
or U11232 (N_11232,N_8311,N_9201);
nand U11233 (N_11233,N_9704,N_8215);
or U11234 (N_11234,N_8405,N_9559);
nand U11235 (N_11235,N_9749,N_9003);
or U11236 (N_11236,N_8246,N_8463);
and U11237 (N_11237,N_9501,N_9556);
xnor U11238 (N_11238,N_9268,N_8328);
or U11239 (N_11239,N_9656,N_8472);
or U11240 (N_11240,N_9094,N_8045);
nand U11241 (N_11241,N_9867,N_8283);
nand U11242 (N_11242,N_8311,N_9741);
nand U11243 (N_11243,N_9071,N_9558);
nand U11244 (N_11244,N_8770,N_8720);
or U11245 (N_11245,N_9753,N_9789);
nor U11246 (N_11246,N_8235,N_9760);
nand U11247 (N_11247,N_9034,N_9740);
and U11248 (N_11248,N_9852,N_9566);
nand U11249 (N_11249,N_9363,N_8802);
nor U11250 (N_11250,N_8560,N_8446);
and U11251 (N_11251,N_8518,N_8625);
nand U11252 (N_11252,N_9844,N_8585);
nand U11253 (N_11253,N_8713,N_8770);
nand U11254 (N_11254,N_9522,N_9451);
nand U11255 (N_11255,N_8180,N_9631);
or U11256 (N_11256,N_8194,N_8356);
or U11257 (N_11257,N_8025,N_8450);
nor U11258 (N_11258,N_8341,N_9051);
or U11259 (N_11259,N_9119,N_8846);
or U11260 (N_11260,N_9435,N_8341);
nor U11261 (N_11261,N_9217,N_8865);
or U11262 (N_11262,N_8334,N_9832);
or U11263 (N_11263,N_8803,N_8752);
nand U11264 (N_11264,N_8646,N_8180);
or U11265 (N_11265,N_8479,N_8642);
nand U11266 (N_11266,N_8816,N_9151);
and U11267 (N_11267,N_9595,N_8560);
nand U11268 (N_11268,N_9181,N_9015);
nand U11269 (N_11269,N_9611,N_8814);
or U11270 (N_11270,N_9683,N_8103);
or U11271 (N_11271,N_9226,N_9316);
nor U11272 (N_11272,N_9719,N_8119);
or U11273 (N_11273,N_8426,N_8646);
nor U11274 (N_11274,N_8415,N_9216);
nor U11275 (N_11275,N_9106,N_8962);
nand U11276 (N_11276,N_8419,N_9109);
or U11277 (N_11277,N_8591,N_8305);
nor U11278 (N_11278,N_9097,N_8480);
and U11279 (N_11279,N_9023,N_8589);
and U11280 (N_11280,N_9075,N_9207);
nor U11281 (N_11281,N_8612,N_8792);
xnor U11282 (N_11282,N_8432,N_9968);
and U11283 (N_11283,N_9080,N_9656);
nand U11284 (N_11284,N_9014,N_8760);
nor U11285 (N_11285,N_9779,N_9599);
or U11286 (N_11286,N_9719,N_9398);
nand U11287 (N_11287,N_9680,N_8265);
or U11288 (N_11288,N_9958,N_8260);
or U11289 (N_11289,N_9349,N_8190);
and U11290 (N_11290,N_9654,N_8132);
nor U11291 (N_11291,N_9761,N_9257);
nor U11292 (N_11292,N_9253,N_9061);
nor U11293 (N_11293,N_9347,N_9645);
nor U11294 (N_11294,N_9962,N_9059);
or U11295 (N_11295,N_8784,N_8222);
nand U11296 (N_11296,N_8257,N_8004);
and U11297 (N_11297,N_9322,N_8566);
nor U11298 (N_11298,N_9324,N_8698);
nand U11299 (N_11299,N_9892,N_9681);
nand U11300 (N_11300,N_8579,N_8995);
or U11301 (N_11301,N_8173,N_9823);
or U11302 (N_11302,N_8612,N_9766);
nand U11303 (N_11303,N_9454,N_8599);
or U11304 (N_11304,N_8038,N_9487);
and U11305 (N_11305,N_8629,N_8730);
and U11306 (N_11306,N_9714,N_8615);
or U11307 (N_11307,N_8555,N_8696);
nor U11308 (N_11308,N_9884,N_9032);
or U11309 (N_11309,N_9488,N_9469);
or U11310 (N_11310,N_8371,N_8502);
nor U11311 (N_11311,N_8636,N_9269);
or U11312 (N_11312,N_8706,N_9413);
and U11313 (N_11313,N_8797,N_8188);
and U11314 (N_11314,N_9642,N_9242);
nand U11315 (N_11315,N_8973,N_9072);
and U11316 (N_11316,N_9503,N_8432);
nor U11317 (N_11317,N_9124,N_8189);
nor U11318 (N_11318,N_8386,N_8496);
or U11319 (N_11319,N_9223,N_8759);
and U11320 (N_11320,N_9812,N_9070);
nand U11321 (N_11321,N_8156,N_8799);
nand U11322 (N_11322,N_9646,N_8844);
nor U11323 (N_11323,N_8264,N_8090);
nor U11324 (N_11324,N_9904,N_8164);
nor U11325 (N_11325,N_8667,N_8042);
or U11326 (N_11326,N_9835,N_9021);
and U11327 (N_11327,N_9973,N_9476);
nand U11328 (N_11328,N_8784,N_9384);
and U11329 (N_11329,N_9164,N_8829);
or U11330 (N_11330,N_8597,N_9108);
nor U11331 (N_11331,N_9340,N_9956);
and U11332 (N_11332,N_9839,N_9688);
or U11333 (N_11333,N_8009,N_8771);
or U11334 (N_11334,N_8955,N_8539);
nand U11335 (N_11335,N_8647,N_9132);
nor U11336 (N_11336,N_8728,N_8033);
or U11337 (N_11337,N_8229,N_8101);
or U11338 (N_11338,N_9433,N_8572);
xor U11339 (N_11339,N_9818,N_8408);
and U11340 (N_11340,N_9785,N_8949);
or U11341 (N_11341,N_8497,N_8755);
and U11342 (N_11342,N_8383,N_8899);
nand U11343 (N_11343,N_9310,N_8804);
and U11344 (N_11344,N_9472,N_8263);
nand U11345 (N_11345,N_9443,N_8394);
or U11346 (N_11346,N_9669,N_8780);
or U11347 (N_11347,N_9240,N_8085);
nor U11348 (N_11348,N_9788,N_9754);
or U11349 (N_11349,N_8900,N_8683);
xor U11350 (N_11350,N_8729,N_9319);
and U11351 (N_11351,N_9638,N_8462);
or U11352 (N_11352,N_8694,N_9470);
nor U11353 (N_11353,N_8055,N_9781);
and U11354 (N_11354,N_9502,N_9886);
and U11355 (N_11355,N_9686,N_8514);
and U11356 (N_11356,N_8151,N_9800);
or U11357 (N_11357,N_9872,N_9683);
nand U11358 (N_11358,N_9819,N_9730);
or U11359 (N_11359,N_9468,N_9301);
or U11360 (N_11360,N_9216,N_8551);
and U11361 (N_11361,N_8856,N_9313);
nand U11362 (N_11362,N_9488,N_9099);
or U11363 (N_11363,N_8196,N_8836);
xnor U11364 (N_11364,N_9535,N_8818);
nor U11365 (N_11365,N_9286,N_9025);
nor U11366 (N_11366,N_8203,N_9462);
or U11367 (N_11367,N_9990,N_9077);
nor U11368 (N_11368,N_9633,N_8467);
and U11369 (N_11369,N_8381,N_8059);
and U11370 (N_11370,N_9642,N_8417);
nor U11371 (N_11371,N_9989,N_8260);
nand U11372 (N_11372,N_9747,N_9840);
or U11373 (N_11373,N_9504,N_8443);
and U11374 (N_11374,N_8724,N_9419);
and U11375 (N_11375,N_9428,N_9477);
nand U11376 (N_11376,N_8165,N_9709);
nor U11377 (N_11377,N_8785,N_9346);
nor U11378 (N_11378,N_8779,N_8867);
nor U11379 (N_11379,N_8515,N_9883);
nand U11380 (N_11380,N_8391,N_8417);
and U11381 (N_11381,N_9418,N_9767);
or U11382 (N_11382,N_9279,N_8026);
nand U11383 (N_11383,N_9627,N_8607);
nand U11384 (N_11384,N_8698,N_9141);
nor U11385 (N_11385,N_8479,N_8766);
and U11386 (N_11386,N_8736,N_8530);
nor U11387 (N_11387,N_8063,N_9989);
nand U11388 (N_11388,N_9348,N_9945);
or U11389 (N_11389,N_9789,N_9291);
and U11390 (N_11390,N_8155,N_8656);
xnor U11391 (N_11391,N_8893,N_9232);
nor U11392 (N_11392,N_9527,N_9378);
and U11393 (N_11393,N_8009,N_8583);
nor U11394 (N_11394,N_8838,N_9110);
or U11395 (N_11395,N_9854,N_8616);
xnor U11396 (N_11396,N_8534,N_8279);
and U11397 (N_11397,N_8367,N_9920);
nor U11398 (N_11398,N_8046,N_9638);
nand U11399 (N_11399,N_8977,N_8469);
and U11400 (N_11400,N_8040,N_8212);
and U11401 (N_11401,N_9080,N_8300);
nand U11402 (N_11402,N_8637,N_9308);
or U11403 (N_11403,N_8764,N_9590);
and U11404 (N_11404,N_9713,N_8253);
and U11405 (N_11405,N_9873,N_8945);
and U11406 (N_11406,N_9988,N_9143);
nand U11407 (N_11407,N_8043,N_9865);
and U11408 (N_11408,N_9584,N_9174);
or U11409 (N_11409,N_9662,N_9357);
and U11410 (N_11410,N_9903,N_8283);
and U11411 (N_11411,N_9683,N_8909);
nor U11412 (N_11412,N_8468,N_9876);
or U11413 (N_11413,N_9478,N_8183);
nor U11414 (N_11414,N_9675,N_8853);
or U11415 (N_11415,N_9684,N_8857);
nand U11416 (N_11416,N_9371,N_9171);
or U11417 (N_11417,N_8817,N_8477);
nand U11418 (N_11418,N_8495,N_8603);
and U11419 (N_11419,N_8055,N_8447);
nor U11420 (N_11420,N_8410,N_9467);
or U11421 (N_11421,N_8596,N_8520);
and U11422 (N_11422,N_8710,N_8997);
or U11423 (N_11423,N_8916,N_8563);
nand U11424 (N_11424,N_9873,N_9325);
nand U11425 (N_11425,N_8566,N_8579);
and U11426 (N_11426,N_8068,N_8462);
nor U11427 (N_11427,N_8692,N_9574);
and U11428 (N_11428,N_8833,N_9054);
nand U11429 (N_11429,N_8217,N_9006);
and U11430 (N_11430,N_9258,N_9777);
nor U11431 (N_11431,N_8542,N_9168);
xnor U11432 (N_11432,N_8556,N_8174);
and U11433 (N_11433,N_8226,N_9122);
nor U11434 (N_11434,N_9515,N_9367);
or U11435 (N_11435,N_8346,N_9604);
nand U11436 (N_11436,N_9735,N_8954);
nand U11437 (N_11437,N_9811,N_8482);
nand U11438 (N_11438,N_8368,N_9931);
and U11439 (N_11439,N_8873,N_9486);
nand U11440 (N_11440,N_9499,N_8124);
nand U11441 (N_11441,N_8435,N_9595);
nor U11442 (N_11442,N_9607,N_9038);
nor U11443 (N_11443,N_8975,N_9725);
nand U11444 (N_11444,N_9865,N_8550);
nor U11445 (N_11445,N_8188,N_8674);
nand U11446 (N_11446,N_9730,N_9084);
or U11447 (N_11447,N_9253,N_9607);
or U11448 (N_11448,N_8948,N_9714);
nor U11449 (N_11449,N_9942,N_9826);
nand U11450 (N_11450,N_9069,N_9745);
and U11451 (N_11451,N_9493,N_9053);
nand U11452 (N_11452,N_8980,N_8804);
or U11453 (N_11453,N_9987,N_8890);
nor U11454 (N_11454,N_8707,N_9998);
nor U11455 (N_11455,N_9323,N_8883);
xor U11456 (N_11456,N_9580,N_9156);
nand U11457 (N_11457,N_8722,N_8426);
and U11458 (N_11458,N_9451,N_8417);
nand U11459 (N_11459,N_8415,N_9816);
nand U11460 (N_11460,N_9407,N_9344);
and U11461 (N_11461,N_9692,N_9886);
and U11462 (N_11462,N_8914,N_8477);
and U11463 (N_11463,N_9777,N_8996);
nand U11464 (N_11464,N_9139,N_8267);
nor U11465 (N_11465,N_9240,N_8585);
or U11466 (N_11466,N_8250,N_8058);
nor U11467 (N_11467,N_9404,N_9185);
and U11468 (N_11468,N_8448,N_9451);
nor U11469 (N_11469,N_8127,N_9533);
or U11470 (N_11470,N_9320,N_9283);
nand U11471 (N_11471,N_9651,N_8578);
nand U11472 (N_11472,N_9404,N_9051);
nand U11473 (N_11473,N_8809,N_8240);
and U11474 (N_11474,N_9097,N_8513);
nor U11475 (N_11475,N_8372,N_9280);
and U11476 (N_11476,N_8333,N_9795);
nand U11477 (N_11477,N_8949,N_8089);
nor U11478 (N_11478,N_9332,N_9701);
and U11479 (N_11479,N_9848,N_9313);
nand U11480 (N_11480,N_9451,N_9610);
or U11481 (N_11481,N_9515,N_9210);
and U11482 (N_11482,N_9868,N_8536);
nor U11483 (N_11483,N_8629,N_8737);
or U11484 (N_11484,N_8387,N_9040);
and U11485 (N_11485,N_9641,N_9992);
and U11486 (N_11486,N_9048,N_8786);
or U11487 (N_11487,N_9259,N_9905);
and U11488 (N_11488,N_8306,N_9627);
and U11489 (N_11489,N_8935,N_9307);
and U11490 (N_11490,N_9115,N_8142);
or U11491 (N_11491,N_9297,N_8238);
nor U11492 (N_11492,N_8313,N_9908);
and U11493 (N_11493,N_9152,N_8987);
nor U11494 (N_11494,N_8436,N_9990);
xnor U11495 (N_11495,N_8757,N_8949);
nand U11496 (N_11496,N_8805,N_8312);
and U11497 (N_11497,N_9615,N_9498);
and U11498 (N_11498,N_9281,N_8954);
or U11499 (N_11499,N_8121,N_9788);
and U11500 (N_11500,N_8046,N_9112);
and U11501 (N_11501,N_8952,N_8346);
nand U11502 (N_11502,N_9199,N_9050);
and U11503 (N_11503,N_9155,N_9328);
nor U11504 (N_11504,N_8864,N_9488);
nor U11505 (N_11505,N_8808,N_8141);
and U11506 (N_11506,N_8861,N_9110);
nand U11507 (N_11507,N_8283,N_8470);
nor U11508 (N_11508,N_9261,N_9933);
nand U11509 (N_11509,N_9305,N_9639);
nor U11510 (N_11510,N_8748,N_8146);
nor U11511 (N_11511,N_9380,N_9217);
and U11512 (N_11512,N_8227,N_9375);
and U11513 (N_11513,N_8419,N_9682);
and U11514 (N_11514,N_9743,N_8235);
nand U11515 (N_11515,N_9469,N_8193);
and U11516 (N_11516,N_8051,N_8220);
or U11517 (N_11517,N_9918,N_8374);
nor U11518 (N_11518,N_8164,N_9423);
or U11519 (N_11519,N_9474,N_9053);
nand U11520 (N_11520,N_9386,N_9672);
nand U11521 (N_11521,N_8996,N_8435);
nor U11522 (N_11522,N_8737,N_8969);
and U11523 (N_11523,N_8808,N_8446);
nand U11524 (N_11524,N_8511,N_9717);
nand U11525 (N_11525,N_9648,N_8461);
and U11526 (N_11526,N_8697,N_8017);
xnor U11527 (N_11527,N_9032,N_8791);
nand U11528 (N_11528,N_8238,N_9466);
nor U11529 (N_11529,N_8618,N_9753);
and U11530 (N_11530,N_9965,N_9876);
and U11531 (N_11531,N_8525,N_9648);
nand U11532 (N_11532,N_8553,N_9882);
nand U11533 (N_11533,N_8647,N_8373);
and U11534 (N_11534,N_8303,N_8389);
or U11535 (N_11535,N_9063,N_9286);
or U11536 (N_11536,N_8305,N_9746);
or U11537 (N_11537,N_9458,N_8336);
or U11538 (N_11538,N_9791,N_8754);
or U11539 (N_11539,N_9126,N_8181);
xnor U11540 (N_11540,N_9270,N_9119);
nor U11541 (N_11541,N_9407,N_9571);
xnor U11542 (N_11542,N_9003,N_8960);
nand U11543 (N_11543,N_9781,N_9302);
nand U11544 (N_11544,N_8537,N_9330);
nand U11545 (N_11545,N_9613,N_9445);
or U11546 (N_11546,N_8619,N_8781);
nor U11547 (N_11547,N_9640,N_9089);
or U11548 (N_11548,N_9978,N_8688);
nor U11549 (N_11549,N_9692,N_9624);
nand U11550 (N_11550,N_8250,N_8930);
and U11551 (N_11551,N_8684,N_9174);
nand U11552 (N_11552,N_9060,N_8496);
xor U11553 (N_11553,N_8419,N_8575);
nand U11554 (N_11554,N_9090,N_8318);
and U11555 (N_11555,N_9262,N_9614);
nor U11556 (N_11556,N_9487,N_9620);
and U11557 (N_11557,N_9379,N_9042);
or U11558 (N_11558,N_9386,N_9373);
nor U11559 (N_11559,N_8954,N_9388);
and U11560 (N_11560,N_9901,N_9126);
or U11561 (N_11561,N_9789,N_9414);
xnor U11562 (N_11562,N_9605,N_8945);
nor U11563 (N_11563,N_9121,N_9744);
nor U11564 (N_11564,N_9114,N_8408);
or U11565 (N_11565,N_9283,N_9209);
nor U11566 (N_11566,N_9801,N_8816);
nor U11567 (N_11567,N_9244,N_9898);
or U11568 (N_11568,N_8984,N_9324);
nor U11569 (N_11569,N_9012,N_9466);
and U11570 (N_11570,N_9918,N_8813);
nand U11571 (N_11571,N_8786,N_8450);
and U11572 (N_11572,N_9595,N_8011);
nand U11573 (N_11573,N_8221,N_8658);
nand U11574 (N_11574,N_9538,N_8741);
or U11575 (N_11575,N_8042,N_8923);
nor U11576 (N_11576,N_9505,N_8824);
nor U11577 (N_11577,N_8682,N_8177);
nor U11578 (N_11578,N_9835,N_8575);
nand U11579 (N_11579,N_8417,N_8443);
nand U11580 (N_11580,N_9072,N_8558);
nand U11581 (N_11581,N_9744,N_9139);
or U11582 (N_11582,N_9475,N_9257);
or U11583 (N_11583,N_9036,N_9733);
nor U11584 (N_11584,N_8905,N_8636);
nor U11585 (N_11585,N_8961,N_8349);
xnor U11586 (N_11586,N_9107,N_9598);
nand U11587 (N_11587,N_9854,N_8521);
nor U11588 (N_11588,N_9074,N_8770);
nand U11589 (N_11589,N_8001,N_8868);
or U11590 (N_11590,N_9401,N_9666);
and U11591 (N_11591,N_8243,N_9392);
nor U11592 (N_11592,N_8804,N_8228);
xor U11593 (N_11593,N_8442,N_8972);
nor U11594 (N_11594,N_9970,N_9964);
nor U11595 (N_11595,N_9706,N_8618);
and U11596 (N_11596,N_9993,N_9685);
nor U11597 (N_11597,N_9945,N_9450);
or U11598 (N_11598,N_9590,N_9597);
nor U11599 (N_11599,N_8458,N_9912);
nor U11600 (N_11600,N_8002,N_9854);
nor U11601 (N_11601,N_8561,N_9045);
and U11602 (N_11602,N_8942,N_9932);
and U11603 (N_11603,N_9894,N_9442);
and U11604 (N_11604,N_9783,N_9852);
nor U11605 (N_11605,N_8907,N_8659);
or U11606 (N_11606,N_8656,N_9882);
or U11607 (N_11607,N_8665,N_8885);
or U11608 (N_11608,N_8738,N_9551);
or U11609 (N_11609,N_8040,N_9047);
or U11610 (N_11610,N_9249,N_9465);
and U11611 (N_11611,N_8123,N_8047);
or U11612 (N_11612,N_9995,N_9250);
nand U11613 (N_11613,N_8422,N_9740);
and U11614 (N_11614,N_8669,N_9184);
nor U11615 (N_11615,N_9376,N_8469);
or U11616 (N_11616,N_9640,N_8421);
nor U11617 (N_11617,N_9156,N_9645);
or U11618 (N_11618,N_9269,N_8815);
nor U11619 (N_11619,N_8616,N_8976);
nor U11620 (N_11620,N_8843,N_9341);
and U11621 (N_11621,N_9366,N_8159);
xor U11622 (N_11622,N_9502,N_8743);
or U11623 (N_11623,N_9432,N_8825);
nor U11624 (N_11624,N_8384,N_9074);
nor U11625 (N_11625,N_9906,N_9925);
or U11626 (N_11626,N_8443,N_8535);
or U11627 (N_11627,N_8748,N_8079);
nand U11628 (N_11628,N_9255,N_8379);
nor U11629 (N_11629,N_8363,N_8437);
or U11630 (N_11630,N_8674,N_9256);
and U11631 (N_11631,N_9586,N_9743);
and U11632 (N_11632,N_9508,N_9419);
and U11633 (N_11633,N_8819,N_9747);
and U11634 (N_11634,N_9607,N_8813);
xnor U11635 (N_11635,N_9246,N_9829);
nand U11636 (N_11636,N_9186,N_8698);
and U11637 (N_11637,N_8270,N_9925);
or U11638 (N_11638,N_9100,N_9161);
and U11639 (N_11639,N_9354,N_9273);
or U11640 (N_11640,N_9023,N_8350);
or U11641 (N_11641,N_8234,N_9193);
and U11642 (N_11642,N_9695,N_8800);
nor U11643 (N_11643,N_9059,N_9176);
nand U11644 (N_11644,N_9765,N_8499);
nand U11645 (N_11645,N_9665,N_8569);
nand U11646 (N_11646,N_8903,N_9431);
and U11647 (N_11647,N_9537,N_9039);
or U11648 (N_11648,N_9690,N_8931);
and U11649 (N_11649,N_8068,N_9605);
and U11650 (N_11650,N_9849,N_8105);
nand U11651 (N_11651,N_9516,N_9593);
and U11652 (N_11652,N_9178,N_9074);
nand U11653 (N_11653,N_9807,N_9573);
and U11654 (N_11654,N_9091,N_9045);
xor U11655 (N_11655,N_8212,N_9698);
or U11656 (N_11656,N_8028,N_8659);
nand U11657 (N_11657,N_8657,N_9792);
nand U11658 (N_11658,N_9185,N_9203);
or U11659 (N_11659,N_9611,N_9451);
and U11660 (N_11660,N_9730,N_9605);
nand U11661 (N_11661,N_8450,N_8338);
nand U11662 (N_11662,N_9882,N_9879);
nor U11663 (N_11663,N_9577,N_9625);
or U11664 (N_11664,N_8020,N_8974);
or U11665 (N_11665,N_8746,N_9925);
nor U11666 (N_11666,N_8429,N_9371);
and U11667 (N_11667,N_8380,N_8427);
or U11668 (N_11668,N_9685,N_8669);
and U11669 (N_11669,N_9928,N_9755);
and U11670 (N_11670,N_8206,N_9704);
or U11671 (N_11671,N_8284,N_9863);
or U11672 (N_11672,N_9223,N_8035);
nand U11673 (N_11673,N_8041,N_8699);
nand U11674 (N_11674,N_8722,N_8240);
or U11675 (N_11675,N_8709,N_9396);
nand U11676 (N_11676,N_8300,N_9534);
or U11677 (N_11677,N_9128,N_9656);
nand U11678 (N_11678,N_8434,N_9542);
nand U11679 (N_11679,N_9554,N_9814);
and U11680 (N_11680,N_8223,N_8033);
or U11681 (N_11681,N_9773,N_8038);
nor U11682 (N_11682,N_9488,N_9981);
and U11683 (N_11683,N_9787,N_9235);
and U11684 (N_11684,N_9109,N_9960);
xor U11685 (N_11685,N_9665,N_8299);
and U11686 (N_11686,N_8246,N_9033);
nand U11687 (N_11687,N_8041,N_8243);
or U11688 (N_11688,N_9407,N_8578);
xnor U11689 (N_11689,N_9229,N_8953);
nor U11690 (N_11690,N_9325,N_8110);
nand U11691 (N_11691,N_8855,N_9968);
nor U11692 (N_11692,N_8331,N_8562);
nand U11693 (N_11693,N_8616,N_9869);
nor U11694 (N_11694,N_8669,N_8845);
and U11695 (N_11695,N_9221,N_8980);
and U11696 (N_11696,N_8055,N_9347);
nor U11697 (N_11697,N_8256,N_9041);
and U11698 (N_11698,N_9357,N_9729);
or U11699 (N_11699,N_9036,N_8342);
and U11700 (N_11700,N_8016,N_9579);
or U11701 (N_11701,N_8877,N_8463);
nand U11702 (N_11702,N_9403,N_8739);
nor U11703 (N_11703,N_8914,N_8212);
or U11704 (N_11704,N_9631,N_8885);
nand U11705 (N_11705,N_9076,N_9065);
and U11706 (N_11706,N_8037,N_8590);
nor U11707 (N_11707,N_8348,N_9006);
nor U11708 (N_11708,N_9338,N_9197);
and U11709 (N_11709,N_8283,N_9815);
nand U11710 (N_11710,N_8829,N_9245);
or U11711 (N_11711,N_8003,N_9260);
or U11712 (N_11712,N_8428,N_9769);
nor U11713 (N_11713,N_9542,N_9258);
xor U11714 (N_11714,N_8483,N_9338);
nor U11715 (N_11715,N_9108,N_8828);
or U11716 (N_11716,N_9864,N_8087);
nor U11717 (N_11717,N_8344,N_9877);
or U11718 (N_11718,N_9633,N_9543);
nor U11719 (N_11719,N_8065,N_9510);
nand U11720 (N_11720,N_9463,N_9831);
nor U11721 (N_11721,N_8922,N_9087);
or U11722 (N_11722,N_8812,N_9667);
or U11723 (N_11723,N_9511,N_9478);
xnor U11724 (N_11724,N_8203,N_9053);
or U11725 (N_11725,N_9738,N_8439);
or U11726 (N_11726,N_9800,N_8520);
nor U11727 (N_11727,N_9742,N_9718);
and U11728 (N_11728,N_9998,N_9940);
and U11729 (N_11729,N_8894,N_9294);
nand U11730 (N_11730,N_8580,N_9827);
nor U11731 (N_11731,N_9727,N_8260);
nand U11732 (N_11732,N_9092,N_8471);
nand U11733 (N_11733,N_9694,N_8603);
or U11734 (N_11734,N_8045,N_8071);
nand U11735 (N_11735,N_9134,N_9262);
nor U11736 (N_11736,N_9870,N_9819);
nor U11737 (N_11737,N_9231,N_8906);
or U11738 (N_11738,N_8691,N_8468);
xor U11739 (N_11739,N_9326,N_8085);
and U11740 (N_11740,N_9758,N_8595);
and U11741 (N_11741,N_9291,N_9575);
and U11742 (N_11742,N_8553,N_9051);
nor U11743 (N_11743,N_8792,N_8085);
and U11744 (N_11744,N_9631,N_8480);
nand U11745 (N_11745,N_9942,N_8775);
nand U11746 (N_11746,N_8060,N_9247);
nand U11747 (N_11747,N_9837,N_9754);
nor U11748 (N_11748,N_9963,N_9806);
and U11749 (N_11749,N_8072,N_8508);
nor U11750 (N_11750,N_9046,N_8560);
and U11751 (N_11751,N_9463,N_8141);
xnor U11752 (N_11752,N_9869,N_9009);
and U11753 (N_11753,N_9951,N_9369);
nor U11754 (N_11754,N_8083,N_8528);
and U11755 (N_11755,N_9936,N_9203);
nand U11756 (N_11756,N_9763,N_9270);
or U11757 (N_11757,N_8352,N_9569);
or U11758 (N_11758,N_9828,N_8880);
nand U11759 (N_11759,N_9474,N_9405);
xnor U11760 (N_11760,N_9648,N_8344);
and U11761 (N_11761,N_8279,N_9776);
or U11762 (N_11762,N_8326,N_9386);
nor U11763 (N_11763,N_9696,N_8518);
or U11764 (N_11764,N_9500,N_8732);
nor U11765 (N_11765,N_9834,N_9059);
and U11766 (N_11766,N_9969,N_9914);
or U11767 (N_11767,N_8312,N_9058);
nand U11768 (N_11768,N_8573,N_8492);
or U11769 (N_11769,N_8328,N_9545);
nor U11770 (N_11770,N_9553,N_9730);
and U11771 (N_11771,N_8805,N_8460);
or U11772 (N_11772,N_9522,N_9021);
nand U11773 (N_11773,N_9889,N_9770);
nand U11774 (N_11774,N_9731,N_8410);
nor U11775 (N_11775,N_9436,N_8252);
and U11776 (N_11776,N_8956,N_8121);
or U11777 (N_11777,N_8697,N_9678);
and U11778 (N_11778,N_9780,N_8779);
nand U11779 (N_11779,N_9689,N_9170);
and U11780 (N_11780,N_8653,N_9769);
or U11781 (N_11781,N_9585,N_8389);
nand U11782 (N_11782,N_9494,N_9340);
nor U11783 (N_11783,N_8533,N_9210);
and U11784 (N_11784,N_9713,N_9671);
nand U11785 (N_11785,N_8352,N_8099);
nand U11786 (N_11786,N_9843,N_8992);
nor U11787 (N_11787,N_9192,N_9189);
xor U11788 (N_11788,N_9521,N_8382);
and U11789 (N_11789,N_8183,N_9081);
nor U11790 (N_11790,N_8148,N_8047);
nand U11791 (N_11791,N_8226,N_8885);
or U11792 (N_11792,N_9940,N_9504);
or U11793 (N_11793,N_8959,N_9442);
and U11794 (N_11794,N_8175,N_8867);
nor U11795 (N_11795,N_9318,N_9376);
nand U11796 (N_11796,N_9309,N_8442);
and U11797 (N_11797,N_9481,N_9299);
nor U11798 (N_11798,N_8822,N_9718);
or U11799 (N_11799,N_8791,N_8984);
or U11800 (N_11800,N_8706,N_8951);
and U11801 (N_11801,N_9813,N_8653);
or U11802 (N_11802,N_9366,N_9249);
or U11803 (N_11803,N_8744,N_9430);
and U11804 (N_11804,N_8089,N_8030);
or U11805 (N_11805,N_8219,N_9083);
nand U11806 (N_11806,N_8328,N_9807);
nand U11807 (N_11807,N_9089,N_8985);
or U11808 (N_11808,N_8276,N_9019);
nand U11809 (N_11809,N_8410,N_8859);
and U11810 (N_11810,N_8020,N_9633);
nor U11811 (N_11811,N_9593,N_9241);
nand U11812 (N_11812,N_8129,N_8142);
nand U11813 (N_11813,N_8893,N_9143);
nand U11814 (N_11814,N_8454,N_9241);
and U11815 (N_11815,N_9243,N_8293);
and U11816 (N_11816,N_9108,N_9189);
nor U11817 (N_11817,N_8679,N_9510);
nor U11818 (N_11818,N_9854,N_9421);
nand U11819 (N_11819,N_8022,N_8835);
nor U11820 (N_11820,N_9461,N_8531);
and U11821 (N_11821,N_8483,N_8863);
nand U11822 (N_11822,N_8114,N_9431);
or U11823 (N_11823,N_9124,N_8015);
nor U11824 (N_11824,N_9032,N_8996);
or U11825 (N_11825,N_8715,N_8672);
or U11826 (N_11826,N_8594,N_9087);
nor U11827 (N_11827,N_9354,N_9258);
nor U11828 (N_11828,N_8183,N_9201);
nor U11829 (N_11829,N_8035,N_8684);
xnor U11830 (N_11830,N_9361,N_8392);
nand U11831 (N_11831,N_8671,N_8928);
nand U11832 (N_11832,N_9663,N_9579);
or U11833 (N_11833,N_8736,N_9424);
or U11834 (N_11834,N_8665,N_9525);
nand U11835 (N_11835,N_8078,N_9830);
nand U11836 (N_11836,N_8715,N_8359);
nor U11837 (N_11837,N_8295,N_8470);
or U11838 (N_11838,N_9692,N_8355);
and U11839 (N_11839,N_8251,N_8783);
nor U11840 (N_11840,N_9437,N_8904);
and U11841 (N_11841,N_9627,N_9805);
or U11842 (N_11842,N_8257,N_8496);
nor U11843 (N_11843,N_8651,N_9491);
or U11844 (N_11844,N_9171,N_9550);
and U11845 (N_11845,N_8882,N_9680);
or U11846 (N_11846,N_9684,N_8898);
or U11847 (N_11847,N_8721,N_8367);
or U11848 (N_11848,N_8450,N_9481);
nand U11849 (N_11849,N_9512,N_9253);
or U11850 (N_11850,N_9187,N_9511);
and U11851 (N_11851,N_8290,N_8925);
or U11852 (N_11852,N_8596,N_8561);
or U11853 (N_11853,N_9708,N_8844);
or U11854 (N_11854,N_9897,N_9028);
nand U11855 (N_11855,N_9258,N_9327);
nand U11856 (N_11856,N_8818,N_9432);
nor U11857 (N_11857,N_9877,N_8022);
or U11858 (N_11858,N_9007,N_9178);
nor U11859 (N_11859,N_9556,N_9598);
or U11860 (N_11860,N_8109,N_8870);
xnor U11861 (N_11861,N_9476,N_8743);
nor U11862 (N_11862,N_9598,N_9372);
and U11863 (N_11863,N_9204,N_9161);
or U11864 (N_11864,N_8910,N_9959);
nor U11865 (N_11865,N_9856,N_8628);
nand U11866 (N_11866,N_9399,N_9045);
nor U11867 (N_11867,N_8914,N_9871);
and U11868 (N_11868,N_9006,N_9152);
nand U11869 (N_11869,N_9051,N_9993);
and U11870 (N_11870,N_8277,N_9411);
nor U11871 (N_11871,N_9815,N_8009);
nand U11872 (N_11872,N_8764,N_9959);
nor U11873 (N_11873,N_9201,N_9022);
nor U11874 (N_11874,N_9950,N_9419);
nor U11875 (N_11875,N_8881,N_9685);
or U11876 (N_11876,N_8355,N_9863);
nand U11877 (N_11877,N_8169,N_8025);
or U11878 (N_11878,N_8709,N_9566);
nor U11879 (N_11879,N_9474,N_8608);
nand U11880 (N_11880,N_8178,N_9949);
nand U11881 (N_11881,N_8795,N_8519);
and U11882 (N_11882,N_9102,N_9079);
and U11883 (N_11883,N_8020,N_9327);
nand U11884 (N_11884,N_9190,N_8090);
nor U11885 (N_11885,N_8911,N_9298);
nor U11886 (N_11886,N_9667,N_8791);
nand U11887 (N_11887,N_8402,N_9932);
nor U11888 (N_11888,N_8371,N_8266);
and U11889 (N_11889,N_8585,N_8834);
or U11890 (N_11890,N_8982,N_9912);
nor U11891 (N_11891,N_9836,N_9430);
and U11892 (N_11892,N_8774,N_8320);
nor U11893 (N_11893,N_8182,N_8328);
nor U11894 (N_11894,N_9766,N_8499);
nor U11895 (N_11895,N_9064,N_9783);
xor U11896 (N_11896,N_9275,N_9745);
nand U11897 (N_11897,N_9827,N_8849);
nand U11898 (N_11898,N_8193,N_8969);
nor U11899 (N_11899,N_8717,N_8284);
and U11900 (N_11900,N_9361,N_8717);
nand U11901 (N_11901,N_9688,N_9289);
and U11902 (N_11902,N_8108,N_8203);
and U11903 (N_11903,N_9188,N_8960);
nor U11904 (N_11904,N_9538,N_9089);
nor U11905 (N_11905,N_9944,N_8399);
nor U11906 (N_11906,N_8981,N_8485);
nand U11907 (N_11907,N_9183,N_8246);
and U11908 (N_11908,N_9570,N_8692);
nand U11909 (N_11909,N_9569,N_8765);
nor U11910 (N_11910,N_8555,N_9510);
nand U11911 (N_11911,N_8109,N_8357);
nand U11912 (N_11912,N_8307,N_8267);
or U11913 (N_11913,N_9989,N_8102);
nor U11914 (N_11914,N_8138,N_9323);
or U11915 (N_11915,N_8021,N_9146);
or U11916 (N_11916,N_8399,N_8647);
nor U11917 (N_11917,N_9432,N_8286);
nand U11918 (N_11918,N_9577,N_8973);
nor U11919 (N_11919,N_8653,N_9315);
nor U11920 (N_11920,N_9241,N_9778);
nand U11921 (N_11921,N_8960,N_9658);
or U11922 (N_11922,N_9633,N_9378);
nand U11923 (N_11923,N_9312,N_9228);
nand U11924 (N_11924,N_9259,N_8672);
or U11925 (N_11925,N_8953,N_9396);
nand U11926 (N_11926,N_8659,N_8385);
or U11927 (N_11927,N_8030,N_9801);
nor U11928 (N_11928,N_9481,N_9515);
nor U11929 (N_11929,N_9783,N_8114);
nand U11930 (N_11930,N_9677,N_8011);
nand U11931 (N_11931,N_8809,N_8576);
xor U11932 (N_11932,N_8524,N_9477);
nand U11933 (N_11933,N_8143,N_9776);
or U11934 (N_11934,N_8196,N_9329);
or U11935 (N_11935,N_9061,N_9494);
and U11936 (N_11936,N_8590,N_8307);
xor U11937 (N_11937,N_8794,N_8058);
nand U11938 (N_11938,N_8296,N_9301);
nor U11939 (N_11939,N_8862,N_8963);
or U11940 (N_11940,N_8865,N_8268);
nor U11941 (N_11941,N_9635,N_8483);
nand U11942 (N_11942,N_9176,N_9867);
and U11943 (N_11943,N_8888,N_9713);
and U11944 (N_11944,N_8706,N_8176);
nor U11945 (N_11945,N_9253,N_8644);
and U11946 (N_11946,N_9307,N_9316);
or U11947 (N_11947,N_9201,N_9398);
nand U11948 (N_11948,N_8499,N_8783);
nor U11949 (N_11949,N_8285,N_9665);
or U11950 (N_11950,N_8551,N_9337);
nor U11951 (N_11951,N_9909,N_9148);
and U11952 (N_11952,N_9165,N_8160);
nor U11953 (N_11953,N_8840,N_9914);
nor U11954 (N_11954,N_9976,N_8443);
or U11955 (N_11955,N_8287,N_9654);
or U11956 (N_11956,N_9870,N_8046);
nor U11957 (N_11957,N_9158,N_9541);
nand U11958 (N_11958,N_9599,N_9789);
nand U11959 (N_11959,N_8194,N_9507);
and U11960 (N_11960,N_8449,N_9460);
nand U11961 (N_11961,N_9874,N_8253);
nor U11962 (N_11962,N_8977,N_8353);
nand U11963 (N_11963,N_9672,N_8549);
and U11964 (N_11964,N_8154,N_8072);
nand U11965 (N_11965,N_8147,N_9457);
and U11966 (N_11966,N_8863,N_9712);
and U11967 (N_11967,N_8141,N_8495);
nand U11968 (N_11968,N_8152,N_8147);
nor U11969 (N_11969,N_9526,N_8474);
nand U11970 (N_11970,N_8225,N_8495);
or U11971 (N_11971,N_9187,N_8043);
nand U11972 (N_11972,N_9501,N_9378);
nand U11973 (N_11973,N_8922,N_9298);
nand U11974 (N_11974,N_8692,N_8107);
nand U11975 (N_11975,N_9267,N_9799);
nor U11976 (N_11976,N_9106,N_8700);
and U11977 (N_11977,N_9165,N_8162);
nor U11978 (N_11978,N_8112,N_8987);
or U11979 (N_11979,N_9127,N_8788);
and U11980 (N_11980,N_8483,N_9892);
xor U11981 (N_11981,N_8622,N_9066);
nand U11982 (N_11982,N_9147,N_8397);
nand U11983 (N_11983,N_8251,N_9289);
nor U11984 (N_11984,N_9374,N_8033);
nand U11985 (N_11985,N_9402,N_8266);
and U11986 (N_11986,N_9660,N_9347);
or U11987 (N_11987,N_8049,N_9000);
nor U11988 (N_11988,N_8045,N_9346);
nand U11989 (N_11989,N_9704,N_8179);
nor U11990 (N_11990,N_9294,N_9174);
or U11991 (N_11991,N_8568,N_8210);
and U11992 (N_11992,N_9105,N_9424);
or U11993 (N_11993,N_8655,N_8121);
nand U11994 (N_11994,N_9371,N_8639);
nand U11995 (N_11995,N_8666,N_9994);
or U11996 (N_11996,N_9198,N_8549);
nand U11997 (N_11997,N_9641,N_8912);
and U11998 (N_11998,N_9091,N_8383);
nor U11999 (N_11999,N_8773,N_9542);
and U12000 (N_12000,N_10421,N_11114);
nand U12001 (N_12001,N_11335,N_10399);
nand U12002 (N_12002,N_10580,N_11530);
nand U12003 (N_12003,N_11087,N_10402);
and U12004 (N_12004,N_10117,N_11359);
or U12005 (N_12005,N_10742,N_10539);
nor U12006 (N_12006,N_10926,N_10959);
nand U12007 (N_12007,N_11216,N_10335);
nor U12008 (N_12008,N_10861,N_11863);
nor U12009 (N_12009,N_10893,N_10288);
nor U12010 (N_12010,N_10990,N_10397);
or U12011 (N_12011,N_11090,N_10406);
or U12012 (N_12012,N_11173,N_11205);
or U12013 (N_12013,N_11720,N_10383);
nand U12014 (N_12014,N_11996,N_11204);
nor U12015 (N_12015,N_10216,N_10964);
or U12016 (N_12016,N_10871,N_11059);
nor U12017 (N_12017,N_10394,N_11372);
or U12018 (N_12018,N_10497,N_10681);
nand U12019 (N_12019,N_10760,N_10365);
or U12020 (N_12020,N_11185,N_10070);
and U12021 (N_12021,N_11903,N_11086);
or U12022 (N_12022,N_10481,N_11180);
nor U12023 (N_12023,N_11941,N_11077);
nand U12024 (N_12024,N_10354,N_10584);
and U12025 (N_12025,N_10029,N_10548);
and U12026 (N_12026,N_11223,N_10302);
nor U12027 (N_12027,N_11315,N_11931);
xor U12028 (N_12028,N_11892,N_11573);
and U12029 (N_12029,N_11475,N_10100);
xnor U12030 (N_12030,N_10518,N_10195);
nand U12031 (N_12031,N_10453,N_11688);
nor U12032 (N_12032,N_11306,N_10155);
nand U12033 (N_12033,N_11511,N_10276);
nand U12034 (N_12034,N_11968,N_10695);
nor U12035 (N_12035,N_11734,N_11435);
nor U12036 (N_12036,N_10436,N_10300);
nand U12037 (N_12037,N_11648,N_10368);
nor U12038 (N_12038,N_11851,N_11444);
nand U12039 (N_12039,N_11091,N_11261);
nor U12040 (N_12040,N_10054,N_10933);
and U12041 (N_12041,N_11760,N_11112);
or U12042 (N_12042,N_10465,N_11754);
or U12043 (N_12043,N_11778,N_10839);
nand U12044 (N_12044,N_11055,N_11982);
nor U12045 (N_12045,N_11886,N_10720);
nor U12046 (N_12046,N_11066,N_11767);
and U12047 (N_12047,N_10133,N_11225);
and U12048 (N_12048,N_11808,N_11345);
nor U12049 (N_12049,N_10255,N_11942);
or U12050 (N_12050,N_11713,N_11743);
or U12051 (N_12051,N_11884,N_11784);
and U12052 (N_12052,N_11718,N_10488);
or U12053 (N_12053,N_11485,N_11780);
and U12054 (N_12054,N_10388,N_11307);
nand U12055 (N_12055,N_11826,N_11341);
nand U12056 (N_12056,N_10956,N_10244);
nor U12057 (N_12057,N_10050,N_10937);
nand U12058 (N_12058,N_11227,N_10150);
xnor U12059 (N_12059,N_11280,N_10200);
or U12060 (N_12060,N_11993,N_10526);
nor U12061 (N_12061,N_11134,N_11148);
and U12062 (N_12062,N_11074,N_10568);
and U12063 (N_12063,N_11505,N_10899);
nor U12064 (N_12064,N_11995,N_10743);
nand U12065 (N_12065,N_11606,N_11024);
nand U12066 (N_12066,N_11735,N_10895);
nand U12067 (N_12067,N_11336,N_10813);
nand U12068 (N_12068,N_10866,N_10361);
nand U12069 (N_12069,N_10753,N_11698);
nand U12070 (N_12070,N_11789,N_11834);
nand U12071 (N_12071,N_11636,N_10787);
nor U12072 (N_12072,N_11226,N_11552);
or U12073 (N_12073,N_10843,N_10545);
nor U12074 (N_12074,N_11289,N_11192);
or U12075 (N_12075,N_11531,N_10731);
nand U12076 (N_12076,N_11125,N_10903);
or U12077 (N_12077,N_10344,N_11326);
xnor U12078 (N_12078,N_10459,N_10651);
nor U12079 (N_12079,N_11130,N_11150);
nor U12080 (N_12080,N_11169,N_10454);
nor U12081 (N_12081,N_11702,N_11913);
nand U12082 (N_12082,N_10359,N_10826);
and U12083 (N_12083,N_10746,N_10706);
or U12084 (N_12084,N_11540,N_11681);
nor U12085 (N_12085,N_11076,N_10414);
or U12086 (N_12086,N_10696,N_11620);
nand U12087 (N_12087,N_11154,N_11382);
nor U12088 (N_12088,N_10233,N_11450);
or U12089 (N_12089,N_10318,N_11253);
nor U12090 (N_12090,N_10814,N_11664);
nand U12091 (N_12091,N_11439,N_11512);
or U12092 (N_12092,N_11237,N_10218);
nor U12093 (N_12093,N_10366,N_11574);
nand U12094 (N_12094,N_11680,N_11413);
and U12095 (N_12095,N_10677,N_11750);
nor U12096 (N_12096,N_11295,N_10351);
nand U12097 (N_12097,N_10081,N_11111);
or U12098 (N_12098,N_11627,N_11194);
nor U12099 (N_12099,N_10786,N_10337);
nand U12100 (N_12100,N_10563,N_10800);
and U12101 (N_12101,N_11417,N_11717);
or U12102 (N_12102,N_10653,N_10795);
and U12103 (N_12103,N_11765,N_11557);
and U12104 (N_12104,N_11605,N_10438);
nor U12105 (N_12105,N_11611,N_10664);
nand U12106 (N_12106,N_11323,N_11166);
nand U12107 (N_12107,N_10562,N_10428);
and U12108 (N_12108,N_10327,N_11570);
nor U12109 (N_12109,N_10816,N_11314);
and U12110 (N_12110,N_11534,N_11036);
or U12111 (N_12111,N_11412,N_11679);
nor U12112 (N_12112,N_10201,N_10080);
and U12113 (N_12113,N_10501,N_10729);
nand U12114 (N_12114,N_11022,N_10531);
and U12115 (N_12115,N_11415,N_10794);
or U12116 (N_12116,N_10851,N_10067);
nand U12117 (N_12117,N_10122,N_11838);
nor U12118 (N_12118,N_10870,N_10745);
or U12119 (N_12119,N_11133,N_11096);
or U12120 (N_12120,N_11689,N_11906);
or U12121 (N_12121,N_10246,N_10534);
and U12122 (N_12122,N_10551,N_10688);
or U12123 (N_12123,N_10510,N_11308);
nor U12124 (N_12124,N_11310,N_11935);
and U12125 (N_12125,N_11350,N_11771);
nand U12126 (N_12126,N_10308,N_10311);
nand U12127 (N_12127,N_10111,N_11468);
nand U12128 (N_12128,N_11398,N_11354);
nand U12129 (N_12129,N_11438,N_10400);
xnor U12130 (N_12130,N_10151,N_11160);
and U12131 (N_12131,N_10396,N_10472);
nor U12132 (N_12132,N_10035,N_11646);
nor U12133 (N_12133,N_10247,N_11951);
and U12134 (N_12134,N_10158,N_11217);
or U12135 (N_12135,N_11487,N_11161);
or U12136 (N_12136,N_10214,N_11203);
nand U12137 (N_12137,N_10382,N_11830);
nand U12138 (N_12138,N_10022,N_10818);
or U12139 (N_12139,N_10528,N_11948);
or U12140 (N_12140,N_11793,N_11279);
nand U12141 (N_12141,N_10102,N_11476);
or U12142 (N_12142,N_10734,N_10628);
nand U12143 (N_12143,N_10636,N_11883);
nand U12144 (N_12144,N_11190,N_11156);
or U12145 (N_12145,N_11955,N_10928);
nand U12146 (N_12146,N_11482,N_10170);
nor U12147 (N_12147,N_11922,N_11973);
nand U12148 (N_12148,N_11019,N_10455);
nand U12149 (N_12149,N_10362,N_11893);
nand U12150 (N_12150,N_10504,N_11804);
and U12151 (N_12151,N_10264,N_11252);
or U12152 (N_12152,N_10585,N_10689);
and U12153 (N_12153,N_10773,N_10521);
nand U12154 (N_12154,N_10714,N_10242);
nor U12155 (N_12155,N_10867,N_10401);
nand U12156 (N_12156,N_10467,N_10908);
nand U12157 (N_12157,N_10916,N_11556);
or U12158 (N_12158,N_10817,N_10702);
and U12159 (N_12159,N_11048,N_11954);
nor U12160 (N_12160,N_10458,N_11590);
xor U12161 (N_12161,N_10630,N_10144);
nor U12162 (N_12162,N_11604,N_10983);
or U12163 (N_12163,N_10321,N_11763);
and U12164 (N_12164,N_10086,N_11854);
xor U12165 (N_12165,N_11183,N_10415);
or U12166 (N_12166,N_11017,N_11168);
nor U12167 (N_12167,N_11891,N_11871);
nor U12168 (N_12168,N_11456,N_11393);
and U12169 (N_12169,N_10046,N_11933);
and U12170 (N_12170,N_10197,N_11785);
or U12171 (N_12171,N_11146,N_10148);
nor U12172 (N_12172,N_10125,N_11554);
nand U12173 (N_12173,N_11281,N_10199);
or U12174 (N_12174,N_11843,N_11312);
and U12175 (N_12175,N_11369,N_10113);
or U12176 (N_12176,N_11016,N_10483);
nand U12177 (N_12177,N_10608,N_10345);
nor U12178 (N_12178,N_11696,N_10373);
nand U12179 (N_12179,N_10303,N_10614);
nor U12180 (N_12180,N_10680,N_11305);
or U12181 (N_12181,N_11008,N_11837);
nand U12182 (N_12182,N_10516,N_11430);
and U12183 (N_12183,N_11943,N_11418);
nor U12184 (N_12184,N_11266,N_11657);
nor U12185 (N_12185,N_11725,N_11451);
and U12186 (N_12186,N_10206,N_11244);
and U12187 (N_12187,N_10685,N_11918);
nand U12188 (N_12188,N_10257,N_11078);
and U12189 (N_12189,N_10727,N_10938);
nor U12190 (N_12190,N_10805,N_11764);
and U12191 (N_12191,N_10767,N_11104);
or U12192 (N_12192,N_11953,N_10434);
xor U12193 (N_12193,N_11729,N_11011);
nor U12194 (N_12194,N_10776,N_10897);
nor U12195 (N_12195,N_10385,N_10073);
or U12196 (N_12196,N_11959,N_10540);
or U12197 (N_12197,N_10477,N_11069);
nor U12198 (N_12198,N_10587,N_11427);
and U12199 (N_12199,N_10644,N_10726);
and U12200 (N_12200,N_10157,N_10326);
nor U12201 (N_12201,N_11902,N_10060);
nor U12202 (N_12202,N_10593,N_10781);
nor U12203 (N_12203,N_10972,N_10995);
nor U12204 (N_12204,N_11888,N_11984);
or U12205 (N_12205,N_11113,N_10053);
or U12206 (N_12206,N_11120,N_10942);
or U12207 (N_12207,N_10845,N_10811);
nand U12208 (N_12208,N_11632,N_11821);
nand U12209 (N_12209,N_10907,N_10156);
and U12210 (N_12210,N_11617,N_11142);
nand U12211 (N_12211,N_11442,N_10292);
or U12212 (N_12212,N_11988,N_10687);
and U12213 (N_12213,N_11409,N_11386);
or U12214 (N_12214,N_10324,N_11625);
and U12215 (N_12215,N_10582,N_11367);
or U12216 (N_12216,N_10087,N_10166);
or U12217 (N_12217,N_10227,N_10096);
or U12218 (N_12218,N_10290,N_10709);
nor U12219 (N_12219,N_10852,N_10850);
or U12220 (N_12220,N_10656,N_10116);
nand U12221 (N_12221,N_10572,N_11517);
nand U12222 (N_12222,N_10014,N_10878);
nand U12223 (N_12223,N_10953,N_10294);
or U12224 (N_12224,N_11296,N_10089);
nor U12225 (N_12225,N_10405,N_10509);
and U12226 (N_12226,N_10925,N_11188);
nor U12227 (N_12227,N_10131,N_11493);
and U12228 (N_12228,N_10554,N_10508);
nand U12229 (N_12229,N_10039,N_10287);
or U12230 (N_12230,N_11304,N_10063);
or U12231 (N_12231,N_11603,N_11164);
nor U12232 (N_12232,N_10493,N_11915);
nand U12233 (N_12233,N_11135,N_11563);
nor U12234 (N_12234,N_11292,N_10639);
and U12235 (N_12235,N_11000,N_10619);
and U12236 (N_12236,N_11018,N_10530);
nor U12237 (N_12237,N_11577,N_11855);
and U12238 (N_12238,N_11660,N_11381);
nand U12239 (N_12239,N_10809,N_11236);
or U12240 (N_12240,N_11348,N_10595);
nand U12241 (N_12241,N_11368,N_11579);
nand U12242 (N_12242,N_10765,N_11123);
xnor U12243 (N_12243,N_10523,N_10346);
nor U12244 (N_12244,N_10419,N_11794);
nand U12245 (N_12245,N_11157,N_10473);
nor U12246 (N_12246,N_11388,N_11737);
or U12247 (N_12247,N_10708,N_10299);
and U12248 (N_12248,N_11116,N_11218);
nand U12249 (N_12249,N_10307,N_10996);
xor U12250 (N_12250,N_11596,N_11525);
or U12251 (N_12251,N_11961,N_11259);
and U12252 (N_12252,N_10954,N_10737);
or U12253 (N_12253,N_10097,N_10234);
xnor U12254 (N_12254,N_10496,N_10934);
nand U12255 (N_12255,N_11582,N_11355);
nor U12256 (N_12256,N_10441,N_11506);
and U12257 (N_12257,N_11706,N_10012);
and U12258 (N_12258,N_11652,N_11520);
nor U12259 (N_12259,N_11469,N_10258);
nand U12260 (N_12260,N_11273,N_10126);
nand U12261 (N_12261,N_11700,N_10780);
nand U12262 (N_12262,N_11044,N_11728);
nand U12263 (N_12263,N_11630,N_10298);
nor U12264 (N_12264,N_11424,N_10537);
nor U12265 (N_12265,N_11472,N_10389);
nor U12266 (N_12266,N_11337,N_11149);
or U12267 (N_12267,N_11846,N_10490);
nand U12268 (N_12268,N_11907,N_11283);
or U12269 (N_12269,N_10789,N_11569);
nand U12270 (N_12270,N_11219,N_10034);
xor U12271 (N_12271,N_10755,N_10691);
nand U12272 (N_12272,N_11053,N_10372);
nand U12273 (N_12273,N_11299,N_11495);
nor U12274 (N_12274,N_10464,N_11587);
nor U12275 (N_12275,N_11802,N_11333);
nor U12276 (N_12276,N_11956,N_11352);
nor U12277 (N_12277,N_11581,N_10770);
nand U12278 (N_12278,N_10295,N_10576);
or U12279 (N_12279,N_10285,N_11421);
and U12280 (N_12280,N_10812,N_10301);
and U12281 (N_12281,N_10910,N_11994);
nand U12282 (N_12282,N_10074,N_11795);
and U12283 (N_12283,N_11980,N_11153);
and U12284 (N_12284,N_10044,N_10643);
nor U12285 (N_12285,N_10169,N_11516);
nand U12286 (N_12286,N_10558,N_11730);
nor U12287 (N_12287,N_10503,N_10618);
nor U12288 (N_12288,N_10579,N_11536);
and U12289 (N_12289,N_11758,N_10777);
or U12290 (N_12290,N_10316,N_10352);
nor U12291 (N_12291,N_10417,N_11810);
or U12292 (N_12292,N_11641,N_10710);
or U12293 (N_12293,N_10976,N_11642);
and U12294 (N_12294,N_10546,N_11356);
nor U12295 (N_12295,N_10693,N_10446);
nand U12296 (N_12296,N_11101,N_11544);
and U12297 (N_12297,N_10888,N_10448);
or U12298 (N_12298,N_11309,N_10048);
nand U12299 (N_12299,N_11080,N_10810);
and U12300 (N_12300,N_11610,N_11110);
or U12301 (N_12301,N_10469,N_11715);
and U12302 (N_12302,N_10457,N_10055);
nor U12303 (N_12303,N_10164,N_11478);
and U12304 (N_12304,N_11499,N_11429);
nor U12305 (N_12305,N_11274,N_11151);
nand U12306 (N_12306,N_10802,N_10369);
and U12307 (N_12307,N_10317,N_10224);
and U12308 (N_12308,N_10191,N_10426);
nor U12309 (N_12309,N_10815,N_11193);
nand U12310 (N_12310,N_11028,N_10784);
and U12311 (N_12311,N_11565,N_10482);
or U12312 (N_12312,N_10274,N_10004);
or U12313 (N_12313,N_10603,N_10371);
and U12314 (N_12314,N_10970,N_11425);
nand U12315 (N_12315,N_10758,N_11402);
nor U12316 (N_12316,N_10842,N_11209);
and U12317 (N_12317,N_10314,N_11376);
and U12318 (N_12318,N_10898,N_11782);
or U12319 (N_12319,N_10532,N_10424);
nand U12320 (N_12320,N_10355,N_10202);
or U12321 (N_12321,N_10387,N_11502);
and U12322 (N_12322,N_10350,N_11242);
nor U12323 (N_12323,N_11944,N_11118);
nand U12324 (N_12324,N_10820,N_11288);
and U12325 (N_12325,N_10284,N_10684);
or U12326 (N_12326,N_11766,N_11026);
nand U12327 (N_12327,N_10890,N_11256);
or U12328 (N_12328,N_10862,N_10975);
or U12329 (N_12329,N_10273,N_10272);
or U12330 (N_12330,N_11033,N_10750);
or U12331 (N_12331,N_10764,N_10236);
or U12332 (N_12332,N_10922,N_10343);
or U12333 (N_12333,N_10184,N_10931);
nand U12334 (N_12334,N_11532,N_10322);
or U12335 (N_12335,N_10038,N_10556);
or U12336 (N_12336,N_11805,N_11929);
nor U12337 (N_12337,N_10023,N_11873);
nor U12338 (N_12338,N_11881,N_10007);
nor U12339 (N_12339,N_10875,N_10120);
and U12340 (N_12340,N_11523,N_11676);
or U12341 (N_12341,N_10849,N_10935);
or U12342 (N_12342,N_10543,N_10686);
and U12343 (N_12343,N_11045,N_10189);
nor U12344 (N_12344,N_10422,N_10574);
and U12345 (N_12345,N_11089,N_10822);
and U12346 (N_12346,N_10803,N_11885);
or U12347 (N_12347,N_11370,N_11790);
or U12348 (N_12348,N_10863,N_11809);
nand U12349 (N_12349,N_10932,N_10586);
or U12350 (N_12350,N_10884,N_10330);
or U12351 (N_12351,N_11270,N_11900);
or U12352 (N_12352,N_11375,N_10183);
nor U12353 (N_12353,N_10245,N_10177);
and U12354 (N_12354,N_11612,N_11938);
nor U12355 (N_12355,N_10635,N_10571);
nand U12356 (N_12356,N_11138,N_10228);
or U12357 (N_12357,N_11965,N_11119);
nand U12358 (N_12358,N_10549,N_10615);
or U12359 (N_12359,N_11094,N_10188);
and U12360 (N_12360,N_10876,N_11990);
nor U12361 (N_12361,N_11063,N_10381);
nor U12362 (N_12362,N_11962,N_10944);
xnor U12363 (N_12363,N_10790,N_11248);
and U12364 (N_12364,N_10957,N_10621);
nand U12365 (N_12365,N_10027,N_10160);
or U12366 (N_12366,N_10041,N_11374);
or U12367 (N_12367,N_10559,N_10847);
and U12368 (N_12368,N_11344,N_10775);
or U12369 (N_12369,N_10315,N_11551);
and U12370 (N_12370,N_10313,N_10210);
nor U12371 (N_12371,N_11377,N_11445);
nor U12372 (N_12372,N_10238,N_11054);
or U12373 (N_12373,N_10834,N_11986);
or U12374 (N_12374,N_10037,N_10798);
or U12375 (N_12375,N_11957,N_10178);
nand U12376 (N_12376,N_10032,N_11342);
nand U12377 (N_12377,N_10143,N_10139);
nor U12378 (N_12378,N_11391,N_11392);
nand U12379 (N_12379,N_11820,N_10506);
nor U12380 (N_12380,N_11842,N_11924);
nand U12381 (N_12381,N_11548,N_10069);
nor U12382 (N_12382,N_11145,N_11201);
or U12383 (N_12383,N_10253,N_11452);
nand U12384 (N_12384,N_11631,N_10989);
and U12385 (N_12385,N_11433,N_11492);
nand U12386 (N_12386,N_10066,N_11067);
nor U12387 (N_12387,N_10565,N_11365);
nand U12388 (N_12388,N_10877,N_10952);
or U12389 (N_12389,N_10728,N_11167);
nor U12390 (N_12390,N_10252,N_10168);
nor U12391 (N_12391,N_10152,N_10768);
nand U12392 (N_12392,N_11539,N_10704);
nor U12393 (N_12393,N_11916,N_11158);
nor U12394 (N_12394,N_10511,N_10736);
and U12395 (N_12395,N_11300,N_10924);
or U12396 (N_12396,N_10021,N_11003);
nand U12397 (N_12397,N_10588,N_11521);
nand U12398 (N_12398,N_10914,N_11635);
or U12399 (N_12399,N_11298,N_11747);
and U12400 (N_12400,N_11649,N_10655);
and U12401 (N_12401,N_10672,N_11231);
nor U12402 (N_12402,N_10207,N_10240);
and U12403 (N_12403,N_10219,N_10075);
nand U12404 (N_12404,N_11165,N_10403);
nor U12405 (N_12405,N_11437,N_11362);
nand U12406 (N_12406,N_11085,N_11419);
nand U12407 (N_12407,N_10262,N_11012);
or U12408 (N_12408,N_10963,N_10320);
and U12409 (N_12409,N_10536,N_10378);
xor U12410 (N_12410,N_11775,N_11013);
or U12411 (N_12411,N_10339,N_11673);
nand U12412 (N_12412,N_11501,N_11366);
or U12413 (N_12413,N_11286,N_11526);
nor U12414 (N_12414,N_11360,N_10648);
and U12415 (N_12415,N_11117,N_11302);
nand U12416 (N_12416,N_10654,N_11489);
nor U12417 (N_12417,N_11602,N_11447);
xor U12418 (N_12418,N_10529,N_11106);
nor U12419 (N_12419,N_10918,N_10443);
nand U12420 (N_12420,N_11220,N_11056);
and U12421 (N_12421,N_10872,N_11853);
and U12422 (N_12422,N_11755,N_10724);
or U12423 (N_12423,N_11509,N_11697);
nand U12424 (N_12424,N_10592,N_10968);
nand U12425 (N_12425,N_11245,N_11249);
and U12426 (N_12426,N_10716,N_10725);
and U12427 (N_12427,N_10541,N_10281);
or U12428 (N_12428,N_11930,N_10987);
nor U12429 (N_12429,N_10208,N_10717);
nand U12430 (N_12430,N_10293,N_11932);
and U12431 (N_12431,N_10106,N_11952);
nand U12432 (N_12432,N_10788,N_10025);
and U12433 (N_12433,N_11254,N_10071);
nand U12434 (N_12434,N_11723,N_10873);
and U12435 (N_12435,N_11172,N_10544);
nor U12436 (N_12436,N_11504,N_10967);
or U12437 (N_12437,N_10675,N_11633);
xnor U12438 (N_12438,N_10594,N_11558);
nand U12439 (N_12439,N_10832,N_11974);
and U12440 (N_12440,N_11265,N_11542);
nand U12441 (N_12441,N_11025,N_10431);
nor U12442 (N_12442,N_11537,N_11757);
or U12443 (N_12443,N_10880,N_10833);
or U12444 (N_12444,N_11410,N_11692);
nand U12445 (N_12445,N_11037,N_10666);
nand U12446 (N_12446,N_11773,N_10182);
nand U12447 (N_12447,N_11650,N_11126);
and U12448 (N_12448,N_10637,N_10147);
and U12449 (N_12449,N_11997,N_10190);
or U12450 (N_12450,N_11816,N_11945);
or U12451 (N_12451,N_10209,N_10740);
nand U12452 (N_12452,N_11867,N_10982);
or U12453 (N_12453,N_11978,N_10946);
nor U12454 (N_12454,N_11030,N_11446);
or U12455 (N_12455,N_10744,N_11890);
and U12456 (N_12456,N_10674,N_10420);
and U12457 (N_12457,N_11599,N_10567);
and U12458 (N_12458,N_10825,N_10485);
nand U12459 (N_12459,N_11494,N_10663);
xnor U12460 (N_12460,N_11670,N_11759);
and U12461 (N_12461,N_10423,N_10163);
nand U12462 (N_12462,N_11600,N_11966);
xor U12463 (N_12463,N_10923,N_11208);
or U12464 (N_12464,N_10578,N_11832);
nor U12465 (N_12465,N_10408,N_11390);
nor U12466 (N_12466,N_11198,N_11562);
or U12467 (N_12467,N_11703,N_11833);
nor U12468 (N_12468,N_10703,N_11290);
or U12469 (N_12469,N_10599,N_11975);
or U12470 (N_12470,N_11958,N_10757);
nor U12471 (N_12471,N_11460,N_11841);
nand U12472 (N_12472,N_10785,N_11082);
nor U12473 (N_12473,N_11385,N_10077);
and U12474 (N_12474,N_11184,N_10965);
and U12475 (N_12475,N_10447,N_11839);
nand U12476 (N_12476,N_11960,N_11812);
xor U12477 (N_12477,N_11009,N_11541);
and U12478 (N_12478,N_10064,N_10006);
or U12479 (N_12479,N_11406,N_11007);
nor U12480 (N_12480,N_10364,N_11250);
nor U12481 (N_12481,N_11387,N_11181);
nand U12482 (N_12482,N_11872,N_10347);
nand U12483 (N_12483,N_11311,N_11238);
and U12484 (N_12484,N_10517,N_10229);
xor U12485 (N_12485,N_11422,N_10193);
nand U12486 (N_12486,N_10623,N_11864);
nor U12487 (N_12487,N_11695,N_11050);
nor U12488 (N_12488,N_11405,N_11338);
nand U12489 (N_12489,N_10409,N_10243);
or U12490 (N_12490,N_11099,N_10642);
or U12491 (N_12491,N_10205,N_11847);
and U12492 (N_12492,N_11484,N_11155);
nand U12493 (N_12493,N_11233,N_11745);
nand U12494 (N_12494,N_11940,N_10484);
nand U12495 (N_12495,N_11860,N_10103);
and U12496 (N_12496,N_10992,N_11132);
nor U12497 (N_12497,N_11399,N_10604);
or U12498 (N_12498,N_10011,N_11187);
nor U12499 (N_12499,N_10124,N_10449);
nor U12500 (N_12500,N_11224,N_11701);
and U12501 (N_12501,N_10348,N_11353);
and U12502 (N_12502,N_11939,N_11685);
nand U12503 (N_12503,N_11403,N_11034);
or U12504 (N_12504,N_10110,N_10913);
or U12505 (N_12505,N_11584,N_10984);
nand U12506 (N_12506,N_10641,N_11210);
nor U12507 (N_12507,N_10804,N_10591);
nor U12508 (N_12508,N_10297,N_11787);
and U12509 (N_12509,N_10991,N_10864);
or U12510 (N_12510,N_11672,N_10036);
nand U12511 (N_12511,N_10042,N_11878);
nand U12512 (N_12512,N_11457,N_11691);
and U12513 (N_12513,N_11733,N_11171);
and U12514 (N_12514,N_10682,N_10017);
nand U12515 (N_12515,N_11144,N_11449);
or U12516 (N_12516,N_11093,N_10429);
nand U12517 (N_12517,N_11947,N_10679);
and U12518 (N_12518,N_10665,N_10392);
nor U12519 (N_12519,N_10263,N_10659);
and U12520 (N_12520,N_10917,N_10001);
or U12521 (N_12521,N_11322,N_11711);
or U12522 (N_12522,N_10280,N_10270);
or U12523 (N_12523,N_11615,N_11919);
or U12524 (N_12524,N_10332,N_10002);
nand U12525 (N_12525,N_10705,N_10404);
and U12526 (N_12526,N_10460,N_11127);
nor U12527 (N_12527,N_11443,N_11396);
or U12528 (N_12528,N_10766,N_11844);
nand U12529 (N_12529,N_11608,N_10052);
nand U12530 (N_12530,N_10265,N_10363);
or U12531 (N_12531,N_11675,N_10222);
nor U12532 (N_12532,N_10829,N_11378);
and U12533 (N_12533,N_10698,N_11719);
nand U12534 (N_12534,N_10719,N_10966);
or U12535 (N_12535,N_10256,N_10225);
nor U12536 (N_12536,N_10629,N_11477);
nor U12537 (N_12537,N_10735,N_11057);
and U12538 (N_12538,N_10853,N_10821);
nand U12539 (N_12539,N_11666,N_10090);
nand U12540 (N_12540,N_11972,N_11420);
or U12541 (N_12541,N_11580,N_10930);
or U12542 (N_12542,N_10779,N_10215);
and U12543 (N_12543,N_11423,N_11967);
and U12544 (N_12544,N_10980,N_10250);
nor U12545 (N_12545,N_10478,N_10323);
xor U12546 (N_12546,N_11320,N_11108);
and U12547 (N_12547,N_10527,N_10159);
nor U12548 (N_12548,N_11683,N_10231);
and U12549 (N_12549,N_10739,N_11065);
nor U12550 (N_12550,N_11428,N_10505);
nor U12551 (N_12551,N_10939,N_10997);
nor U12552 (N_12552,N_11411,N_11467);
nand U12553 (N_12553,N_11490,N_10699);
and U12554 (N_12554,N_10919,N_10911);
nor U12555 (N_12555,N_11277,N_11800);
nand U12556 (N_12556,N_10783,N_10386);
nor U12557 (N_12557,N_11936,N_11928);
nor U12558 (N_12558,N_10683,N_10678);
nor U12559 (N_12559,N_10756,N_11107);
and U12560 (N_12560,N_11591,N_11147);
and U12561 (N_12561,N_11303,N_10226);
or U12562 (N_12562,N_10439,N_11278);
nand U12563 (N_12563,N_10487,N_11176);
xnor U12564 (N_12564,N_11213,N_10198);
or U12565 (N_12565,N_11682,N_11197);
nor U12566 (N_12566,N_11232,N_11538);
nand U12567 (N_12567,N_10092,N_11578);
nor U12568 (N_12568,N_10566,N_11098);
nand U12569 (N_12569,N_11693,N_11079);
and U12570 (N_12570,N_11550,N_10083);
and U12571 (N_12571,N_11006,N_11749);
and U12572 (N_12572,N_11199,N_10161);
or U12573 (N_12573,N_10652,N_11870);
or U12574 (N_12574,N_11561,N_11647);
or U12575 (N_12575,N_10988,N_11251);
or U12576 (N_12576,N_10831,N_10435);
nand U12577 (N_12577,N_11051,N_11638);
xnor U12578 (N_12578,N_11607,N_11257);
nand U12579 (N_12579,N_10416,N_11704);
nor U12580 (N_12580,N_10486,N_10432);
nor U12581 (N_12581,N_10223,N_11408);
and U12582 (N_12582,N_11555,N_11985);
nand U12583 (N_12583,N_11268,N_10374);
and U12584 (N_12584,N_11513,N_11849);
nand U12585 (N_12585,N_11895,N_10154);
or U12586 (N_12586,N_11897,N_11178);
and U12587 (N_12587,N_10393,N_10310);
xor U12588 (N_12588,N_10752,N_10146);
nor U12589 (N_12589,N_11340,N_11207);
xor U12590 (N_12590,N_10412,N_11215);
and U12591 (N_12591,N_11777,N_10627);
xor U12592 (N_12592,N_11364,N_10577);
xor U12593 (N_12593,N_10634,N_11246);
and U12594 (N_12594,N_11927,N_10016);
nand U12595 (N_12595,N_10093,N_11708);
or U12596 (N_12596,N_10806,N_10974);
or U12597 (N_12597,N_10261,N_10552);
and U12598 (N_12598,N_10512,N_10379);
nand U12599 (N_12599,N_10879,N_11015);
nand U12600 (N_12600,N_11979,N_11568);
nand U12601 (N_12601,N_11357,N_11686);
and U12602 (N_12602,N_11609,N_11170);
nor U12603 (N_12603,N_11141,N_11038);
xor U12604 (N_12604,N_10305,N_10462);
or U12605 (N_12605,N_10172,N_10936);
or U12606 (N_12606,N_10519,N_10370);
nor U12607 (N_12607,N_10165,N_11061);
xnor U12608 (N_12608,N_11002,N_11819);
nand U12609 (N_12609,N_11035,N_11243);
or U12610 (N_12610,N_11920,N_11619);
and U12611 (N_12611,N_11262,N_11815);
or U12612 (N_12612,N_11799,N_11291);
nand U12613 (N_12613,N_10841,N_11371);
nand U12614 (N_12614,N_11572,N_10241);
nand U12615 (N_12615,N_10865,N_10277);
or U12616 (N_12616,N_11546,N_10993);
nand U12617 (N_12617,N_11879,N_10221);
nand U12618 (N_12618,N_11200,N_11926);
nor U12619 (N_12619,N_11383,N_11182);
nand U12620 (N_12620,N_10945,N_11914);
nor U12621 (N_12621,N_10555,N_11507);
or U12622 (N_12622,N_11005,N_11852);
and U12623 (N_12623,N_11159,N_10542);
nor U12624 (N_12624,N_11571,N_11347);
nand U12625 (N_12625,N_10848,N_11690);
or U12626 (N_12626,N_10480,N_10333);
and U12627 (N_12627,N_11239,N_10440);
nor U12628 (N_12628,N_11732,N_10430);
or U12629 (N_12629,N_11070,N_10660);
xor U12630 (N_12630,N_10749,N_11643);
nor U12631 (N_12631,N_11097,N_11162);
or U12632 (N_12632,N_11716,N_11740);
or U12633 (N_12633,N_11589,N_11214);
or U12634 (N_12634,N_11373,N_11121);
and U12635 (N_12635,N_10960,N_10380);
nand U12636 (N_12636,N_10823,N_11901);
and U12637 (N_12637,N_10561,N_11742);
or U12638 (N_12638,N_10858,N_11075);
nor U12639 (N_12639,N_11276,N_10762);
nand U12640 (N_12640,N_10882,N_11414);
nor U12641 (N_12641,N_11329,N_11228);
nor U12642 (N_12642,N_11317,N_11859);
nand U12643 (N_12643,N_11598,N_10723);
nor U12644 (N_12644,N_11510,N_10410);
xnor U12645 (N_12645,N_10010,N_10732);
nor U12646 (N_12646,N_10874,N_10961);
or U12647 (N_12647,N_11434,N_11593);
xnor U12648 (N_12648,N_11684,N_11894);
nand U12649 (N_12649,N_10738,N_10107);
nor U12650 (N_12650,N_11746,N_10260);
or U12651 (N_12651,N_10610,N_11547);
nor U12652 (N_12652,N_10793,N_10994);
nand U12653 (N_12653,N_11896,N_10840);
and U12654 (N_12654,N_11659,N_10329);
or U12655 (N_12655,N_10179,N_11977);
xor U12656 (N_12656,N_10611,N_11235);
or U12657 (N_12657,N_10140,N_11103);
and U12658 (N_12658,N_10638,N_10949);
nand U12659 (N_12659,N_10837,N_10915);
or U12660 (N_12660,N_11508,N_11575);
xnor U12661 (N_12661,N_11395,N_10792);
xnor U12662 (N_12662,N_11062,N_11436);
or U12663 (N_12663,N_11721,N_11191);
or U12664 (N_12664,N_11905,N_10887);
nor U12665 (N_12665,N_11349,N_10033);
nor U12666 (N_12666,N_11152,N_10058);
nand U12667 (N_12667,N_10220,N_11710);
nor U12668 (N_12668,N_10072,N_11241);
nand U12669 (N_12669,N_10217,N_11828);
or U12670 (N_12670,N_11470,N_11663);
or U12671 (N_12671,N_10068,N_10962);
nand U12672 (N_12672,N_10112,N_10338);
nand U12673 (N_12673,N_10707,N_10570);
and U12674 (N_12674,N_10921,N_10525);
and U12675 (N_12675,N_11753,N_11923);
nor U12676 (N_12676,N_11678,N_10134);
and U12677 (N_12677,N_11744,N_10203);
nand U12678 (N_12678,N_11515,N_11705);
nor U12679 (N_12679,N_11752,N_10912);
or U12680 (N_12680,N_11665,N_10977);
nor U12681 (N_12681,N_10141,N_10082);
nand U12682 (N_12682,N_10173,N_10712);
and U12683 (N_12683,N_11328,N_11109);
or U12684 (N_12684,N_10751,N_11762);
nand U12685 (N_12685,N_10411,N_11865);
nand U12686 (N_12686,N_11084,N_10008);
and U12687 (N_12687,N_10661,N_11862);
or U12688 (N_12688,N_11488,N_10859);
nor U12689 (N_12689,N_10137,N_10617);
nand U12690 (N_12690,N_10132,N_10407);
or U12691 (N_12691,N_10088,N_11327);
nand U12692 (N_12692,N_10824,N_10883);
and U12693 (N_12693,N_10662,N_10747);
or U12694 (N_12694,N_10413,N_11594);
or U12695 (N_12695,N_10328,N_10266);
or U12696 (N_12696,N_10979,N_11644);
nand U12697 (N_12697,N_11671,N_11313);
or U12698 (N_12698,N_11461,N_11628);
nor U12699 (N_12699,N_10341,N_11321);
or U12700 (N_12700,N_11840,N_11882);
and U12701 (N_12701,N_11346,N_11731);
or U12702 (N_12702,N_10631,N_10836);
nor U12703 (N_12703,N_11950,N_10005);
nand U12704 (N_12704,N_11661,N_11818);
nand U12705 (N_12705,N_10492,N_11836);
or U12706 (N_12706,N_11272,N_11426);
or U12707 (N_12707,N_11397,N_11001);
nor U12708 (N_12708,N_10626,N_10676);
nand U12709 (N_12709,N_10024,N_11528);
or U12710 (N_12710,N_11480,N_11964);
nor U12711 (N_12711,N_10955,N_10940);
xor U12712 (N_12712,N_11824,N_11806);
nor U12713 (N_12713,N_10569,N_10797);
and U12714 (N_12714,N_10251,N_11140);
nor U12715 (N_12715,N_10835,N_11856);
nor U12716 (N_12716,N_10985,N_10331);
or U12717 (N_12717,N_10375,N_10204);
nand U12718 (N_12718,N_11634,N_11284);
or U12719 (N_12719,N_10900,N_10186);
or U12720 (N_12720,N_10607,N_11042);
nor U12721 (N_12721,N_11937,N_10466);
nand U12722 (N_12722,N_10358,N_11827);
nor U12723 (N_12723,N_11814,N_11549);
and U12724 (N_12724,N_10282,N_10948);
nor U12725 (N_12725,N_11791,N_10239);
and U12726 (N_12726,N_10101,N_10056);
nand U12727 (N_12727,N_10043,N_10763);
nand U12728 (N_12728,N_11769,N_11068);
and U12729 (N_12729,N_11293,N_11564);
or U12730 (N_12730,N_11081,N_11898);
nand U12731 (N_12731,N_10442,N_11621);
or U12732 (N_12732,N_11043,N_11263);
or U12733 (N_12733,N_11294,N_11921);
nor U12734 (N_12734,N_10095,N_11518);
nor U12735 (N_12735,N_11004,N_11404);
nand U12736 (N_12736,N_10646,N_11058);
nand U12737 (N_12737,N_11783,N_11275);
or U12738 (N_12738,N_11014,N_11825);
and U12739 (N_12739,N_10754,N_11234);
nor U12740 (N_12740,N_10869,N_10180);
or U12741 (N_12741,N_10119,N_11835);
nor U12742 (N_12742,N_10774,N_11786);
nand U12743 (N_12743,N_11285,N_11674);
or U12744 (N_12744,N_10547,N_11908);
nand U12745 (N_12745,N_11072,N_11831);
or U12746 (N_12746,N_10769,N_10601);
and U12747 (N_12747,N_10461,N_10377);
nand U12748 (N_12748,N_11687,N_10135);
nor U12749 (N_12749,N_11458,N_10468);
nor U12750 (N_12750,N_11361,N_11726);
and U12751 (N_12751,N_11911,N_11131);
nor U12752 (N_12752,N_11622,N_10085);
or U12753 (N_12753,N_11522,N_11500);
nand U12754 (N_12754,N_11529,N_11654);
xnor U12755 (N_12755,N_11032,N_10078);
or U12756 (N_12756,N_11020,N_11662);
nor U12757 (N_12757,N_10718,N_10590);
nand U12758 (N_12758,N_10136,N_11560);
nand U12759 (N_12759,N_10500,N_11999);
nand U12760 (N_12760,N_10550,N_11400);
or U12761 (N_12761,N_10065,N_11543);
nor U12762 (N_12762,N_11064,N_11866);
and U12763 (N_12763,N_11768,N_10061);
or U12764 (N_12764,N_10020,N_11060);
xnor U12765 (N_12765,N_10782,N_10697);
and U12766 (N_12766,N_10971,N_11023);
and U12767 (N_12767,N_11533,N_11868);
or U12768 (N_12768,N_10892,N_10606);
nor U12769 (N_12769,N_10951,N_11230);
nand U12770 (N_12770,N_10437,N_11637);
or U12771 (N_12771,N_11904,N_11202);
nor U12772 (N_12772,N_10583,N_11021);
nor U12773 (N_12773,N_11401,N_10367);
nand U12774 (N_12774,N_11453,N_10084);
or U12775 (N_12775,N_11229,N_10213);
nand U12776 (N_12776,N_10452,N_11124);
nor U12777 (N_12777,N_10271,N_11597);
or U12778 (N_12778,N_10881,N_11206);
xnor U12779 (N_12779,N_10444,N_11128);
nand U12780 (N_12780,N_10167,N_10830);
xnor U12781 (N_12781,N_10248,N_11455);
and U12782 (N_12782,N_11137,N_10309);
and U12783 (N_12783,N_11189,N_10819);
nand U12784 (N_12784,N_11240,N_10856);
and U12785 (N_12785,N_10973,N_11432);
and U12786 (N_12786,N_11576,N_11798);
nand U12787 (N_12787,N_11796,N_10609);
nor U12788 (N_12788,N_10633,N_11822);
nor U12789 (N_12789,N_10495,N_11491);
nor U12790 (N_12790,N_11624,N_11811);
or U12791 (N_12791,N_10491,N_11027);
or U12792 (N_12792,N_10799,N_10909);
and U12793 (N_12793,N_11334,N_10384);
or U12794 (N_12794,N_10259,N_11788);
or U12795 (N_12795,N_10612,N_10575);
and U12796 (N_12796,N_10722,N_11917);
nand U12797 (N_12797,N_11514,N_11774);
or U12798 (N_12798,N_11524,N_10129);
nand U12799 (N_12799,N_10771,N_11613);
nand U12800 (N_12800,N_11971,N_11739);
nor U12801 (N_12801,N_10115,N_10855);
nor U12802 (N_12802,N_10433,N_11588);
nor U12803 (N_12803,N_11105,N_10857);
or U12804 (N_12804,N_10941,N_10057);
nand U12805 (N_12805,N_10425,N_10109);
and U12806 (N_12806,N_11845,N_10499);
and U12807 (N_12807,N_11496,N_11875);
nand U12808 (N_12808,N_10502,N_11221);
and U12809 (N_12809,N_10885,N_10376);
nor U12810 (N_12810,N_11179,N_10476);
and U12811 (N_12811,N_10846,N_10650);
nand U12812 (N_12812,N_11324,N_11981);
and U12813 (N_12813,N_10049,N_10616);
and U12814 (N_12814,N_11761,N_11260);
nand U12815 (N_12815,N_11503,N_11462);
nand U12816 (N_12816,N_10153,N_10009);
and U12817 (N_12817,N_10360,N_11946);
xnor U12818 (N_12818,N_11876,N_11473);
and U12819 (N_12819,N_10232,N_10560);
nand U12820 (N_12820,N_11163,N_10645);
or U12821 (N_12821,N_10690,N_11709);
nand U12822 (N_12822,N_11770,N_11651);
nand U12823 (N_12823,N_11618,N_11083);
and U12824 (N_12824,N_11351,N_11553);
or U12825 (N_12825,N_10827,N_10319);
and U12826 (N_12826,N_11100,N_10657);
or U12827 (N_12827,N_11463,N_10114);
or U12828 (N_12828,N_11748,N_10185);
nor U12829 (N_12829,N_10533,N_11407);
and U12830 (N_12830,N_11416,N_11498);
nor U12831 (N_12831,N_11175,N_11655);
and U12832 (N_12832,N_10721,N_10958);
nand U12833 (N_12833,N_10451,N_10427);
and U12834 (N_12834,N_10597,N_10235);
nor U12835 (N_12835,N_10669,N_11316);
nor U12836 (N_12836,N_10950,N_10489);
nor U12837 (N_12837,N_10108,N_10589);
xor U12838 (N_12838,N_11653,N_11858);
and U12839 (N_12839,N_10647,N_10171);
nand U12840 (N_12840,N_10920,N_11195);
nand U12841 (N_12841,N_11586,N_11949);
and U12842 (N_12842,N_10450,N_11925);
nor U12843 (N_12843,N_11889,N_11139);
and U12844 (N_12844,N_10130,N_10291);
nand U12845 (N_12845,N_10602,N_10999);
and U12846 (N_12846,N_10927,N_10620);
xor U12847 (N_12847,N_11143,N_10860);
nor U12848 (N_12848,N_10494,N_11092);
nor U12849 (N_12849,N_11136,N_11566);
nor U12850 (N_12850,N_11694,N_10418);
nand U12851 (N_12851,N_10145,N_10981);
xnor U12852 (N_12852,N_11724,N_11330);
nand U12853 (N_12853,N_10013,N_11850);
and U12854 (N_12854,N_10475,N_11115);
nor U12855 (N_12855,N_11073,N_10237);
and U12856 (N_12856,N_10479,N_11332);
and U12857 (N_12857,N_10667,N_10162);
and U12858 (N_12858,N_10671,N_10514);
nor U12859 (N_12859,N_11102,N_10187);
or U12860 (N_12860,N_10398,N_11722);
nand U12861 (N_12861,N_11358,N_10943);
or U12862 (N_12862,N_11269,N_11987);
or U12863 (N_12863,N_11813,N_11595);
nand U12864 (N_12864,N_10613,N_11714);
nor U12865 (N_12865,N_11431,N_10349);
xor U12866 (N_12866,N_11331,N_10828);
and U12867 (N_12867,N_11088,N_10456);
and U12868 (N_12868,N_11049,N_11247);
and U12869 (N_12869,N_10269,N_10868);
or U12870 (N_12870,N_11874,N_10498);
nor U12871 (N_12871,N_10573,N_10535);
xnor U12872 (N_12872,N_11640,N_10929);
nor U12873 (N_12873,N_10118,N_10047);
nor U12874 (N_12874,N_11601,N_10254);
and U12875 (N_12875,N_11668,N_11177);
nor U12876 (N_12876,N_10028,N_10513);
and U12877 (N_12877,N_10854,N_10336);
nor U12878 (N_12878,N_10700,N_11545);
or U12879 (N_12879,N_10211,N_11122);
nor U12880 (N_12880,N_10286,N_10031);
or U12881 (N_12881,N_10279,N_11989);
or U12882 (N_12882,N_10658,N_11029);
and U12883 (N_12883,N_10051,N_11497);
nor U12884 (N_12884,N_10894,N_11095);
and U12885 (N_12885,N_11040,N_10711);
nand U12886 (N_12886,N_10306,N_11880);
nor U12887 (N_12887,N_10947,N_11471);
nor U12888 (N_12888,N_10230,N_11912);
and U12889 (N_12889,N_11585,N_10249);
and U12890 (N_12890,N_10896,N_11998);
or U12891 (N_12891,N_10015,N_10212);
nor U12892 (N_12892,N_10905,N_10515);
nor U12893 (N_12893,N_10470,N_11325);
nand U12894 (N_12894,N_11707,N_10391);
and U12895 (N_12895,N_11267,N_10445);
nand U12896 (N_12896,N_10390,N_10901);
and U12897 (N_12897,N_11474,N_10557);
or U12898 (N_12898,N_11535,N_10507);
and U12899 (N_12899,N_10670,N_11301);
nand U12900 (N_12900,N_10000,N_10127);
and U12901 (N_12901,N_11129,N_11869);
or U12902 (N_12902,N_11756,N_11807);
nor U12903 (N_12903,N_10018,N_11297);
or U12904 (N_12904,N_11817,N_11801);
and U12905 (N_12905,N_10673,N_11465);
and U12906 (N_12906,N_11629,N_11010);
and U12907 (N_12907,N_11441,N_10149);
or U12908 (N_12908,N_10003,N_11031);
nand U12909 (N_12909,N_10045,N_11741);
and U12910 (N_12910,N_10340,N_10889);
and U12911 (N_12911,N_10059,N_10701);
nor U12912 (N_12912,N_11466,N_11712);
nor U12913 (N_12913,N_11047,N_10761);
and U12914 (N_12914,N_10395,N_11623);
or U12915 (N_12915,N_11264,N_11751);
nor U12916 (N_12916,N_10759,N_10694);
nor U12917 (N_12917,N_10296,N_10353);
nor U12918 (N_12918,N_10019,N_10463);
nand U12919 (N_12919,N_11389,N_11258);
and U12920 (N_12920,N_11899,N_10121);
and U12921 (N_12921,N_10625,N_11727);
or U12922 (N_12922,N_10891,N_10098);
nor U12923 (N_12923,N_10342,N_11963);
nor U12924 (N_12924,N_10356,N_11339);
or U12925 (N_12925,N_10801,N_10474);
or U12926 (N_12926,N_11519,N_11486);
or U12927 (N_12927,N_10062,N_10778);
nor U12928 (N_12928,N_10128,N_11196);
xnor U12929 (N_12929,N_11909,N_11211);
and U12930 (N_12930,N_10192,N_10267);
nor U12931 (N_12931,N_11991,N_11343);
and U12932 (N_12932,N_11440,N_11861);
nor U12933 (N_12933,N_11394,N_10138);
or U12934 (N_12934,N_11287,N_11992);
and U12935 (N_12935,N_10076,N_10904);
nor U12936 (N_12936,N_10030,N_10986);
or U12937 (N_12937,N_10194,N_10796);
and U12938 (N_12938,N_10807,N_11567);
nand U12939 (N_12939,N_11448,N_10564);
nor U12940 (N_12940,N_10312,N_11614);
and U12941 (N_12941,N_11667,N_10174);
nor U12942 (N_12942,N_10632,N_11848);
nand U12943 (N_12943,N_10791,N_11626);
nor U12944 (N_12944,N_10275,N_11699);
and U12945 (N_12945,N_11039,N_11363);
nand U12946 (N_12946,N_10176,N_10520);
nor U12947 (N_12947,N_10091,N_10906);
nand U12948 (N_12948,N_10553,N_10079);
or U12949 (N_12949,N_11592,N_11583);
xnor U12950 (N_12950,N_10713,N_10094);
nand U12951 (N_12951,N_11803,N_10886);
nand U12952 (N_12952,N_10538,N_11222);
nand U12953 (N_12953,N_11379,N_10902);
or U12954 (N_12954,N_11479,N_10471);
or U12955 (N_12955,N_11639,N_10524);
and U12956 (N_12956,N_11736,N_11823);
nor U12957 (N_12957,N_10624,N_10175);
nor U12958 (N_12958,N_11464,N_11934);
nor U12959 (N_12959,N_11384,N_10998);
nand U12960 (N_12960,N_11656,N_10741);
or U12961 (N_12961,N_11046,N_11071);
nand U12962 (N_12962,N_11255,N_10099);
nor U12963 (N_12963,N_11459,N_11857);
nor U12964 (N_12964,N_11481,N_11527);
nor U12965 (N_12965,N_11779,N_10123);
or U12966 (N_12966,N_11174,N_11776);
and U12967 (N_12967,N_11483,N_10598);
or U12968 (N_12968,N_11616,N_10581);
nand U12969 (N_12969,N_11677,N_11976);
nand U12970 (N_12970,N_11887,N_10622);
nor U12971 (N_12971,N_11877,N_10748);
and U12972 (N_12972,N_10596,N_10649);
nand U12973 (N_12973,N_10357,N_10334);
xor U12974 (N_12974,N_10325,N_10692);
or U12975 (N_12975,N_10978,N_10522);
nand U12976 (N_12976,N_11658,N_10142);
nand U12977 (N_12977,N_11318,N_11380);
or U12978 (N_12978,N_11319,N_11829);
nor U12979 (N_12979,N_11282,N_11738);
or U12980 (N_12980,N_11212,N_10772);
nor U12981 (N_12981,N_11645,N_11792);
xnor U12982 (N_12982,N_10181,N_10304);
and U12983 (N_12983,N_10283,N_10026);
and U12984 (N_12984,N_11983,N_10733);
or U12985 (N_12985,N_11969,N_10278);
and U12986 (N_12986,N_10969,N_10668);
and U12987 (N_12987,N_11772,N_10808);
nor U12988 (N_12988,N_10268,N_10715);
xnor U12989 (N_12989,N_11669,N_10040);
nor U12990 (N_12990,N_10105,N_11781);
and U12991 (N_12991,N_10605,N_11186);
nand U12992 (N_12992,N_11052,N_11271);
nand U12993 (N_12993,N_10730,N_10104);
or U12994 (N_12994,N_11797,N_11910);
nor U12995 (N_12995,N_10640,N_10844);
or U12996 (N_12996,N_10196,N_10600);
and U12997 (N_12997,N_11559,N_11970);
and U12998 (N_12998,N_10838,N_11041);
nand U12999 (N_12999,N_11454,N_10289);
and U13000 (N_13000,N_10412,N_10527);
nand U13001 (N_13001,N_10960,N_10025);
or U13002 (N_13002,N_11482,N_10142);
and U13003 (N_13003,N_11504,N_11524);
and U13004 (N_13004,N_10670,N_11481);
or U13005 (N_13005,N_11778,N_11148);
or U13006 (N_13006,N_10539,N_11774);
nand U13007 (N_13007,N_11337,N_11495);
nor U13008 (N_13008,N_11038,N_10728);
xnor U13009 (N_13009,N_10776,N_11554);
or U13010 (N_13010,N_11351,N_10635);
and U13011 (N_13011,N_10326,N_10500);
nor U13012 (N_13012,N_11704,N_11414);
nand U13013 (N_13013,N_10690,N_11590);
nand U13014 (N_13014,N_11441,N_10375);
nor U13015 (N_13015,N_11126,N_10820);
or U13016 (N_13016,N_10833,N_11258);
nand U13017 (N_13017,N_10388,N_10398);
nor U13018 (N_13018,N_11628,N_11604);
and U13019 (N_13019,N_10020,N_11221);
nand U13020 (N_13020,N_10525,N_10441);
and U13021 (N_13021,N_11169,N_11154);
or U13022 (N_13022,N_11219,N_11676);
or U13023 (N_13023,N_11444,N_11865);
and U13024 (N_13024,N_11834,N_11219);
nor U13025 (N_13025,N_10744,N_10135);
or U13026 (N_13026,N_11273,N_11628);
xnor U13027 (N_13027,N_11648,N_10164);
nor U13028 (N_13028,N_10212,N_10563);
nand U13029 (N_13029,N_11452,N_11435);
nor U13030 (N_13030,N_10877,N_10269);
and U13031 (N_13031,N_10503,N_11694);
or U13032 (N_13032,N_10467,N_11179);
and U13033 (N_13033,N_10544,N_11652);
nor U13034 (N_13034,N_11073,N_11123);
xnor U13035 (N_13035,N_11475,N_10571);
nor U13036 (N_13036,N_10094,N_11482);
and U13037 (N_13037,N_10668,N_10815);
nor U13038 (N_13038,N_10097,N_10430);
nor U13039 (N_13039,N_11976,N_10153);
and U13040 (N_13040,N_10171,N_11974);
or U13041 (N_13041,N_10406,N_11005);
nand U13042 (N_13042,N_11494,N_11106);
nor U13043 (N_13043,N_10216,N_10139);
nand U13044 (N_13044,N_11379,N_10119);
nor U13045 (N_13045,N_10422,N_11945);
nand U13046 (N_13046,N_11462,N_10507);
or U13047 (N_13047,N_11224,N_11908);
or U13048 (N_13048,N_11286,N_11711);
nor U13049 (N_13049,N_11625,N_11658);
nor U13050 (N_13050,N_10240,N_11350);
nand U13051 (N_13051,N_10649,N_10206);
nand U13052 (N_13052,N_10309,N_10212);
nor U13053 (N_13053,N_11930,N_11376);
or U13054 (N_13054,N_11913,N_10343);
and U13055 (N_13055,N_10049,N_10067);
or U13056 (N_13056,N_11913,N_10114);
and U13057 (N_13057,N_10814,N_10713);
and U13058 (N_13058,N_11981,N_10606);
nand U13059 (N_13059,N_10110,N_10398);
or U13060 (N_13060,N_10709,N_11151);
nor U13061 (N_13061,N_11374,N_11589);
nor U13062 (N_13062,N_11688,N_10492);
and U13063 (N_13063,N_11396,N_10999);
and U13064 (N_13064,N_11944,N_11675);
nor U13065 (N_13065,N_10653,N_11583);
or U13066 (N_13066,N_11704,N_10774);
nor U13067 (N_13067,N_10631,N_10281);
and U13068 (N_13068,N_10458,N_11721);
nand U13069 (N_13069,N_11116,N_10563);
nor U13070 (N_13070,N_10042,N_11490);
and U13071 (N_13071,N_11144,N_10436);
nor U13072 (N_13072,N_11234,N_11145);
nand U13073 (N_13073,N_10619,N_10245);
nor U13074 (N_13074,N_11268,N_10026);
or U13075 (N_13075,N_11893,N_10457);
and U13076 (N_13076,N_10297,N_11713);
nor U13077 (N_13077,N_10304,N_10425);
and U13078 (N_13078,N_11884,N_10735);
and U13079 (N_13079,N_10597,N_10056);
or U13080 (N_13080,N_10134,N_11777);
and U13081 (N_13081,N_10735,N_11895);
nor U13082 (N_13082,N_11069,N_10853);
or U13083 (N_13083,N_11608,N_10722);
and U13084 (N_13084,N_11810,N_11332);
nor U13085 (N_13085,N_10002,N_11446);
or U13086 (N_13086,N_10031,N_11812);
or U13087 (N_13087,N_11407,N_10832);
or U13088 (N_13088,N_11541,N_11900);
or U13089 (N_13089,N_10430,N_10477);
nand U13090 (N_13090,N_11065,N_11557);
or U13091 (N_13091,N_11574,N_10026);
and U13092 (N_13092,N_10754,N_11315);
nand U13093 (N_13093,N_10969,N_11095);
nand U13094 (N_13094,N_11168,N_11981);
or U13095 (N_13095,N_10776,N_10793);
and U13096 (N_13096,N_11807,N_10799);
nor U13097 (N_13097,N_10709,N_10533);
nand U13098 (N_13098,N_10112,N_11075);
or U13099 (N_13099,N_10106,N_10552);
and U13100 (N_13100,N_11779,N_10854);
nand U13101 (N_13101,N_10454,N_10603);
nor U13102 (N_13102,N_10434,N_11828);
or U13103 (N_13103,N_10205,N_11660);
nand U13104 (N_13104,N_11370,N_10372);
or U13105 (N_13105,N_11197,N_10801);
and U13106 (N_13106,N_11028,N_10675);
and U13107 (N_13107,N_11812,N_11922);
nor U13108 (N_13108,N_11878,N_11790);
or U13109 (N_13109,N_10065,N_10623);
nand U13110 (N_13110,N_11652,N_10913);
nor U13111 (N_13111,N_11202,N_11739);
nor U13112 (N_13112,N_11029,N_11180);
or U13113 (N_13113,N_10078,N_10902);
and U13114 (N_13114,N_10895,N_11685);
nor U13115 (N_13115,N_10424,N_11707);
and U13116 (N_13116,N_10294,N_11281);
nand U13117 (N_13117,N_10439,N_10744);
and U13118 (N_13118,N_10010,N_10795);
nand U13119 (N_13119,N_10424,N_10219);
nand U13120 (N_13120,N_11483,N_10930);
nand U13121 (N_13121,N_11774,N_10315);
nand U13122 (N_13122,N_11115,N_11738);
or U13123 (N_13123,N_10069,N_10461);
or U13124 (N_13124,N_11241,N_10789);
nand U13125 (N_13125,N_11839,N_11613);
nand U13126 (N_13126,N_10856,N_11774);
and U13127 (N_13127,N_11348,N_10482);
and U13128 (N_13128,N_11074,N_10129);
or U13129 (N_13129,N_10136,N_11274);
nor U13130 (N_13130,N_10377,N_10960);
nand U13131 (N_13131,N_10119,N_10714);
or U13132 (N_13132,N_10317,N_11424);
nor U13133 (N_13133,N_11900,N_11433);
and U13134 (N_13134,N_10710,N_10916);
nor U13135 (N_13135,N_10279,N_10734);
nor U13136 (N_13136,N_10622,N_10820);
or U13137 (N_13137,N_10515,N_10650);
nand U13138 (N_13138,N_10203,N_11434);
nand U13139 (N_13139,N_11791,N_11241);
and U13140 (N_13140,N_11341,N_10507);
and U13141 (N_13141,N_11403,N_10558);
nor U13142 (N_13142,N_11036,N_11278);
or U13143 (N_13143,N_10305,N_11573);
nand U13144 (N_13144,N_11545,N_11568);
and U13145 (N_13145,N_11566,N_11265);
or U13146 (N_13146,N_11085,N_11653);
and U13147 (N_13147,N_10281,N_11199);
nor U13148 (N_13148,N_11050,N_10900);
or U13149 (N_13149,N_11147,N_11778);
and U13150 (N_13150,N_11569,N_10879);
and U13151 (N_13151,N_10902,N_10874);
or U13152 (N_13152,N_10827,N_10065);
nand U13153 (N_13153,N_10233,N_11919);
and U13154 (N_13154,N_11371,N_11140);
or U13155 (N_13155,N_10606,N_10841);
nand U13156 (N_13156,N_10591,N_11760);
and U13157 (N_13157,N_11571,N_11053);
nand U13158 (N_13158,N_11474,N_11599);
nor U13159 (N_13159,N_11406,N_11526);
and U13160 (N_13160,N_11336,N_11014);
nor U13161 (N_13161,N_10456,N_10493);
or U13162 (N_13162,N_10880,N_10289);
nand U13163 (N_13163,N_10689,N_10786);
or U13164 (N_13164,N_10421,N_11913);
nor U13165 (N_13165,N_10325,N_11932);
nand U13166 (N_13166,N_10698,N_11803);
and U13167 (N_13167,N_11546,N_10554);
or U13168 (N_13168,N_11489,N_10275);
nor U13169 (N_13169,N_10333,N_10384);
nand U13170 (N_13170,N_10436,N_11097);
or U13171 (N_13171,N_11688,N_11983);
and U13172 (N_13172,N_10590,N_11956);
nor U13173 (N_13173,N_11235,N_10898);
or U13174 (N_13174,N_10101,N_10656);
nor U13175 (N_13175,N_10157,N_10302);
and U13176 (N_13176,N_11965,N_10348);
xnor U13177 (N_13177,N_11987,N_10717);
or U13178 (N_13178,N_11145,N_11063);
nor U13179 (N_13179,N_10853,N_11614);
or U13180 (N_13180,N_10909,N_10580);
or U13181 (N_13181,N_10225,N_10358);
and U13182 (N_13182,N_10560,N_10596);
nand U13183 (N_13183,N_10620,N_11924);
and U13184 (N_13184,N_11460,N_10251);
nor U13185 (N_13185,N_10865,N_11540);
nor U13186 (N_13186,N_10633,N_10806);
nand U13187 (N_13187,N_10599,N_10140);
nand U13188 (N_13188,N_10006,N_11394);
or U13189 (N_13189,N_10543,N_11077);
and U13190 (N_13190,N_10560,N_11076);
nor U13191 (N_13191,N_10700,N_10683);
nand U13192 (N_13192,N_11294,N_11301);
and U13193 (N_13193,N_11515,N_10274);
nor U13194 (N_13194,N_11463,N_10966);
nand U13195 (N_13195,N_11215,N_11402);
nand U13196 (N_13196,N_10101,N_11942);
nand U13197 (N_13197,N_10935,N_10195);
and U13198 (N_13198,N_10507,N_10476);
nand U13199 (N_13199,N_11578,N_10133);
or U13200 (N_13200,N_10906,N_10395);
nand U13201 (N_13201,N_11717,N_11868);
or U13202 (N_13202,N_10396,N_11348);
nand U13203 (N_13203,N_10818,N_11516);
or U13204 (N_13204,N_11855,N_10855);
nor U13205 (N_13205,N_10656,N_11516);
nor U13206 (N_13206,N_10484,N_11954);
nand U13207 (N_13207,N_11388,N_10094);
and U13208 (N_13208,N_11926,N_10952);
nor U13209 (N_13209,N_11210,N_10279);
nor U13210 (N_13210,N_11035,N_10821);
nor U13211 (N_13211,N_11749,N_10399);
nand U13212 (N_13212,N_10863,N_10986);
and U13213 (N_13213,N_11407,N_11519);
nor U13214 (N_13214,N_10993,N_10326);
nand U13215 (N_13215,N_10471,N_10938);
xor U13216 (N_13216,N_11470,N_11081);
nand U13217 (N_13217,N_11252,N_11355);
or U13218 (N_13218,N_11224,N_11322);
nand U13219 (N_13219,N_11144,N_10637);
and U13220 (N_13220,N_11679,N_10600);
nor U13221 (N_13221,N_11998,N_10197);
or U13222 (N_13222,N_11166,N_11183);
or U13223 (N_13223,N_11934,N_11660);
or U13224 (N_13224,N_11549,N_11081);
and U13225 (N_13225,N_10820,N_10362);
or U13226 (N_13226,N_10719,N_10730);
nor U13227 (N_13227,N_11412,N_11114);
and U13228 (N_13228,N_10145,N_11745);
nand U13229 (N_13229,N_11847,N_11986);
and U13230 (N_13230,N_10510,N_11190);
or U13231 (N_13231,N_10176,N_10480);
nand U13232 (N_13232,N_11200,N_10585);
nor U13233 (N_13233,N_11424,N_10615);
nor U13234 (N_13234,N_11209,N_11557);
or U13235 (N_13235,N_11113,N_10020);
xnor U13236 (N_13236,N_10041,N_11973);
or U13237 (N_13237,N_11579,N_10528);
or U13238 (N_13238,N_11809,N_10598);
nand U13239 (N_13239,N_11161,N_11433);
or U13240 (N_13240,N_10873,N_10458);
nand U13241 (N_13241,N_10049,N_11827);
or U13242 (N_13242,N_11641,N_10048);
and U13243 (N_13243,N_10270,N_11203);
and U13244 (N_13244,N_11772,N_11472);
nand U13245 (N_13245,N_10200,N_11974);
nand U13246 (N_13246,N_10807,N_10137);
nand U13247 (N_13247,N_10202,N_11747);
nand U13248 (N_13248,N_11016,N_10353);
or U13249 (N_13249,N_10610,N_11499);
and U13250 (N_13250,N_10438,N_11032);
nand U13251 (N_13251,N_11942,N_11828);
nor U13252 (N_13252,N_11955,N_11176);
or U13253 (N_13253,N_11261,N_11950);
and U13254 (N_13254,N_11093,N_10433);
or U13255 (N_13255,N_10984,N_10696);
nor U13256 (N_13256,N_11909,N_11189);
and U13257 (N_13257,N_11626,N_10220);
nand U13258 (N_13258,N_10669,N_10322);
xnor U13259 (N_13259,N_10776,N_11446);
or U13260 (N_13260,N_11204,N_11746);
nand U13261 (N_13261,N_11779,N_10736);
and U13262 (N_13262,N_11948,N_11688);
nor U13263 (N_13263,N_11429,N_11569);
nor U13264 (N_13264,N_10536,N_11754);
and U13265 (N_13265,N_11997,N_11194);
or U13266 (N_13266,N_10106,N_11980);
nor U13267 (N_13267,N_10252,N_10178);
xor U13268 (N_13268,N_11909,N_10030);
xnor U13269 (N_13269,N_10764,N_10681);
nor U13270 (N_13270,N_11619,N_10923);
or U13271 (N_13271,N_10618,N_10565);
nand U13272 (N_13272,N_10050,N_11329);
nor U13273 (N_13273,N_11658,N_10811);
nor U13274 (N_13274,N_10673,N_11015);
nor U13275 (N_13275,N_10839,N_10339);
nand U13276 (N_13276,N_11800,N_10680);
or U13277 (N_13277,N_11916,N_10241);
and U13278 (N_13278,N_10484,N_10229);
nor U13279 (N_13279,N_11778,N_11238);
and U13280 (N_13280,N_10865,N_11405);
or U13281 (N_13281,N_10215,N_11600);
nand U13282 (N_13282,N_10130,N_10389);
nand U13283 (N_13283,N_10308,N_10381);
nand U13284 (N_13284,N_10382,N_10645);
nand U13285 (N_13285,N_10309,N_11188);
or U13286 (N_13286,N_10413,N_11751);
nor U13287 (N_13287,N_11685,N_10591);
nor U13288 (N_13288,N_10005,N_11725);
and U13289 (N_13289,N_10161,N_10279);
or U13290 (N_13290,N_11135,N_11584);
or U13291 (N_13291,N_10670,N_11462);
or U13292 (N_13292,N_11035,N_11260);
nand U13293 (N_13293,N_11628,N_10932);
nor U13294 (N_13294,N_10849,N_11030);
nor U13295 (N_13295,N_10346,N_11896);
or U13296 (N_13296,N_11563,N_10247);
or U13297 (N_13297,N_11969,N_10959);
or U13298 (N_13298,N_10425,N_11213);
and U13299 (N_13299,N_11812,N_10075);
and U13300 (N_13300,N_11192,N_11170);
or U13301 (N_13301,N_11244,N_11141);
or U13302 (N_13302,N_11772,N_11823);
nor U13303 (N_13303,N_10960,N_10753);
and U13304 (N_13304,N_11254,N_10105);
or U13305 (N_13305,N_11796,N_10390);
or U13306 (N_13306,N_11078,N_11622);
and U13307 (N_13307,N_11398,N_10007);
and U13308 (N_13308,N_10665,N_11011);
nor U13309 (N_13309,N_10196,N_10177);
nor U13310 (N_13310,N_11240,N_11346);
nor U13311 (N_13311,N_11561,N_11638);
and U13312 (N_13312,N_10663,N_10841);
nor U13313 (N_13313,N_11823,N_11428);
and U13314 (N_13314,N_10399,N_10240);
nor U13315 (N_13315,N_11131,N_11379);
nand U13316 (N_13316,N_10959,N_11804);
nand U13317 (N_13317,N_10154,N_10384);
and U13318 (N_13318,N_10258,N_11757);
nor U13319 (N_13319,N_10628,N_10330);
nor U13320 (N_13320,N_10990,N_10352);
and U13321 (N_13321,N_10209,N_10257);
or U13322 (N_13322,N_10758,N_11712);
nand U13323 (N_13323,N_10013,N_11945);
nor U13324 (N_13324,N_11920,N_10759);
or U13325 (N_13325,N_11554,N_10182);
and U13326 (N_13326,N_11826,N_11054);
or U13327 (N_13327,N_10993,N_10278);
nand U13328 (N_13328,N_10426,N_10454);
and U13329 (N_13329,N_10117,N_11895);
nor U13330 (N_13330,N_10653,N_10942);
nand U13331 (N_13331,N_11426,N_11838);
or U13332 (N_13332,N_10796,N_10072);
and U13333 (N_13333,N_10717,N_11400);
nand U13334 (N_13334,N_10907,N_10189);
or U13335 (N_13335,N_10807,N_10996);
nand U13336 (N_13336,N_10979,N_11249);
or U13337 (N_13337,N_10905,N_11401);
or U13338 (N_13338,N_10798,N_10512);
and U13339 (N_13339,N_11062,N_11156);
or U13340 (N_13340,N_10167,N_11484);
and U13341 (N_13341,N_11777,N_11861);
nor U13342 (N_13342,N_11662,N_10515);
and U13343 (N_13343,N_11404,N_11212);
or U13344 (N_13344,N_11584,N_10545);
nor U13345 (N_13345,N_11876,N_10251);
or U13346 (N_13346,N_10951,N_10773);
nor U13347 (N_13347,N_10091,N_11780);
nor U13348 (N_13348,N_10318,N_10031);
or U13349 (N_13349,N_10356,N_10988);
nand U13350 (N_13350,N_10548,N_10653);
and U13351 (N_13351,N_10422,N_10312);
nor U13352 (N_13352,N_10937,N_10625);
and U13353 (N_13353,N_11057,N_11936);
and U13354 (N_13354,N_10233,N_11260);
nor U13355 (N_13355,N_11737,N_10469);
nor U13356 (N_13356,N_11711,N_10195);
nor U13357 (N_13357,N_10014,N_11768);
nor U13358 (N_13358,N_11530,N_11577);
nor U13359 (N_13359,N_10801,N_10653);
or U13360 (N_13360,N_11283,N_11639);
nand U13361 (N_13361,N_11092,N_10813);
and U13362 (N_13362,N_10692,N_11383);
and U13363 (N_13363,N_10944,N_10917);
xnor U13364 (N_13364,N_11061,N_10179);
or U13365 (N_13365,N_10407,N_10704);
and U13366 (N_13366,N_10672,N_11686);
nor U13367 (N_13367,N_10207,N_11126);
and U13368 (N_13368,N_10215,N_10290);
nor U13369 (N_13369,N_11236,N_11730);
nand U13370 (N_13370,N_11515,N_11721);
or U13371 (N_13371,N_10204,N_11369);
nand U13372 (N_13372,N_11322,N_10082);
nand U13373 (N_13373,N_11453,N_11401);
nand U13374 (N_13374,N_11128,N_11094);
and U13375 (N_13375,N_11766,N_10426);
nand U13376 (N_13376,N_10450,N_11208);
or U13377 (N_13377,N_10303,N_11515);
and U13378 (N_13378,N_11260,N_11967);
or U13379 (N_13379,N_11469,N_10511);
nor U13380 (N_13380,N_10811,N_10723);
nand U13381 (N_13381,N_11401,N_11113);
nor U13382 (N_13382,N_11122,N_10351);
and U13383 (N_13383,N_10515,N_10458);
or U13384 (N_13384,N_11442,N_11297);
nand U13385 (N_13385,N_11206,N_11542);
and U13386 (N_13386,N_11103,N_11374);
or U13387 (N_13387,N_11549,N_11899);
nor U13388 (N_13388,N_10471,N_10654);
nand U13389 (N_13389,N_10670,N_11683);
or U13390 (N_13390,N_10656,N_11975);
nand U13391 (N_13391,N_11824,N_10861);
nand U13392 (N_13392,N_10572,N_10557);
nand U13393 (N_13393,N_11219,N_10906);
and U13394 (N_13394,N_10684,N_10742);
or U13395 (N_13395,N_11433,N_10487);
or U13396 (N_13396,N_10290,N_11860);
nand U13397 (N_13397,N_10925,N_11756);
nor U13398 (N_13398,N_11602,N_10008);
or U13399 (N_13399,N_10992,N_11431);
and U13400 (N_13400,N_11253,N_10312);
nor U13401 (N_13401,N_11593,N_11519);
or U13402 (N_13402,N_11024,N_11419);
nor U13403 (N_13403,N_10762,N_10107);
nor U13404 (N_13404,N_11280,N_11087);
nor U13405 (N_13405,N_11093,N_10894);
nand U13406 (N_13406,N_11664,N_10271);
and U13407 (N_13407,N_10034,N_10846);
or U13408 (N_13408,N_10890,N_10709);
or U13409 (N_13409,N_11650,N_11859);
or U13410 (N_13410,N_10046,N_10856);
nand U13411 (N_13411,N_10359,N_10602);
and U13412 (N_13412,N_11813,N_10811);
nor U13413 (N_13413,N_11940,N_11326);
nand U13414 (N_13414,N_11583,N_11912);
and U13415 (N_13415,N_11973,N_10270);
nor U13416 (N_13416,N_10177,N_10623);
or U13417 (N_13417,N_10302,N_11830);
nand U13418 (N_13418,N_10451,N_10253);
nor U13419 (N_13419,N_10390,N_10768);
and U13420 (N_13420,N_11934,N_10403);
nor U13421 (N_13421,N_11092,N_10627);
nand U13422 (N_13422,N_10025,N_10571);
nor U13423 (N_13423,N_10617,N_11889);
nand U13424 (N_13424,N_10886,N_10004);
or U13425 (N_13425,N_10859,N_11584);
and U13426 (N_13426,N_10217,N_10782);
and U13427 (N_13427,N_10938,N_11461);
nor U13428 (N_13428,N_10680,N_11448);
and U13429 (N_13429,N_10631,N_11712);
nand U13430 (N_13430,N_11481,N_10456);
nand U13431 (N_13431,N_11622,N_11256);
nand U13432 (N_13432,N_10542,N_11180);
nor U13433 (N_13433,N_11962,N_10966);
nor U13434 (N_13434,N_11321,N_10475);
nand U13435 (N_13435,N_11691,N_11774);
nor U13436 (N_13436,N_11254,N_10195);
and U13437 (N_13437,N_10128,N_10561);
nor U13438 (N_13438,N_11461,N_11340);
and U13439 (N_13439,N_11458,N_11711);
and U13440 (N_13440,N_10585,N_10810);
nand U13441 (N_13441,N_11498,N_11927);
nor U13442 (N_13442,N_11358,N_11604);
and U13443 (N_13443,N_11848,N_11805);
nor U13444 (N_13444,N_11066,N_11201);
nand U13445 (N_13445,N_10928,N_10293);
nand U13446 (N_13446,N_10628,N_11812);
nand U13447 (N_13447,N_10184,N_10152);
or U13448 (N_13448,N_11552,N_11510);
nand U13449 (N_13449,N_11328,N_11429);
nor U13450 (N_13450,N_11244,N_11430);
and U13451 (N_13451,N_11513,N_11975);
nor U13452 (N_13452,N_11083,N_11465);
nor U13453 (N_13453,N_11170,N_11988);
and U13454 (N_13454,N_11557,N_10099);
nor U13455 (N_13455,N_10815,N_10757);
and U13456 (N_13456,N_11759,N_11835);
nor U13457 (N_13457,N_11077,N_11473);
or U13458 (N_13458,N_10677,N_10149);
nand U13459 (N_13459,N_10528,N_10050);
and U13460 (N_13460,N_11191,N_10780);
nor U13461 (N_13461,N_11941,N_11812);
nand U13462 (N_13462,N_11835,N_10888);
nor U13463 (N_13463,N_11015,N_11105);
nor U13464 (N_13464,N_10109,N_11835);
nor U13465 (N_13465,N_10696,N_10317);
or U13466 (N_13466,N_11599,N_10802);
and U13467 (N_13467,N_10886,N_10332);
nand U13468 (N_13468,N_11152,N_10957);
or U13469 (N_13469,N_10706,N_11018);
nand U13470 (N_13470,N_11075,N_11028);
and U13471 (N_13471,N_11103,N_10828);
and U13472 (N_13472,N_11444,N_10316);
and U13473 (N_13473,N_11849,N_11735);
nand U13474 (N_13474,N_11102,N_11647);
and U13475 (N_13475,N_10739,N_10801);
or U13476 (N_13476,N_10146,N_11726);
or U13477 (N_13477,N_10900,N_10539);
or U13478 (N_13478,N_10639,N_10777);
and U13479 (N_13479,N_11906,N_11457);
xor U13480 (N_13480,N_11471,N_10042);
or U13481 (N_13481,N_10060,N_10670);
nand U13482 (N_13482,N_11309,N_11084);
nor U13483 (N_13483,N_10728,N_10959);
nor U13484 (N_13484,N_10143,N_10862);
and U13485 (N_13485,N_10071,N_11635);
nand U13486 (N_13486,N_10116,N_11153);
or U13487 (N_13487,N_11808,N_11633);
nand U13488 (N_13488,N_11378,N_10294);
or U13489 (N_13489,N_11430,N_11403);
or U13490 (N_13490,N_10898,N_11770);
nor U13491 (N_13491,N_10916,N_10610);
and U13492 (N_13492,N_10786,N_10963);
nor U13493 (N_13493,N_11317,N_11283);
nor U13494 (N_13494,N_11422,N_11058);
or U13495 (N_13495,N_11102,N_10312);
or U13496 (N_13496,N_11281,N_11563);
nand U13497 (N_13497,N_11923,N_11725);
and U13498 (N_13498,N_10486,N_10510);
nor U13499 (N_13499,N_11898,N_10433);
nand U13500 (N_13500,N_11459,N_10058);
nand U13501 (N_13501,N_11073,N_10656);
or U13502 (N_13502,N_11042,N_10115);
nor U13503 (N_13503,N_10568,N_11827);
nand U13504 (N_13504,N_11839,N_11106);
nor U13505 (N_13505,N_10745,N_11450);
nor U13506 (N_13506,N_10050,N_10270);
or U13507 (N_13507,N_11614,N_11937);
or U13508 (N_13508,N_10875,N_10370);
nor U13509 (N_13509,N_11080,N_10117);
nor U13510 (N_13510,N_10052,N_11160);
nor U13511 (N_13511,N_11141,N_10092);
and U13512 (N_13512,N_11530,N_10679);
or U13513 (N_13513,N_10671,N_10743);
or U13514 (N_13514,N_10843,N_11965);
and U13515 (N_13515,N_10358,N_10976);
and U13516 (N_13516,N_11200,N_10235);
xnor U13517 (N_13517,N_10611,N_11919);
or U13518 (N_13518,N_11110,N_11186);
or U13519 (N_13519,N_10420,N_11672);
nand U13520 (N_13520,N_11866,N_10325);
or U13521 (N_13521,N_10781,N_11864);
and U13522 (N_13522,N_11029,N_10981);
xor U13523 (N_13523,N_11770,N_11591);
nor U13524 (N_13524,N_11177,N_11309);
and U13525 (N_13525,N_11371,N_11800);
nand U13526 (N_13526,N_11366,N_11763);
and U13527 (N_13527,N_10385,N_11058);
and U13528 (N_13528,N_11788,N_10459);
nand U13529 (N_13529,N_11617,N_11732);
nand U13530 (N_13530,N_11454,N_11372);
and U13531 (N_13531,N_10934,N_10878);
or U13532 (N_13532,N_11923,N_11971);
nand U13533 (N_13533,N_11949,N_10190);
xor U13534 (N_13534,N_10360,N_10131);
or U13535 (N_13535,N_11181,N_10947);
nor U13536 (N_13536,N_11174,N_10020);
nand U13537 (N_13537,N_11082,N_11383);
nor U13538 (N_13538,N_10164,N_10991);
nand U13539 (N_13539,N_11439,N_10721);
nor U13540 (N_13540,N_10382,N_11425);
and U13541 (N_13541,N_10282,N_10183);
and U13542 (N_13542,N_10746,N_10895);
nor U13543 (N_13543,N_11860,N_11172);
nor U13544 (N_13544,N_10024,N_10515);
nor U13545 (N_13545,N_10285,N_11561);
or U13546 (N_13546,N_10560,N_10511);
or U13547 (N_13547,N_10718,N_10414);
nor U13548 (N_13548,N_10977,N_10850);
or U13549 (N_13549,N_11880,N_11294);
nor U13550 (N_13550,N_11652,N_11548);
nor U13551 (N_13551,N_10558,N_10595);
or U13552 (N_13552,N_10403,N_11661);
nand U13553 (N_13553,N_10094,N_11803);
nand U13554 (N_13554,N_10954,N_11131);
nor U13555 (N_13555,N_11986,N_10254);
nor U13556 (N_13556,N_11130,N_10184);
nand U13557 (N_13557,N_10503,N_10262);
and U13558 (N_13558,N_10041,N_10494);
xnor U13559 (N_13559,N_10791,N_11451);
nand U13560 (N_13560,N_10112,N_10987);
nor U13561 (N_13561,N_11853,N_11530);
or U13562 (N_13562,N_10646,N_10556);
and U13563 (N_13563,N_11524,N_10932);
and U13564 (N_13564,N_10474,N_11513);
nand U13565 (N_13565,N_11541,N_11350);
nor U13566 (N_13566,N_10545,N_10342);
and U13567 (N_13567,N_10360,N_10860);
and U13568 (N_13568,N_10241,N_11284);
nand U13569 (N_13569,N_10744,N_10297);
or U13570 (N_13570,N_10589,N_11990);
nor U13571 (N_13571,N_10154,N_10899);
nor U13572 (N_13572,N_11126,N_10311);
nor U13573 (N_13573,N_11020,N_10814);
nor U13574 (N_13574,N_11792,N_10318);
nor U13575 (N_13575,N_10739,N_11620);
and U13576 (N_13576,N_10145,N_11207);
and U13577 (N_13577,N_11563,N_11699);
or U13578 (N_13578,N_11900,N_11371);
nand U13579 (N_13579,N_10157,N_10520);
or U13580 (N_13580,N_10268,N_10922);
nand U13581 (N_13581,N_11108,N_11316);
or U13582 (N_13582,N_10325,N_10028);
or U13583 (N_13583,N_10507,N_10554);
and U13584 (N_13584,N_11134,N_11172);
nor U13585 (N_13585,N_10081,N_11177);
nand U13586 (N_13586,N_10781,N_11620);
and U13587 (N_13587,N_11189,N_10138);
or U13588 (N_13588,N_11138,N_11177);
and U13589 (N_13589,N_10743,N_10165);
or U13590 (N_13590,N_10374,N_11373);
nand U13591 (N_13591,N_11332,N_11013);
or U13592 (N_13592,N_10836,N_11306);
nor U13593 (N_13593,N_11263,N_10947);
nand U13594 (N_13594,N_11709,N_10856);
nand U13595 (N_13595,N_10919,N_10190);
and U13596 (N_13596,N_11399,N_11798);
nand U13597 (N_13597,N_11480,N_11273);
and U13598 (N_13598,N_10779,N_11978);
nor U13599 (N_13599,N_11765,N_11780);
and U13600 (N_13600,N_11932,N_11241);
nor U13601 (N_13601,N_11019,N_10895);
nand U13602 (N_13602,N_10386,N_10620);
nor U13603 (N_13603,N_11207,N_11449);
and U13604 (N_13604,N_11978,N_11662);
and U13605 (N_13605,N_10374,N_10205);
or U13606 (N_13606,N_10747,N_11667);
or U13607 (N_13607,N_10827,N_11748);
and U13608 (N_13608,N_10838,N_10112);
and U13609 (N_13609,N_11248,N_11880);
nor U13610 (N_13610,N_10429,N_11450);
and U13611 (N_13611,N_10167,N_11416);
nand U13612 (N_13612,N_10446,N_10066);
or U13613 (N_13613,N_11361,N_10535);
nor U13614 (N_13614,N_10695,N_11700);
nor U13615 (N_13615,N_11116,N_11800);
and U13616 (N_13616,N_11064,N_10666);
nand U13617 (N_13617,N_10391,N_10637);
nand U13618 (N_13618,N_10806,N_11942);
nor U13619 (N_13619,N_10043,N_11128);
and U13620 (N_13620,N_11764,N_10171);
nor U13621 (N_13621,N_11947,N_11627);
or U13622 (N_13622,N_10562,N_10054);
and U13623 (N_13623,N_11062,N_11052);
or U13624 (N_13624,N_11043,N_11904);
xor U13625 (N_13625,N_11300,N_10544);
and U13626 (N_13626,N_11227,N_10189);
and U13627 (N_13627,N_10887,N_10687);
nand U13628 (N_13628,N_11550,N_10081);
and U13629 (N_13629,N_10539,N_10125);
or U13630 (N_13630,N_10783,N_11523);
nor U13631 (N_13631,N_11392,N_11096);
nand U13632 (N_13632,N_10989,N_10793);
nand U13633 (N_13633,N_11002,N_11076);
nand U13634 (N_13634,N_11745,N_11937);
and U13635 (N_13635,N_11498,N_10576);
and U13636 (N_13636,N_11676,N_10609);
or U13637 (N_13637,N_11611,N_11729);
or U13638 (N_13638,N_11368,N_11133);
nor U13639 (N_13639,N_10493,N_10864);
nand U13640 (N_13640,N_11580,N_10358);
nor U13641 (N_13641,N_10075,N_10267);
and U13642 (N_13642,N_11640,N_11925);
and U13643 (N_13643,N_10610,N_11825);
and U13644 (N_13644,N_11509,N_10438);
or U13645 (N_13645,N_11853,N_11465);
and U13646 (N_13646,N_10319,N_10009);
or U13647 (N_13647,N_10040,N_10655);
nor U13648 (N_13648,N_10711,N_11156);
nand U13649 (N_13649,N_11320,N_10219);
or U13650 (N_13650,N_11552,N_11593);
and U13651 (N_13651,N_10944,N_10778);
nor U13652 (N_13652,N_11635,N_10420);
and U13653 (N_13653,N_10375,N_10583);
nor U13654 (N_13654,N_11093,N_10700);
nand U13655 (N_13655,N_10540,N_11162);
or U13656 (N_13656,N_11086,N_10114);
nand U13657 (N_13657,N_11108,N_11965);
nor U13658 (N_13658,N_10523,N_11184);
nand U13659 (N_13659,N_11649,N_11995);
nand U13660 (N_13660,N_10262,N_11094);
and U13661 (N_13661,N_10654,N_10603);
nor U13662 (N_13662,N_10456,N_10559);
or U13663 (N_13663,N_10423,N_11056);
and U13664 (N_13664,N_11435,N_10077);
or U13665 (N_13665,N_10231,N_10676);
nand U13666 (N_13666,N_11607,N_10242);
and U13667 (N_13667,N_10515,N_10114);
and U13668 (N_13668,N_10637,N_11734);
nand U13669 (N_13669,N_10157,N_11543);
and U13670 (N_13670,N_11994,N_11937);
nand U13671 (N_13671,N_10501,N_10968);
and U13672 (N_13672,N_11768,N_11810);
or U13673 (N_13673,N_10571,N_11368);
nand U13674 (N_13674,N_10802,N_11800);
or U13675 (N_13675,N_10581,N_10660);
nand U13676 (N_13676,N_11595,N_10323);
nor U13677 (N_13677,N_11420,N_10470);
nand U13678 (N_13678,N_11808,N_10965);
nand U13679 (N_13679,N_10851,N_11132);
nand U13680 (N_13680,N_10558,N_10138);
and U13681 (N_13681,N_11188,N_11976);
or U13682 (N_13682,N_11672,N_11771);
nand U13683 (N_13683,N_11487,N_11690);
nand U13684 (N_13684,N_10707,N_11254);
nand U13685 (N_13685,N_10261,N_11015);
or U13686 (N_13686,N_11530,N_10838);
and U13687 (N_13687,N_11853,N_11804);
nand U13688 (N_13688,N_11590,N_11879);
or U13689 (N_13689,N_11582,N_11017);
nor U13690 (N_13690,N_10045,N_11393);
or U13691 (N_13691,N_11871,N_11396);
nand U13692 (N_13692,N_10818,N_11653);
nand U13693 (N_13693,N_10090,N_10109);
and U13694 (N_13694,N_10586,N_11931);
and U13695 (N_13695,N_11970,N_10099);
or U13696 (N_13696,N_11699,N_10055);
nor U13697 (N_13697,N_10452,N_11775);
and U13698 (N_13698,N_10842,N_10573);
nor U13699 (N_13699,N_11401,N_10236);
nand U13700 (N_13700,N_11070,N_10970);
or U13701 (N_13701,N_10354,N_11561);
nor U13702 (N_13702,N_10606,N_11398);
nor U13703 (N_13703,N_10190,N_11133);
nor U13704 (N_13704,N_11777,N_11143);
nor U13705 (N_13705,N_11791,N_11581);
nor U13706 (N_13706,N_11415,N_10403);
nand U13707 (N_13707,N_11274,N_10031);
nand U13708 (N_13708,N_10272,N_10970);
nand U13709 (N_13709,N_11480,N_11911);
or U13710 (N_13710,N_10112,N_10004);
and U13711 (N_13711,N_10650,N_10599);
xnor U13712 (N_13712,N_11259,N_11543);
nor U13713 (N_13713,N_11530,N_10122);
xnor U13714 (N_13714,N_10785,N_11887);
nor U13715 (N_13715,N_11148,N_11776);
nor U13716 (N_13716,N_10298,N_11146);
nand U13717 (N_13717,N_11969,N_10744);
xnor U13718 (N_13718,N_11542,N_11497);
nor U13719 (N_13719,N_10302,N_11624);
and U13720 (N_13720,N_10611,N_10366);
and U13721 (N_13721,N_10253,N_11095);
nor U13722 (N_13722,N_11484,N_11636);
xnor U13723 (N_13723,N_10392,N_11400);
or U13724 (N_13724,N_11193,N_10324);
nand U13725 (N_13725,N_10125,N_10413);
nand U13726 (N_13726,N_10766,N_11972);
xnor U13727 (N_13727,N_10220,N_10338);
nand U13728 (N_13728,N_11661,N_11461);
nand U13729 (N_13729,N_10867,N_11418);
and U13730 (N_13730,N_11299,N_11831);
nand U13731 (N_13731,N_10477,N_11653);
and U13732 (N_13732,N_11998,N_10566);
xor U13733 (N_13733,N_11334,N_11279);
xor U13734 (N_13734,N_11612,N_10979);
and U13735 (N_13735,N_10864,N_11485);
nor U13736 (N_13736,N_11228,N_11963);
or U13737 (N_13737,N_10956,N_10616);
or U13738 (N_13738,N_10996,N_11868);
nand U13739 (N_13739,N_10715,N_11808);
nand U13740 (N_13740,N_10771,N_11450);
or U13741 (N_13741,N_11616,N_10701);
or U13742 (N_13742,N_11868,N_10700);
or U13743 (N_13743,N_11300,N_10561);
and U13744 (N_13744,N_10746,N_10477);
or U13745 (N_13745,N_10683,N_10273);
nor U13746 (N_13746,N_11646,N_10146);
and U13747 (N_13747,N_10444,N_11387);
nand U13748 (N_13748,N_11176,N_10725);
xor U13749 (N_13749,N_11558,N_11674);
or U13750 (N_13750,N_10102,N_11589);
nand U13751 (N_13751,N_10393,N_11212);
xnor U13752 (N_13752,N_10019,N_11010);
nand U13753 (N_13753,N_11314,N_10320);
nor U13754 (N_13754,N_10591,N_11026);
or U13755 (N_13755,N_10025,N_10436);
nor U13756 (N_13756,N_11906,N_10848);
nand U13757 (N_13757,N_10240,N_11892);
or U13758 (N_13758,N_10041,N_10226);
nand U13759 (N_13759,N_11950,N_11013);
and U13760 (N_13760,N_10232,N_11391);
or U13761 (N_13761,N_11607,N_11609);
xnor U13762 (N_13762,N_10043,N_11182);
nor U13763 (N_13763,N_10722,N_10039);
or U13764 (N_13764,N_10720,N_11371);
nor U13765 (N_13765,N_11542,N_10734);
nor U13766 (N_13766,N_11178,N_10014);
and U13767 (N_13767,N_10438,N_10214);
nor U13768 (N_13768,N_11420,N_11937);
or U13769 (N_13769,N_10686,N_10636);
nor U13770 (N_13770,N_11747,N_10016);
nand U13771 (N_13771,N_11752,N_11462);
nand U13772 (N_13772,N_11996,N_11710);
and U13773 (N_13773,N_11137,N_10793);
or U13774 (N_13774,N_11359,N_11268);
nand U13775 (N_13775,N_11358,N_11533);
nor U13776 (N_13776,N_11443,N_10728);
nand U13777 (N_13777,N_11900,N_11860);
or U13778 (N_13778,N_11388,N_11273);
or U13779 (N_13779,N_10046,N_11807);
nor U13780 (N_13780,N_11486,N_11203);
xnor U13781 (N_13781,N_10576,N_10387);
and U13782 (N_13782,N_10400,N_10281);
nor U13783 (N_13783,N_11270,N_11771);
and U13784 (N_13784,N_10199,N_10054);
and U13785 (N_13785,N_10304,N_10649);
nand U13786 (N_13786,N_10368,N_11702);
nor U13787 (N_13787,N_10291,N_11671);
and U13788 (N_13788,N_11871,N_10466);
nand U13789 (N_13789,N_10643,N_10680);
and U13790 (N_13790,N_11241,N_11849);
or U13791 (N_13791,N_11775,N_11682);
xor U13792 (N_13792,N_11293,N_10825);
xnor U13793 (N_13793,N_11007,N_10169);
xnor U13794 (N_13794,N_10451,N_11258);
and U13795 (N_13795,N_10475,N_10447);
nor U13796 (N_13796,N_11392,N_10950);
and U13797 (N_13797,N_10581,N_10343);
nor U13798 (N_13798,N_11768,N_10171);
and U13799 (N_13799,N_11791,N_10348);
nand U13800 (N_13800,N_11556,N_10608);
and U13801 (N_13801,N_10757,N_11646);
nand U13802 (N_13802,N_11944,N_11936);
and U13803 (N_13803,N_11517,N_11758);
nor U13804 (N_13804,N_11088,N_10469);
and U13805 (N_13805,N_10064,N_10631);
nand U13806 (N_13806,N_10988,N_11903);
and U13807 (N_13807,N_11229,N_10340);
or U13808 (N_13808,N_11352,N_10333);
and U13809 (N_13809,N_10906,N_11135);
and U13810 (N_13810,N_11093,N_11669);
nand U13811 (N_13811,N_10526,N_10421);
and U13812 (N_13812,N_10397,N_11023);
or U13813 (N_13813,N_10444,N_11784);
or U13814 (N_13814,N_10167,N_11388);
or U13815 (N_13815,N_11874,N_11022);
nand U13816 (N_13816,N_10282,N_11898);
and U13817 (N_13817,N_11934,N_11272);
or U13818 (N_13818,N_11033,N_11501);
nor U13819 (N_13819,N_11022,N_11965);
nor U13820 (N_13820,N_10273,N_11996);
nor U13821 (N_13821,N_10486,N_10667);
nor U13822 (N_13822,N_10144,N_10860);
nor U13823 (N_13823,N_11990,N_10853);
nor U13824 (N_13824,N_11086,N_11487);
or U13825 (N_13825,N_10322,N_10825);
nand U13826 (N_13826,N_10520,N_10982);
and U13827 (N_13827,N_10770,N_10599);
or U13828 (N_13828,N_11874,N_10121);
nand U13829 (N_13829,N_10678,N_11458);
nand U13830 (N_13830,N_10619,N_10282);
nor U13831 (N_13831,N_11237,N_10560);
or U13832 (N_13832,N_10651,N_11398);
or U13833 (N_13833,N_11734,N_10887);
or U13834 (N_13834,N_11649,N_10800);
nand U13835 (N_13835,N_11633,N_11001);
nand U13836 (N_13836,N_10427,N_11429);
and U13837 (N_13837,N_11506,N_10162);
and U13838 (N_13838,N_11210,N_10164);
nand U13839 (N_13839,N_11172,N_10001);
nand U13840 (N_13840,N_10413,N_11933);
nor U13841 (N_13841,N_10686,N_10504);
and U13842 (N_13842,N_11903,N_11500);
and U13843 (N_13843,N_11373,N_11298);
xnor U13844 (N_13844,N_11742,N_11612);
nor U13845 (N_13845,N_11413,N_10481);
nor U13846 (N_13846,N_11092,N_11666);
nand U13847 (N_13847,N_10315,N_10707);
or U13848 (N_13848,N_11071,N_10622);
or U13849 (N_13849,N_10108,N_10723);
nor U13850 (N_13850,N_11736,N_11078);
xor U13851 (N_13851,N_11300,N_10746);
or U13852 (N_13852,N_10923,N_11454);
nand U13853 (N_13853,N_10171,N_10741);
nand U13854 (N_13854,N_11088,N_10246);
or U13855 (N_13855,N_11153,N_10855);
or U13856 (N_13856,N_11111,N_10285);
and U13857 (N_13857,N_10197,N_11250);
nand U13858 (N_13858,N_11751,N_10456);
nand U13859 (N_13859,N_10239,N_10798);
or U13860 (N_13860,N_10365,N_10622);
and U13861 (N_13861,N_10899,N_11789);
nor U13862 (N_13862,N_11592,N_10600);
nand U13863 (N_13863,N_11436,N_10104);
nand U13864 (N_13864,N_10896,N_10789);
nor U13865 (N_13865,N_10324,N_10587);
and U13866 (N_13866,N_11492,N_10780);
or U13867 (N_13867,N_10374,N_10942);
nor U13868 (N_13868,N_11733,N_10104);
and U13869 (N_13869,N_10492,N_10255);
or U13870 (N_13870,N_10875,N_10754);
nand U13871 (N_13871,N_10766,N_11411);
nand U13872 (N_13872,N_11326,N_10701);
and U13873 (N_13873,N_10495,N_10812);
nor U13874 (N_13874,N_11712,N_11046);
or U13875 (N_13875,N_10312,N_10568);
and U13876 (N_13876,N_10513,N_10564);
nor U13877 (N_13877,N_10058,N_10170);
and U13878 (N_13878,N_10967,N_10868);
or U13879 (N_13879,N_11247,N_11510);
xnor U13880 (N_13880,N_11833,N_10104);
and U13881 (N_13881,N_10275,N_11832);
and U13882 (N_13882,N_11991,N_10396);
and U13883 (N_13883,N_10592,N_10935);
nor U13884 (N_13884,N_11767,N_11336);
nand U13885 (N_13885,N_10880,N_11586);
nand U13886 (N_13886,N_10233,N_10976);
or U13887 (N_13887,N_11711,N_10362);
nand U13888 (N_13888,N_11555,N_11667);
or U13889 (N_13889,N_11728,N_10289);
nor U13890 (N_13890,N_11728,N_11928);
nand U13891 (N_13891,N_10415,N_11412);
nand U13892 (N_13892,N_11644,N_10674);
xnor U13893 (N_13893,N_11515,N_11133);
and U13894 (N_13894,N_11551,N_11993);
and U13895 (N_13895,N_10960,N_10249);
nand U13896 (N_13896,N_10261,N_10522);
and U13897 (N_13897,N_11525,N_10531);
xnor U13898 (N_13898,N_11084,N_10477);
nand U13899 (N_13899,N_10271,N_11736);
nor U13900 (N_13900,N_10884,N_10044);
nor U13901 (N_13901,N_10867,N_11282);
nand U13902 (N_13902,N_10411,N_10055);
nor U13903 (N_13903,N_11499,N_11288);
nor U13904 (N_13904,N_10975,N_11996);
and U13905 (N_13905,N_11968,N_10694);
nor U13906 (N_13906,N_10304,N_11601);
xnor U13907 (N_13907,N_10843,N_10340);
and U13908 (N_13908,N_10586,N_10903);
nand U13909 (N_13909,N_10087,N_11463);
and U13910 (N_13910,N_11110,N_10039);
nand U13911 (N_13911,N_10160,N_10649);
nor U13912 (N_13912,N_11756,N_11865);
nand U13913 (N_13913,N_11899,N_10440);
nand U13914 (N_13914,N_10046,N_11459);
nand U13915 (N_13915,N_11132,N_11463);
nand U13916 (N_13916,N_11708,N_11005);
nand U13917 (N_13917,N_11009,N_10560);
nand U13918 (N_13918,N_10183,N_10629);
or U13919 (N_13919,N_10310,N_10790);
or U13920 (N_13920,N_11904,N_11289);
nand U13921 (N_13921,N_10276,N_11540);
and U13922 (N_13922,N_11571,N_11144);
nor U13923 (N_13923,N_10538,N_11936);
and U13924 (N_13924,N_10992,N_11648);
nor U13925 (N_13925,N_10468,N_10264);
nand U13926 (N_13926,N_11680,N_10740);
xor U13927 (N_13927,N_10776,N_11614);
and U13928 (N_13928,N_11815,N_11545);
nor U13929 (N_13929,N_10461,N_10919);
and U13930 (N_13930,N_10812,N_10859);
nand U13931 (N_13931,N_10950,N_11117);
or U13932 (N_13932,N_11214,N_11812);
or U13933 (N_13933,N_11859,N_11912);
nor U13934 (N_13934,N_10603,N_10163);
nor U13935 (N_13935,N_11705,N_10977);
or U13936 (N_13936,N_10438,N_10832);
and U13937 (N_13937,N_10161,N_10137);
nand U13938 (N_13938,N_10621,N_11831);
and U13939 (N_13939,N_10390,N_10949);
and U13940 (N_13940,N_10731,N_10981);
or U13941 (N_13941,N_11591,N_10625);
or U13942 (N_13942,N_10465,N_11482);
or U13943 (N_13943,N_11805,N_11451);
nor U13944 (N_13944,N_11636,N_11093);
and U13945 (N_13945,N_10042,N_10290);
or U13946 (N_13946,N_10506,N_10842);
nand U13947 (N_13947,N_11897,N_10377);
or U13948 (N_13948,N_11088,N_11541);
nand U13949 (N_13949,N_11134,N_11417);
nor U13950 (N_13950,N_11478,N_10102);
and U13951 (N_13951,N_10825,N_10448);
or U13952 (N_13952,N_11770,N_11613);
nor U13953 (N_13953,N_10329,N_11367);
nand U13954 (N_13954,N_10549,N_10653);
or U13955 (N_13955,N_11773,N_10835);
or U13956 (N_13956,N_11496,N_10525);
and U13957 (N_13957,N_11619,N_10678);
nand U13958 (N_13958,N_11651,N_10959);
and U13959 (N_13959,N_10082,N_10666);
or U13960 (N_13960,N_11505,N_10270);
or U13961 (N_13961,N_11597,N_10085);
nor U13962 (N_13962,N_10710,N_11727);
nor U13963 (N_13963,N_10608,N_10291);
nor U13964 (N_13964,N_11482,N_10431);
or U13965 (N_13965,N_11419,N_10442);
or U13966 (N_13966,N_10113,N_11953);
and U13967 (N_13967,N_11672,N_11026);
or U13968 (N_13968,N_11615,N_11605);
nor U13969 (N_13969,N_10978,N_10520);
nor U13970 (N_13970,N_11231,N_11546);
and U13971 (N_13971,N_11694,N_10382);
nor U13972 (N_13972,N_10559,N_10902);
nor U13973 (N_13973,N_11039,N_10036);
or U13974 (N_13974,N_10615,N_10922);
and U13975 (N_13975,N_10133,N_11226);
nand U13976 (N_13976,N_10818,N_10704);
nor U13977 (N_13977,N_10318,N_10951);
nand U13978 (N_13978,N_10598,N_10241);
and U13979 (N_13979,N_10112,N_11207);
or U13980 (N_13980,N_10298,N_10226);
or U13981 (N_13981,N_11988,N_10977);
or U13982 (N_13982,N_11465,N_10479);
and U13983 (N_13983,N_11880,N_11206);
or U13984 (N_13984,N_10942,N_10874);
nand U13985 (N_13985,N_11208,N_10333);
nand U13986 (N_13986,N_10323,N_10140);
or U13987 (N_13987,N_10512,N_10874);
nor U13988 (N_13988,N_11705,N_10900);
or U13989 (N_13989,N_11384,N_10616);
and U13990 (N_13990,N_10047,N_11694);
nand U13991 (N_13991,N_11444,N_10338);
or U13992 (N_13992,N_11622,N_11229);
and U13993 (N_13993,N_11171,N_10074);
nor U13994 (N_13994,N_10162,N_11651);
or U13995 (N_13995,N_11304,N_11786);
or U13996 (N_13996,N_10814,N_10358);
or U13997 (N_13997,N_10450,N_10130);
nand U13998 (N_13998,N_11928,N_10710);
nor U13999 (N_13999,N_11078,N_11126);
and U14000 (N_14000,N_13168,N_12467);
nand U14001 (N_14001,N_13285,N_12487);
and U14002 (N_14002,N_12660,N_12578);
and U14003 (N_14003,N_13846,N_12858);
and U14004 (N_14004,N_12838,N_13666);
and U14005 (N_14005,N_13665,N_12241);
and U14006 (N_14006,N_12419,N_13271);
nor U14007 (N_14007,N_13693,N_12523);
nand U14008 (N_14008,N_12230,N_12281);
nand U14009 (N_14009,N_12205,N_12980);
or U14010 (N_14010,N_12129,N_12007);
nor U14011 (N_14011,N_12783,N_13197);
nor U14012 (N_14012,N_13106,N_12184);
nor U14013 (N_14013,N_13873,N_13681);
nor U14014 (N_14014,N_13630,N_12508);
nand U14015 (N_14015,N_12801,N_13986);
and U14016 (N_14016,N_13469,N_13415);
and U14017 (N_14017,N_12163,N_13974);
and U14018 (N_14018,N_12485,N_13350);
or U14019 (N_14019,N_12320,N_13939);
nor U14020 (N_14020,N_13572,N_13828);
and U14021 (N_14021,N_12152,N_12536);
or U14022 (N_14022,N_12628,N_12583);
xnor U14023 (N_14023,N_13375,N_12438);
and U14024 (N_14024,N_13321,N_12121);
nand U14025 (N_14025,N_13006,N_13839);
nand U14026 (N_14026,N_12107,N_13274);
nand U14027 (N_14027,N_12826,N_13752);
nor U14028 (N_14028,N_12340,N_12076);
nor U14029 (N_14029,N_13998,N_12940);
nand U14030 (N_14030,N_12224,N_13568);
or U14031 (N_14031,N_13475,N_12965);
nand U14032 (N_14032,N_13709,N_13025);
and U14033 (N_14033,N_12469,N_13161);
and U14034 (N_14034,N_12183,N_12564);
and U14035 (N_14035,N_12011,N_13169);
or U14036 (N_14036,N_13145,N_12910);
or U14037 (N_14037,N_12461,N_12203);
nand U14038 (N_14038,N_13157,N_12214);
nor U14039 (N_14039,N_13774,N_12410);
nand U14040 (N_14040,N_13509,N_12997);
nor U14041 (N_14041,N_12913,N_13719);
nor U14042 (N_14042,N_12266,N_13066);
nand U14043 (N_14043,N_12159,N_13635);
nor U14044 (N_14044,N_13857,N_12416);
and U14045 (N_14045,N_12135,N_13526);
and U14046 (N_14046,N_13007,N_13311);
nor U14047 (N_14047,N_13448,N_12894);
nand U14048 (N_14048,N_13990,N_12659);
nor U14049 (N_14049,N_12324,N_13551);
or U14050 (N_14050,N_12992,N_12365);
and U14051 (N_14051,N_12207,N_12930);
nor U14052 (N_14052,N_13439,N_13513);
and U14053 (N_14053,N_12932,N_12554);
or U14054 (N_14054,N_13332,N_13878);
or U14055 (N_14055,N_13250,N_13421);
nand U14056 (N_14056,N_13139,N_12552);
or U14057 (N_14057,N_13823,N_12982);
nand U14058 (N_14058,N_12532,N_12585);
nor U14059 (N_14059,N_12069,N_13540);
or U14060 (N_14060,N_12041,N_12002);
nor U14061 (N_14061,N_13686,N_13435);
nor U14062 (N_14062,N_13026,N_12791);
or U14063 (N_14063,N_13201,N_13278);
nand U14064 (N_14064,N_12644,N_13223);
and U14065 (N_14065,N_13347,N_13362);
and U14066 (N_14066,N_13517,N_13736);
nand U14067 (N_14067,N_13726,N_13104);
or U14068 (N_14068,N_12465,N_12026);
nor U14069 (N_14069,N_13877,N_12453);
or U14070 (N_14070,N_12722,N_12418);
or U14071 (N_14071,N_12983,N_12031);
nor U14072 (N_14072,N_12223,N_13874);
nand U14073 (N_14073,N_12912,N_12767);
and U14074 (N_14074,N_13324,N_13925);
or U14075 (N_14075,N_13902,N_13587);
and U14076 (N_14076,N_12387,N_12968);
or U14077 (N_14077,N_13987,N_12926);
nand U14078 (N_14078,N_13247,N_12609);
or U14079 (N_14079,N_13956,N_13651);
and U14080 (N_14080,N_12287,N_13705);
and U14081 (N_14081,N_13413,N_12384);
nand U14082 (N_14082,N_13335,N_13267);
or U14083 (N_14083,N_12662,N_12579);
and U14084 (N_14084,N_12586,N_13617);
nand U14085 (N_14085,N_13804,N_13391);
and U14086 (N_14086,N_12004,N_12924);
and U14087 (N_14087,N_12096,N_13944);
xnor U14088 (N_14088,N_13239,N_13156);
and U14089 (N_14089,N_13142,N_13782);
nor U14090 (N_14090,N_12678,N_13794);
or U14091 (N_14091,N_13009,N_13395);
nor U14092 (N_14092,N_13042,N_12078);
or U14093 (N_14093,N_13253,N_12015);
nor U14094 (N_14094,N_12298,N_13141);
nand U14095 (N_14095,N_13124,N_12423);
nor U14096 (N_14096,N_13543,N_13763);
or U14097 (N_14097,N_12909,N_12645);
nor U14098 (N_14098,N_12428,N_13240);
nor U14099 (N_14099,N_12219,N_13359);
nand U14100 (N_14100,N_12346,N_13904);
or U14101 (N_14101,N_13633,N_12988);
and U14102 (N_14102,N_13649,N_13401);
or U14103 (N_14103,N_13638,N_12040);
and U14104 (N_14104,N_12702,N_13843);
or U14105 (N_14105,N_12788,N_12496);
or U14106 (N_14106,N_13631,N_12058);
nand U14107 (N_14107,N_12921,N_13648);
and U14108 (N_14108,N_12671,N_12746);
and U14109 (N_14109,N_13748,N_13487);
nand U14110 (N_14110,N_13099,N_12378);
or U14111 (N_14111,N_12080,N_13716);
or U14112 (N_14112,N_12302,N_12769);
or U14113 (N_14113,N_13871,N_13653);
and U14114 (N_14114,N_13833,N_12394);
and U14115 (N_14115,N_12435,N_12313);
or U14116 (N_14116,N_13452,N_12179);
nor U14117 (N_14117,N_12970,N_12650);
or U14118 (N_14118,N_12310,N_13030);
nand U14119 (N_14119,N_13641,N_12082);
nand U14120 (N_14120,N_12484,N_12326);
nand U14121 (N_14121,N_12314,N_13714);
nor U14122 (N_14122,N_13056,N_12831);
and U14123 (N_14123,N_13863,N_12717);
or U14124 (N_14124,N_12683,N_13268);
or U14125 (N_14125,N_12665,N_13565);
and U14126 (N_14126,N_12631,N_12502);
nor U14127 (N_14127,N_13672,N_12399);
and U14128 (N_14128,N_12236,N_13972);
nand U14129 (N_14129,N_13118,N_13047);
nand U14130 (N_14130,N_13144,N_12268);
nor U14131 (N_14131,N_12425,N_13573);
and U14132 (N_14132,N_13095,N_12250);
nand U14133 (N_14133,N_13241,N_13701);
and U14134 (N_14134,N_13928,N_12088);
nor U14135 (N_14135,N_13130,N_13361);
nor U14136 (N_14136,N_12882,N_12760);
nand U14137 (N_14137,N_13230,N_12775);
and U14138 (N_14138,N_13964,N_13249);
xor U14139 (N_14139,N_13154,N_13343);
nand U14140 (N_14140,N_12692,N_12871);
and U14141 (N_14141,N_12251,N_12466);
and U14142 (N_14142,N_12866,N_12855);
nor U14143 (N_14143,N_13379,N_12696);
and U14144 (N_14144,N_12613,N_12931);
nand U14145 (N_14145,N_12701,N_12049);
and U14146 (N_14146,N_12402,N_12571);
nor U14147 (N_14147,N_13720,N_13861);
and U14148 (N_14148,N_12807,N_12259);
nand U14149 (N_14149,N_13504,N_13731);
nor U14150 (N_14150,N_12663,N_12307);
nor U14151 (N_14151,N_13766,N_13708);
or U14152 (N_14152,N_13780,N_13417);
nand U14153 (N_14153,N_13847,N_12883);
nor U14154 (N_14154,N_12772,N_12367);
or U14155 (N_14155,N_13005,N_12561);
and U14156 (N_14156,N_13536,N_12518);
nand U14157 (N_14157,N_13560,N_13165);
and U14158 (N_14158,N_13880,N_13446);
or U14159 (N_14159,N_13498,N_13398);
and U14160 (N_14160,N_13558,N_12857);
or U14161 (N_14161,N_12208,N_13325);
and U14162 (N_14162,N_13741,N_12569);
nand U14163 (N_14163,N_12906,N_12110);
nand U14164 (N_14164,N_13858,N_13341);
or U14165 (N_14165,N_12376,N_12967);
or U14166 (N_14166,N_12265,N_13367);
nor U14167 (N_14167,N_12549,N_12584);
or U14168 (N_14168,N_13897,N_13948);
nand U14169 (N_14169,N_13835,N_13349);
and U14170 (N_14170,N_12424,N_13955);
nor U14171 (N_14171,N_13945,N_13192);
or U14172 (N_14172,N_12094,N_13967);
nor U14173 (N_14173,N_13221,N_12289);
nand U14174 (N_14174,N_12710,N_12821);
or U14175 (N_14175,N_12407,N_12217);
and U14176 (N_14176,N_12155,N_13205);
nor U14177 (N_14177,N_13992,N_13302);
and U14178 (N_14178,N_12477,N_13832);
or U14179 (N_14179,N_13266,N_13979);
nor U14180 (N_14180,N_13935,N_12182);
nor U14181 (N_14181,N_13834,N_13055);
and U14182 (N_14182,N_12503,N_12512);
or U14183 (N_14183,N_12869,N_12386);
and U14184 (N_14184,N_13788,N_12032);
nand U14185 (N_14185,N_12859,N_13771);
or U14186 (N_14186,N_12351,N_12133);
nand U14187 (N_14187,N_12501,N_12447);
and U14188 (N_14188,N_12150,N_13258);
nand U14189 (N_14189,N_13508,N_13661);
and U14190 (N_14190,N_12872,N_12669);
or U14191 (N_14191,N_12934,N_13209);
and U14192 (N_14192,N_12491,N_12830);
nand U14193 (N_14193,N_13767,N_12140);
or U14194 (N_14194,N_12810,N_13358);
nand U14195 (N_14195,N_13200,N_13078);
nor U14196 (N_14196,N_12846,N_13773);
or U14197 (N_14197,N_13203,N_12328);
or U14198 (N_14198,N_12527,N_13346);
or U14199 (N_14199,N_13123,N_13461);
and U14200 (N_14200,N_13533,N_12488);
and U14201 (N_14201,N_12691,N_12733);
or U14202 (N_14202,N_13656,N_13314);
nor U14203 (N_14203,N_13876,N_12030);
nor U14204 (N_14204,N_13229,N_13495);
nand U14205 (N_14205,N_13769,N_13962);
nand U14206 (N_14206,N_13381,N_12668);
nand U14207 (N_14207,N_13447,N_13492);
or U14208 (N_14208,N_13580,N_13330);
and U14209 (N_14209,N_12961,N_13818);
nor U14210 (N_14210,N_12945,N_13566);
nor U14211 (N_14211,N_13232,N_13569);
or U14212 (N_14212,N_12739,N_12306);
nor U14213 (N_14213,N_13520,N_13762);
nand U14214 (N_14214,N_12889,N_13400);
or U14215 (N_14215,N_12437,N_13930);
or U14216 (N_14216,N_12162,N_12500);
nor U14217 (N_14217,N_13734,N_12044);
and U14218 (N_14218,N_12835,N_13462);
and U14219 (N_14219,N_12641,N_13018);
and U14220 (N_14220,N_12526,N_13844);
nor U14221 (N_14221,N_12867,N_13336);
nand U14222 (N_14222,N_13899,N_12212);
and U14223 (N_14223,N_12101,N_12918);
nand U14224 (N_14224,N_12610,N_13942);
nor U14225 (N_14225,N_12352,N_13724);
nand U14226 (N_14226,N_12687,N_12765);
and U14227 (N_14227,N_12379,N_12812);
and U14228 (N_14228,N_13171,N_13685);
and U14229 (N_14229,N_13021,N_12881);
or U14230 (N_14230,N_12793,N_13723);
and U14231 (N_14231,N_12543,N_12548);
and U14232 (N_14232,N_13778,N_13973);
and U14233 (N_14233,N_12027,N_12618);
or U14234 (N_14234,N_12256,N_12242);
nor U14235 (N_14235,N_12648,N_13922);
nand U14236 (N_14236,N_13084,N_12651);
or U14237 (N_14237,N_12122,N_13254);
and U14238 (N_14238,N_13014,N_12361);
nor U14239 (N_14239,N_12360,N_13147);
and U14240 (N_14240,N_13287,N_13135);
nor U14241 (N_14241,N_12401,N_12167);
and U14242 (N_14242,N_13585,N_12270);
nor U14243 (N_14243,N_13372,N_12299);
and U14244 (N_14244,N_12226,N_13989);
nand U14245 (N_14245,N_13996,N_12837);
or U14246 (N_14246,N_12095,N_12892);
and U14247 (N_14247,N_12750,N_13983);
nor U14248 (N_14248,N_12814,N_13327);
nor U14249 (N_14249,N_13750,N_13959);
nor U14250 (N_14250,N_12354,N_12252);
nand U14251 (N_14251,N_13614,N_13176);
and U14252 (N_14252,N_13418,N_13451);
nor U14253 (N_14253,N_12600,N_12161);
xor U14254 (N_14254,N_12245,N_12603);
nor U14255 (N_14255,N_13597,N_13860);
or U14256 (N_14256,N_12178,N_12852);
and U14257 (N_14257,N_12994,N_13488);
nor U14258 (N_14258,N_12590,N_12978);
or U14259 (N_14259,N_13288,N_12398);
nor U14260 (N_14260,N_12559,N_12827);
nand U14261 (N_14261,N_13999,N_13941);
xnor U14262 (N_14262,N_13320,N_12470);
and U14263 (N_14263,N_13202,N_12781);
or U14264 (N_14264,N_12938,N_12146);
or U14265 (N_14265,N_12865,N_12596);
or U14266 (N_14266,N_12165,N_13473);
and U14267 (N_14267,N_12235,N_13991);
or U14268 (N_14268,N_13337,N_13982);
and U14269 (N_14269,N_12192,N_13669);
nand U14270 (N_14270,N_13386,N_12933);
or U14271 (N_14271,N_12958,N_12396);
and U14272 (N_14272,N_13465,N_13545);
nand U14273 (N_14273,N_13663,N_13235);
nand U14274 (N_14274,N_12278,N_12318);
and U14275 (N_14275,N_12064,N_13383);
and U14276 (N_14276,N_12305,N_13182);
nor U14277 (N_14277,N_13515,N_13091);
nor U14278 (N_14278,N_12533,N_12370);
nand U14279 (N_14279,N_13131,N_12777);
or U14280 (N_14280,N_13215,N_13261);
nand U14281 (N_14281,N_12634,N_13622);
and U14282 (N_14282,N_12332,N_12341);
nor U14283 (N_14283,N_13525,N_13159);
or U14284 (N_14284,N_12137,N_12694);
or U14285 (N_14285,N_12363,N_12144);
nand U14286 (N_14286,N_13751,N_12499);
and U14287 (N_14287,N_12276,N_12815);
or U14288 (N_14288,N_12718,N_13152);
nand U14289 (N_14289,N_12339,N_12462);
and U14290 (N_14290,N_13830,N_12784);
and U14291 (N_14291,N_12254,N_13694);
xor U14292 (N_14292,N_12685,N_12563);
or U14293 (N_14293,N_13153,N_12822);
nor U14294 (N_14294,N_13073,N_13997);
nand U14295 (N_14295,N_13053,N_13183);
nor U14296 (N_14296,N_13424,N_13329);
and U14297 (N_14297,N_13419,N_13514);
or U14298 (N_14298,N_12151,N_13707);
or U14299 (N_14299,N_13017,N_12130);
nor U14300 (N_14300,N_12464,N_13623);
or U14301 (N_14301,N_12751,N_13920);
nor U14302 (N_14302,N_12357,N_12322);
and U14303 (N_14303,N_12025,N_13554);
xor U14304 (N_14304,N_12635,N_12333);
or U14305 (N_14305,N_13425,N_13326);
nand U14306 (N_14306,N_13076,N_12656);
or U14307 (N_14307,N_12755,N_13575);
nor U14308 (N_14308,N_13454,N_12525);
or U14309 (N_14309,N_12055,N_12029);
or U14310 (N_14310,N_12917,N_13932);
nand U14311 (N_14311,N_12412,N_13339);
nand U14312 (N_14312,N_13069,N_13862);
or U14313 (N_14313,N_13746,N_13164);
nand U14314 (N_14314,N_13770,N_13364);
and U14315 (N_14315,N_12483,N_12726);
or U14316 (N_14316,N_12863,N_12524);
nor U14317 (N_14317,N_12492,N_13529);
nand U14318 (N_14318,N_13696,N_12850);
xnor U14319 (N_14319,N_12759,N_12991);
or U14320 (N_14320,N_13836,N_13260);
or U14321 (N_14321,N_12316,N_13033);
or U14322 (N_14322,N_12482,N_12218);
and U14323 (N_14323,N_12275,N_13371);
and U14324 (N_14324,N_13946,N_12787);
nor U14325 (N_14325,N_13096,N_13423);
and U14326 (N_14326,N_13875,N_12575);
nor U14327 (N_14327,N_13411,N_12238);
nor U14328 (N_14328,N_13039,N_12989);
nand U14329 (N_14329,N_12607,N_13115);
nand U14330 (N_14330,N_13518,N_13786);
and U14331 (N_14331,N_12890,N_13032);
nand U14332 (N_14332,N_13270,N_13706);
or U14333 (N_14333,N_12427,N_13403);
nor U14334 (N_14334,N_13604,N_13521);
nand U14335 (N_14335,N_12854,N_12381);
and U14336 (N_14336,N_12626,N_13754);
or U14337 (N_14337,N_13747,N_13976);
and U14338 (N_14338,N_12056,N_12795);
nand U14339 (N_14339,N_13655,N_13679);
nand U14340 (N_14340,N_13743,N_12836);
or U14341 (N_14341,N_13023,N_13660);
nand U14342 (N_14342,N_12369,N_13695);
xor U14343 (N_14343,N_12046,N_13943);
or U14344 (N_14344,N_13645,N_12963);
and U14345 (N_14345,N_13698,N_12560);
or U14346 (N_14346,N_12506,N_12808);
or U14347 (N_14347,N_12504,N_12581);
nor U14348 (N_14348,N_12068,N_13703);
nand U14349 (N_14349,N_12720,N_12842);
or U14350 (N_14350,N_12061,N_13700);
and U14351 (N_14351,N_12415,N_13310);
or U14352 (N_14352,N_13281,N_13909);
and U14353 (N_14353,N_12681,N_13355);
or U14354 (N_14354,N_12463,N_13378);
nor U14355 (N_14355,N_12849,N_12020);
nand U14356 (N_14356,N_13108,N_12771);
and U14357 (N_14357,N_12098,N_13792);
and U14358 (N_14358,N_12215,N_12422);
and U14359 (N_14359,N_12077,N_12293);
or U14360 (N_14360,N_13246,N_12630);
or U14361 (N_14361,N_13965,N_13603);
nor U14362 (N_14362,N_13901,N_13284);
nor U14363 (N_14363,N_13632,N_12962);
and U14364 (N_14364,N_12149,N_12105);
or U14365 (N_14365,N_12706,N_12716);
or U14366 (N_14366,N_12887,N_13801);
and U14367 (N_14367,N_13166,N_12377);
nand U14368 (N_14368,N_12216,N_12738);
nand U14369 (N_14369,N_13499,N_13412);
or U14370 (N_14370,N_12132,N_13644);
or U14371 (N_14371,N_13426,N_13789);
nor U14372 (N_14372,N_12770,N_13598);
or U14373 (N_14373,N_13718,N_13231);
and U14374 (N_14374,N_13879,N_13405);
xor U14375 (N_14375,N_12799,N_13890);
nand U14376 (N_14376,N_12395,N_13579);
nand U14377 (N_14377,N_13757,N_13065);
and U14378 (N_14378,N_13502,N_13307);
nor U14379 (N_14379,N_12478,N_12517);
nor U14380 (N_14380,N_13036,N_12951);
or U14381 (N_14381,N_12201,N_12421);
and U14382 (N_14382,N_13552,N_13211);
and U14383 (N_14383,N_13984,N_12390);
or U14384 (N_14384,N_12373,N_12019);
nand U14385 (N_14385,N_13228,N_13564);
and U14386 (N_14386,N_13352,N_13016);
nor U14387 (N_14387,N_13480,N_12338);
nand U14388 (N_14388,N_12345,N_13429);
or U14389 (N_14389,N_13914,N_13697);
nand U14390 (N_14390,N_13344,N_13460);
nand U14391 (N_14391,N_13810,N_13092);
or U14392 (N_14392,N_13219,N_12953);
nor U14393 (N_14393,N_13980,N_13994);
nand U14394 (N_14394,N_12944,N_12284);
nand U14395 (N_14395,N_13822,N_13220);
or U14396 (N_14396,N_13713,N_13969);
nand U14397 (N_14397,N_13402,N_12870);
or U14398 (N_14398,N_12344,N_12868);
and U14399 (N_14399,N_12758,N_13272);
and U14400 (N_14400,N_12556,N_12100);
nor U14401 (N_14401,N_12113,N_13783);
or U14402 (N_14402,N_13600,N_13082);
nor U14403 (N_14403,N_12493,N_12452);
or U14404 (N_14404,N_13732,N_13257);
nand U14405 (N_14405,N_12138,N_13457);
and U14406 (N_14406,N_12035,N_13584);
and U14407 (N_14407,N_12375,N_13855);
or U14408 (N_14408,N_12257,N_12763);
nor U14409 (N_14409,N_12005,N_12160);
nand U14410 (N_14410,N_12898,N_12582);
nor U14411 (N_14411,N_12321,N_13629);
nand U14412 (N_14412,N_13608,N_13808);
nor U14413 (N_14413,N_13127,N_12615);
or U14414 (N_14414,N_12774,N_12737);
nand U14415 (N_14415,N_13276,N_12756);
nor U14416 (N_14416,N_13592,N_13472);
nand U14417 (N_14417,N_12239,N_13385);
nor U14418 (N_14418,N_12145,N_12187);
and U14419 (N_14419,N_13668,N_13952);
and U14420 (N_14420,N_12206,N_12286);
nand U14421 (N_14421,N_13640,N_12253);
or U14422 (N_14422,N_12602,N_12118);
or U14423 (N_14423,N_12195,N_13134);
and U14424 (N_14424,N_13895,N_12786);
nor U14425 (N_14425,N_12747,N_12742);
and U14426 (N_14426,N_12877,N_12010);
nand U14427 (N_14427,N_13885,N_13081);
nor U14428 (N_14428,N_13802,N_12862);
nand U14429 (N_14429,N_12768,N_12753);
and U14430 (N_14430,N_12573,N_13158);
nand U14431 (N_14431,N_12511,N_12444);
nand U14432 (N_14432,N_12083,N_13322);
or U14433 (N_14433,N_12903,N_12432);
and U14434 (N_14434,N_12522,N_12975);
or U14435 (N_14435,N_13305,N_13530);
nor U14436 (N_14436,N_13599,N_13132);
nor U14437 (N_14437,N_12211,N_13671);
or U14438 (N_14438,N_12516,N_12247);
nand U14439 (N_14439,N_13328,N_12309);
or U14440 (N_14440,N_13527,N_12127);
nor U14441 (N_14441,N_13816,N_12947);
nor U14442 (N_14442,N_13667,N_13392);
or U14443 (N_14443,N_13826,N_13259);
or U14444 (N_14444,N_12404,N_12034);
and U14445 (N_14445,N_12723,N_12673);
nand U14446 (N_14446,N_13298,N_13122);
and U14447 (N_14447,N_13294,N_12530);
and U14448 (N_14448,N_12780,N_13044);
and U14449 (N_14449,N_12655,N_13756);
nor U14450 (N_14450,N_12979,N_13831);
nor U14451 (N_14451,N_12012,N_13620);
xnor U14452 (N_14452,N_12244,N_13216);
or U14453 (N_14453,N_13471,N_12383);
nor U14454 (N_14454,N_13315,N_13683);
nor U14455 (N_14455,N_12411,N_12606);
and U14456 (N_14456,N_13576,N_12672);
nor U14457 (N_14457,N_13796,N_13547);
or U14458 (N_14458,N_12841,N_12181);
nand U14459 (N_14459,N_12153,N_12649);
or U14460 (N_14460,N_12601,N_12697);
and U14461 (N_14461,N_12764,N_13674);
and U14462 (N_14462,N_13699,N_12274);
or U14463 (N_14463,N_12355,N_13595);
nand U14464 (N_14464,N_12232,N_12816);
or U14465 (N_14465,N_13704,N_13478);
nor U14466 (N_14466,N_12176,N_13582);
or U14467 (N_14467,N_13761,N_12893);
or U14468 (N_14468,N_12292,N_12368);
nor U14469 (N_14469,N_13865,N_12534);
or U14470 (N_14470,N_13848,N_12426);
and U14471 (N_14471,N_13390,N_12175);
or U14472 (N_14472,N_12169,N_12013);
nor U14473 (N_14473,N_12874,N_12018);
nor U14474 (N_14474,N_13290,N_12599);
or U14475 (N_14475,N_12562,N_12999);
nand U14476 (N_14476,N_13279,N_13970);
or U14477 (N_14477,N_13217,N_13243);
or U14478 (N_14478,N_12342,N_12695);
nand U14479 (N_14479,N_13966,N_12356);
nor U14480 (N_14480,N_13126,N_12897);
and U14481 (N_14481,N_13917,N_12172);
nor U14482 (N_14482,N_13366,N_13975);
nor U14483 (N_14483,N_13926,N_12228);
nor U14484 (N_14484,N_13434,N_13179);
nand U14485 (N_14485,N_13800,N_12832);
and U14486 (N_14486,N_12762,N_13275);
and U14487 (N_14487,N_13170,N_12164);
and U14488 (N_14488,N_12014,N_13758);
or U14489 (N_14489,N_13299,N_12661);
nand U14490 (N_14490,N_13357,N_13483);
or U14491 (N_14491,N_13040,N_12053);
and U14492 (N_14492,N_12006,N_12984);
and U14493 (N_14493,N_12577,N_12824);
xor U14494 (N_14494,N_12490,N_12120);
nor U14495 (N_14495,N_12246,N_12269);
nor U14496 (N_14496,N_13851,N_13181);
xnor U14497 (N_14497,N_13577,N_12108);
nand U14498 (N_14498,N_13236,N_13376);
and U14499 (N_14499,N_12704,N_13531);
or U14500 (N_14500,N_13721,N_12594);
nand U14501 (N_14501,N_12380,N_13618);
nor U14502 (N_14502,N_13803,N_13397);
nand U14503 (N_14503,N_12705,N_12900);
nor U14504 (N_14504,N_13760,N_13121);
or U14505 (N_14505,N_13059,N_12388);
nor U14506 (N_14506,N_12896,N_13195);
and U14507 (N_14507,N_13918,N_13348);
nor U14508 (N_14508,N_13870,N_12180);
nor U14509 (N_14509,N_13916,N_13610);
and U14510 (N_14510,N_13884,N_12986);
nor U14511 (N_14511,N_13430,N_12093);
nand U14512 (N_14512,N_13555,N_12899);
or U14513 (N_14513,N_12147,N_13072);
nand U14514 (N_14514,N_12358,N_13813);
xnor U14515 (N_14515,N_13553,N_13812);
and U14516 (N_14516,N_13226,N_12173);
nand U14517 (N_14517,N_12675,N_12204);
nand U14518 (N_14518,N_12392,N_12553);
nand U14519 (N_14519,N_13109,N_12680);
or U14520 (N_14520,N_12170,N_12519);
and U14521 (N_14521,N_13467,N_13840);
nor U14522 (N_14522,N_12017,N_12497);
or U14523 (N_14523,N_12789,N_13048);
and U14524 (N_14524,N_13459,N_13012);
nand U14525 (N_14525,N_12263,N_12194);
and U14526 (N_14526,N_13814,N_12325);
or U14527 (N_14527,N_12636,N_13008);
xor U14528 (N_14528,N_12457,N_13180);
and U14529 (N_14529,N_12956,N_12022);
and U14530 (N_14530,N_13837,N_12290);
and U14531 (N_14531,N_13938,N_12486);
nand U14532 (N_14532,N_13850,N_13208);
or U14533 (N_14533,N_13589,N_13896);
or U14534 (N_14534,N_13729,N_13297);
and U14535 (N_14535,N_12288,N_12752);
nor U14536 (N_14536,N_12740,N_12796);
nand U14537 (N_14537,N_12168,N_13609);
nor U14538 (N_14538,N_12067,N_13416);
nand U14539 (N_14539,N_13510,N_12736);
nor U14540 (N_14540,N_12699,N_12608);
or U14541 (N_14541,N_13887,N_12943);
and U14542 (N_14542,N_13245,N_12729);
and U14543 (N_14543,N_12389,N_13308);
or U14544 (N_14544,N_13331,N_12627);
nor U14545 (N_14545,N_12529,N_13541);
or U14546 (N_14546,N_13913,N_12901);
or U14547 (N_14547,N_12703,N_12198);
nand U14548 (N_14548,N_13643,N_13316);
and U14549 (N_14549,N_13881,N_12923);
nor U14550 (N_14550,N_13995,N_12301);
nor U14551 (N_14551,N_13639,N_12948);
nand U14552 (N_14552,N_13776,N_13912);
xor U14553 (N_14553,N_12191,N_12126);
or U14554 (N_14554,N_13854,N_12928);
or U14555 (N_14555,N_13503,N_13002);
nand U14556 (N_14556,N_13606,N_12277);
or U14557 (N_14557,N_12714,N_12942);
or U14558 (N_14558,N_12875,N_13440);
nand U14559 (N_14559,N_13849,N_13041);
nand U14560 (N_14560,N_12657,N_12479);
nand U14561 (N_14561,N_13485,N_13781);
xor U14562 (N_14562,N_12079,N_13000);
nor U14563 (N_14563,N_13301,N_13466);
nand U14564 (N_14564,N_13470,N_13433);
nand U14565 (N_14565,N_13049,N_12790);
or U14566 (N_14566,N_12036,N_13712);
nor U14567 (N_14567,N_12063,N_13866);
nand U14568 (N_14568,N_12220,N_12589);
xnor U14569 (N_14569,N_13688,N_13252);
nor U14570 (N_14570,N_13523,N_13657);
nand U14571 (N_14571,N_13934,N_13950);
or U14572 (N_14572,N_12234,N_12177);
nand U14573 (N_14573,N_12513,N_12920);
nand U14574 (N_14574,N_12397,N_12713);
nor U14575 (N_14575,N_12449,N_12674);
xnor U14576 (N_14576,N_12653,N_12474);
nor U14577 (N_14577,N_12123,N_12915);
nor U14578 (N_14578,N_12642,N_12454);
and U14579 (N_14579,N_13151,N_12828);
and U14580 (N_14580,N_12558,N_12757);
nor U14581 (N_14581,N_13450,N_13054);
nor U14582 (N_14582,N_13393,N_12337);
nand U14583 (N_14583,N_13787,N_13199);
nor U14584 (N_14584,N_12853,N_13213);
nor U14585 (N_14585,N_12054,N_13711);
nand U14586 (N_14586,N_12825,N_13027);
nor U14587 (N_14587,N_12335,N_12319);
nand U14588 (N_14588,N_12766,N_12851);
and U14589 (N_14589,N_12124,N_12919);
and U14590 (N_14590,N_12735,N_12185);
or U14591 (N_14591,N_13951,N_12102);
nor U14592 (N_14592,N_13841,N_12542);
nor U14593 (N_14593,N_12861,N_12433);
and U14594 (N_14594,N_12878,N_13024);
or U14595 (N_14595,N_13993,N_13586);
and U14596 (N_14596,N_13805,N_13856);
and U14597 (N_14597,N_13627,N_13702);
or U14598 (N_14598,N_12544,N_12570);
or U14599 (N_14599,N_12408,N_13210);
and U14600 (N_14600,N_12834,N_13692);
or U14601 (N_14601,N_13689,N_12291);
or U14602 (N_14602,N_12406,N_12249);
or U14603 (N_14603,N_13728,N_13512);
or U14604 (N_14604,N_12640,N_12413);
and U14605 (N_14605,N_13981,N_12000);
nor U14606 (N_14606,N_13029,N_12450);
or U14607 (N_14607,N_12954,N_13162);
and U14608 (N_14608,N_13280,N_13571);
or U14609 (N_14609,N_13143,N_12860);
nor U14610 (N_14610,N_13915,N_13759);
or U14611 (N_14611,N_12231,N_13742);
or U14612 (N_14612,N_13494,N_12654);
and U14613 (N_14613,N_13458,N_12595);
or U14614 (N_14614,N_12847,N_12621);
or U14615 (N_14615,N_13407,N_13167);
and U14616 (N_14616,N_13957,N_13406);
nand U14617 (N_14617,N_12964,N_13825);
and U14618 (N_14618,N_13624,N_12028);
and U14619 (N_14619,N_13768,N_13105);
or U14620 (N_14620,N_13085,N_12403);
or U14621 (N_14621,N_13368,N_12065);
and U14622 (N_14622,N_13562,N_13206);
nand U14623 (N_14623,N_12604,N_13684);
nor U14624 (N_14624,N_13790,N_12666);
nor U14625 (N_14625,N_13737,N_13111);
nand U14626 (N_14626,N_13043,N_12317);
nor U14627 (N_14627,N_13262,N_12261);
and U14628 (N_14628,N_12873,N_12264);
and U14629 (N_14629,N_13534,N_12876);
nand U14630 (N_14630,N_12131,N_12633);
and U14631 (N_14631,N_12073,N_13538);
xnor U14632 (N_14632,N_13738,N_13384);
xnor U14633 (N_14633,N_12950,N_13616);
and U14634 (N_14634,N_13273,N_13615);
or U14635 (N_14635,N_13227,N_13650);
xnor U14636 (N_14636,N_13034,N_13497);
nand U14637 (N_14637,N_13125,N_13893);
and U14638 (N_14638,N_13612,N_12071);
nor U14639 (N_14639,N_13178,N_12436);
nand U14640 (N_14640,N_12547,N_13455);
nand U14641 (N_14641,N_12844,N_12473);
xor U14642 (N_14642,N_13978,N_13086);
or U14643 (N_14643,N_12248,N_13468);
or U14644 (N_14644,N_12086,N_13408);
nand U14645 (N_14645,N_12537,N_12619);
and U14646 (N_14646,N_13177,N_12304);
nand U14647 (N_14647,N_12362,N_12001);
nor U14648 (N_14648,N_12374,N_13730);
or U14649 (N_14649,N_12743,N_13590);
and U14650 (N_14650,N_12611,N_13404);
or U14651 (N_14651,N_12985,N_13333);
nor U14652 (N_14652,N_12895,N_13593);
and U14653 (N_14653,N_13882,N_12353);
or U14654 (N_14654,N_13140,N_12545);
or U14655 (N_14655,N_13785,N_12455);
nor U14656 (N_14656,N_12243,N_12442);
or U14657 (N_14657,N_12202,N_12282);
nand U14658 (N_14658,N_13581,N_12143);
and U14659 (N_14659,N_12712,N_12057);
nor U14660 (N_14660,N_12535,N_12623);
and U14661 (N_14661,N_13292,N_12748);
nand U14662 (N_14662,N_13464,N_12916);
and U14663 (N_14663,N_13570,N_12476);
and U14664 (N_14664,N_12688,N_13443);
nand U14665 (N_14665,N_12431,N_13775);
nor U14666 (N_14666,N_13908,N_12708);
and U14667 (N_14667,N_12038,N_13432);
or U14668 (N_14668,N_13764,N_12744);
nand U14669 (N_14669,N_13037,N_12498);
nor U14670 (N_14670,N_13382,N_13093);
nand U14671 (N_14671,N_12188,N_13437);
nor U14672 (N_14672,N_13845,N_13351);
nor U14673 (N_14673,N_13251,N_12272);
nand U14674 (N_14674,N_12489,N_13340);
nor U14675 (N_14675,N_12089,N_12295);
nand U14676 (N_14676,N_13658,N_12097);
or U14677 (N_14677,N_12798,N_12114);
nor U14678 (N_14678,N_13119,N_12009);
nor U14679 (N_14679,N_13755,N_13185);
or U14680 (N_14680,N_13463,N_12062);
nand U14681 (N_14681,N_12166,N_12066);
and U14682 (N_14682,N_13486,N_13677);
or U14683 (N_14683,N_13516,N_13690);
and U14684 (N_14684,N_13410,N_13652);
nand U14685 (N_14685,N_13654,N_12620);
nand U14686 (N_14686,N_12136,N_12514);
or U14687 (N_14687,N_12134,N_13634);
and U14688 (N_14688,N_12255,N_12084);
nor U14689 (N_14689,N_12990,N_13365);
and U14690 (N_14690,N_12521,N_13422);
nand U14691 (N_14691,N_13559,N_13753);
and U14692 (N_14692,N_13815,N_13662);
nor U14693 (N_14693,N_13772,N_13594);
nor U14694 (N_14694,N_12052,N_12125);
nand U14695 (N_14695,N_12813,N_12441);
or U14696 (N_14696,N_13088,N_13196);
and U14697 (N_14697,N_13601,N_13636);
nor U14698 (N_14698,N_13050,N_13524);
or U14699 (N_14699,N_12567,N_13449);
or U14700 (N_14700,N_12572,N_12949);
nor U14701 (N_14701,N_13493,N_13563);
or U14702 (N_14702,N_12664,N_13637);
nand U14703 (N_14703,N_13682,N_13283);
or U14704 (N_14704,N_13149,N_13838);
and U14705 (N_14705,N_13484,N_12409);
and U14706 (N_14706,N_12686,N_12331);
nor U14707 (N_14707,N_12271,N_13621);
nor U14708 (N_14708,N_12315,N_13172);
nand U14709 (N_14709,N_13811,N_13160);
and U14710 (N_14710,N_12460,N_13872);
and U14711 (N_14711,N_13557,N_12300);
nor U14712 (N_14712,N_12580,N_13146);
or U14713 (N_14713,N_13074,N_13377);
and U14714 (N_14714,N_12612,N_13456);
or U14715 (N_14715,N_12043,N_12154);
xor U14716 (N_14716,N_13710,N_13820);
and U14717 (N_14717,N_12481,N_13175);
nor U14718 (N_14718,N_12196,N_12364);
and U14719 (N_14719,N_13101,N_12914);
nand U14720 (N_14720,N_13063,N_12797);
or U14721 (N_14721,N_12366,N_12646);
or U14722 (N_14722,N_13356,N_12109);
nor U14723 (N_14723,N_13868,N_13607);
or U14724 (N_14724,N_13296,N_12042);
xnor U14725 (N_14725,N_13481,N_13222);
or U14726 (N_14726,N_12509,N_12959);
or U14727 (N_14727,N_12528,N_13988);
nand U14728 (N_14728,N_13374,N_12565);
or U14729 (N_14729,N_12539,N_13256);
and U14730 (N_14730,N_12385,N_12864);
nor U14731 (N_14731,N_13799,N_12566);
nand U14732 (N_14732,N_13057,N_12142);
and U14733 (N_14733,N_13626,N_13903);
nand U14734 (N_14734,N_13113,N_13052);
nor U14735 (N_14735,N_12260,N_13548);
and U14736 (N_14736,N_12856,N_12116);
nor U14737 (N_14737,N_13323,N_12280);
and U14738 (N_14738,N_12727,N_13338);
nand U14739 (N_14739,N_13100,N_13441);
and U14740 (N_14740,N_13490,N_12792);
nand U14741 (N_14741,N_13479,N_12617);
nor U14742 (N_14742,N_13295,N_12707);
or U14743 (N_14743,N_13075,N_12778);
nand U14744 (N_14744,N_12805,N_12800);
nand U14745 (N_14745,N_12059,N_12391);
or U14746 (N_14746,N_12885,N_12724);
nor U14747 (N_14747,N_12818,N_13907);
and U14748 (N_14748,N_12520,N_12719);
nor U14749 (N_14749,N_13237,N_13539);
or U14750 (N_14750,N_12106,N_12343);
or U14751 (N_14751,N_12622,N_12741);
nand U14752 (N_14752,N_12996,N_12085);
nand U14753 (N_14753,N_13186,N_12475);
nor U14754 (N_14754,N_12731,N_12957);
xor U14755 (N_14755,N_13574,N_13954);
and U14756 (N_14756,N_12393,N_12471);
nand U14757 (N_14757,N_13807,N_13137);
or U14758 (N_14758,N_13038,N_13958);
nor U14759 (N_14759,N_13387,N_13605);
or U14760 (N_14760,N_13817,N_13136);
or U14761 (N_14761,N_13189,N_13675);
and U14762 (N_14762,N_13242,N_12051);
nor U14763 (N_14763,N_12715,N_13013);
nand U14764 (N_14764,N_12658,N_12285);
or U14765 (N_14765,N_13507,N_13544);
nor U14766 (N_14766,N_12888,N_13098);
nor U14767 (N_14767,N_12540,N_13691);
nor U14768 (N_14768,N_12946,N_12803);
and U14769 (N_14769,N_13342,N_12448);
nor U14770 (N_14770,N_13898,N_13212);
and U14771 (N_14771,N_12199,N_12451);
nor U14772 (N_14772,N_12682,N_13353);
or U14773 (N_14773,N_12210,N_13264);
xnor U14774 (N_14774,N_13673,N_13567);
and U14775 (N_14775,N_13960,N_12927);
nor U14776 (N_14776,N_12848,N_12952);
and U14777 (N_14777,N_12977,N_12405);
nand U14778 (N_14778,N_13427,N_12443);
or U14779 (N_14779,N_13313,N_13546);
nor U14780 (N_14780,N_13791,N_12336);
and U14781 (N_14781,N_13797,N_12128);
nor U14782 (N_14782,N_13318,N_12117);
or U14783 (N_14783,N_12976,N_12922);
nor U14784 (N_14784,N_13070,N_13596);
and U14785 (N_14785,N_12221,N_13373);
nand U14786 (N_14786,N_12969,N_12939);
nor U14787 (N_14787,N_13233,N_12823);
nand U14788 (N_14788,N_12839,N_12267);
nand U14789 (N_14789,N_13064,N_12531);
and U14790 (N_14790,N_13004,N_13354);
nand U14791 (N_14791,N_12400,N_12625);
or U14792 (N_14792,N_13911,N_13187);
nand U14793 (N_14793,N_13046,N_13619);
or U14794 (N_14794,N_13438,N_13319);
nor U14795 (N_14795,N_12785,N_13798);
and U14796 (N_14796,N_12229,N_12709);
nor U14797 (N_14797,N_13282,N_13806);
xnor U14798 (N_14798,N_13080,N_12222);
nand U14799 (N_14799,N_12884,N_13399);
nand U14800 (N_14800,N_13784,N_13071);
nor U14801 (N_14801,N_13910,N_12190);
and U14802 (N_14802,N_12891,N_12700);
nand U14803 (N_14803,N_12074,N_12782);
and U14804 (N_14804,N_13103,N_13511);
or U14805 (N_14805,N_12732,N_12639);
or U14806 (N_14806,N_12941,N_13937);
nor U14807 (N_14807,N_12200,N_13923);
nand U14808 (N_14808,N_12279,N_13188);
or U14809 (N_14809,N_13889,N_13010);
nand U14810 (N_14810,N_12186,N_13953);
or U14811 (N_14811,N_13061,N_13090);
nand U14812 (N_14812,N_13117,N_12225);
nor U14813 (N_14813,N_12981,N_12227);
and U14814 (N_14814,N_13409,N_13924);
nor U14815 (N_14815,N_13089,N_13022);
nor U14816 (N_14816,N_12294,N_12624);
or U14817 (N_14817,N_13853,N_12845);
nor U14818 (N_14818,N_13864,N_12330);
or U14819 (N_14819,N_13277,N_13163);
xor U14820 (N_14820,N_12629,N_13148);
and U14821 (N_14821,N_12139,N_12303);
nor U14822 (N_14822,N_13225,N_13001);
nor U14823 (N_14823,N_13128,N_12698);
and U14824 (N_14824,N_12037,N_12417);
nand U14825 (N_14825,N_12327,N_12574);
nor U14826 (N_14826,N_12987,N_13528);
nor U14827 (N_14827,N_12904,N_12843);
and U14828 (N_14828,N_13501,N_12045);
or U14829 (N_14829,N_12016,N_12480);
or U14830 (N_14830,N_13133,N_13428);
nor U14831 (N_14831,N_12262,N_12157);
or U14832 (N_14832,N_13060,N_12779);
nor U14833 (N_14833,N_12430,N_13611);
or U14834 (N_14834,N_13491,N_13191);
nor U14835 (N_14835,N_13370,N_13112);
nand U14836 (N_14836,N_12446,N_12047);
nor U14837 (N_14837,N_12907,N_12197);
nor U14838 (N_14838,N_12972,N_13476);
nand U14839 (N_14839,N_12515,N_12081);
nor U14840 (N_14840,N_13028,N_13900);
nand U14841 (N_14841,N_12806,N_13224);
and U14842 (N_14842,N_12754,N_12911);
nor U14843 (N_14843,N_13602,N_13204);
nand U14844 (N_14844,N_13613,N_12557);
nor U14845 (N_14845,N_13094,N_12350);
nand U14846 (N_14846,N_12060,N_12935);
or U14847 (N_14847,N_13248,N_13985);
nor U14848 (N_14848,N_13888,N_13207);
or U14849 (N_14849,N_12329,N_13727);
nor U14850 (N_14850,N_13031,N_13214);
and U14851 (N_14851,N_13929,N_12880);
nor U14852 (N_14852,N_13363,N_13345);
or U14853 (N_14853,N_13255,N_13646);
and U14854 (N_14854,N_13369,N_12677);
and U14855 (N_14855,N_13150,N_13535);
nand U14856 (N_14856,N_12308,N_12749);
nand U14857 (N_14857,N_13676,N_13809);
or U14858 (N_14858,N_13444,N_13765);
nand U14859 (N_14859,N_13289,N_13194);
xnor U14860 (N_14860,N_12679,N_13110);
or U14861 (N_14861,N_13869,N_13414);
nor U14862 (N_14862,N_12008,N_12745);
nand U14863 (N_14863,N_13174,N_12349);
nand U14864 (N_14864,N_13793,N_12273);
nand U14865 (N_14865,N_13442,N_13129);
and U14866 (N_14866,N_13733,N_13474);
or U14867 (N_14867,N_12734,N_12546);
nor U14868 (N_14868,N_12616,N_12297);
nor U14869 (N_14869,N_12111,N_12156);
nor U14870 (N_14870,N_13919,N_12382);
nor U14871 (N_14871,N_13067,N_13380);
or U14872 (N_14872,N_13715,N_12296);
nand U14873 (N_14873,N_12023,N_13931);
or U14874 (N_14874,N_12761,N_12439);
and U14875 (N_14875,N_12725,N_13303);
nand U14876 (N_14876,N_13334,N_13360);
nor U14877 (N_14877,N_13051,N_13522);
nand U14878 (N_14878,N_13735,N_12936);
nand U14879 (N_14879,N_13819,N_12039);
or U14880 (N_14880,N_13218,N_12024);
nand U14881 (N_14881,N_12359,N_12598);
nand U14882 (N_14882,N_12588,N_13827);
nand U14883 (N_14883,N_13628,N_13961);
nand U14884 (N_14884,N_13453,N_12960);
nand U14885 (N_14885,N_12112,N_12075);
xnor U14886 (N_14886,N_13678,N_12614);
xnor U14887 (N_14887,N_12587,N_12494);
nand U14888 (N_14888,N_12092,N_12647);
and U14889 (N_14889,N_12551,N_13542);
or U14890 (N_14890,N_12937,N_12905);
and U14891 (N_14891,N_13198,N_12240);
nand U14892 (N_14892,N_12721,N_13963);
or U14893 (N_14893,N_12652,N_12070);
or U14894 (N_14894,N_12643,N_12141);
nand U14895 (N_14895,N_13725,N_12171);
or U14896 (N_14896,N_13120,N_13389);
and U14897 (N_14897,N_12879,N_13949);
and U14898 (N_14898,N_13114,N_12033);
nand U14899 (N_14899,N_12148,N_13906);
nand U14900 (N_14900,N_13291,N_12811);
nor U14901 (N_14901,N_13500,N_12458);
nand U14902 (N_14902,N_12237,N_12495);
or U14903 (N_14903,N_13583,N_13482);
or U14904 (N_14904,N_12819,N_13269);
and U14905 (N_14905,N_12820,N_12817);
nor U14906 (N_14906,N_13561,N_13821);
or U14907 (N_14907,N_12048,N_13647);
or U14908 (N_14908,N_12468,N_12804);
nor U14909 (N_14909,N_13779,N_12115);
and U14910 (N_14910,N_13940,N_12311);
nand U14911 (N_14911,N_12445,N_13933);
and U14912 (N_14912,N_12676,N_12103);
and U14913 (N_14913,N_13537,N_12158);
and U14914 (N_14914,N_13744,N_13062);
or U14915 (N_14915,N_12050,N_13077);
nand U14916 (N_14916,N_12605,N_13777);
and U14917 (N_14917,N_12902,N_12925);
nand U14918 (N_14918,N_12993,N_12420);
nand U14919 (N_14919,N_12995,N_12728);
or U14920 (N_14920,N_12693,N_12119);
nand U14921 (N_14921,N_12334,N_12091);
and U14922 (N_14922,N_13293,N_13396);
xor U14923 (N_14923,N_12773,N_12638);
nand U14924 (N_14924,N_13859,N_12213);
and U14925 (N_14925,N_13489,N_13977);
xor U14926 (N_14926,N_13588,N_13107);
nand U14927 (N_14927,N_12555,N_12632);
nor U14928 (N_14928,N_13852,N_12684);
nand U14929 (N_14929,N_13886,N_13436);
nor U14930 (N_14930,N_13011,N_13306);
and U14931 (N_14931,N_13687,N_12711);
or U14932 (N_14932,N_13717,N_13102);
nor U14933 (N_14933,N_12929,N_12472);
and U14934 (N_14934,N_13019,N_13921);
nor U14935 (N_14935,N_12829,N_12689);
nor U14936 (N_14936,N_13971,N_13947);
or U14937 (N_14937,N_12456,N_12510);
nor U14938 (N_14938,N_12072,N_13905);
and U14939 (N_14939,N_12347,N_13193);
nand U14940 (N_14940,N_13578,N_13087);
xor U14941 (N_14941,N_12258,N_13388);
nand U14942 (N_14942,N_13892,N_12802);
and U14943 (N_14943,N_13968,N_13625);
nor U14944 (N_14944,N_12087,N_12090);
nor U14945 (N_14945,N_13234,N_12973);
and U14946 (N_14946,N_12833,N_13015);
nor U14947 (N_14947,N_12886,N_13003);
nand U14948 (N_14948,N_13312,N_13317);
or U14949 (N_14949,N_12440,N_13184);
and U14950 (N_14950,N_12966,N_13155);
nand U14951 (N_14951,N_13506,N_12459);
nor U14952 (N_14952,N_12312,N_13286);
or U14953 (N_14953,N_13829,N_12597);
or U14954 (N_14954,N_12809,N_12550);
and U14955 (N_14955,N_12323,N_12730);
nor U14956 (N_14956,N_13477,N_13739);
xor U14957 (N_14957,N_13035,N_13263);
or U14958 (N_14958,N_13083,N_13173);
nand U14959 (N_14959,N_12003,N_13309);
or U14960 (N_14960,N_13549,N_13722);
and U14961 (N_14961,N_12667,N_13680);
nor U14962 (N_14962,N_13420,N_12593);
nor U14963 (N_14963,N_12955,N_13058);
nor U14964 (N_14964,N_12576,N_13936);
and U14965 (N_14965,N_12209,N_12974);
and U14966 (N_14966,N_13795,N_12908);
nand U14967 (N_14967,N_13664,N_12507);
nand U14968 (N_14968,N_13244,N_12541);
and U14969 (N_14969,N_13045,N_13591);
or U14970 (N_14970,N_12193,N_12794);
and U14971 (N_14971,N_13238,N_13519);
or U14972 (N_14972,N_12690,N_13505);
nand U14973 (N_14973,N_13138,N_12670);
and U14974 (N_14974,N_13894,N_13824);
nor U14975 (N_14975,N_13431,N_13642);
nor U14976 (N_14976,N_13445,N_13304);
or U14977 (N_14977,N_13867,N_12538);
and U14978 (N_14978,N_13265,N_13532);
and U14979 (N_14979,N_12840,N_13556);
nor U14980 (N_14980,N_13190,N_13300);
nand U14981 (N_14981,N_13496,N_12776);
nand U14982 (N_14982,N_12434,N_12971);
and U14983 (N_14983,N_13927,N_13883);
or U14984 (N_14984,N_13020,N_13394);
and U14985 (N_14985,N_12021,N_13079);
and U14986 (N_14986,N_13670,N_12371);
and U14987 (N_14987,N_13891,N_12099);
nor U14988 (N_14988,N_13749,N_13116);
nor U14989 (N_14989,N_12104,N_12283);
and U14990 (N_14990,N_13097,N_13740);
nand U14991 (N_14991,N_12637,N_12189);
nor U14992 (N_14992,N_12591,N_12998);
or U14993 (N_14993,N_12568,N_13550);
nor U14994 (N_14994,N_12174,N_12505);
or U14995 (N_14995,N_12372,N_13068);
nand U14996 (N_14996,N_13745,N_12233);
nand U14997 (N_14997,N_12429,N_13842);
nand U14998 (N_14998,N_12592,N_12348);
nand U14999 (N_14999,N_12414,N_13659);
and U15000 (N_15000,N_13344,N_12642);
nor U15001 (N_15001,N_13172,N_13098);
xnor U15002 (N_15002,N_13507,N_13002);
nand U15003 (N_15003,N_12558,N_12340);
nand U15004 (N_15004,N_13600,N_12845);
xnor U15005 (N_15005,N_13060,N_12204);
and U15006 (N_15006,N_13496,N_12033);
and U15007 (N_15007,N_13046,N_13227);
or U15008 (N_15008,N_12246,N_13136);
nor U15009 (N_15009,N_13145,N_13638);
or U15010 (N_15010,N_12752,N_12122);
nor U15011 (N_15011,N_12488,N_13647);
or U15012 (N_15012,N_12377,N_13218);
nor U15013 (N_15013,N_12490,N_13874);
nor U15014 (N_15014,N_12761,N_12668);
and U15015 (N_15015,N_12542,N_13713);
nand U15016 (N_15016,N_13297,N_12785);
or U15017 (N_15017,N_12727,N_13198);
or U15018 (N_15018,N_12452,N_12249);
and U15019 (N_15019,N_13657,N_13490);
nor U15020 (N_15020,N_13932,N_13712);
nor U15021 (N_15021,N_12568,N_12062);
nor U15022 (N_15022,N_12969,N_13816);
and U15023 (N_15023,N_13958,N_13332);
and U15024 (N_15024,N_12030,N_12123);
nor U15025 (N_15025,N_12943,N_13778);
nor U15026 (N_15026,N_12693,N_12227);
nand U15027 (N_15027,N_13637,N_12535);
and U15028 (N_15028,N_13170,N_13611);
and U15029 (N_15029,N_12856,N_13298);
and U15030 (N_15030,N_13678,N_12874);
nand U15031 (N_15031,N_12916,N_12301);
xor U15032 (N_15032,N_13478,N_13769);
or U15033 (N_15033,N_12777,N_13434);
and U15034 (N_15034,N_12161,N_13288);
or U15035 (N_15035,N_12438,N_13374);
or U15036 (N_15036,N_13804,N_12216);
or U15037 (N_15037,N_13374,N_12397);
or U15038 (N_15038,N_12497,N_13873);
or U15039 (N_15039,N_12900,N_13043);
nor U15040 (N_15040,N_12364,N_12630);
and U15041 (N_15041,N_13689,N_12868);
nor U15042 (N_15042,N_13134,N_13103);
and U15043 (N_15043,N_13214,N_12857);
and U15044 (N_15044,N_13502,N_12065);
or U15045 (N_15045,N_13552,N_13694);
or U15046 (N_15046,N_12352,N_13843);
nand U15047 (N_15047,N_12880,N_13064);
nor U15048 (N_15048,N_13883,N_13447);
or U15049 (N_15049,N_13226,N_13802);
nand U15050 (N_15050,N_13074,N_13186);
or U15051 (N_15051,N_13721,N_13750);
or U15052 (N_15052,N_12507,N_13541);
nand U15053 (N_15053,N_13766,N_12602);
nand U15054 (N_15054,N_12126,N_13834);
nand U15055 (N_15055,N_13514,N_13746);
nor U15056 (N_15056,N_12788,N_13729);
and U15057 (N_15057,N_12233,N_12258);
and U15058 (N_15058,N_13091,N_12524);
xor U15059 (N_15059,N_12114,N_12843);
or U15060 (N_15060,N_13866,N_12918);
and U15061 (N_15061,N_12646,N_13017);
nor U15062 (N_15062,N_12488,N_13255);
nor U15063 (N_15063,N_12812,N_12604);
nor U15064 (N_15064,N_13556,N_13756);
and U15065 (N_15065,N_13341,N_13380);
or U15066 (N_15066,N_13913,N_13849);
nor U15067 (N_15067,N_12423,N_13006);
and U15068 (N_15068,N_12530,N_12896);
nor U15069 (N_15069,N_13369,N_13496);
nand U15070 (N_15070,N_12939,N_12314);
or U15071 (N_15071,N_13589,N_13709);
or U15072 (N_15072,N_13306,N_13690);
and U15073 (N_15073,N_13400,N_12624);
and U15074 (N_15074,N_13411,N_13006);
and U15075 (N_15075,N_12264,N_13022);
nand U15076 (N_15076,N_12874,N_13700);
or U15077 (N_15077,N_12404,N_12993);
and U15078 (N_15078,N_13239,N_13215);
and U15079 (N_15079,N_12220,N_12369);
and U15080 (N_15080,N_12817,N_13730);
nor U15081 (N_15081,N_12541,N_13135);
nor U15082 (N_15082,N_12573,N_12219);
nand U15083 (N_15083,N_13759,N_12230);
nor U15084 (N_15084,N_12105,N_12583);
nor U15085 (N_15085,N_13975,N_12120);
or U15086 (N_15086,N_13462,N_13749);
or U15087 (N_15087,N_12739,N_13872);
nand U15088 (N_15088,N_13343,N_12084);
or U15089 (N_15089,N_12915,N_12066);
or U15090 (N_15090,N_13209,N_13211);
xnor U15091 (N_15091,N_13174,N_13394);
nor U15092 (N_15092,N_12513,N_12400);
or U15093 (N_15093,N_12015,N_13840);
and U15094 (N_15094,N_13891,N_13594);
nor U15095 (N_15095,N_13419,N_12181);
and U15096 (N_15096,N_12590,N_12235);
xnor U15097 (N_15097,N_12411,N_12481);
and U15098 (N_15098,N_13608,N_13329);
and U15099 (N_15099,N_13356,N_13671);
or U15100 (N_15100,N_12591,N_13545);
and U15101 (N_15101,N_12609,N_12482);
nor U15102 (N_15102,N_12971,N_13887);
nor U15103 (N_15103,N_12287,N_13240);
nor U15104 (N_15104,N_12455,N_12803);
and U15105 (N_15105,N_12695,N_13455);
or U15106 (N_15106,N_12766,N_12717);
nor U15107 (N_15107,N_12576,N_12979);
or U15108 (N_15108,N_12938,N_12449);
nor U15109 (N_15109,N_13279,N_12600);
nor U15110 (N_15110,N_13757,N_12763);
or U15111 (N_15111,N_12599,N_12886);
and U15112 (N_15112,N_12064,N_12102);
or U15113 (N_15113,N_12922,N_13364);
nand U15114 (N_15114,N_13975,N_13701);
nand U15115 (N_15115,N_12577,N_13562);
and U15116 (N_15116,N_13433,N_13948);
nor U15117 (N_15117,N_13783,N_12997);
and U15118 (N_15118,N_12902,N_12784);
nor U15119 (N_15119,N_13803,N_13477);
or U15120 (N_15120,N_13333,N_12335);
and U15121 (N_15121,N_12550,N_12803);
nor U15122 (N_15122,N_13435,N_12924);
nand U15123 (N_15123,N_13452,N_12053);
nand U15124 (N_15124,N_12959,N_12812);
and U15125 (N_15125,N_12947,N_12428);
nand U15126 (N_15126,N_13520,N_13343);
or U15127 (N_15127,N_13864,N_13349);
or U15128 (N_15128,N_12287,N_13257);
and U15129 (N_15129,N_13865,N_13464);
nand U15130 (N_15130,N_12711,N_13485);
or U15131 (N_15131,N_12310,N_13672);
nand U15132 (N_15132,N_12942,N_13496);
nor U15133 (N_15133,N_12709,N_12554);
nor U15134 (N_15134,N_12416,N_13259);
or U15135 (N_15135,N_12088,N_12478);
nand U15136 (N_15136,N_13171,N_13479);
nor U15137 (N_15137,N_13153,N_12866);
and U15138 (N_15138,N_12581,N_13491);
or U15139 (N_15139,N_12177,N_12332);
and U15140 (N_15140,N_13744,N_12325);
or U15141 (N_15141,N_12918,N_13089);
or U15142 (N_15142,N_12515,N_12823);
and U15143 (N_15143,N_13667,N_13200);
and U15144 (N_15144,N_12506,N_13793);
and U15145 (N_15145,N_13276,N_12499);
nand U15146 (N_15146,N_12476,N_13767);
and U15147 (N_15147,N_12334,N_13886);
nand U15148 (N_15148,N_12105,N_12298);
and U15149 (N_15149,N_13529,N_13498);
nor U15150 (N_15150,N_13616,N_13743);
or U15151 (N_15151,N_13970,N_13611);
or U15152 (N_15152,N_13700,N_12198);
and U15153 (N_15153,N_13460,N_12056);
nand U15154 (N_15154,N_12923,N_12209);
nor U15155 (N_15155,N_13590,N_12561);
nor U15156 (N_15156,N_12941,N_13870);
nand U15157 (N_15157,N_12997,N_13836);
nand U15158 (N_15158,N_12959,N_12183);
nor U15159 (N_15159,N_13902,N_13038);
nor U15160 (N_15160,N_13334,N_12543);
and U15161 (N_15161,N_12331,N_13947);
xor U15162 (N_15162,N_12354,N_13016);
and U15163 (N_15163,N_13123,N_13524);
xor U15164 (N_15164,N_13837,N_13005);
and U15165 (N_15165,N_13404,N_13904);
nand U15166 (N_15166,N_13634,N_12170);
nor U15167 (N_15167,N_13775,N_12573);
nor U15168 (N_15168,N_13100,N_13991);
nand U15169 (N_15169,N_13957,N_12699);
nand U15170 (N_15170,N_13043,N_13774);
nor U15171 (N_15171,N_12407,N_13723);
nor U15172 (N_15172,N_12256,N_13136);
and U15173 (N_15173,N_13688,N_12541);
nor U15174 (N_15174,N_12613,N_13380);
nand U15175 (N_15175,N_13162,N_12096);
or U15176 (N_15176,N_12014,N_12821);
or U15177 (N_15177,N_12667,N_13888);
and U15178 (N_15178,N_13672,N_12351);
nor U15179 (N_15179,N_12767,N_12421);
and U15180 (N_15180,N_13899,N_12640);
and U15181 (N_15181,N_13431,N_12129);
and U15182 (N_15182,N_12833,N_12628);
and U15183 (N_15183,N_12344,N_12479);
or U15184 (N_15184,N_12076,N_12807);
or U15185 (N_15185,N_12464,N_12274);
nor U15186 (N_15186,N_13055,N_13301);
nand U15187 (N_15187,N_13795,N_12917);
or U15188 (N_15188,N_12129,N_12307);
and U15189 (N_15189,N_12608,N_12581);
nand U15190 (N_15190,N_13197,N_12856);
nor U15191 (N_15191,N_12106,N_13542);
nor U15192 (N_15192,N_13858,N_13930);
nor U15193 (N_15193,N_13703,N_13662);
xnor U15194 (N_15194,N_12630,N_13742);
nand U15195 (N_15195,N_12283,N_13219);
or U15196 (N_15196,N_12620,N_13478);
nand U15197 (N_15197,N_13332,N_12601);
and U15198 (N_15198,N_12398,N_13868);
nand U15199 (N_15199,N_12131,N_13415);
and U15200 (N_15200,N_12690,N_12397);
or U15201 (N_15201,N_12836,N_13683);
or U15202 (N_15202,N_13000,N_13390);
and U15203 (N_15203,N_13639,N_12944);
or U15204 (N_15204,N_12756,N_12288);
or U15205 (N_15205,N_12236,N_13092);
nand U15206 (N_15206,N_13550,N_12530);
nor U15207 (N_15207,N_12687,N_12728);
and U15208 (N_15208,N_12231,N_13212);
nor U15209 (N_15209,N_13632,N_13126);
or U15210 (N_15210,N_13525,N_12599);
or U15211 (N_15211,N_13628,N_13942);
nor U15212 (N_15212,N_13293,N_12896);
nor U15213 (N_15213,N_12163,N_13921);
nor U15214 (N_15214,N_12405,N_12097);
or U15215 (N_15215,N_13132,N_13812);
nor U15216 (N_15216,N_13231,N_13769);
xnor U15217 (N_15217,N_13037,N_12012);
or U15218 (N_15218,N_13385,N_13608);
and U15219 (N_15219,N_12190,N_12095);
or U15220 (N_15220,N_13726,N_13348);
nor U15221 (N_15221,N_13969,N_13196);
or U15222 (N_15222,N_12211,N_12188);
and U15223 (N_15223,N_12135,N_13437);
nor U15224 (N_15224,N_13771,N_12967);
and U15225 (N_15225,N_12862,N_12027);
nand U15226 (N_15226,N_12240,N_13049);
nand U15227 (N_15227,N_13762,N_13179);
or U15228 (N_15228,N_12047,N_12260);
or U15229 (N_15229,N_13498,N_12824);
or U15230 (N_15230,N_13039,N_13308);
nor U15231 (N_15231,N_12463,N_13888);
nor U15232 (N_15232,N_13978,N_13510);
or U15233 (N_15233,N_12942,N_13688);
or U15234 (N_15234,N_12323,N_12356);
nor U15235 (N_15235,N_12638,N_13964);
or U15236 (N_15236,N_13384,N_13804);
or U15237 (N_15237,N_13156,N_12718);
and U15238 (N_15238,N_13808,N_13352);
and U15239 (N_15239,N_12467,N_12445);
and U15240 (N_15240,N_12288,N_13074);
nand U15241 (N_15241,N_12924,N_13966);
nand U15242 (N_15242,N_12132,N_13832);
and U15243 (N_15243,N_13059,N_12044);
nor U15244 (N_15244,N_13897,N_13920);
nand U15245 (N_15245,N_12474,N_12172);
or U15246 (N_15246,N_12618,N_12303);
or U15247 (N_15247,N_13523,N_13599);
or U15248 (N_15248,N_13522,N_12215);
or U15249 (N_15249,N_13015,N_12476);
or U15250 (N_15250,N_12916,N_13263);
nor U15251 (N_15251,N_13443,N_13996);
nand U15252 (N_15252,N_12376,N_13494);
xor U15253 (N_15253,N_12732,N_12171);
or U15254 (N_15254,N_13395,N_13022);
nor U15255 (N_15255,N_12176,N_13139);
nand U15256 (N_15256,N_13750,N_13259);
nor U15257 (N_15257,N_12589,N_12384);
and U15258 (N_15258,N_12440,N_13052);
nand U15259 (N_15259,N_12531,N_12703);
nor U15260 (N_15260,N_13579,N_13333);
xor U15261 (N_15261,N_13792,N_13346);
and U15262 (N_15262,N_12380,N_13477);
or U15263 (N_15263,N_13185,N_13037);
nor U15264 (N_15264,N_12488,N_13874);
nor U15265 (N_15265,N_12230,N_13189);
or U15266 (N_15266,N_13022,N_13873);
or U15267 (N_15267,N_13370,N_13990);
nor U15268 (N_15268,N_13203,N_13015);
nor U15269 (N_15269,N_13691,N_13276);
nor U15270 (N_15270,N_12296,N_12336);
or U15271 (N_15271,N_12699,N_13304);
nand U15272 (N_15272,N_13127,N_12545);
and U15273 (N_15273,N_12345,N_13717);
nor U15274 (N_15274,N_13295,N_13836);
nor U15275 (N_15275,N_13743,N_13440);
nor U15276 (N_15276,N_12898,N_12674);
nand U15277 (N_15277,N_12063,N_13733);
and U15278 (N_15278,N_13994,N_12304);
and U15279 (N_15279,N_12253,N_12878);
nor U15280 (N_15280,N_13183,N_13490);
xnor U15281 (N_15281,N_12814,N_13031);
nor U15282 (N_15282,N_13343,N_12584);
nand U15283 (N_15283,N_13392,N_12391);
and U15284 (N_15284,N_12094,N_13494);
and U15285 (N_15285,N_12292,N_12857);
and U15286 (N_15286,N_13331,N_13479);
nor U15287 (N_15287,N_13905,N_12067);
nor U15288 (N_15288,N_12324,N_13882);
nor U15289 (N_15289,N_12795,N_12858);
nor U15290 (N_15290,N_12476,N_13640);
or U15291 (N_15291,N_13340,N_13765);
nand U15292 (N_15292,N_12175,N_13703);
nor U15293 (N_15293,N_12213,N_13552);
and U15294 (N_15294,N_13431,N_13634);
nor U15295 (N_15295,N_13302,N_13058);
nand U15296 (N_15296,N_12580,N_12545);
nand U15297 (N_15297,N_13732,N_12066);
or U15298 (N_15298,N_13732,N_12309);
nand U15299 (N_15299,N_13213,N_13779);
nor U15300 (N_15300,N_13508,N_12940);
or U15301 (N_15301,N_12161,N_13840);
nand U15302 (N_15302,N_13720,N_13765);
and U15303 (N_15303,N_12759,N_13440);
nor U15304 (N_15304,N_13753,N_12401);
or U15305 (N_15305,N_12071,N_12199);
and U15306 (N_15306,N_13415,N_13741);
xnor U15307 (N_15307,N_13484,N_12926);
nand U15308 (N_15308,N_12807,N_12941);
nand U15309 (N_15309,N_13490,N_12056);
and U15310 (N_15310,N_13620,N_12618);
nand U15311 (N_15311,N_13881,N_13306);
nor U15312 (N_15312,N_12856,N_12656);
and U15313 (N_15313,N_13699,N_12216);
and U15314 (N_15314,N_13908,N_12052);
or U15315 (N_15315,N_13714,N_13257);
nand U15316 (N_15316,N_12564,N_12429);
and U15317 (N_15317,N_13576,N_13512);
nand U15318 (N_15318,N_12936,N_12501);
nand U15319 (N_15319,N_13934,N_13479);
and U15320 (N_15320,N_12021,N_12788);
nand U15321 (N_15321,N_13339,N_13318);
nand U15322 (N_15322,N_13336,N_12375);
or U15323 (N_15323,N_12387,N_13818);
and U15324 (N_15324,N_13686,N_13915);
or U15325 (N_15325,N_12814,N_13114);
nand U15326 (N_15326,N_13046,N_12709);
and U15327 (N_15327,N_12809,N_13024);
nand U15328 (N_15328,N_13332,N_12276);
or U15329 (N_15329,N_13453,N_12703);
nor U15330 (N_15330,N_12956,N_13452);
and U15331 (N_15331,N_12378,N_12981);
and U15332 (N_15332,N_13926,N_13772);
and U15333 (N_15333,N_13422,N_13989);
nor U15334 (N_15334,N_13436,N_13218);
nor U15335 (N_15335,N_12592,N_13600);
nand U15336 (N_15336,N_13811,N_12168);
or U15337 (N_15337,N_13025,N_12191);
nand U15338 (N_15338,N_12529,N_13029);
and U15339 (N_15339,N_12173,N_13654);
nand U15340 (N_15340,N_12925,N_12053);
nand U15341 (N_15341,N_13369,N_12697);
or U15342 (N_15342,N_13818,N_13967);
nand U15343 (N_15343,N_13830,N_12205);
and U15344 (N_15344,N_12862,N_13542);
nor U15345 (N_15345,N_12766,N_13556);
nand U15346 (N_15346,N_13612,N_12548);
nand U15347 (N_15347,N_12659,N_13144);
and U15348 (N_15348,N_12266,N_12619);
and U15349 (N_15349,N_13095,N_13398);
nor U15350 (N_15350,N_12729,N_13233);
or U15351 (N_15351,N_13307,N_13613);
nor U15352 (N_15352,N_12161,N_13308);
nand U15353 (N_15353,N_13190,N_12944);
and U15354 (N_15354,N_13584,N_13211);
or U15355 (N_15355,N_13797,N_13825);
nand U15356 (N_15356,N_13732,N_13881);
or U15357 (N_15357,N_13409,N_13688);
or U15358 (N_15358,N_13421,N_13271);
nor U15359 (N_15359,N_12981,N_12008);
or U15360 (N_15360,N_13941,N_12339);
or U15361 (N_15361,N_13756,N_12381);
nor U15362 (N_15362,N_12730,N_13000);
and U15363 (N_15363,N_12625,N_12146);
nor U15364 (N_15364,N_12281,N_12339);
nor U15365 (N_15365,N_13064,N_13504);
nand U15366 (N_15366,N_12501,N_12111);
and U15367 (N_15367,N_13951,N_13346);
or U15368 (N_15368,N_13790,N_12734);
nand U15369 (N_15369,N_12447,N_12913);
or U15370 (N_15370,N_13168,N_12256);
nand U15371 (N_15371,N_13158,N_13922);
and U15372 (N_15372,N_12213,N_13341);
and U15373 (N_15373,N_12648,N_13707);
and U15374 (N_15374,N_12880,N_13222);
nor U15375 (N_15375,N_13559,N_13940);
and U15376 (N_15376,N_12856,N_12610);
nor U15377 (N_15377,N_12782,N_13410);
nand U15378 (N_15378,N_13770,N_12025);
and U15379 (N_15379,N_12847,N_12002);
nor U15380 (N_15380,N_12574,N_12001);
or U15381 (N_15381,N_13202,N_13810);
and U15382 (N_15382,N_12395,N_12316);
or U15383 (N_15383,N_13412,N_12226);
or U15384 (N_15384,N_13622,N_12123);
nor U15385 (N_15385,N_13490,N_13168);
nand U15386 (N_15386,N_13978,N_13498);
nand U15387 (N_15387,N_12410,N_12626);
nor U15388 (N_15388,N_13450,N_12098);
nor U15389 (N_15389,N_13373,N_13340);
nand U15390 (N_15390,N_13344,N_12374);
nor U15391 (N_15391,N_12880,N_13156);
or U15392 (N_15392,N_13108,N_13422);
and U15393 (N_15393,N_12546,N_12148);
or U15394 (N_15394,N_12892,N_13621);
and U15395 (N_15395,N_12900,N_13683);
nand U15396 (N_15396,N_13058,N_12959);
nand U15397 (N_15397,N_13753,N_13712);
or U15398 (N_15398,N_12788,N_12388);
or U15399 (N_15399,N_12780,N_13968);
and U15400 (N_15400,N_12591,N_13441);
or U15401 (N_15401,N_13702,N_12045);
nor U15402 (N_15402,N_12726,N_13899);
nand U15403 (N_15403,N_13391,N_13365);
and U15404 (N_15404,N_13550,N_12489);
nand U15405 (N_15405,N_13884,N_13930);
xor U15406 (N_15406,N_13083,N_13769);
nand U15407 (N_15407,N_13163,N_13219);
or U15408 (N_15408,N_12005,N_13883);
or U15409 (N_15409,N_13337,N_13170);
or U15410 (N_15410,N_13957,N_12150);
nand U15411 (N_15411,N_12449,N_13742);
nand U15412 (N_15412,N_13084,N_13010);
xor U15413 (N_15413,N_12171,N_13601);
xor U15414 (N_15414,N_12253,N_13213);
or U15415 (N_15415,N_13942,N_12521);
and U15416 (N_15416,N_12510,N_12317);
and U15417 (N_15417,N_12162,N_13393);
or U15418 (N_15418,N_13640,N_12282);
or U15419 (N_15419,N_12827,N_13378);
nand U15420 (N_15420,N_13328,N_13284);
and U15421 (N_15421,N_12453,N_13128);
nor U15422 (N_15422,N_13624,N_13518);
or U15423 (N_15423,N_12733,N_13263);
nor U15424 (N_15424,N_13862,N_13513);
nor U15425 (N_15425,N_13207,N_12995);
or U15426 (N_15426,N_12585,N_13620);
nand U15427 (N_15427,N_12564,N_12723);
and U15428 (N_15428,N_12280,N_13719);
nor U15429 (N_15429,N_13420,N_13225);
nand U15430 (N_15430,N_13160,N_13137);
or U15431 (N_15431,N_12198,N_12102);
and U15432 (N_15432,N_12924,N_12266);
and U15433 (N_15433,N_13524,N_12659);
nor U15434 (N_15434,N_13946,N_12608);
and U15435 (N_15435,N_12577,N_13347);
and U15436 (N_15436,N_12405,N_12981);
nor U15437 (N_15437,N_12389,N_13224);
or U15438 (N_15438,N_13319,N_13840);
or U15439 (N_15439,N_13543,N_13716);
nor U15440 (N_15440,N_12482,N_13911);
and U15441 (N_15441,N_12462,N_13154);
nand U15442 (N_15442,N_13463,N_12605);
nand U15443 (N_15443,N_13044,N_12730);
or U15444 (N_15444,N_12797,N_12543);
nand U15445 (N_15445,N_13735,N_12900);
nand U15446 (N_15446,N_13125,N_12841);
nor U15447 (N_15447,N_13743,N_12055);
and U15448 (N_15448,N_13057,N_13977);
and U15449 (N_15449,N_13990,N_13010);
and U15450 (N_15450,N_12086,N_13978);
nor U15451 (N_15451,N_13242,N_13789);
or U15452 (N_15452,N_12896,N_13340);
nand U15453 (N_15453,N_12815,N_13311);
nor U15454 (N_15454,N_12353,N_12323);
nand U15455 (N_15455,N_13264,N_12894);
and U15456 (N_15456,N_12378,N_12197);
nor U15457 (N_15457,N_13179,N_13604);
nand U15458 (N_15458,N_13050,N_13829);
nand U15459 (N_15459,N_12294,N_13765);
nand U15460 (N_15460,N_13462,N_12216);
nor U15461 (N_15461,N_13699,N_12807);
nand U15462 (N_15462,N_12425,N_13320);
and U15463 (N_15463,N_12612,N_13695);
nor U15464 (N_15464,N_12203,N_13648);
and U15465 (N_15465,N_12492,N_12123);
nor U15466 (N_15466,N_13889,N_12061);
or U15467 (N_15467,N_12389,N_12804);
nor U15468 (N_15468,N_12547,N_13808);
nand U15469 (N_15469,N_13372,N_13434);
xor U15470 (N_15470,N_12441,N_12859);
nand U15471 (N_15471,N_13968,N_13111);
or U15472 (N_15472,N_12804,N_12486);
and U15473 (N_15473,N_12522,N_13585);
nor U15474 (N_15474,N_12489,N_12731);
and U15475 (N_15475,N_12078,N_12679);
nand U15476 (N_15476,N_13204,N_13358);
and U15477 (N_15477,N_13639,N_13683);
xnor U15478 (N_15478,N_13919,N_13429);
and U15479 (N_15479,N_13943,N_13099);
nor U15480 (N_15480,N_13714,N_12328);
and U15481 (N_15481,N_13031,N_12370);
and U15482 (N_15482,N_12257,N_12275);
and U15483 (N_15483,N_13819,N_12959);
or U15484 (N_15484,N_13387,N_13012);
nand U15485 (N_15485,N_13056,N_13357);
nand U15486 (N_15486,N_12794,N_12666);
nand U15487 (N_15487,N_13229,N_13696);
nor U15488 (N_15488,N_13161,N_13905);
or U15489 (N_15489,N_12011,N_12801);
or U15490 (N_15490,N_13997,N_12267);
nand U15491 (N_15491,N_12107,N_12743);
nor U15492 (N_15492,N_12915,N_13000);
xnor U15493 (N_15493,N_13084,N_12519);
nor U15494 (N_15494,N_13554,N_12662);
nand U15495 (N_15495,N_12776,N_12791);
and U15496 (N_15496,N_13865,N_13240);
or U15497 (N_15497,N_13045,N_12013);
nand U15498 (N_15498,N_12215,N_13861);
and U15499 (N_15499,N_12665,N_13196);
or U15500 (N_15500,N_13654,N_12791);
nand U15501 (N_15501,N_12037,N_13739);
or U15502 (N_15502,N_12479,N_13888);
xnor U15503 (N_15503,N_13396,N_12759);
nor U15504 (N_15504,N_13559,N_13700);
nand U15505 (N_15505,N_13094,N_13392);
nor U15506 (N_15506,N_13915,N_12515);
and U15507 (N_15507,N_13064,N_12734);
nand U15508 (N_15508,N_13815,N_12339);
xor U15509 (N_15509,N_12471,N_12840);
nor U15510 (N_15510,N_12008,N_12590);
xor U15511 (N_15511,N_12287,N_13284);
nor U15512 (N_15512,N_12270,N_12661);
nor U15513 (N_15513,N_13469,N_13878);
or U15514 (N_15514,N_13229,N_13634);
and U15515 (N_15515,N_12960,N_12307);
and U15516 (N_15516,N_13648,N_13206);
nand U15517 (N_15517,N_12719,N_13430);
xor U15518 (N_15518,N_12716,N_13817);
or U15519 (N_15519,N_13873,N_13563);
and U15520 (N_15520,N_13181,N_12120);
nor U15521 (N_15521,N_12293,N_12186);
and U15522 (N_15522,N_13594,N_12311);
and U15523 (N_15523,N_13717,N_13842);
and U15524 (N_15524,N_12614,N_12482);
nand U15525 (N_15525,N_12555,N_13496);
nand U15526 (N_15526,N_12027,N_13961);
and U15527 (N_15527,N_12567,N_13626);
and U15528 (N_15528,N_12434,N_12594);
nor U15529 (N_15529,N_12881,N_12662);
or U15530 (N_15530,N_12936,N_12737);
nand U15531 (N_15531,N_13977,N_13982);
or U15532 (N_15532,N_12135,N_13095);
nand U15533 (N_15533,N_13078,N_12609);
nor U15534 (N_15534,N_12851,N_13797);
and U15535 (N_15535,N_13466,N_12249);
and U15536 (N_15536,N_12276,N_12845);
nand U15537 (N_15537,N_13701,N_12941);
or U15538 (N_15538,N_12353,N_12343);
or U15539 (N_15539,N_12143,N_12090);
nor U15540 (N_15540,N_13994,N_12253);
xor U15541 (N_15541,N_13382,N_12850);
or U15542 (N_15542,N_12815,N_13701);
and U15543 (N_15543,N_12200,N_13813);
nand U15544 (N_15544,N_12613,N_13426);
and U15545 (N_15545,N_12021,N_13284);
xnor U15546 (N_15546,N_13432,N_12404);
or U15547 (N_15547,N_13292,N_13375);
and U15548 (N_15548,N_12148,N_13936);
or U15549 (N_15549,N_13379,N_12764);
and U15550 (N_15550,N_12395,N_12562);
nor U15551 (N_15551,N_12756,N_13634);
nand U15552 (N_15552,N_12012,N_13668);
or U15553 (N_15553,N_12820,N_12823);
xnor U15554 (N_15554,N_13856,N_12608);
nand U15555 (N_15555,N_13751,N_13276);
nand U15556 (N_15556,N_12932,N_13528);
or U15557 (N_15557,N_12369,N_13408);
nor U15558 (N_15558,N_12844,N_12178);
nor U15559 (N_15559,N_12011,N_13965);
or U15560 (N_15560,N_13463,N_13296);
nor U15561 (N_15561,N_12490,N_12654);
or U15562 (N_15562,N_12038,N_12283);
and U15563 (N_15563,N_13525,N_13611);
nor U15564 (N_15564,N_12094,N_13294);
and U15565 (N_15565,N_13524,N_12021);
nand U15566 (N_15566,N_13448,N_12487);
and U15567 (N_15567,N_13262,N_13477);
nand U15568 (N_15568,N_13749,N_12406);
xor U15569 (N_15569,N_13256,N_12632);
and U15570 (N_15570,N_13955,N_12596);
nand U15571 (N_15571,N_13574,N_12903);
and U15572 (N_15572,N_13955,N_12845);
nor U15573 (N_15573,N_13604,N_13210);
and U15574 (N_15574,N_12306,N_13358);
nor U15575 (N_15575,N_12719,N_13192);
nand U15576 (N_15576,N_13597,N_13981);
or U15577 (N_15577,N_13828,N_13522);
and U15578 (N_15578,N_13549,N_13181);
nor U15579 (N_15579,N_12140,N_13003);
and U15580 (N_15580,N_12708,N_13356);
nand U15581 (N_15581,N_12389,N_12229);
nand U15582 (N_15582,N_12104,N_12444);
nand U15583 (N_15583,N_12553,N_13422);
nor U15584 (N_15584,N_12210,N_13008);
xnor U15585 (N_15585,N_12614,N_13611);
and U15586 (N_15586,N_13424,N_13190);
nor U15587 (N_15587,N_13311,N_13620);
nor U15588 (N_15588,N_12336,N_13137);
nand U15589 (N_15589,N_12972,N_13159);
nor U15590 (N_15590,N_13995,N_12507);
xor U15591 (N_15591,N_13875,N_13805);
and U15592 (N_15592,N_12049,N_13933);
nor U15593 (N_15593,N_12182,N_12312);
nor U15594 (N_15594,N_13853,N_13791);
nand U15595 (N_15595,N_12441,N_12408);
and U15596 (N_15596,N_12833,N_12112);
or U15597 (N_15597,N_12013,N_13908);
or U15598 (N_15598,N_13281,N_13969);
or U15599 (N_15599,N_13229,N_12547);
nor U15600 (N_15600,N_12793,N_12714);
nor U15601 (N_15601,N_13342,N_13669);
or U15602 (N_15602,N_12015,N_12813);
and U15603 (N_15603,N_12925,N_12649);
or U15604 (N_15604,N_12359,N_12805);
or U15605 (N_15605,N_13842,N_12682);
and U15606 (N_15606,N_13623,N_12787);
or U15607 (N_15607,N_13433,N_13618);
nand U15608 (N_15608,N_13581,N_13569);
or U15609 (N_15609,N_13821,N_13897);
nor U15610 (N_15610,N_12353,N_13976);
xor U15611 (N_15611,N_12656,N_13703);
or U15612 (N_15612,N_12911,N_13873);
nor U15613 (N_15613,N_13244,N_13368);
nor U15614 (N_15614,N_13937,N_12492);
and U15615 (N_15615,N_12013,N_12089);
nor U15616 (N_15616,N_12750,N_13985);
or U15617 (N_15617,N_12990,N_13711);
or U15618 (N_15618,N_13836,N_13578);
nand U15619 (N_15619,N_13756,N_12356);
nand U15620 (N_15620,N_12900,N_13581);
nand U15621 (N_15621,N_13349,N_12123);
nand U15622 (N_15622,N_12635,N_12402);
and U15623 (N_15623,N_12979,N_12126);
and U15624 (N_15624,N_13279,N_13655);
and U15625 (N_15625,N_13992,N_12396);
and U15626 (N_15626,N_13706,N_13036);
and U15627 (N_15627,N_13012,N_13013);
and U15628 (N_15628,N_12213,N_12592);
or U15629 (N_15629,N_12101,N_13521);
nor U15630 (N_15630,N_13664,N_13599);
nor U15631 (N_15631,N_13063,N_13303);
nor U15632 (N_15632,N_12654,N_12333);
nand U15633 (N_15633,N_12494,N_12730);
and U15634 (N_15634,N_13088,N_12452);
nand U15635 (N_15635,N_12727,N_13674);
or U15636 (N_15636,N_13404,N_12501);
nor U15637 (N_15637,N_12873,N_13320);
nand U15638 (N_15638,N_13382,N_13499);
or U15639 (N_15639,N_13110,N_13741);
or U15640 (N_15640,N_12505,N_12150);
nand U15641 (N_15641,N_12175,N_13405);
and U15642 (N_15642,N_13642,N_13719);
and U15643 (N_15643,N_13801,N_12695);
nor U15644 (N_15644,N_13911,N_13101);
nand U15645 (N_15645,N_12614,N_12775);
nor U15646 (N_15646,N_12472,N_12431);
nor U15647 (N_15647,N_12706,N_13529);
nor U15648 (N_15648,N_12463,N_13250);
or U15649 (N_15649,N_13785,N_13486);
nor U15650 (N_15650,N_13710,N_13031);
and U15651 (N_15651,N_12102,N_12250);
and U15652 (N_15652,N_12997,N_13953);
or U15653 (N_15653,N_12060,N_12685);
and U15654 (N_15654,N_13094,N_12039);
or U15655 (N_15655,N_13747,N_12500);
nor U15656 (N_15656,N_12955,N_13786);
nor U15657 (N_15657,N_13670,N_12254);
nand U15658 (N_15658,N_12131,N_13255);
nor U15659 (N_15659,N_12736,N_12268);
nor U15660 (N_15660,N_13401,N_12572);
and U15661 (N_15661,N_12009,N_12951);
nor U15662 (N_15662,N_12425,N_12903);
nor U15663 (N_15663,N_13878,N_12616);
nand U15664 (N_15664,N_12434,N_12683);
and U15665 (N_15665,N_13320,N_12102);
or U15666 (N_15666,N_13952,N_12153);
and U15667 (N_15667,N_13429,N_12352);
and U15668 (N_15668,N_12332,N_13554);
nand U15669 (N_15669,N_12524,N_13566);
nor U15670 (N_15670,N_13382,N_13904);
nor U15671 (N_15671,N_12038,N_13184);
and U15672 (N_15672,N_12828,N_13803);
and U15673 (N_15673,N_12630,N_13761);
and U15674 (N_15674,N_13804,N_13182);
nor U15675 (N_15675,N_12771,N_13376);
or U15676 (N_15676,N_13322,N_13213);
nor U15677 (N_15677,N_13357,N_13758);
nor U15678 (N_15678,N_12246,N_13847);
or U15679 (N_15679,N_12172,N_12840);
xor U15680 (N_15680,N_12873,N_12781);
nor U15681 (N_15681,N_12072,N_13819);
or U15682 (N_15682,N_12149,N_12326);
nand U15683 (N_15683,N_12064,N_12852);
and U15684 (N_15684,N_13222,N_12453);
and U15685 (N_15685,N_12928,N_12319);
or U15686 (N_15686,N_12020,N_12730);
nor U15687 (N_15687,N_13196,N_13677);
and U15688 (N_15688,N_13499,N_13916);
or U15689 (N_15689,N_12707,N_13081);
and U15690 (N_15690,N_13135,N_13547);
nand U15691 (N_15691,N_13981,N_12422);
or U15692 (N_15692,N_13462,N_13521);
nor U15693 (N_15693,N_12839,N_13010);
nor U15694 (N_15694,N_13499,N_13142);
or U15695 (N_15695,N_12709,N_12914);
and U15696 (N_15696,N_12877,N_13044);
nand U15697 (N_15697,N_12964,N_12352);
and U15698 (N_15698,N_13898,N_13093);
or U15699 (N_15699,N_12465,N_13883);
nor U15700 (N_15700,N_13442,N_12410);
and U15701 (N_15701,N_12349,N_12546);
nand U15702 (N_15702,N_12354,N_13750);
nor U15703 (N_15703,N_12972,N_13908);
and U15704 (N_15704,N_12410,N_13658);
nand U15705 (N_15705,N_12502,N_13589);
or U15706 (N_15706,N_12015,N_13173);
nand U15707 (N_15707,N_12851,N_12631);
xor U15708 (N_15708,N_13959,N_13917);
nor U15709 (N_15709,N_13479,N_13279);
and U15710 (N_15710,N_12593,N_12355);
or U15711 (N_15711,N_13554,N_12476);
nor U15712 (N_15712,N_12994,N_13043);
or U15713 (N_15713,N_13749,N_13133);
or U15714 (N_15714,N_12473,N_12451);
or U15715 (N_15715,N_13524,N_13052);
nor U15716 (N_15716,N_13657,N_13293);
and U15717 (N_15717,N_13026,N_13202);
or U15718 (N_15718,N_13768,N_13243);
or U15719 (N_15719,N_13536,N_12730);
nand U15720 (N_15720,N_12302,N_13846);
and U15721 (N_15721,N_12310,N_13611);
nand U15722 (N_15722,N_13192,N_13148);
and U15723 (N_15723,N_13922,N_13476);
or U15724 (N_15724,N_13363,N_13199);
nor U15725 (N_15725,N_12840,N_13931);
and U15726 (N_15726,N_13323,N_12945);
nor U15727 (N_15727,N_13954,N_12549);
nor U15728 (N_15728,N_12860,N_12336);
nand U15729 (N_15729,N_13518,N_12970);
nand U15730 (N_15730,N_13239,N_13388);
nor U15731 (N_15731,N_12406,N_13411);
or U15732 (N_15732,N_13931,N_13228);
nor U15733 (N_15733,N_13609,N_13638);
and U15734 (N_15734,N_13662,N_12031);
nor U15735 (N_15735,N_13762,N_12057);
nand U15736 (N_15736,N_13760,N_12975);
or U15737 (N_15737,N_13480,N_13242);
or U15738 (N_15738,N_12418,N_12871);
and U15739 (N_15739,N_13824,N_13725);
nand U15740 (N_15740,N_12980,N_13455);
nand U15741 (N_15741,N_13513,N_13011);
and U15742 (N_15742,N_12416,N_13545);
and U15743 (N_15743,N_13202,N_13920);
and U15744 (N_15744,N_12588,N_12203);
or U15745 (N_15745,N_12154,N_12460);
xnor U15746 (N_15746,N_12024,N_13594);
or U15747 (N_15747,N_13707,N_13612);
nand U15748 (N_15748,N_13472,N_13107);
nand U15749 (N_15749,N_12792,N_12228);
nor U15750 (N_15750,N_13828,N_12940);
xor U15751 (N_15751,N_13617,N_13078);
and U15752 (N_15752,N_12475,N_13171);
or U15753 (N_15753,N_13713,N_13421);
nand U15754 (N_15754,N_13974,N_12050);
and U15755 (N_15755,N_12078,N_12911);
or U15756 (N_15756,N_13196,N_13977);
nand U15757 (N_15757,N_12746,N_13024);
nand U15758 (N_15758,N_13737,N_12109);
and U15759 (N_15759,N_12452,N_13335);
xnor U15760 (N_15760,N_13001,N_13656);
nor U15761 (N_15761,N_13075,N_13660);
or U15762 (N_15762,N_12566,N_12201);
or U15763 (N_15763,N_12776,N_13698);
or U15764 (N_15764,N_13101,N_12666);
nand U15765 (N_15765,N_13224,N_13263);
and U15766 (N_15766,N_13206,N_12418);
and U15767 (N_15767,N_13778,N_13752);
and U15768 (N_15768,N_13648,N_13976);
xor U15769 (N_15769,N_13102,N_13030);
or U15770 (N_15770,N_12246,N_13604);
and U15771 (N_15771,N_13510,N_13579);
and U15772 (N_15772,N_12699,N_12541);
and U15773 (N_15773,N_12853,N_12091);
nor U15774 (N_15774,N_12723,N_12577);
nand U15775 (N_15775,N_12836,N_13062);
and U15776 (N_15776,N_12230,N_13932);
nor U15777 (N_15777,N_12016,N_12384);
or U15778 (N_15778,N_12794,N_13207);
and U15779 (N_15779,N_12507,N_13977);
and U15780 (N_15780,N_13484,N_12124);
nand U15781 (N_15781,N_13880,N_12040);
nand U15782 (N_15782,N_12931,N_12497);
nor U15783 (N_15783,N_12247,N_13206);
nor U15784 (N_15784,N_13034,N_13133);
nor U15785 (N_15785,N_12946,N_12909);
nor U15786 (N_15786,N_13692,N_13170);
nor U15787 (N_15787,N_12922,N_13903);
nor U15788 (N_15788,N_12485,N_13904);
or U15789 (N_15789,N_13530,N_13032);
or U15790 (N_15790,N_12131,N_12564);
nand U15791 (N_15791,N_12223,N_12449);
or U15792 (N_15792,N_13068,N_13613);
nand U15793 (N_15793,N_12438,N_12099);
or U15794 (N_15794,N_12276,N_12967);
nor U15795 (N_15795,N_12336,N_13798);
nor U15796 (N_15796,N_13234,N_13757);
nor U15797 (N_15797,N_12204,N_12991);
and U15798 (N_15798,N_13866,N_12614);
nor U15799 (N_15799,N_12188,N_12099);
or U15800 (N_15800,N_13935,N_13714);
and U15801 (N_15801,N_13733,N_12018);
and U15802 (N_15802,N_13839,N_13013);
nor U15803 (N_15803,N_12798,N_12868);
or U15804 (N_15804,N_13052,N_12146);
or U15805 (N_15805,N_12292,N_12255);
and U15806 (N_15806,N_13635,N_13481);
nor U15807 (N_15807,N_12531,N_12844);
nor U15808 (N_15808,N_12596,N_12654);
nor U15809 (N_15809,N_13039,N_13096);
nor U15810 (N_15810,N_13091,N_13437);
or U15811 (N_15811,N_12871,N_13278);
and U15812 (N_15812,N_12232,N_13985);
nand U15813 (N_15813,N_13191,N_13619);
nand U15814 (N_15814,N_12276,N_12185);
or U15815 (N_15815,N_12110,N_12372);
nor U15816 (N_15816,N_13178,N_13924);
and U15817 (N_15817,N_12949,N_12588);
or U15818 (N_15818,N_12374,N_12221);
nand U15819 (N_15819,N_12506,N_13255);
or U15820 (N_15820,N_13562,N_12058);
or U15821 (N_15821,N_13700,N_12891);
or U15822 (N_15822,N_12886,N_13939);
and U15823 (N_15823,N_12554,N_12490);
and U15824 (N_15824,N_13715,N_13845);
or U15825 (N_15825,N_12466,N_12958);
nand U15826 (N_15826,N_12261,N_12712);
nand U15827 (N_15827,N_13778,N_13641);
and U15828 (N_15828,N_12812,N_12569);
nand U15829 (N_15829,N_12416,N_12478);
nand U15830 (N_15830,N_12157,N_13945);
nor U15831 (N_15831,N_12817,N_13117);
and U15832 (N_15832,N_13709,N_13741);
nand U15833 (N_15833,N_13391,N_12052);
nor U15834 (N_15834,N_13898,N_13796);
or U15835 (N_15835,N_12378,N_13302);
xor U15836 (N_15836,N_12222,N_13964);
or U15837 (N_15837,N_13771,N_12274);
nand U15838 (N_15838,N_13428,N_13413);
and U15839 (N_15839,N_12713,N_13425);
nand U15840 (N_15840,N_12803,N_13086);
or U15841 (N_15841,N_12376,N_12449);
nand U15842 (N_15842,N_13368,N_12995);
nor U15843 (N_15843,N_13535,N_12245);
and U15844 (N_15844,N_13538,N_12006);
nand U15845 (N_15845,N_12277,N_12378);
and U15846 (N_15846,N_13275,N_12074);
and U15847 (N_15847,N_12577,N_12093);
and U15848 (N_15848,N_12190,N_12549);
and U15849 (N_15849,N_12439,N_12716);
and U15850 (N_15850,N_13811,N_13622);
nand U15851 (N_15851,N_13204,N_12973);
nor U15852 (N_15852,N_13760,N_13233);
and U15853 (N_15853,N_12434,N_13897);
xor U15854 (N_15854,N_13965,N_12617);
and U15855 (N_15855,N_13130,N_12098);
or U15856 (N_15856,N_12436,N_13968);
nor U15857 (N_15857,N_13651,N_13593);
and U15858 (N_15858,N_13288,N_12971);
nor U15859 (N_15859,N_13822,N_13055);
nor U15860 (N_15860,N_12744,N_12355);
and U15861 (N_15861,N_13717,N_13229);
nand U15862 (N_15862,N_12955,N_13682);
nor U15863 (N_15863,N_12744,N_13629);
nor U15864 (N_15864,N_13902,N_12993);
nand U15865 (N_15865,N_13046,N_12603);
or U15866 (N_15866,N_13810,N_12305);
nand U15867 (N_15867,N_13475,N_13566);
xnor U15868 (N_15868,N_12372,N_12289);
or U15869 (N_15869,N_13973,N_13579);
nand U15870 (N_15870,N_12310,N_12973);
and U15871 (N_15871,N_13836,N_13623);
nor U15872 (N_15872,N_12664,N_12931);
nor U15873 (N_15873,N_13232,N_12551);
nand U15874 (N_15874,N_12255,N_12725);
or U15875 (N_15875,N_13763,N_12622);
xnor U15876 (N_15876,N_12734,N_13949);
nand U15877 (N_15877,N_13073,N_12418);
or U15878 (N_15878,N_12607,N_12936);
nor U15879 (N_15879,N_12031,N_13943);
nand U15880 (N_15880,N_12036,N_12225);
nand U15881 (N_15881,N_12021,N_12723);
or U15882 (N_15882,N_12510,N_12926);
nor U15883 (N_15883,N_12425,N_12342);
and U15884 (N_15884,N_12180,N_13518);
nor U15885 (N_15885,N_13188,N_13990);
nand U15886 (N_15886,N_12358,N_13986);
nor U15887 (N_15887,N_13218,N_12922);
or U15888 (N_15888,N_12148,N_12092);
or U15889 (N_15889,N_13887,N_12590);
and U15890 (N_15890,N_12994,N_13660);
nor U15891 (N_15891,N_12294,N_13746);
nand U15892 (N_15892,N_12219,N_13841);
xnor U15893 (N_15893,N_12142,N_13326);
or U15894 (N_15894,N_13145,N_13560);
nor U15895 (N_15895,N_13630,N_13895);
or U15896 (N_15896,N_13628,N_13151);
and U15897 (N_15897,N_13819,N_13284);
and U15898 (N_15898,N_12359,N_13616);
or U15899 (N_15899,N_12722,N_12591);
and U15900 (N_15900,N_12185,N_13031);
nor U15901 (N_15901,N_13856,N_13774);
and U15902 (N_15902,N_12177,N_12024);
nand U15903 (N_15903,N_12053,N_13278);
or U15904 (N_15904,N_13401,N_13772);
nor U15905 (N_15905,N_12735,N_13264);
or U15906 (N_15906,N_13243,N_12243);
nand U15907 (N_15907,N_13145,N_12810);
nand U15908 (N_15908,N_12893,N_13668);
xnor U15909 (N_15909,N_13239,N_13976);
or U15910 (N_15910,N_13039,N_13393);
and U15911 (N_15911,N_12408,N_12222);
nor U15912 (N_15912,N_13104,N_13420);
or U15913 (N_15913,N_13044,N_12529);
or U15914 (N_15914,N_12069,N_13142);
and U15915 (N_15915,N_12124,N_12900);
nor U15916 (N_15916,N_12148,N_12387);
nand U15917 (N_15917,N_12511,N_12086);
nand U15918 (N_15918,N_13227,N_13267);
and U15919 (N_15919,N_13583,N_12202);
and U15920 (N_15920,N_12016,N_12497);
and U15921 (N_15921,N_13391,N_12413);
and U15922 (N_15922,N_12456,N_12613);
or U15923 (N_15923,N_13210,N_13023);
nor U15924 (N_15924,N_13583,N_12970);
nor U15925 (N_15925,N_13127,N_12552);
or U15926 (N_15926,N_13789,N_12995);
and U15927 (N_15927,N_12928,N_12110);
nor U15928 (N_15928,N_12012,N_12422);
nor U15929 (N_15929,N_12436,N_12390);
nor U15930 (N_15930,N_12329,N_13160);
nand U15931 (N_15931,N_13335,N_13420);
or U15932 (N_15932,N_12218,N_13963);
nor U15933 (N_15933,N_12214,N_12243);
nand U15934 (N_15934,N_13628,N_12864);
xnor U15935 (N_15935,N_12011,N_12126);
and U15936 (N_15936,N_12473,N_13984);
or U15937 (N_15937,N_13743,N_12385);
and U15938 (N_15938,N_13544,N_12296);
and U15939 (N_15939,N_12088,N_12425);
nand U15940 (N_15940,N_13234,N_12013);
and U15941 (N_15941,N_12037,N_12173);
or U15942 (N_15942,N_12222,N_12307);
nand U15943 (N_15943,N_12199,N_12495);
and U15944 (N_15944,N_13113,N_12300);
and U15945 (N_15945,N_13700,N_12292);
or U15946 (N_15946,N_13813,N_13496);
nor U15947 (N_15947,N_12349,N_12941);
and U15948 (N_15948,N_12823,N_12302);
or U15949 (N_15949,N_13821,N_12299);
and U15950 (N_15950,N_12798,N_13819);
nor U15951 (N_15951,N_13768,N_13760);
and U15952 (N_15952,N_13964,N_13676);
and U15953 (N_15953,N_13151,N_13216);
nand U15954 (N_15954,N_12706,N_13523);
nand U15955 (N_15955,N_13813,N_12001);
or U15956 (N_15956,N_12946,N_13695);
nand U15957 (N_15957,N_12307,N_13724);
and U15958 (N_15958,N_12652,N_12492);
and U15959 (N_15959,N_13520,N_13486);
xor U15960 (N_15960,N_12106,N_13810);
and U15961 (N_15961,N_12658,N_13453);
or U15962 (N_15962,N_13668,N_12726);
xor U15963 (N_15963,N_13404,N_13196);
and U15964 (N_15964,N_13576,N_13677);
nand U15965 (N_15965,N_12985,N_13624);
nand U15966 (N_15966,N_13363,N_12550);
nand U15967 (N_15967,N_13629,N_13818);
and U15968 (N_15968,N_12455,N_13862);
nor U15969 (N_15969,N_12926,N_13444);
or U15970 (N_15970,N_13742,N_13400);
nand U15971 (N_15971,N_13545,N_12939);
nor U15972 (N_15972,N_12877,N_12721);
or U15973 (N_15973,N_12825,N_12787);
or U15974 (N_15974,N_12167,N_12675);
and U15975 (N_15975,N_13346,N_13857);
xnor U15976 (N_15976,N_13052,N_12486);
or U15977 (N_15977,N_12508,N_12353);
or U15978 (N_15978,N_12737,N_13208);
nand U15979 (N_15979,N_13473,N_12158);
and U15980 (N_15980,N_12406,N_12917);
and U15981 (N_15981,N_12736,N_13809);
and U15982 (N_15982,N_13306,N_13966);
nor U15983 (N_15983,N_12527,N_13918);
and U15984 (N_15984,N_13296,N_12227);
nand U15985 (N_15985,N_12907,N_13049);
or U15986 (N_15986,N_12776,N_13069);
or U15987 (N_15987,N_13428,N_13635);
and U15988 (N_15988,N_13380,N_12020);
or U15989 (N_15989,N_12563,N_13991);
and U15990 (N_15990,N_13023,N_12464);
and U15991 (N_15991,N_12403,N_12888);
nand U15992 (N_15992,N_13393,N_13408);
nor U15993 (N_15993,N_13984,N_13672);
nand U15994 (N_15994,N_13755,N_12899);
and U15995 (N_15995,N_13245,N_12656);
nor U15996 (N_15996,N_13541,N_13212);
nand U15997 (N_15997,N_13438,N_12672);
or U15998 (N_15998,N_12114,N_13563);
nor U15999 (N_15999,N_12356,N_13441);
nand U16000 (N_16000,N_15211,N_15387);
or U16001 (N_16001,N_15988,N_15359);
nor U16002 (N_16002,N_15701,N_14819);
or U16003 (N_16003,N_14280,N_14856);
nand U16004 (N_16004,N_14468,N_15605);
nor U16005 (N_16005,N_14992,N_15782);
and U16006 (N_16006,N_15669,N_14885);
nand U16007 (N_16007,N_15149,N_15552);
and U16008 (N_16008,N_14096,N_14424);
nand U16009 (N_16009,N_15096,N_14516);
nand U16010 (N_16010,N_15586,N_14886);
nand U16011 (N_16011,N_15421,N_14167);
nand U16012 (N_16012,N_15826,N_15792);
and U16013 (N_16013,N_14095,N_14942);
nor U16014 (N_16014,N_14683,N_15884);
nand U16015 (N_16015,N_15021,N_14928);
or U16016 (N_16016,N_14050,N_14228);
and U16017 (N_16017,N_14475,N_14590);
nand U16018 (N_16018,N_14694,N_14234);
or U16019 (N_16019,N_15070,N_14481);
nand U16020 (N_16020,N_15194,N_14699);
nor U16021 (N_16021,N_14571,N_14966);
nor U16022 (N_16022,N_15079,N_15896);
nor U16023 (N_16023,N_15001,N_15136);
nor U16024 (N_16024,N_15921,N_15502);
nand U16025 (N_16025,N_14727,N_14472);
nand U16026 (N_16026,N_15542,N_15963);
nor U16027 (N_16027,N_14852,N_14408);
xor U16028 (N_16028,N_15187,N_14011);
or U16029 (N_16029,N_14193,N_14977);
and U16030 (N_16030,N_14687,N_15532);
nand U16031 (N_16031,N_14250,N_14213);
nor U16032 (N_16032,N_15870,N_14373);
nor U16033 (N_16033,N_14238,N_15695);
or U16034 (N_16034,N_14645,N_14256);
nand U16035 (N_16035,N_14696,N_15318);
and U16036 (N_16036,N_15959,N_15095);
nand U16037 (N_16037,N_14765,N_15843);
nand U16038 (N_16038,N_14367,N_15992);
and U16039 (N_16039,N_14340,N_14496);
or U16040 (N_16040,N_15683,N_14638);
or U16041 (N_16041,N_15232,N_14337);
and U16042 (N_16042,N_15508,N_15202);
and U16043 (N_16043,N_14537,N_15269);
nor U16044 (N_16044,N_14515,N_14031);
nand U16045 (N_16045,N_14394,N_15799);
and U16046 (N_16046,N_15590,N_14166);
and U16047 (N_16047,N_15611,N_15007);
nor U16048 (N_16048,N_15419,N_14872);
nand U16049 (N_16049,N_15214,N_15009);
nand U16050 (N_16050,N_14319,N_14118);
and U16051 (N_16051,N_15958,N_15395);
nand U16052 (N_16052,N_14538,N_15371);
or U16053 (N_16053,N_14438,N_14579);
or U16054 (N_16054,N_15282,N_15533);
and U16055 (N_16055,N_14415,N_14439);
and U16056 (N_16056,N_14907,N_14176);
nand U16057 (N_16057,N_14999,N_14321);
nand U16058 (N_16058,N_14491,N_14123);
nor U16059 (N_16059,N_15497,N_15706);
or U16060 (N_16060,N_14422,N_14851);
and U16061 (N_16061,N_14072,N_15505);
nand U16062 (N_16062,N_14704,N_15373);
nand U16063 (N_16063,N_14099,N_14655);
nand U16064 (N_16064,N_14542,N_15957);
nor U16065 (N_16065,N_15711,N_14157);
nor U16066 (N_16066,N_14062,N_14376);
nor U16067 (N_16067,N_14676,N_15939);
or U16068 (N_16068,N_14806,N_14890);
nor U16069 (N_16069,N_15818,N_14633);
nor U16070 (N_16070,N_15610,N_15769);
and U16071 (N_16071,N_15338,N_14086);
or U16072 (N_16072,N_15727,N_15721);
and U16073 (N_16073,N_14188,N_14114);
and U16074 (N_16074,N_15834,N_15735);
nand U16075 (N_16075,N_15372,N_15573);
and U16076 (N_16076,N_14345,N_14018);
and U16077 (N_16077,N_14764,N_15265);
or U16078 (N_16078,N_14378,N_15644);
nor U16079 (N_16079,N_15556,N_15544);
nor U16080 (N_16080,N_15844,N_15239);
or U16081 (N_16081,N_15408,N_14656);
or U16082 (N_16082,N_14414,N_14453);
or U16083 (N_16083,N_15821,N_15245);
and U16084 (N_16084,N_14117,N_15115);
nor U16085 (N_16085,N_15829,N_15615);
nor U16086 (N_16086,N_15926,N_14503);
or U16087 (N_16087,N_15109,N_14776);
nor U16088 (N_16088,N_14845,N_14254);
nor U16089 (N_16089,N_15734,N_14181);
xnor U16090 (N_16090,N_14901,N_14292);
or U16091 (N_16091,N_14494,N_14930);
or U16092 (N_16092,N_15308,N_15920);
or U16093 (N_16093,N_14330,N_14665);
and U16094 (N_16094,N_14941,N_15567);
nand U16095 (N_16095,N_14070,N_15437);
nor U16096 (N_16096,N_14785,N_15041);
nand U16097 (N_16097,N_14214,N_14544);
nor U16098 (N_16098,N_15512,N_14893);
nor U16099 (N_16099,N_14354,N_14342);
nor U16100 (N_16100,N_14952,N_14803);
and U16101 (N_16101,N_14305,N_15268);
and U16102 (N_16102,N_15349,N_15463);
nor U16103 (N_16103,N_14358,N_14150);
or U16104 (N_16104,N_15401,N_15306);
and U16105 (N_16105,N_15496,N_14641);
and U16106 (N_16106,N_15962,N_15072);
and U16107 (N_16107,N_14149,N_15598);
or U16108 (N_16108,N_15277,N_14388);
nand U16109 (N_16109,N_15775,N_14458);
or U16110 (N_16110,N_15777,N_15218);
nand U16111 (N_16111,N_14637,N_15723);
or U16112 (N_16112,N_14860,N_15872);
or U16113 (N_16113,N_14836,N_14314);
nand U16114 (N_16114,N_15370,N_14680);
and U16115 (N_16115,N_15725,N_15259);
nand U16116 (N_16116,N_15112,N_15916);
or U16117 (N_16117,N_14457,N_14362);
and U16118 (N_16118,N_14713,N_14377);
or U16119 (N_16119,N_14034,N_14584);
nor U16120 (N_16120,N_14627,N_15581);
nor U16121 (N_16121,N_14846,N_14546);
nand U16122 (N_16122,N_14366,N_14406);
or U16123 (N_16123,N_15594,N_15032);
or U16124 (N_16124,N_14834,N_14141);
and U16125 (N_16125,N_14582,N_15653);
nor U16126 (N_16126,N_15886,N_14842);
nand U16127 (N_16127,N_15716,N_14707);
nand U16128 (N_16128,N_15694,N_14751);
nand U16129 (N_16129,N_14081,N_14074);
or U16130 (N_16130,N_14547,N_14235);
and U16131 (N_16131,N_14772,N_15092);
or U16132 (N_16132,N_15182,N_14790);
nand U16133 (N_16133,N_15297,N_15976);
or U16134 (N_16134,N_14083,N_14614);
or U16135 (N_16135,N_14716,N_14116);
or U16136 (N_16136,N_15430,N_15828);
and U16137 (N_16137,N_14393,N_14989);
or U16138 (N_16138,N_14705,N_15473);
and U16139 (N_16139,N_15053,N_15179);
and U16140 (N_16140,N_14489,N_14626);
or U16141 (N_16141,N_14786,N_14636);
or U16142 (N_16142,N_14476,N_14525);
nand U16143 (N_16143,N_14741,N_15833);
nor U16144 (N_16144,N_14051,N_14658);
nand U16145 (N_16145,N_15944,N_15196);
nor U16146 (N_16146,N_15666,N_15368);
nor U16147 (N_16147,N_14243,N_14490);
xnor U16148 (N_16148,N_14389,N_15974);
nand U16149 (N_16149,N_15912,N_14024);
and U16150 (N_16150,N_15504,N_15804);
and U16151 (N_16151,N_14442,N_14121);
or U16152 (N_16152,N_15914,N_14770);
or U16153 (N_16153,N_14210,N_14561);
and U16154 (N_16154,N_14762,N_14313);
or U16155 (N_16155,N_14281,N_15099);
or U16156 (N_16156,N_15341,N_14302);
nor U16157 (N_16157,N_14621,N_15948);
nor U16158 (N_16158,N_14372,N_15907);
and U16159 (N_16159,N_15641,N_14355);
or U16160 (N_16160,N_14905,N_15241);
or U16161 (N_16161,N_15759,N_14267);
nor U16162 (N_16162,N_14653,N_14271);
nand U16163 (N_16163,N_15073,N_14833);
nor U16164 (N_16164,N_14146,N_15130);
and U16165 (N_16165,N_14369,N_14264);
nor U16166 (N_16166,N_14237,N_15464);
nor U16167 (N_16167,N_15671,N_15290);
nor U16168 (N_16168,N_14242,N_15493);
or U16169 (N_16169,N_14165,N_15819);
and U16170 (N_16170,N_14087,N_14784);
and U16171 (N_16171,N_15856,N_14756);
and U16172 (N_16172,N_14335,N_14016);
nand U16173 (N_16173,N_14822,N_15173);
or U16174 (N_16174,N_15044,N_15322);
nor U16175 (N_16175,N_15619,N_15517);
nor U16176 (N_16176,N_15082,N_15050);
nor U16177 (N_16177,N_15979,N_15090);
nand U16178 (N_16178,N_14192,N_14898);
or U16179 (N_16179,N_14502,N_14606);
or U16180 (N_16180,N_15681,N_15474);
or U16181 (N_16181,N_14059,N_15745);
or U16182 (N_16182,N_14216,N_14576);
nand U16183 (N_16183,N_14331,N_15452);
nand U16184 (N_16184,N_14743,N_14451);
or U16185 (N_16185,N_14965,N_14049);
nand U16186 (N_16186,N_15761,N_14748);
and U16187 (N_16187,N_15147,N_14398);
or U16188 (N_16188,N_14385,N_14041);
nor U16189 (N_16189,N_14077,N_15283);
or U16190 (N_16190,N_14275,N_15319);
or U16191 (N_16191,N_14100,N_14792);
nor U16192 (N_16192,N_14040,N_15812);
nand U16193 (N_16193,N_15097,N_15927);
nand U16194 (N_16194,N_15540,N_14509);
nor U16195 (N_16195,N_15750,N_14679);
nor U16196 (N_16196,N_14558,N_15783);
nand U16197 (N_16197,N_15732,N_15191);
nor U16198 (N_16198,N_15647,N_14556);
nand U16199 (N_16199,N_15295,N_15918);
and U16200 (N_16200,N_15840,N_15230);
nand U16201 (N_16201,N_15402,N_15913);
or U16202 (N_16202,N_14329,N_14974);
nor U16203 (N_16203,N_15140,N_14831);
and U16204 (N_16204,N_15728,N_14519);
xor U16205 (N_16205,N_14171,N_14353);
or U16206 (N_16206,N_15827,N_14071);
or U16207 (N_16207,N_15094,N_15879);
xor U16208 (N_16208,N_14858,N_14828);
nand U16209 (N_16209,N_15609,N_14501);
and U16210 (N_16210,N_15863,N_14948);
or U16211 (N_16211,N_14168,N_15171);
nand U16212 (N_16212,N_15026,N_14971);
nor U16213 (N_16213,N_14585,N_15847);
or U16214 (N_16214,N_14409,N_15674);
or U16215 (N_16215,N_15722,N_15465);
nand U16216 (N_16216,N_15961,N_14722);
or U16217 (N_16217,N_15867,N_14597);
nor U16218 (N_16218,N_14418,N_15085);
nand U16219 (N_16219,N_15760,N_15928);
or U16220 (N_16220,N_15225,N_15541);
or U16221 (N_16221,N_15579,N_14425);
nor U16222 (N_16222,N_15547,N_14957);
nor U16223 (N_16223,N_14443,N_15880);
nor U16224 (N_16224,N_14032,N_15312);
nand U16225 (N_16225,N_15990,N_15687);
nor U16226 (N_16226,N_15289,N_14937);
nor U16227 (N_16227,N_15231,N_15328);
nor U16228 (N_16228,N_15688,N_15816);
nor U16229 (N_16229,N_14747,N_14742);
nor U16230 (N_16230,N_15849,N_15400);
nand U16231 (N_16231,N_15931,N_14437);
nor U16232 (N_16232,N_15601,N_14460);
and U16233 (N_16233,N_15864,N_14285);
xor U16234 (N_16234,N_14586,N_14924);
or U16235 (N_16235,N_15158,N_15443);
or U16236 (N_16236,N_15924,N_15790);
nor U16237 (N_16237,N_14844,N_14545);
or U16238 (N_16238,N_15055,N_15820);
nor U16239 (N_16239,N_15845,N_15117);
nor U16240 (N_16240,N_14944,N_15146);
or U16241 (N_16241,N_15654,N_15565);
nor U16242 (N_16242,N_14308,N_15578);
or U16243 (N_16243,N_14820,N_15235);
and U16244 (N_16244,N_14970,N_15684);
nor U16245 (N_16245,N_15530,N_14867);
nor U16246 (N_16246,N_14950,N_14604);
nand U16247 (N_16247,N_14246,N_14144);
nor U16248 (N_16248,N_15252,N_14396);
or U16249 (N_16249,N_15257,N_14904);
nand U16250 (N_16250,N_15686,N_14498);
and U16251 (N_16251,N_14122,N_15281);
or U16252 (N_16252,N_14675,N_14916);
nand U16253 (N_16253,N_14093,N_15878);
or U16254 (N_16254,N_14701,N_15755);
and U16255 (N_16255,N_15071,N_15538);
and U16256 (N_16256,N_14972,N_15923);
and U16257 (N_16257,N_15985,N_15134);
nor U16258 (N_16258,N_15469,N_14463);
nor U16259 (N_16259,N_15301,N_15510);
and U16260 (N_16260,N_14286,N_14789);
or U16261 (N_16261,N_15160,N_14883);
and U16262 (N_16262,N_15919,N_14471);
nor U16263 (N_16263,N_15893,N_14288);
nand U16264 (N_16264,N_15868,N_14467);
nand U16265 (N_16265,N_15577,N_15608);
and U16266 (N_16266,N_14344,N_15993);
nand U16267 (N_16267,N_15574,N_15904);
and U16268 (N_16268,N_15410,N_15851);
nand U16269 (N_16269,N_15059,N_15120);
nor U16270 (N_16270,N_14779,N_14877);
nor U16271 (N_16271,N_15270,N_15910);
nand U16272 (N_16272,N_15456,N_15320);
nand U16273 (N_16273,N_14283,N_15063);
or U16274 (N_16274,N_15661,N_14732);
or U16275 (N_16275,N_14771,N_15651);
nand U16276 (N_16276,N_15899,N_15405);
nor U16277 (N_16277,N_14129,N_14124);
nand U16278 (N_16278,N_14925,N_14349);
or U16279 (N_16279,N_14777,N_14401);
nor U16280 (N_16280,N_15162,N_15936);
nand U16281 (N_16281,N_15221,N_15718);
or U16282 (N_16282,N_14397,N_14220);
nor U16283 (N_16283,N_15704,N_15881);
or U16284 (N_16284,N_14013,N_14829);
and U16285 (N_16285,N_15922,N_14801);
nor U16286 (N_16286,N_15639,N_15814);
and U16287 (N_16287,N_15104,N_15213);
and U16288 (N_16288,N_14706,N_14015);
nand U16289 (N_16289,N_15066,N_15087);
or U16290 (N_16290,N_14486,N_14350);
nand U16291 (N_16291,N_14588,N_14363);
nand U16292 (N_16292,N_15485,N_14560);
nand U16293 (N_16293,N_15444,N_15431);
or U16294 (N_16294,N_14681,N_15305);
nor U16295 (N_16295,N_14581,N_14686);
nor U16296 (N_16296,N_14474,N_14399);
xor U16297 (N_16297,N_14044,N_14339);
and U16298 (N_16298,N_14336,N_14382);
nor U16299 (N_16299,N_14642,N_14236);
or U16300 (N_16300,N_14324,N_14441);
nor U16301 (N_16301,N_15930,N_14026);
or U16302 (N_16302,N_15111,N_15825);
and U16303 (N_16303,N_14333,N_14697);
and U16304 (N_16304,N_15757,N_14030);
nor U16305 (N_16305,N_15702,N_14624);
or U16306 (N_16306,N_15786,N_15911);
and U16307 (N_16307,N_15207,N_14110);
nand U16308 (N_16308,N_15486,N_14673);
nor U16309 (N_16309,N_15388,N_14360);
and U16310 (N_16310,N_14229,N_15472);
and U16311 (N_16311,N_15815,N_15057);
or U16312 (N_16312,N_15744,N_15709);
and U16313 (N_16313,N_14029,N_15568);
nor U16314 (N_16314,N_14282,N_15185);
and U16315 (N_16315,N_14569,N_14461);
nand U16316 (N_16316,N_14370,N_14631);
or U16317 (N_16317,N_15503,N_14555);
or U16318 (N_16318,N_14787,N_15470);
nand U16319 (N_16319,N_15429,N_14714);
nand U16320 (N_16320,N_15204,N_14793);
nor U16321 (N_16321,N_14809,N_15972);
or U16322 (N_16322,N_15475,N_14808);
and U16323 (N_16323,N_15733,N_15700);
and U16324 (N_16324,N_14311,N_14493);
or U16325 (N_16325,N_15135,N_14734);
nor U16326 (N_16326,N_14570,N_14497);
nor U16327 (N_16327,N_14152,N_14611);
or U16328 (N_16328,N_14618,N_15352);
or U16329 (N_16329,N_15738,N_14287);
nor U16330 (N_16330,N_15038,N_15521);
nor U16331 (N_16331,N_14534,N_15527);
nand U16332 (N_16332,N_14866,N_14137);
nand U16333 (N_16333,N_15593,N_14207);
or U16334 (N_16334,N_14812,N_15752);
nand U16335 (N_16335,N_15435,N_14274);
or U16336 (N_16336,N_15383,N_14774);
nor U16337 (N_16337,N_14954,N_14573);
nand U16338 (N_16338,N_15676,N_15137);
nor U16339 (N_16339,N_14303,N_15652);
or U16340 (N_16340,N_15366,N_15874);
and U16341 (N_16341,N_14723,N_15340);
nand U16342 (N_16342,N_14036,N_15679);
and U16343 (N_16343,N_14884,N_14514);
nand U16344 (N_16344,N_14297,N_14536);
and U16345 (N_16345,N_15536,N_14580);
nand U16346 (N_16346,N_14693,N_14064);
or U16347 (N_16347,N_14427,N_15380);
nand U16348 (N_16348,N_15758,N_15584);
nor U16349 (N_16349,N_14109,N_14383);
or U16350 (N_16350,N_15524,N_14089);
xor U16351 (N_16351,N_15048,N_15570);
and U16352 (N_16352,N_15580,N_15168);
nand U16353 (N_16353,N_15222,N_15363);
nor U16354 (N_16354,N_15005,N_14245);
or U16355 (N_16355,N_14426,N_14719);
and U16356 (N_16356,N_15302,N_14200);
nand U16357 (N_16357,N_15069,N_15300);
nor U16358 (N_16358,N_15596,N_15663);
xnor U16359 (N_16359,N_14518,N_15587);
or U16360 (N_16360,N_14753,N_14273);
or U16361 (N_16361,N_15217,N_14252);
nor U16362 (N_16362,N_14768,N_15244);
nor U16363 (N_16363,N_14865,N_14020);
nor U16364 (N_16364,N_14177,N_15309);
nor U16365 (N_16365,N_14932,N_15238);
nor U16366 (N_16366,N_15646,N_15223);
nand U16367 (N_16367,N_15736,N_14241);
nor U16368 (N_16368,N_14419,N_15551);
and U16369 (N_16369,N_15088,N_15811);
and U16370 (N_16370,N_14724,N_15209);
xor U16371 (N_16371,N_15386,N_15873);
nor U16372 (N_16372,N_14215,N_15550);
and U16373 (N_16373,N_14730,N_15049);
nand U16374 (N_16374,N_14539,N_15315);
and U16375 (N_16375,N_15479,N_14470);
nor U16376 (N_16376,N_15025,N_15501);
and U16377 (N_16377,N_14002,N_14182);
or U16378 (N_16378,N_15802,N_15737);
nor U16379 (N_16379,N_14959,N_14183);
nor U16380 (N_16380,N_14446,N_15106);
nor U16381 (N_16381,N_14454,N_15665);
nor U16382 (N_16382,N_14630,N_15176);
nor U16383 (N_16383,N_15977,N_15292);
nor U16384 (N_16384,N_14507,N_14379);
and U16385 (N_16385,N_15835,N_14140);
and U16386 (N_16386,N_15477,N_15638);
and U16387 (N_16387,N_14592,N_14386);
nand U16388 (N_16388,N_14943,N_14299);
or U16389 (N_16389,N_15822,N_14767);
or U16390 (N_16390,N_14484,N_15618);
and U16391 (N_16391,N_15433,N_14270);
or U16392 (N_16392,N_15076,N_15582);
and U16393 (N_16393,N_14535,N_14158);
and U16394 (N_16394,N_15678,N_15288);
and U16395 (N_16395,N_15384,N_15086);
nand U16396 (N_16396,N_14084,N_15746);
or U16397 (N_16397,N_14102,N_14700);
nand U16398 (N_16398,N_15743,N_15519);
and U16399 (N_16399,N_15170,N_15215);
nand U16400 (N_16400,N_15101,N_15513);
nor U16401 (N_16401,N_15999,N_14375);
and U16402 (N_16402,N_14849,N_14896);
or U16403 (N_16403,N_14847,N_14825);
or U16404 (N_16404,N_15626,N_15789);
nor U16405 (N_16405,N_15973,N_14961);
nor U16406 (N_16406,N_14411,N_14143);
and U16407 (N_16407,N_14310,N_14304);
xnor U16408 (N_16408,N_15773,N_14757);
nand U16409 (N_16409,N_15707,N_15107);
nor U16410 (N_16410,N_15397,N_14483);
nor U16411 (N_16411,N_15129,N_15377);
and U16412 (N_16412,N_14052,N_15330);
and U16413 (N_16413,N_14880,N_14987);
nand U16414 (N_16414,N_15051,N_15817);
or U16415 (N_16415,N_15188,N_14692);
nand U16416 (N_16416,N_15762,N_14445);
nor U16417 (N_16417,N_15422,N_15607);
or U16418 (N_16418,N_14039,N_15374);
and U16419 (N_16419,N_14563,N_14224);
nor U16420 (N_16420,N_14783,N_15986);
and U16421 (N_16421,N_15020,N_15237);
or U16422 (N_16422,N_14218,N_15122);
or U16423 (N_16423,N_15585,N_15242);
and U16424 (N_16424,N_14400,N_15848);
and U16425 (N_16425,N_14998,N_15576);
xor U16426 (N_16426,N_14205,N_15157);
nand U16427 (N_16427,N_15591,N_15764);
or U16428 (N_16428,N_15656,N_15836);
or U16429 (N_16429,N_15018,N_14802);
or U16430 (N_16430,N_15569,N_15857);
nor U16431 (N_16431,N_14583,N_14249);
nand U16432 (N_16432,N_15393,N_14529);
or U16433 (N_16433,N_15362,N_14047);
or U16434 (N_16434,N_14824,N_15226);
nor U16435 (N_16435,N_14392,N_15036);
and U16436 (N_16436,N_14332,N_14668);
nor U16437 (N_16437,N_15945,N_15901);
or U16438 (N_16438,N_14870,N_15997);
nand U16439 (N_16439,N_15633,N_14485);
or U16440 (N_16440,N_14019,N_14874);
and U16441 (N_16441,N_15796,N_15813);
or U16442 (N_16442,N_15390,N_14639);
nand U16443 (N_16443,N_15455,N_14664);
nand U16444 (N_16444,N_14796,N_15778);
nand U16445 (N_16445,N_14301,N_15592);
xnor U16446 (N_16446,N_14853,N_14195);
nor U16447 (N_16447,N_15518,N_14919);
and U16448 (N_16448,N_15407,N_15554);
nand U16449 (N_16449,N_14951,N_14007);
nor U16450 (N_16450,N_15186,N_14568);
nand U16451 (N_16451,N_15313,N_14455);
nand U16452 (N_16452,N_14773,N_15030);
nor U16453 (N_16453,N_14648,N_15299);
nand U16454 (N_16454,N_15680,N_15915);
or U16455 (N_16455,N_15011,N_14891);
or U16456 (N_16456,N_15730,N_14293);
nor U16457 (N_16457,N_14126,N_15648);
nand U16458 (N_16458,N_14995,N_15278);
nand U16459 (N_16459,N_14174,N_15181);
nand U16460 (N_16460,N_14107,N_14384);
nand U16461 (N_16461,N_15537,N_15102);
nand U16462 (N_16462,N_14922,N_15358);
nor U16463 (N_16463,N_14320,N_14488);
or U16464 (N_16464,N_14564,N_14230);
or U16465 (N_16465,N_15756,N_14403);
and U16466 (N_16466,N_15047,N_14108);
nand U16467 (N_16467,N_14088,N_15753);
nor U16468 (N_16468,N_14659,N_15285);
nand U16469 (N_16469,N_15449,N_15091);
nor U16470 (N_16470,N_14428,N_15877);
nand U16471 (N_16471,N_15143,N_15507);
nor U16472 (N_16472,N_14878,N_15529);
nand U16473 (N_16473,N_15258,N_14465);
and U16474 (N_16474,N_15776,N_14404);
xor U16475 (N_16475,N_15982,N_14436);
or U16476 (N_16476,N_14873,N_15515);
nor U16477 (N_16477,N_15394,N_15523);
or U16478 (N_16478,N_15621,N_15131);
or U16479 (N_16479,N_14986,N_14410);
nor U16480 (N_16480,N_14717,N_15858);
and U16481 (N_16481,N_14832,N_15327);
or U16482 (N_16482,N_15126,N_15832);
or U16483 (N_16483,N_15052,N_14910);
nor U16484 (N_16484,N_15412,N_15046);
nor U16485 (N_16485,N_14835,N_15511);
nand U16486 (N_16486,N_15314,N_14348);
nor U16487 (N_16487,N_14155,N_14855);
xor U16488 (N_16488,N_15634,N_15494);
nand U16489 (N_16489,N_14456,N_15480);
and U16490 (N_16490,N_14008,N_14841);
nor U16491 (N_16491,N_15121,N_14625);
nand U16492 (N_16492,N_15212,N_15650);
nand U16493 (N_16493,N_14938,N_14608);
nor U16494 (N_16494,N_15772,N_14993);
or U16495 (N_16495,N_14931,N_15291);
nand U16496 (N_16496,N_14253,N_15206);
or U16497 (N_16497,N_14949,N_14861);
or U16498 (N_16498,N_14232,N_14450);
nor U16499 (N_16499,N_15113,N_15024);
or U16500 (N_16500,N_14487,N_15148);
or U16501 (N_16501,N_15561,N_15434);
nor U16502 (N_16502,N_15342,N_15017);
nor U16503 (N_16503,N_14021,N_14712);
and U16504 (N_16504,N_15078,N_15749);
and U16505 (N_16505,N_14615,N_15898);
nor U16506 (N_16506,N_15253,N_14429);
or U16507 (N_16507,N_14978,N_15027);
or U16508 (N_16508,N_14685,N_14565);
nor U16509 (N_16509,N_15854,N_15951);
nand U16510 (N_16510,N_14374,N_14657);
nor U16511 (N_16511,N_15446,N_14698);
nand U16512 (N_16512,N_15953,N_15411);
nand U16513 (N_16513,N_14201,N_15768);
nand U16514 (N_16514,N_14524,N_15062);
nand U16515 (N_16515,N_14097,N_14887);
nand U16516 (N_16516,N_15203,N_15145);
or U16517 (N_16517,N_14927,N_15360);
and U16518 (N_16518,N_14721,N_15629);
nor U16519 (N_16519,N_15399,N_14127);
or U16520 (N_16520,N_14973,N_14120);
and U16521 (N_16521,N_14823,N_15975);
nand U16522 (N_16522,N_15487,N_14368);
nand U16523 (N_16523,N_14164,N_15458);
nor U16524 (N_16524,N_15454,N_15575);
nand U16525 (N_16525,N_15141,N_14520);
nor U16526 (N_16526,N_15229,N_15876);
nand U16527 (N_16527,N_14058,N_15809);
nor U16528 (N_16528,N_15166,N_14112);
and U16529 (N_16529,N_14710,N_14364);
or U16530 (N_16530,N_14602,N_14262);
or U16531 (N_16531,N_14170,N_14654);
nand U16532 (N_16532,N_14447,N_14900);
nand U16533 (N_16533,N_15682,N_15114);
nor U16534 (N_16534,N_14130,N_14616);
and U16535 (N_16535,N_15897,N_15555);
nand U16536 (N_16536,N_15672,N_15557);
and U16537 (N_16537,N_15946,N_15740);
nor U16538 (N_16538,N_14781,N_14325);
nand U16539 (N_16539,N_14480,N_14632);
and U16540 (N_16540,N_15488,N_14996);
nor U16541 (N_16541,N_15793,N_14327);
and U16542 (N_16542,N_15635,N_14562);
or U16543 (N_16543,N_14198,N_15869);
or U16544 (N_16544,N_15224,N_15438);
nor U16545 (N_16545,N_14433,N_15810);
or U16546 (N_16546,N_15178,N_15075);
nand U16547 (N_16547,N_14955,N_15273);
nor U16548 (N_16548,N_15664,N_15779);
nand U16549 (N_16549,N_15325,N_14227);
and U16550 (N_16550,N_14209,N_15348);
and U16551 (N_16551,N_14111,N_15506);
nor U16552 (N_16552,N_15420,N_15193);
or U16553 (N_16553,N_15139,N_15572);
xor U16554 (N_16554,N_15000,N_15673);
nor U16555 (N_16555,N_15056,N_14926);
nor U16556 (N_16556,N_15860,N_15697);
nand U16557 (N_16557,N_15124,N_14035);
nor U16558 (N_16558,N_15003,N_15566);
or U16559 (N_16559,N_14380,N_15406);
nor U16560 (N_16560,N_14259,N_14466);
or U16561 (N_16561,N_15531,N_14014);
nand U16562 (N_16562,N_15805,N_15043);
and U16563 (N_16563,N_14733,N_15184);
and U16564 (N_16564,N_15441,N_15606);
nand U16565 (N_16565,N_15205,N_15724);
nand U16566 (N_16566,N_14543,N_15905);
nand U16567 (N_16567,N_14541,N_15637);
nand U16568 (N_16568,N_14755,N_14033);
or U16569 (N_16569,N_14042,N_14260);
and U16570 (N_16570,N_14479,N_14752);
or U16571 (N_16571,N_14964,N_14997);
or U16572 (N_16572,N_15264,N_15228);
nor U16573 (N_16573,N_14945,N_15996);
and U16574 (N_16574,N_14431,N_15365);
nand U16575 (N_16575,N_15233,N_15970);
xor U16576 (N_16576,N_15144,N_15190);
nor U16577 (N_16577,N_14612,N_14899);
and U16578 (N_16578,N_14395,N_15770);
or U16579 (N_16579,N_14343,N_14391);
nor U16580 (N_16580,N_15266,N_14290);
nand U16581 (N_16581,N_14903,N_15478);
and U16582 (N_16582,N_15116,N_15560);
or U16583 (N_16583,N_14532,N_14605);
nand U16584 (N_16584,N_14045,N_14827);
nand U16585 (N_16585,N_15199,N_14889);
nor U16586 (N_16586,N_14263,N_15462);
or U16587 (N_16587,N_14156,N_14702);
and U16588 (N_16588,N_14745,N_14814);
and U16589 (N_16589,N_14859,N_15317);
xor U16590 (N_16590,N_15098,N_15016);
nand U16591 (N_16591,N_15333,N_14004);
nand U16592 (N_16592,N_15984,N_14635);
or U16593 (N_16593,N_15807,N_14718);
or U16594 (N_16594,N_14173,N_14038);
nor U16595 (N_16595,N_14760,N_14323);
nor U16596 (N_16596,N_14691,N_15516);
and U16597 (N_16597,N_14918,N_15528);
or U16598 (N_16598,N_14761,N_14749);
and U16599 (N_16599,N_14794,N_15364);
nand U16600 (N_16600,N_14620,N_15423);
xor U16601 (N_16601,N_15457,N_15917);
nor U16602 (N_16602,N_15622,N_14417);
or U16603 (N_16603,N_15938,N_15632);
nor U16604 (N_16604,N_14028,N_14651);
nand U16605 (N_16605,N_14548,N_15903);
and U16606 (N_16606,N_15599,N_15447);
nand U16607 (N_16607,N_15389,N_14206);
and U16608 (N_16608,N_15785,N_14085);
nand U16609 (N_16609,N_14566,N_15061);
and U16610 (N_16610,N_15471,N_14600);
or U16611 (N_16611,N_14800,N_14508);
and U16612 (N_16612,N_14115,N_14482);
nor U16613 (N_16613,N_14082,N_14758);
nand U16614 (N_16614,N_15483,N_15035);
and U16615 (N_16615,N_14985,N_14868);
nand U16616 (N_16616,N_14278,N_14261);
nand U16617 (N_16617,N_14079,N_14821);
nor U16618 (N_16618,N_15719,N_14247);
and U16619 (N_16619,N_15426,N_14356);
nor U16620 (N_16620,N_15495,N_15801);
and U16621 (N_16621,N_14607,N_14994);
nor U16622 (N_16622,N_14135,N_15624);
nor U16623 (N_16623,N_15304,N_14172);
or U16624 (N_16624,N_14405,N_14908);
nand U16625 (N_16625,N_14850,N_15693);
or U16626 (N_16626,N_14430,N_14272);
nand U16627 (N_16627,N_14005,N_15118);
nor U16628 (N_16628,N_15991,N_15128);
and U16629 (N_16629,N_14359,N_15439);
nand U16630 (N_16630,N_15885,N_15795);
xnor U16631 (N_16631,N_15164,N_15971);
nand U16632 (N_16632,N_14574,N_14906);
and U16633 (N_16633,N_15823,N_15889);
or U16634 (N_16634,N_15156,N_15655);
and U16635 (N_16635,N_14688,N_15602);
and U16636 (N_16636,N_15274,N_15453);
and U16637 (N_16637,N_15645,N_14969);
or U16638 (N_16638,N_15369,N_15033);
and U16639 (N_16639,N_15460,N_15381);
and U16640 (N_16640,N_15246,N_15074);
nor U16641 (N_16641,N_15806,N_15105);
and U16642 (N_16642,N_14980,N_14352);
nor U16643 (N_16643,N_14813,N_15932);
nand U16644 (N_16644,N_14775,N_15200);
nand U16645 (N_16645,N_14737,N_15824);
nand U16646 (N_16646,N_15326,N_15028);
and U16647 (N_16647,N_15323,N_14983);
xor U16648 (N_16648,N_15353,N_14025);
nand U16649 (N_16649,N_14240,N_14958);
nand U16650 (N_16650,N_14258,N_15416);
and U16651 (N_16651,N_15334,N_14805);
nand U16652 (N_16652,N_15631,N_15459);
or U16653 (N_16653,N_15771,N_14142);
nand U16654 (N_16654,N_14662,N_14098);
nand U16655 (N_16655,N_14953,N_14202);
nand U16656 (N_16656,N_15262,N_15690);
or U16657 (N_16657,N_14512,N_14478);
nor U16658 (N_16658,N_15925,N_15013);
and U16659 (N_16659,N_15023,N_15685);
and U16660 (N_16660,N_14554,N_15800);
nand U16661 (N_16661,N_15391,N_14416);
nor U16662 (N_16662,N_14709,N_15831);
and U16663 (N_16663,N_15691,N_14551);
and U16664 (N_16664,N_15689,N_14736);
or U16665 (N_16665,N_14371,N_14334);
nand U16666 (N_16666,N_14559,N_15859);
or U16667 (N_16667,N_14991,N_14268);
or U16668 (N_16668,N_15077,N_15748);
nor U16669 (N_16669,N_14046,N_14711);
or U16670 (N_16670,N_14092,N_14589);
or U16671 (N_16671,N_14361,N_15553);
and U16672 (N_16672,N_14567,N_14423);
nand U16673 (N_16673,N_14009,N_15174);
nand U16674 (N_16674,N_15279,N_15514);
or U16675 (N_16675,N_15436,N_14807);
and U16676 (N_16676,N_15249,N_14477);
nand U16677 (N_16677,N_14434,N_14432);
or U16678 (N_16678,N_15649,N_15165);
nand U16679 (N_16679,N_14090,N_15337);
nand U16680 (N_16680,N_15367,N_15361);
and U16681 (N_16681,N_15219,N_14136);
nor U16682 (N_16682,N_14552,N_14412);
or U16683 (N_16683,N_14864,N_15031);
and U16684 (N_16684,N_14613,N_14672);
nand U16685 (N_16685,N_14682,N_15583);
or U16686 (N_16686,N_14075,N_15351);
or U16687 (N_16687,N_15509,N_15084);
and U16688 (N_16688,N_15243,N_15883);
nor U16689 (N_16689,N_14990,N_15588);
nor U16690 (N_16690,N_15699,N_14186);
or U16691 (N_16691,N_14294,N_14289);
or U16692 (N_16692,N_15029,N_15335);
and U16693 (N_16693,N_14799,N_15929);
and U16694 (N_16694,N_14644,N_14162);
nor U16695 (N_16695,N_15154,N_14381);
nand U16696 (N_16696,N_14138,N_14725);
nand U16697 (N_16697,N_14739,N_15960);
xnor U16698 (N_16698,N_15255,N_14043);
and U16699 (N_16699,N_14068,N_15852);
or U16700 (N_16700,N_14413,N_15280);
and U16701 (N_16701,N_15415,N_14306);
and U16702 (N_16702,N_15628,N_15339);
and U16703 (N_16703,N_15103,N_15267);
xor U16704 (N_16704,N_14871,N_14816);
nor U16705 (N_16705,N_14940,N_14357);
and U16706 (N_16706,N_14277,N_14731);
nor U16707 (N_16707,N_15100,N_15355);
or U16708 (N_16708,N_14911,N_14139);
nand U16709 (N_16709,N_15172,N_15955);
nand U16710 (N_16710,N_15943,N_15981);
or U16711 (N_16711,N_15451,N_15571);
nand U16712 (N_16712,N_15808,N_14175);
or U16713 (N_16713,N_14572,N_15636);
nor U16714 (N_16714,N_15175,N_15022);
or U16715 (N_16715,N_14557,N_15167);
nor U16716 (N_16716,N_14609,N_14968);
nand U16717 (N_16717,N_14640,N_14128);
or U16718 (N_16718,N_14328,N_15006);
nor U16719 (N_16719,N_15747,N_15791);
nor U16720 (N_16720,N_14132,N_14528);
nor U16721 (N_16721,N_14595,N_15956);
and U16722 (N_16722,N_14628,N_14862);
xor U16723 (N_16723,N_14915,N_15888);
and U16724 (N_16724,N_15350,N_15549);
nand U16725 (N_16725,N_15132,N_14750);
or U16726 (N_16726,N_15316,N_15546);
or U16727 (N_16727,N_14677,N_14511);
nor U16728 (N_16728,N_14798,N_14650);
nor U16729 (N_16729,N_14326,N_15713);
or U16730 (N_16730,N_15272,N_14875);
and U16731 (N_16731,N_15763,N_14056);
nor U16732 (N_16732,N_14500,N_15534);
or U16733 (N_16733,N_15989,N_14876);
and U16734 (N_16734,N_15548,N_15484);
and U16735 (N_16735,N_15428,N_14226);
or U16736 (N_16736,N_15712,N_15965);
nor U16737 (N_16737,N_15662,N_15286);
and U16738 (N_16738,N_15346,N_14791);
and U16739 (N_16739,N_14929,N_15675);
nor U16740 (N_16740,N_14674,N_15490);
and U16741 (N_16741,N_14239,N_14178);
or U16742 (N_16742,N_14670,N_14449);
and U16743 (N_16743,N_15015,N_15742);
and U16744 (N_16744,N_14023,N_15396);
or U16745 (N_16745,N_14145,N_14053);
nand U16746 (N_16746,N_15949,N_15336);
and U16747 (N_16747,N_15163,N_14963);
nand U16748 (N_16748,N_14817,N_14473);
nand U16749 (N_16749,N_15293,N_14048);
nand U16750 (N_16750,N_15123,N_15002);
and U16751 (N_16751,N_14153,N_14222);
nor U16752 (N_16752,N_15138,N_14550);
nor U16753 (N_16753,N_14810,N_14204);
nor U16754 (N_16754,N_15612,N_15660);
nor U16755 (N_16755,N_14440,N_15425);
nor U16756 (N_16756,N_14840,N_15110);
nand U16757 (N_16757,N_14661,N_15220);
nand U16758 (N_16758,N_14495,N_14818);
nor U16759 (N_16759,N_14131,N_15717);
and U16760 (N_16760,N_14882,N_15210);
nand U16761 (N_16761,N_15375,N_14854);
nor U16762 (N_16762,N_14001,N_15589);
and U16763 (N_16763,N_15535,N_15766);
and U16764 (N_16764,N_15276,N_14312);
xnor U16765 (N_16765,N_15838,N_14257);
nand U16766 (N_16766,N_15875,N_14462);
and U16767 (N_16767,N_15489,N_14499);
or U16768 (N_16768,N_14151,N_14012);
and U16769 (N_16769,N_14055,N_15754);
nor U16770 (N_16770,N_15842,N_14284);
or U16771 (N_16771,N_14935,N_14577);
nor U16772 (N_16772,N_15227,N_14838);
or U16773 (N_16773,N_15376,N_15658);
or U16774 (N_16774,N_15448,N_15417);
and U16775 (N_16775,N_14251,N_14255);
and U16776 (N_16776,N_15714,N_15710);
and U16777 (N_16777,N_14895,N_15385);
or U16778 (N_16778,N_14623,N_15781);
nor U16779 (N_16779,N_15189,N_15354);
nand U16780 (N_16780,N_14469,N_15153);
and U16781 (N_16781,N_14351,N_15617);
nand U16782 (N_16782,N_14067,N_15564);
nand U16783 (N_16783,N_15155,N_15620);
nand U16784 (N_16784,N_15404,N_14671);
nor U16785 (N_16785,N_15392,N_14982);
or U16786 (N_16786,N_15964,N_15500);
and U16787 (N_16787,N_15287,N_15332);
or U16788 (N_16788,N_15846,N_15739);
and U16789 (N_16789,N_14599,N_14106);
nor U16790 (N_16790,N_15934,N_15837);
nor U16791 (N_16791,N_15698,N_15787);
and U16792 (N_16792,N_15201,N_14811);
or U16793 (N_16793,N_14506,N_14402);
nand U16794 (N_16794,N_14217,N_15980);
and U16795 (N_16795,N_15520,N_14160);
and U16796 (N_16796,N_14522,N_15558);
nand U16797 (N_16797,N_15169,N_15119);
nor U16798 (N_16798,N_15108,N_15696);
nor U16799 (N_16799,N_14603,N_14523);
and U16800 (N_16800,N_14103,N_14452);
or U16801 (N_16801,N_14596,N_15195);
and U16802 (N_16802,N_15933,N_14594);
or U16803 (N_16803,N_15794,N_14909);
nand U16804 (N_16804,N_15866,N_15461);
nand U16805 (N_16805,N_14746,N_14830);
nand U16806 (N_16806,N_14869,N_14265);
nand U16807 (N_16807,N_14988,N_15941);
nand U16808 (N_16808,N_14269,N_15068);
and U16809 (N_16809,N_15040,N_14649);
or U16810 (N_16810,N_15720,N_14060);
or U16811 (N_16811,N_15797,N_15378);
nand U16812 (N_16812,N_14912,N_15627);
xnor U16813 (N_16813,N_14769,N_15667);
nand U16814 (N_16814,N_15198,N_14184);
nand U16815 (N_16815,N_15468,N_15726);
nor U16816 (N_16816,N_14307,N_14956);
nand U16817 (N_16817,N_14587,N_14735);
and U16818 (N_16818,N_14540,N_14652);
nor U16819 (N_16819,N_14318,N_15356);
nor U16820 (N_16820,N_15331,N_15251);
nand U16821 (N_16821,N_15019,N_14598);
nand U16822 (N_16822,N_15967,N_15382);
nor U16823 (N_16823,N_14464,N_15784);
nor U16824 (N_16824,N_15256,N_15294);
nand U16825 (N_16825,N_14902,N_14967);
nand U16826 (N_16826,N_15543,N_15892);
and U16827 (N_16827,N_15424,N_14161);
nand U16828 (N_16828,N_14387,N_14421);
nand U16829 (N_16829,N_15481,N_14897);
and U16830 (N_16830,N_15642,N_14211);
nor U16831 (N_16831,N_14133,N_15234);
nor U16832 (N_16832,N_14815,N_14179);
or U16833 (N_16833,N_14892,N_14420);
nand U16834 (N_16834,N_15900,N_14322);
or U16835 (N_16835,N_15254,N_15871);
or U16836 (N_16836,N_14578,N_14521);
and U16837 (N_16837,N_15659,N_15780);
and U16838 (N_16838,N_15159,N_15054);
and U16839 (N_16839,N_14231,N_15064);
or U16840 (N_16840,N_14720,N_15216);
or U16841 (N_16841,N_15597,N_14169);
nand U16842 (N_16842,N_15357,N_14766);
nand U16843 (N_16843,N_15952,N_15142);
and U16844 (N_16844,N_14148,N_14754);
nor U16845 (N_16845,N_15995,N_15906);
and U16846 (N_16846,N_14505,N_14795);
and U16847 (N_16847,N_15409,N_14689);
and U16848 (N_16848,N_14197,N_14076);
or U16849 (N_16849,N_15894,N_15751);
or U16850 (N_16850,N_15539,N_15014);
or U16851 (N_16851,N_15125,N_14296);
or U16852 (N_16852,N_14448,N_15307);
nor U16853 (N_16853,N_14510,N_15640);
and U16854 (N_16854,N_15731,N_14894);
nor U16855 (N_16855,N_14300,N_14740);
nor U16856 (N_16856,N_14728,N_15670);
nand U16857 (N_16857,N_15298,N_15705);
nor U16858 (N_16858,N_14444,N_14667);
and U16859 (N_16859,N_14622,N_14459);
or U16860 (N_16860,N_15152,N_15321);
nand U16861 (N_16861,N_14888,N_15347);
and U16862 (N_16862,N_15060,N_14061);
and U16863 (N_16863,N_14843,N_14017);
or U16864 (N_16864,N_15008,N_14684);
nor U16865 (N_16865,N_14839,N_14591);
nand U16866 (N_16866,N_15850,N_15522);
nand U16867 (N_16867,N_14960,N_14962);
and U16868 (N_16868,N_14203,N_14782);
nand U16869 (N_16869,N_14189,N_14920);
or U16870 (N_16870,N_14703,N_14341);
nor U16871 (N_16871,N_14276,N_15127);
or U16872 (N_16872,N_14134,N_15998);
nand U16873 (N_16873,N_14212,N_14936);
xor U16874 (N_16874,N_15865,N_15545);
and U16875 (N_16875,N_14914,N_14780);
or U16876 (N_16876,N_14125,N_14695);
or U16877 (N_16877,N_15089,N_14837);
nand U16878 (N_16878,N_15183,N_15729);
nor U16879 (N_16879,N_14857,N_14526);
nor U16880 (N_16880,N_15311,N_14549);
and U16881 (N_16881,N_15613,N_15492);
nor U16882 (N_16882,N_15427,N_15668);
xnor U16883 (N_16883,N_15954,N_14933);
nand U16884 (N_16884,N_14517,N_14979);
and U16885 (N_16885,N_14163,N_14003);
nor U16886 (N_16886,N_14848,N_15440);
xor U16887 (N_16887,N_15765,N_14390);
or U16888 (N_16888,N_15630,N_14027);
and U16889 (N_16889,N_15862,N_15498);
nor U16890 (N_16890,N_14913,N_15432);
nand U16891 (N_16891,N_14073,N_14154);
nand U16892 (N_16892,N_14194,N_14726);
or U16893 (N_16893,N_15476,N_14984);
nor U16894 (N_16894,N_14317,N_15379);
nor U16895 (N_16895,N_15093,N_14863);
or U16896 (N_16896,N_15208,N_14663);
or U16897 (N_16897,N_14069,N_15616);
or U16898 (N_16898,N_14346,N_15841);
or U16899 (N_16899,N_15677,N_15788);
nand U16900 (N_16900,N_15467,N_15414);
nor U16901 (N_16901,N_14223,N_15065);
nor U16902 (N_16902,N_14006,N_14101);
and U16903 (N_16903,N_15345,N_14881);
and U16904 (N_16904,N_14678,N_15983);
or U16905 (N_16905,N_14921,N_14619);
and U16906 (N_16906,N_14492,N_15969);
or U16907 (N_16907,N_14666,N_14879);
or U16908 (N_16908,N_14646,N_15703);
nor U16909 (N_16909,N_15909,N_15908);
xor U16910 (N_16910,N_15887,N_14010);
nor U16911 (N_16911,N_15798,N_15855);
nand U16912 (N_16912,N_15271,N_15942);
and U16913 (N_16913,N_15526,N_14338);
or U16914 (N_16914,N_15987,N_14298);
xor U16915 (N_16915,N_14187,N_15275);
or U16916 (N_16916,N_14593,N_15150);
nor U16917 (N_16917,N_14199,N_14078);
nand U16918 (N_16918,N_14660,N_15491);
or U16919 (N_16919,N_14744,N_15767);
or U16920 (N_16920,N_14000,N_15261);
nor U16921 (N_16921,N_14669,N_15197);
nor U16922 (N_16922,N_15296,N_15010);
or U16923 (N_16923,N_14266,N_15853);
nor U16924 (N_16924,N_15418,N_14185);
and U16925 (N_16925,N_14946,N_14054);
or U16926 (N_16926,N_14037,N_15708);
nand U16927 (N_16927,N_14738,N_15248);
xnor U16928 (N_16928,N_15643,N_14647);
nand U16929 (N_16929,N_14113,N_15978);
or U16930 (N_16930,N_15250,N_15861);
nand U16931 (N_16931,N_15525,N_14105);
or U16932 (N_16932,N_14610,N_15466);
nor U16933 (N_16933,N_15882,N_15803);
nand U16934 (N_16934,N_15042,N_15966);
or U16935 (N_16935,N_15004,N_14066);
nor U16936 (N_16936,N_14309,N_15595);
or U16937 (N_16937,N_15559,N_14365);
or U16938 (N_16938,N_14248,N_14022);
or U16939 (N_16939,N_15413,N_14094);
nand U16940 (N_16940,N_14981,N_14407);
or U16941 (N_16941,N_14826,N_14601);
nor U16942 (N_16942,N_15830,N_15310);
or U16943 (N_16943,N_14190,N_15895);
or U16944 (N_16944,N_14196,N_14065);
and U16945 (N_16945,N_14091,N_14759);
and U16946 (N_16946,N_15600,N_15994);
or U16947 (N_16947,N_14527,N_14690);
nand U16948 (N_16948,N_15240,N_14221);
or U16949 (N_16949,N_15324,N_14708);
and U16950 (N_16950,N_15657,N_14923);
or U16951 (N_16951,N_15839,N_14788);
and U16952 (N_16952,N_14208,N_14233);
and U16953 (N_16953,N_14643,N_15450);
nor U16954 (N_16954,N_15482,N_15058);
or U16955 (N_16955,N_15034,N_15614);
nor U16956 (N_16956,N_14080,N_15177);
nand U16957 (N_16957,N_14147,N_14316);
nor U16958 (N_16958,N_14533,N_14513);
nand U16959 (N_16959,N_15192,N_15442);
or U16960 (N_16960,N_14315,N_15604);
nor U16961 (N_16961,N_15263,N_14975);
nor U16962 (N_16962,N_14763,N_14797);
nand U16963 (N_16963,N_15890,N_15083);
and U16964 (N_16964,N_15133,N_14939);
and U16965 (N_16965,N_15398,N_14976);
or U16966 (N_16966,N_14180,N_15303);
nor U16967 (N_16967,N_15940,N_14225);
nand U16968 (N_16968,N_15343,N_14104);
nand U16969 (N_16969,N_14531,N_14191);
nor U16970 (N_16970,N_15741,N_14634);
nand U16971 (N_16971,N_15247,N_14291);
or U16972 (N_16972,N_15161,N_14917);
and U16973 (N_16973,N_14804,N_15067);
nor U16974 (N_16974,N_14347,N_15603);
nor U16975 (N_16975,N_15692,N_15623);
nand U16976 (N_16976,N_14279,N_15445);
or U16977 (N_16977,N_15344,N_14617);
or U16978 (N_16978,N_14295,N_15715);
nand U16979 (N_16979,N_14119,N_15950);
nand U16980 (N_16980,N_14729,N_14934);
nand U16981 (N_16981,N_15891,N_15947);
xor U16982 (N_16982,N_14629,N_15625);
and U16983 (N_16983,N_15937,N_14715);
nand U16984 (N_16984,N_15081,N_15080);
nand U16985 (N_16985,N_15499,N_15037);
and U16986 (N_16986,N_15968,N_15045);
nand U16987 (N_16987,N_14778,N_14057);
nand U16988 (N_16988,N_14435,N_15562);
nor U16989 (N_16989,N_15902,N_14159);
and U16990 (N_16990,N_15403,N_15935);
or U16991 (N_16991,N_14244,N_15180);
nor U16992 (N_16992,N_14063,N_15329);
nor U16993 (N_16993,N_15012,N_15151);
or U16994 (N_16994,N_14530,N_15236);
xor U16995 (N_16995,N_14947,N_15260);
and U16996 (N_16996,N_14504,N_14575);
nor U16997 (N_16997,N_15039,N_15563);
and U16998 (N_16998,N_15774,N_14553);
and U16999 (N_16999,N_15284,N_14219);
or U17000 (N_17000,N_14787,N_14471);
nor U17001 (N_17001,N_15897,N_15006);
or U17002 (N_17002,N_15771,N_14138);
xnor U17003 (N_17003,N_15896,N_14998);
nand U17004 (N_17004,N_14212,N_15008);
and U17005 (N_17005,N_15719,N_14438);
and U17006 (N_17006,N_15998,N_15988);
and U17007 (N_17007,N_15154,N_15490);
nand U17008 (N_17008,N_14853,N_15761);
and U17009 (N_17009,N_14165,N_15225);
nand U17010 (N_17010,N_15618,N_14582);
nor U17011 (N_17011,N_15090,N_15195);
nand U17012 (N_17012,N_14301,N_15059);
xor U17013 (N_17013,N_15924,N_15706);
nand U17014 (N_17014,N_15348,N_15650);
and U17015 (N_17015,N_14475,N_14653);
nand U17016 (N_17016,N_14439,N_14108);
or U17017 (N_17017,N_15862,N_14123);
and U17018 (N_17018,N_14660,N_15364);
and U17019 (N_17019,N_14280,N_14428);
and U17020 (N_17020,N_15488,N_14748);
nand U17021 (N_17021,N_15271,N_15669);
nand U17022 (N_17022,N_14263,N_14080);
nor U17023 (N_17023,N_15344,N_15634);
and U17024 (N_17024,N_15953,N_14533);
and U17025 (N_17025,N_14881,N_14403);
or U17026 (N_17026,N_15531,N_14527);
or U17027 (N_17027,N_15881,N_15402);
or U17028 (N_17028,N_15859,N_15598);
and U17029 (N_17029,N_14827,N_15541);
nand U17030 (N_17030,N_15846,N_15007);
nand U17031 (N_17031,N_15160,N_15868);
nor U17032 (N_17032,N_15826,N_14720);
or U17033 (N_17033,N_14776,N_15789);
and U17034 (N_17034,N_15378,N_14235);
and U17035 (N_17035,N_15593,N_14681);
nor U17036 (N_17036,N_15493,N_14395);
or U17037 (N_17037,N_15334,N_15179);
and U17038 (N_17038,N_15389,N_15362);
nor U17039 (N_17039,N_15640,N_15727);
or U17040 (N_17040,N_15839,N_14751);
or U17041 (N_17041,N_15873,N_14936);
nor U17042 (N_17042,N_14554,N_15315);
nand U17043 (N_17043,N_14172,N_14200);
and U17044 (N_17044,N_15109,N_15296);
and U17045 (N_17045,N_15846,N_14146);
or U17046 (N_17046,N_15308,N_14343);
and U17047 (N_17047,N_14591,N_15416);
and U17048 (N_17048,N_14628,N_14510);
nor U17049 (N_17049,N_15771,N_14063);
and U17050 (N_17050,N_14753,N_15670);
nor U17051 (N_17051,N_14536,N_15111);
nor U17052 (N_17052,N_15069,N_15859);
and U17053 (N_17053,N_15758,N_14888);
or U17054 (N_17054,N_15947,N_14238);
or U17055 (N_17055,N_15469,N_15966);
nand U17056 (N_17056,N_14607,N_15812);
and U17057 (N_17057,N_14361,N_15616);
or U17058 (N_17058,N_14154,N_14397);
and U17059 (N_17059,N_15706,N_15328);
xnor U17060 (N_17060,N_15534,N_14326);
and U17061 (N_17061,N_15690,N_15881);
or U17062 (N_17062,N_15984,N_15779);
or U17063 (N_17063,N_15374,N_14061);
nand U17064 (N_17064,N_14435,N_15823);
or U17065 (N_17065,N_15352,N_15958);
nand U17066 (N_17066,N_14344,N_15809);
and U17067 (N_17067,N_14512,N_14661);
xnor U17068 (N_17068,N_15540,N_14448);
nand U17069 (N_17069,N_14627,N_14522);
and U17070 (N_17070,N_15723,N_14497);
and U17071 (N_17071,N_14018,N_15535);
nand U17072 (N_17072,N_15883,N_15230);
or U17073 (N_17073,N_15290,N_14480);
and U17074 (N_17074,N_14743,N_15900);
xnor U17075 (N_17075,N_14334,N_15910);
nor U17076 (N_17076,N_14112,N_15734);
nor U17077 (N_17077,N_14130,N_15507);
nand U17078 (N_17078,N_15618,N_14794);
or U17079 (N_17079,N_14389,N_15472);
and U17080 (N_17080,N_14502,N_15495);
nand U17081 (N_17081,N_14682,N_14573);
nand U17082 (N_17082,N_14820,N_14537);
and U17083 (N_17083,N_14802,N_15212);
nor U17084 (N_17084,N_14911,N_15633);
nor U17085 (N_17085,N_14832,N_15127);
or U17086 (N_17086,N_14983,N_14879);
nor U17087 (N_17087,N_15034,N_14164);
nand U17088 (N_17088,N_14089,N_15335);
nand U17089 (N_17089,N_15635,N_14361);
nand U17090 (N_17090,N_15495,N_14053);
nor U17091 (N_17091,N_15350,N_14947);
nor U17092 (N_17092,N_15318,N_14511);
and U17093 (N_17093,N_14245,N_15305);
nor U17094 (N_17094,N_15528,N_15297);
or U17095 (N_17095,N_14530,N_15945);
nand U17096 (N_17096,N_15817,N_14495);
nor U17097 (N_17097,N_14731,N_15320);
and U17098 (N_17098,N_15882,N_15306);
or U17099 (N_17099,N_15435,N_15328);
or U17100 (N_17100,N_15288,N_15836);
or U17101 (N_17101,N_15351,N_15673);
nor U17102 (N_17102,N_14300,N_14597);
or U17103 (N_17103,N_15018,N_14386);
nor U17104 (N_17104,N_15042,N_14405);
and U17105 (N_17105,N_14297,N_14454);
and U17106 (N_17106,N_15100,N_15837);
or U17107 (N_17107,N_14567,N_15305);
and U17108 (N_17108,N_15365,N_15967);
nand U17109 (N_17109,N_14005,N_15566);
nand U17110 (N_17110,N_15575,N_15466);
nand U17111 (N_17111,N_15892,N_14769);
nand U17112 (N_17112,N_14191,N_14646);
nor U17113 (N_17113,N_14661,N_15791);
or U17114 (N_17114,N_14733,N_14760);
nand U17115 (N_17115,N_15965,N_15806);
nand U17116 (N_17116,N_15079,N_15536);
and U17117 (N_17117,N_14872,N_15875);
nor U17118 (N_17118,N_14155,N_15507);
nand U17119 (N_17119,N_15687,N_14490);
and U17120 (N_17120,N_14573,N_14030);
nor U17121 (N_17121,N_14030,N_14918);
nand U17122 (N_17122,N_15210,N_15778);
nor U17123 (N_17123,N_15900,N_14514);
nand U17124 (N_17124,N_15104,N_15566);
and U17125 (N_17125,N_14930,N_14196);
nor U17126 (N_17126,N_14947,N_15077);
nor U17127 (N_17127,N_14943,N_14253);
nor U17128 (N_17128,N_14770,N_15067);
nand U17129 (N_17129,N_14281,N_15281);
nor U17130 (N_17130,N_15461,N_14475);
nand U17131 (N_17131,N_15839,N_14772);
nor U17132 (N_17132,N_15909,N_15709);
nor U17133 (N_17133,N_14206,N_15249);
nand U17134 (N_17134,N_15531,N_15558);
nand U17135 (N_17135,N_15040,N_15708);
nand U17136 (N_17136,N_14257,N_14576);
or U17137 (N_17137,N_14973,N_14415);
nand U17138 (N_17138,N_15102,N_14403);
nor U17139 (N_17139,N_14185,N_14511);
nor U17140 (N_17140,N_14052,N_14996);
nor U17141 (N_17141,N_14803,N_14598);
nor U17142 (N_17142,N_14746,N_15636);
and U17143 (N_17143,N_14024,N_14005);
or U17144 (N_17144,N_14081,N_15765);
nor U17145 (N_17145,N_15381,N_14502);
and U17146 (N_17146,N_15719,N_14610);
or U17147 (N_17147,N_14186,N_14402);
or U17148 (N_17148,N_14987,N_15505);
and U17149 (N_17149,N_14583,N_14150);
and U17150 (N_17150,N_15844,N_15101);
or U17151 (N_17151,N_14317,N_15732);
or U17152 (N_17152,N_15817,N_14858);
and U17153 (N_17153,N_14437,N_14868);
or U17154 (N_17154,N_15937,N_14740);
or U17155 (N_17155,N_15708,N_15241);
nand U17156 (N_17156,N_15803,N_15787);
nor U17157 (N_17157,N_14987,N_14587);
nand U17158 (N_17158,N_14040,N_14312);
nor U17159 (N_17159,N_15547,N_14989);
or U17160 (N_17160,N_15537,N_14859);
nor U17161 (N_17161,N_14239,N_14454);
nor U17162 (N_17162,N_15191,N_15206);
nand U17163 (N_17163,N_15906,N_14334);
nand U17164 (N_17164,N_15621,N_15833);
and U17165 (N_17165,N_14410,N_15642);
nor U17166 (N_17166,N_15547,N_14392);
and U17167 (N_17167,N_15501,N_15655);
and U17168 (N_17168,N_14338,N_14845);
nor U17169 (N_17169,N_15384,N_14088);
or U17170 (N_17170,N_14750,N_15399);
and U17171 (N_17171,N_14556,N_15697);
nor U17172 (N_17172,N_14376,N_15657);
and U17173 (N_17173,N_14824,N_14309);
or U17174 (N_17174,N_14144,N_15707);
or U17175 (N_17175,N_14908,N_15954);
nor U17176 (N_17176,N_15954,N_14046);
nor U17177 (N_17177,N_15186,N_15939);
nor U17178 (N_17178,N_14052,N_15899);
nor U17179 (N_17179,N_14528,N_15684);
nor U17180 (N_17180,N_15679,N_14717);
nor U17181 (N_17181,N_15267,N_15860);
nand U17182 (N_17182,N_14404,N_15054);
and U17183 (N_17183,N_14655,N_14478);
nand U17184 (N_17184,N_14790,N_14380);
or U17185 (N_17185,N_14581,N_15505);
or U17186 (N_17186,N_14231,N_14230);
xnor U17187 (N_17187,N_14721,N_15962);
nand U17188 (N_17188,N_14811,N_14566);
nand U17189 (N_17189,N_15623,N_15215);
nor U17190 (N_17190,N_14900,N_14054);
or U17191 (N_17191,N_14820,N_15371);
nor U17192 (N_17192,N_15767,N_14668);
xor U17193 (N_17193,N_15006,N_15694);
nor U17194 (N_17194,N_14290,N_14594);
nand U17195 (N_17195,N_14625,N_15660);
nor U17196 (N_17196,N_14681,N_15274);
nand U17197 (N_17197,N_14924,N_14369);
nor U17198 (N_17198,N_14491,N_15649);
nand U17199 (N_17199,N_14944,N_14148);
nand U17200 (N_17200,N_14454,N_14571);
nor U17201 (N_17201,N_14770,N_14662);
and U17202 (N_17202,N_15835,N_14492);
nand U17203 (N_17203,N_14478,N_14918);
or U17204 (N_17204,N_14301,N_15157);
nor U17205 (N_17205,N_14899,N_15274);
nor U17206 (N_17206,N_15851,N_15707);
nand U17207 (N_17207,N_14840,N_14468);
or U17208 (N_17208,N_15826,N_15595);
and U17209 (N_17209,N_14468,N_14922);
nand U17210 (N_17210,N_15046,N_14581);
nand U17211 (N_17211,N_15381,N_15571);
and U17212 (N_17212,N_15184,N_14820);
and U17213 (N_17213,N_15147,N_15141);
nor U17214 (N_17214,N_14549,N_15226);
and U17215 (N_17215,N_15324,N_14328);
xnor U17216 (N_17216,N_14408,N_15646);
and U17217 (N_17217,N_15729,N_14199);
nand U17218 (N_17218,N_14570,N_15044);
nor U17219 (N_17219,N_15189,N_15014);
or U17220 (N_17220,N_14127,N_15080);
or U17221 (N_17221,N_15827,N_15584);
nand U17222 (N_17222,N_15642,N_15630);
nand U17223 (N_17223,N_14558,N_15525);
or U17224 (N_17224,N_15796,N_15237);
nor U17225 (N_17225,N_15785,N_14672);
nand U17226 (N_17226,N_15212,N_14837);
nor U17227 (N_17227,N_15466,N_14788);
and U17228 (N_17228,N_14749,N_15034);
nand U17229 (N_17229,N_14748,N_14287);
nor U17230 (N_17230,N_14958,N_14843);
nand U17231 (N_17231,N_15669,N_14075);
and U17232 (N_17232,N_14356,N_15508);
nor U17233 (N_17233,N_15099,N_15130);
and U17234 (N_17234,N_15285,N_14693);
xnor U17235 (N_17235,N_15015,N_15487);
nand U17236 (N_17236,N_15481,N_15697);
nor U17237 (N_17237,N_15547,N_14795);
or U17238 (N_17238,N_15372,N_14738);
nor U17239 (N_17239,N_14155,N_14438);
and U17240 (N_17240,N_15824,N_14641);
nor U17241 (N_17241,N_14052,N_15935);
nand U17242 (N_17242,N_14371,N_14606);
or U17243 (N_17243,N_14426,N_14507);
and U17244 (N_17244,N_15009,N_14297);
or U17245 (N_17245,N_14785,N_15613);
and U17246 (N_17246,N_14312,N_15839);
nor U17247 (N_17247,N_15169,N_15595);
or U17248 (N_17248,N_14064,N_15694);
and U17249 (N_17249,N_14255,N_14054);
nor U17250 (N_17250,N_15868,N_14646);
nand U17251 (N_17251,N_14349,N_14599);
or U17252 (N_17252,N_14025,N_14194);
nor U17253 (N_17253,N_15052,N_14189);
xor U17254 (N_17254,N_15597,N_14353);
nand U17255 (N_17255,N_15872,N_14213);
and U17256 (N_17256,N_15467,N_15152);
nand U17257 (N_17257,N_15142,N_14574);
nand U17258 (N_17258,N_15167,N_14464);
nor U17259 (N_17259,N_15299,N_15011);
nor U17260 (N_17260,N_15447,N_14691);
or U17261 (N_17261,N_15098,N_14379);
and U17262 (N_17262,N_14703,N_15692);
nand U17263 (N_17263,N_15846,N_15729);
nor U17264 (N_17264,N_14059,N_14153);
or U17265 (N_17265,N_15595,N_14005);
nor U17266 (N_17266,N_14032,N_15572);
or U17267 (N_17267,N_14819,N_14196);
nand U17268 (N_17268,N_15822,N_14707);
or U17269 (N_17269,N_15998,N_15873);
or U17270 (N_17270,N_15843,N_15056);
or U17271 (N_17271,N_14734,N_15557);
or U17272 (N_17272,N_15493,N_15282);
and U17273 (N_17273,N_14125,N_14005);
or U17274 (N_17274,N_14855,N_15632);
and U17275 (N_17275,N_15529,N_15905);
xor U17276 (N_17276,N_15127,N_15721);
or U17277 (N_17277,N_14747,N_15512);
nand U17278 (N_17278,N_15983,N_14506);
nand U17279 (N_17279,N_15279,N_15915);
or U17280 (N_17280,N_14372,N_14773);
or U17281 (N_17281,N_15746,N_14860);
nor U17282 (N_17282,N_14919,N_14527);
nor U17283 (N_17283,N_14319,N_15656);
and U17284 (N_17284,N_15300,N_14647);
or U17285 (N_17285,N_14802,N_14160);
or U17286 (N_17286,N_14472,N_14941);
or U17287 (N_17287,N_14423,N_14228);
and U17288 (N_17288,N_14379,N_15084);
or U17289 (N_17289,N_15965,N_14390);
nand U17290 (N_17290,N_14321,N_15641);
and U17291 (N_17291,N_15450,N_14026);
xnor U17292 (N_17292,N_14308,N_15278);
nand U17293 (N_17293,N_14437,N_15867);
or U17294 (N_17294,N_14141,N_14369);
nand U17295 (N_17295,N_15900,N_15090);
or U17296 (N_17296,N_14361,N_14855);
or U17297 (N_17297,N_14911,N_14816);
nand U17298 (N_17298,N_14582,N_15525);
and U17299 (N_17299,N_14089,N_14760);
nor U17300 (N_17300,N_14681,N_14116);
and U17301 (N_17301,N_14320,N_15316);
nand U17302 (N_17302,N_15968,N_15515);
and U17303 (N_17303,N_15035,N_15410);
nor U17304 (N_17304,N_15705,N_14662);
and U17305 (N_17305,N_14850,N_14196);
and U17306 (N_17306,N_14255,N_15520);
nor U17307 (N_17307,N_14577,N_15234);
or U17308 (N_17308,N_14871,N_15174);
and U17309 (N_17309,N_15675,N_15921);
or U17310 (N_17310,N_14445,N_14307);
nor U17311 (N_17311,N_14373,N_14409);
and U17312 (N_17312,N_15749,N_15359);
nor U17313 (N_17313,N_14295,N_14165);
or U17314 (N_17314,N_15667,N_14147);
nand U17315 (N_17315,N_15813,N_14358);
nand U17316 (N_17316,N_14503,N_14511);
and U17317 (N_17317,N_15959,N_14413);
and U17318 (N_17318,N_14827,N_14127);
and U17319 (N_17319,N_14711,N_14013);
nand U17320 (N_17320,N_15002,N_15367);
nor U17321 (N_17321,N_15389,N_15368);
nand U17322 (N_17322,N_15640,N_15490);
or U17323 (N_17323,N_15491,N_15753);
and U17324 (N_17324,N_14328,N_14667);
or U17325 (N_17325,N_15750,N_15800);
or U17326 (N_17326,N_14324,N_14538);
and U17327 (N_17327,N_14127,N_14809);
nor U17328 (N_17328,N_15054,N_14331);
and U17329 (N_17329,N_15165,N_14934);
and U17330 (N_17330,N_14725,N_15383);
nor U17331 (N_17331,N_15042,N_15682);
nor U17332 (N_17332,N_15154,N_14891);
nor U17333 (N_17333,N_15395,N_15241);
nor U17334 (N_17334,N_14510,N_14147);
and U17335 (N_17335,N_15336,N_15359);
nand U17336 (N_17336,N_14142,N_15811);
or U17337 (N_17337,N_15065,N_15025);
nor U17338 (N_17338,N_15912,N_14911);
nand U17339 (N_17339,N_14658,N_15157);
and U17340 (N_17340,N_14270,N_14003);
or U17341 (N_17341,N_15202,N_15705);
nand U17342 (N_17342,N_14556,N_14495);
nor U17343 (N_17343,N_15477,N_15495);
or U17344 (N_17344,N_14397,N_15187);
or U17345 (N_17345,N_15061,N_15667);
and U17346 (N_17346,N_14788,N_14868);
and U17347 (N_17347,N_15002,N_14636);
or U17348 (N_17348,N_14379,N_14636);
or U17349 (N_17349,N_14097,N_14827);
and U17350 (N_17350,N_14392,N_15459);
or U17351 (N_17351,N_15124,N_14633);
nand U17352 (N_17352,N_14453,N_15457);
or U17353 (N_17353,N_14348,N_14897);
xor U17354 (N_17354,N_15422,N_15269);
nor U17355 (N_17355,N_14629,N_15518);
and U17356 (N_17356,N_15473,N_15110);
nand U17357 (N_17357,N_15705,N_15058);
and U17358 (N_17358,N_14384,N_15982);
or U17359 (N_17359,N_14133,N_15641);
and U17360 (N_17360,N_14685,N_15678);
or U17361 (N_17361,N_14992,N_14695);
and U17362 (N_17362,N_15343,N_14747);
and U17363 (N_17363,N_14878,N_14414);
nor U17364 (N_17364,N_15885,N_14241);
or U17365 (N_17365,N_15986,N_14566);
or U17366 (N_17366,N_14024,N_14955);
nor U17367 (N_17367,N_15194,N_15943);
and U17368 (N_17368,N_15441,N_15066);
and U17369 (N_17369,N_14586,N_14858);
and U17370 (N_17370,N_14016,N_14214);
xnor U17371 (N_17371,N_14156,N_15471);
nand U17372 (N_17372,N_15160,N_14682);
xnor U17373 (N_17373,N_15332,N_14729);
and U17374 (N_17374,N_14968,N_14820);
nor U17375 (N_17375,N_15618,N_14394);
or U17376 (N_17376,N_14485,N_15038);
or U17377 (N_17377,N_15420,N_14941);
nor U17378 (N_17378,N_15923,N_14718);
or U17379 (N_17379,N_14259,N_15360);
nand U17380 (N_17380,N_14964,N_15085);
or U17381 (N_17381,N_15837,N_14851);
nor U17382 (N_17382,N_15257,N_15360);
nand U17383 (N_17383,N_15399,N_14122);
nor U17384 (N_17384,N_15179,N_14361);
or U17385 (N_17385,N_14412,N_15802);
nand U17386 (N_17386,N_14774,N_15765);
or U17387 (N_17387,N_14408,N_14121);
nor U17388 (N_17388,N_14248,N_14611);
nor U17389 (N_17389,N_14491,N_15056);
nor U17390 (N_17390,N_14097,N_14625);
or U17391 (N_17391,N_15298,N_14488);
or U17392 (N_17392,N_15200,N_15416);
nand U17393 (N_17393,N_15349,N_14760);
and U17394 (N_17394,N_15311,N_15640);
or U17395 (N_17395,N_14240,N_15535);
or U17396 (N_17396,N_15290,N_15890);
or U17397 (N_17397,N_14618,N_15439);
nor U17398 (N_17398,N_15904,N_14839);
nor U17399 (N_17399,N_14506,N_15938);
nor U17400 (N_17400,N_15550,N_15995);
or U17401 (N_17401,N_15801,N_14832);
and U17402 (N_17402,N_15609,N_14554);
nand U17403 (N_17403,N_14857,N_15799);
or U17404 (N_17404,N_15033,N_15658);
nor U17405 (N_17405,N_15772,N_14286);
or U17406 (N_17406,N_15641,N_15883);
xnor U17407 (N_17407,N_15544,N_15506);
nand U17408 (N_17408,N_14174,N_14585);
and U17409 (N_17409,N_15968,N_14091);
nand U17410 (N_17410,N_15529,N_14121);
nand U17411 (N_17411,N_15632,N_14905);
and U17412 (N_17412,N_14970,N_15126);
and U17413 (N_17413,N_15347,N_14091);
or U17414 (N_17414,N_14750,N_14451);
and U17415 (N_17415,N_14866,N_15583);
nand U17416 (N_17416,N_15921,N_15382);
nand U17417 (N_17417,N_14969,N_15686);
or U17418 (N_17418,N_15709,N_14886);
xnor U17419 (N_17419,N_14406,N_15212);
and U17420 (N_17420,N_15522,N_14062);
and U17421 (N_17421,N_14517,N_14742);
nor U17422 (N_17422,N_14804,N_14813);
and U17423 (N_17423,N_15642,N_15918);
nor U17424 (N_17424,N_14421,N_14040);
and U17425 (N_17425,N_14739,N_15498);
or U17426 (N_17426,N_14945,N_14761);
nand U17427 (N_17427,N_14459,N_14307);
nand U17428 (N_17428,N_14397,N_14895);
and U17429 (N_17429,N_15534,N_15332);
or U17430 (N_17430,N_15807,N_14953);
xor U17431 (N_17431,N_15779,N_14456);
and U17432 (N_17432,N_14627,N_14330);
nand U17433 (N_17433,N_15800,N_14500);
nand U17434 (N_17434,N_15452,N_14051);
or U17435 (N_17435,N_15913,N_15064);
nor U17436 (N_17436,N_14050,N_14877);
nand U17437 (N_17437,N_14397,N_14400);
nand U17438 (N_17438,N_15337,N_14249);
or U17439 (N_17439,N_14389,N_14985);
nand U17440 (N_17440,N_15397,N_14542);
and U17441 (N_17441,N_15223,N_15194);
nor U17442 (N_17442,N_15746,N_14458);
and U17443 (N_17443,N_14916,N_15847);
nand U17444 (N_17444,N_15681,N_14134);
nand U17445 (N_17445,N_14937,N_15128);
and U17446 (N_17446,N_15365,N_15233);
and U17447 (N_17447,N_14419,N_15324);
nor U17448 (N_17448,N_15450,N_14361);
nor U17449 (N_17449,N_14521,N_14255);
or U17450 (N_17450,N_15286,N_14732);
nor U17451 (N_17451,N_14732,N_15986);
or U17452 (N_17452,N_14245,N_15878);
or U17453 (N_17453,N_15963,N_15203);
or U17454 (N_17454,N_15402,N_15093);
nand U17455 (N_17455,N_14569,N_15349);
or U17456 (N_17456,N_14064,N_14702);
or U17457 (N_17457,N_14980,N_15413);
and U17458 (N_17458,N_15363,N_14531);
nor U17459 (N_17459,N_15389,N_15083);
or U17460 (N_17460,N_14266,N_14026);
nor U17461 (N_17461,N_14431,N_14999);
and U17462 (N_17462,N_15424,N_15633);
or U17463 (N_17463,N_15238,N_15908);
or U17464 (N_17464,N_14877,N_15945);
or U17465 (N_17465,N_14592,N_15823);
or U17466 (N_17466,N_15600,N_15897);
and U17467 (N_17467,N_14188,N_15367);
nor U17468 (N_17468,N_15869,N_14751);
and U17469 (N_17469,N_15781,N_14003);
nand U17470 (N_17470,N_15415,N_14658);
nand U17471 (N_17471,N_14206,N_14428);
or U17472 (N_17472,N_14464,N_14891);
and U17473 (N_17473,N_14189,N_14465);
and U17474 (N_17474,N_14956,N_14925);
or U17475 (N_17475,N_15205,N_15941);
nand U17476 (N_17476,N_15439,N_15689);
and U17477 (N_17477,N_14716,N_15913);
nor U17478 (N_17478,N_14727,N_14797);
xnor U17479 (N_17479,N_15989,N_15465);
and U17480 (N_17480,N_14404,N_14150);
nand U17481 (N_17481,N_14574,N_14212);
nand U17482 (N_17482,N_14919,N_14865);
or U17483 (N_17483,N_15326,N_14882);
and U17484 (N_17484,N_14075,N_15056);
nand U17485 (N_17485,N_15436,N_14459);
nor U17486 (N_17486,N_14260,N_14939);
nor U17487 (N_17487,N_15610,N_15492);
or U17488 (N_17488,N_14678,N_14734);
nand U17489 (N_17489,N_14891,N_15249);
nor U17490 (N_17490,N_15941,N_14621);
nor U17491 (N_17491,N_15958,N_14625);
and U17492 (N_17492,N_15784,N_15541);
nor U17493 (N_17493,N_15218,N_15733);
nor U17494 (N_17494,N_15214,N_15983);
or U17495 (N_17495,N_14134,N_15132);
nand U17496 (N_17496,N_15356,N_14990);
nor U17497 (N_17497,N_15162,N_15009);
or U17498 (N_17498,N_15338,N_15563);
nor U17499 (N_17499,N_15958,N_14470);
nand U17500 (N_17500,N_14860,N_15424);
nor U17501 (N_17501,N_15630,N_14391);
or U17502 (N_17502,N_14850,N_15043);
nand U17503 (N_17503,N_14092,N_14420);
nor U17504 (N_17504,N_14329,N_15881);
nand U17505 (N_17505,N_14112,N_15562);
xnor U17506 (N_17506,N_14044,N_14816);
or U17507 (N_17507,N_15946,N_14786);
nand U17508 (N_17508,N_14083,N_14865);
and U17509 (N_17509,N_14106,N_14190);
or U17510 (N_17510,N_14545,N_14582);
or U17511 (N_17511,N_14714,N_15670);
nor U17512 (N_17512,N_15912,N_14788);
nand U17513 (N_17513,N_14591,N_15391);
and U17514 (N_17514,N_14857,N_15225);
and U17515 (N_17515,N_15542,N_14091);
nand U17516 (N_17516,N_15354,N_14903);
or U17517 (N_17517,N_15043,N_15021);
xor U17518 (N_17518,N_15391,N_14907);
and U17519 (N_17519,N_14955,N_14972);
or U17520 (N_17520,N_14937,N_14350);
and U17521 (N_17521,N_14719,N_15591);
nor U17522 (N_17522,N_14265,N_15410);
nand U17523 (N_17523,N_14646,N_15446);
and U17524 (N_17524,N_15429,N_14866);
or U17525 (N_17525,N_15791,N_14861);
or U17526 (N_17526,N_15818,N_15379);
nor U17527 (N_17527,N_14652,N_15753);
nand U17528 (N_17528,N_14311,N_14354);
nand U17529 (N_17529,N_15556,N_15657);
nor U17530 (N_17530,N_14355,N_15155);
nand U17531 (N_17531,N_14316,N_15446);
and U17532 (N_17532,N_14670,N_15699);
and U17533 (N_17533,N_14240,N_15844);
or U17534 (N_17534,N_15570,N_14483);
nor U17535 (N_17535,N_14164,N_14623);
and U17536 (N_17536,N_15991,N_15379);
nand U17537 (N_17537,N_15571,N_14143);
nor U17538 (N_17538,N_15287,N_14287);
and U17539 (N_17539,N_14163,N_15800);
or U17540 (N_17540,N_14535,N_14820);
and U17541 (N_17541,N_15658,N_15877);
nor U17542 (N_17542,N_14410,N_15236);
xor U17543 (N_17543,N_15747,N_15479);
nor U17544 (N_17544,N_14559,N_15757);
nor U17545 (N_17545,N_15846,N_15228);
nor U17546 (N_17546,N_14739,N_14655);
nand U17547 (N_17547,N_14278,N_14243);
nand U17548 (N_17548,N_15963,N_15424);
nand U17549 (N_17549,N_14787,N_15227);
and U17550 (N_17550,N_15683,N_14952);
nor U17551 (N_17551,N_15221,N_15320);
xor U17552 (N_17552,N_15969,N_14662);
nand U17553 (N_17553,N_14551,N_14075);
or U17554 (N_17554,N_15940,N_15577);
and U17555 (N_17555,N_15280,N_14486);
and U17556 (N_17556,N_15863,N_15843);
nand U17557 (N_17557,N_14327,N_14735);
or U17558 (N_17558,N_14176,N_15188);
nor U17559 (N_17559,N_14233,N_14928);
and U17560 (N_17560,N_14540,N_14817);
or U17561 (N_17561,N_14810,N_14344);
and U17562 (N_17562,N_15900,N_14364);
nor U17563 (N_17563,N_15304,N_15460);
or U17564 (N_17564,N_15453,N_14633);
nor U17565 (N_17565,N_15773,N_15951);
or U17566 (N_17566,N_15639,N_15056);
or U17567 (N_17567,N_15555,N_14124);
nand U17568 (N_17568,N_15934,N_15807);
nor U17569 (N_17569,N_15699,N_14218);
nand U17570 (N_17570,N_14692,N_14455);
or U17571 (N_17571,N_15889,N_15878);
or U17572 (N_17572,N_14111,N_14928);
and U17573 (N_17573,N_15482,N_15295);
nand U17574 (N_17574,N_15252,N_14491);
nand U17575 (N_17575,N_14893,N_15727);
nand U17576 (N_17576,N_14116,N_15958);
nand U17577 (N_17577,N_15306,N_14532);
or U17578 (N_17578,N_14776,N_14292);
nand U17579 (N_17579,N_15136,N_15543);
nor U17580 (N_17580,N_15048,N_15642);
and U17581 (N_17581,N_15764,N_15867);
nor U17582 (N_17582,N_15161,N_14103);
nand U17583 (N_17583,N_15028,N_15867);
or U17584 (N_17584,N_14515,N_15302);
or U17585 (N_17585,N_14427,N_15549);
nand U17586 (N_17586,N_14116,N_14069);
or U17587 (N_17587,N_14877,N_15199);
nor U17588 (N_17588,N_15134,N_15449);
nor U17589 (N_17589,N_14058,N_15643);
and U17590 (N_17590,N_15991,N_14525);
xor U17591 (N_17591,N_14958,N_15688);
and U17592 (N_17592,N_15817,N_14065);
nand U17593 (N_17593,N_14618,N_14101);
or U17594 (N_17594,N_14307,N_14389);
xnor U17595 (N_17595,N_14361,N_15819);
nand U17596 (N_17596,N_15076,N_14204);
nor U17597 (N_17597,N_14882,N_14340);
nand U17598 (N_17598,N_15221,N_14303);
and U17599 (N_17599,N_14094,N_15202);
or U17600 (N_17600,N_14681,N_15396);
nor U17601 (N_17601,N_15047,N_14720);
and U17602 (N_17602,N_15330,N_15206);
or U17603 (N_17603,N_14544,N_15633);
nand U17604 (N_17604,N_15904,N_14948);
or U17605 (N_17605,N_15710,N_14298);
nor U17606 (N_17606,N_14400,N_15822);
and U17607 (N_17607,N_15348,N_15493);
nor U17608 (N_17608,N_15369,N_14932);
and U17609 (N_17609,N_15217,N_14212);
nor U17610 (N_17610,N_14108,N_15443);
nor U17611 (N_17611,N_15426,N_15969);
or U17612 (N_17612,N_15290,N_14350);
nor U17613 (N_17613,N_14009,N_14454);
nand U17614 (N_17614,N_14847,N_15293);
and U17615 (N_17615,N_15027,N_15938);
nor U17616 (N_17616,N_14354,N_14809);
and U17617 (N_17617,N_14686,N_15688);
nand U17618 (N_17618,N_15023,N_15598);
and U17619 (N_17619,N_14386,N_14510);
or U17620 (N_17620,N_14310,N_15011);
nor U17621 (N_17621,N_15977,N_14179);
nand U17622 (N_17622,N_14388,N_15511);
nor U17623 (N_17623,N_14193,N_15595);
or U17624 (N_17624,N_15048,N_15437);
nor U17625 (N_17625,N_15459,N_14697);
and U17626 (N_17626,N_15792,N_14464);
nand U17627 (N_17627,N_15001,N_14393);
and U17628 (N_17628,N_14600,N_14245);
nand U17629 (N_17629,N_14847,N_15287);
or U17630 (N_17630,N_14621,N_14422);
nand U17631 (N_17631,N_14394,N_14744);
nand U17632 (N_17632,N_14836,N_14947);
nor U17633 (N_17633,N_15273,N_15937);
nand U17634 (N_17634,N_15129,N_14889);
or U17635 (N_17635,N_15641,N_14625);
nor U17636 (N_17636,N_15813,N_14661);
nor U17637 (N_17637,N_14954,N_14894);
and U17638 (N_17638,N_15969,N_15820);
nor U17639 (N_17639,N_14745,N_15488);
and U17640 (N_17640,N_14869,N_15128);
and U17641 (N_17641,N_14755,N_14560);
and U17642 (N_17642,N_15542,N_15729);
and U17643 (N_17643,N_14016,N_15440);
and U17644 (N_17644,N_15196,N_15555);
and U17645 (N_17645,N_14406,N_14691);
or U17646 (N_17646,N_14746,N_14507);
nor U17647 (N_17647,N_14173,N_15386);
nand U17648 (N_17648,N_14270,N_15021);
and U17649 (N_17649,N_14897,N_15501);
or U17650 (N_17650,N_15368,N_15382);
nor U17651 (N_17651,N_15197,N_15404);
nand U17652 (N_17652,N_15998,N_15452);
nand U17653 (N_17653,N_14539,N_15015);
nor U17654 (N_17654,N_15854,N_14772);
nand U17655 (N_17655,N_14209,N_14107);
nand U17656 (N_17656,N_15869,N_15358);
nand U17657 (N_17657,N_14626,N_14050);
or U17658 (N_17658,N_15127,N_15547);
or U17659 (N_17659,N_14851,N_15061);
or U17660 (N_17660,N_14163,N_15663);
nand U17661 (N_17661,N_14476,N_14026);
xor U17662 (N_17662,N_15193,N_15335);
nand U17663 (N_17663,N_15348,N_14027);
and U17664 (N_17664,N_15724,N_15327);
nor U17665 (N_17665,N_15168,N_15750);
nor U17666 (N_17666,N_15268,N_14087);
and U17667 (N_17667,N_15602,N_14490);
and U17668 (N_17668,N_15092,N_14447);
nand U17669 (N_17669,N_15137,N_15304);
or U17670 (N_17670,N_14548,N_14302);
or U17671 (N_17671,N_14008,N_15998);
xnor U17672 (N_17672,N_15139,N_15058);
and U17673 (N_17673,N_15978,N_14322);
or U17674 (N_17674,N_15194,N_14010);
nor U17675 (N_17675,N_15504,N_14153);
xnor U17676 (N_17676,N_15951,N_14438);
and U17677 (N_17677,N_15986,N_14011);
and U17678 (N_17678,N_15882,N_14475);
or U17679 (N_17679,N_15712,N_14572);
nand U17680 (N_17680,N_15401,N_14122);
or U17681 (N_17681,N_14691,N_14476);
and U17682 (N_17682,N_14863,N_15963);
or U17683 (N_17683,N_15359,N_15846);
or U17684 (N_17684,N_14935,N_15786);
nor U17685 (N_17685,N_15954,N_14538);
and U17686 (N_17686,N_14223,N_14380);
nand U17687 (N_17687,N_15938,N_14210);
nor U17688 (N_17688,N_15423,N_15030);
nor U17689 (N_17689,N_15062,N_15567);
or U17690 (N_17690,N_14346,N_14842);
and U17691 (N_17691,N_14529,N_15804);
or U17692 (N_17692,N_15119,N_15567);
and U17693 (N_17693,N_15985,N_15635);
nor U17694 (N_17694,N_15382,N_14795);
and U17695 (N_17695,N_14516,N_15039);
nor U17696 (N_17696,N_14177,N_15595);
nand U17697 (N_17697,N_14858,N_14533);
or U17698 (N_17698,N_14113,N_15604);
or U17699 (N_17699,N_15145,N_14173);
nand U17700 (N_17700,N_14885,N_15776);
nor U17701 (N_17701,N_15977,N_14242);
and U17702 (N_17702,N_14134,N_14642);
nand U17703 (N_17703,N_14322,N_15030);
and U17704 (N_17704,N_15014,N_14836);
and U17705 (N_17705,N_15121,N_15946);
and U17706 (N_17706,N_14205,N_15647);
or U17707 (N_17707,N_15018,N_14685);
nand U17708 (N_17708,N_15475,N_14054);
nand U17709 (N_17709,N_15043,N_14250);
or U17710 (N_17710,N_14318,N_15614);
or U17711 (N_17711,N_15607,N_15651);
nand U17712 (N_17712,N_15184,N_14299);
nand U17713 (N_17713,N_15884,N_14867);
and U17714 (N_17714,N_14509,N_15350);
and U17715 (N_17715,N_15445,N_15500);
nor U17716 (N_17716,N_14415,N_14134);
or U17717 (N_17717,N_15518,N_14963);
nand U17718 (N_17718,N_15648,N_15738);
or U17719 (N_17719,N_14329,N_14408);
nand U17720 (N_17720,N_15018,N_14943);
xor U17721 (N_17721,N_15344,N_14805);
nor U17722 (N_17722,N_15679,N_15826);
and U17723 (N_17723,N_14095,N_15345);
nand U17724 (N_17724,N_15488,N_14740);
xor U17725 (N_17725,N_14002,N_15371);
or U17726 (N_17726,N_14623,N_14342);
and U17727 (N_17727,N_15597,N_15758);
nand U17728 (N_17728,N_14044,N_15083);
nand U17729 (N_17729,N_15735,N_15747);
or U17730 (N_17730,N_15887,N_14951);
and U17731 (N_17731,N_15259,N_14276);
xor U17732 (N_17732,N_14083,N_15793);
nand U17733 (N_17733,N_14187,N_15062);
and U17734 (N_17734,N_14685,N_15661);
and U17735 (N_17735,N_14768,N_14817);
and U17736 (N_17736,N_14547,N_14414);
nand U17737 (N_17737,N_14759,N_14503);
and U17738 (N_17738,N_14464,N_14315);
nand U17739 (N_17739,N_14319,N_14747);
or U17740 (N_17740,N_14800,N_15146);
and U17741 (N_17741,N_14382,N_15063);
or U17742 (N_17742,N_14676,N_14440);
nor U17743 (N_17743,N_14120,N_14611);
nor U17744 (N_17744,N_15785,N_14776);
nor U17745 (N_17745,N_15549,N_15957);
and U17746 (N_17746,N_14756,N_14129);
or U17747 (N_17747,N_15696,N_14535);
nand U17748 (N_17748,N_14159,N_14574);
and U17749 (N_17749,N_14700,N_15738);
nand U17750 (N_17750,N_15275,N_15131);
nand U17751 (N_17751,N_15993,N_15669);
and U17752 (N_17752,N_15900,N_15096);
and U17753 (N_17753,N_14365,N_15126);
and U17754 (N_17754,N_14219,N_15350);
or U17755 (N_17755,N_15060,N_14533);
or U17756 (N_17756,N_14092,N_14382);
nor U17757 (N_17757,N_14270,N_14595);
or U17758 (N_17758,N_15843,N_15245);
nand U17759 (N_17759,N_15290,N_14111);
nand U17760 (N_17760,N_14156,N_15336);
and U17761 (N_17761,N_14763,N_15664);
nor U17762 (N_17762,N_15571,N_15762);
or U17763 (N_17763,N_15130,N_15483);
nor U17764 (N_17764,N_15854,N_14768);
nand U17765 (N_17765,N_15442,N_15090);
nand U17766 (N_17766,N_15042,N_14610);
or U17767 (N_17767,N_15280,N_14407);
nand U17768 (N_17768,N_14302,N_14567);
nand U17769 (N_17769,N_15295,N_15322);
and U17770 (N_17770,N_15948,N_15410);
and U17771 (N_17771,N_15968,N_14574);
and U17772 (N_17772,N_14898,N_15309);
nor U17773 (N_17773,N_15035,N_14947);
nand U17774 (N_17774,N_14333,N_15444);
nand U17775 (N_17775,N_14084,N_14761);
nor U17776 (N_17776,N_15743,N_15827);
or U17777 (N_17777,N_14330,N_14470);
nor U17778 (N_17778,N_14119,N_15420);
nor U17779 (N_17779,N_15573,N_14610);
and U17780 (N_17780,N_14826,N_15030);
or U17781 (N_17781,N_15386,N_15165);
and U17782 (N_17782,N_15876,N_15616);
nor U17783 (N_17783,N_14934,N_14353);
nor U17784 (N_17784,N_15276,N_14559);
nand U17785 (N_17785,N_15187,N_15899);
or U17786 (N_17786,N_15498,N_14560);
or U17787 (N_17787,N_15709,N_15713);
and U17788 (N_17788,N_15267,N_14522);
or U17789 (N_17789,N_14741,N_14218);
or U17790 (N_17790,N_14247,N_14905);
or U17791 (N_17791,N_15980,N_15073);
nand U17792 (N_17792,N_15653,N_15924);
nand U17793 (N_17793,N_15853,N_15053);
nand U17794 (N_17794,N_14145,N_14916);
and U17795 (N_17795,N_15788,N_14307);
or U17796 (N_17796,N_15954,N_15856);
xnor U17797 (N_17797,N_15633,N_14996);
and U17798 (N_17798,N_15622,N_15360);
nand U17799 (N_17799,N_15780,N_14939);
or U17800 (N_17800,N_14441,N_15965);
or U17801 (N_17801,N_14826,N_14882);
and U17802 (N_17802,N_15176,N_14901);
nor U17803 (N_17803,N_15992,N_15707);
nand U17804 (N_17804,N_14314,N_14196);
or U17805 (N_17805,N_14486,N_14224);
nor U17806 (N_17806,N_15790,N_14747);
or U17807 (N_17807,N_15374,N_14411);
and U17808 (N_17808,N_14214,N_15766);
or U17809 (N_17809,N_15747,N_15192);
or U17810 (N_17810,N_14611,N_15584);
nand U17811 (N_17811,N_14757,N_14874);
or U17812 (N_17812,N_14836,N_15854);
or U17813 (N_17813,N_15066,N_15680);
nand U17814 (N_17814,N_14629,N_15504);
nand U17815 (N_17815,N_15263,N_14433);
nand U17816 (N_17816,N_15052,N_15657);
nand U17817 (N_17817,N_14320,N_15332);
xor U17818 (N_17818,N_14307,N_14494);
nor U17819 (N_17819,N_15686,N_14138);
nand U17820 (N_17820,N_15113,N_15261);
nor U17821 (N_17821,N_14066,N_15526);
and U17822 (N_17822,N_14368,N_15571);
nand U17823 (N_17823,N_15997,N_14131);
or U17824 (N_17824,N_15764,N_15925);
nand U17825 (N_17825,N_15423,N_14530);
and U17826 (N_17826,N_14226,N_15980);
nand U17827 (N_17827,N_15916,N_15982);
or U17828 (N_17828,N_14301,N_15306);
or U17829 (N_17829,N_15495,N_15839);
or U17830 (N_17830,N_14709,N_14797);
nor U17831 (N_17831,N_15981,N_14974);
or U17832 (N_17832,N_14254,N_15095);
nand U17833 (N_17833,N_14523,N_14631);
nand U17834 (N_17834,N_15087,N_15580);
or U17835 (N_17835,N_15168,N_14748);
and U17836 (N_17836,N_14656,N_15714);
nand U17837 (N_17837,N_14516,N_15226);
or U17838 (N_17838,N_15765,N_15068);
nor U17839 (N_17839,N_15819,N_15192);
nand U17840 (N_17840,N_15349,N_14862);
and U17841 (N_17841,N_15547,N_14250);
nand U17842 (N_17842,N_14985,N_14581);
nand U17843 (N_17843,N_14677,N_15173);
nor U17844 (N_17844,N_14639,N_15160);
nor U17845 (N_17845,N_14818,N_15280);
xor U17846 (N_17846,N_15689,N_15644);
nand U17847 (N_17847,N_15211,N_14099);
nor U17848 (N_17848,N_15608,N_14605);
nand U17849 (N_17849,N_15125,N_14879);
nor U17850 (N_17850,N_15210,N_14234);
and U17851 (N_17851,N_15674,N_15148);
nand U17852 (N_17852,N_14273,N_14043);
and U17853 (N_17853,N_14882,N_15953);
nand U17854 (N_17854,N_14000,N_14101);
and U17855 (N_17855,N_14296,N_14892);
nand U17856 (N_17856,N_15195,N_15777);
or U17857 (N_17857,N_14901,N_14090);
and U17858 (N_17858,N_14114,N_15217);
nor U17859 (N_17859,N_15123,N_14195);
nor U17860 (N_17860,N_14783,N_15703);
and U17861 (N_17861,N_15576,N_15917);
nor U17862 (N_17862,N_14065,N_14035);
or U17863 (N_17863,N_14319,N_15845);
and U17864 (N_17864,N_15417,N_15585);
nand U17865 (N_17865,N_14765,N_14419);
nand U17866 (N_17866,N_14070,N_14093);
xor U17867 (N_17867,N_14490,N_14801);
nor U17868 (N_17868,N_15824,N_15265);
or U17869 (N_17869,N_14219,N_15954);
nand U17870 (N_17870,N_14133,N_14364);
nand U17871 (N_17871,N_15291,N_14134);
nand U17872 (N_17872,N_14690,N_15027);
and U17873 (N_17873,N_14392,N_14758);
and U17874 (N_17874,N_15979,N_14982);
nand U17875 (N_17875,N_14259,N_15658);
and U17876 (N_17876,N_15769,N_14315);
nand U17877 (N_17877,N_15352,N_15687);
nor U17878 (N_17878,N_15386,N_15245);
nor U17879 (N_17879,N_14664,N_14026);
nand U17880 (N_17880,N_15330,N_15307);
xnor U17881 (N_17881,N_15310,N_15908);
nand U17882 (N_17882,N_14867,N_15894);
or U17883 (N_17883,N_14801,N_15863);
nor U17884 (N_17884,N_14808,N_15830);
or U17885 (N_17885,N_14475,N_15048);
and U17886 (N_17886,N_14668,N_14729);
nand U17887 (N_17887,N_15799,N_15882);
and U17888 (N_17888,N_14643,N_14794);
nand U17889 (N_17889,N_14655,N_14314);
or U17890 (N_17890,N_14827,N_15567);
nor U17891 (N_17891,N_14350,N_15404);
nand U17892 (N_17892,N_14137,N_15634);
nand U17893 (N_17893,N_15377,N_14158);
nor U17894 (N_17894,N_15522,N_14850);
nand U17895 (N_17895,N_15901,N_15813);
and U17896 (N_17896,N_14318,N_14648);
and U17897 (N_17897,N_15526,N_14522);
nand U17898 (N_17898,N_15880,N_14169);
nand U17899 (N_17899,N_14592,N_14090);
nor U17900 (N_17900,N_14204,N_14607);
and U17901 (N_17901,N_15308,N_14963);
or U17902 (N_17902,N_15189,N_14687);
nor U17903 (N_17903,N_15381,N_14233);
nor U17904 (N_17904,N_15455,N_15100);
or U17905 (N_17905,N_14179,N_15314);
and U17906 (N_17906,N_14697,N_14180);
and U17907 (N_17907,N_14527,N_14460);
and U17908 (N_17908,N_14786,N_14339);
nor U17909 (N_17909,N_15646,N_14442);
and U17910 (N_17910,N_14739,N_14062);
and U17911 (N_17911,N_15269,N_15270);
and U17912 (N_17912,N_15793,N_15713);
or U17913 (N_17913,N_15359,N_14981);
or U17914 (N_17914,N_14136,N_14095);
nand U17915 (N_17915,N_15604,N_14200);
nand U17916 (N_17916,N_14263,N_14975);
or U17917 (N_17917,N_14838,N_15223);
or U17918 (N_17918,N_15069,N_15910);
nand U17919 (N_17919,N_14809,N_14031);
nand U17920 (N_17920,N_15343,N_14622);
and U17921 (N_17921,N_14188,N_14372);
nand U17922 (N_17922,N_14255,N_15900);
and U17923 (N_17923,N_14762,N_15968);
nor U17924 (N_17924,N_14238,N_14016);
nand U17925 (N_17925,N_15553,N_14219);
or U17926 (N_17926,N_14995,N_15910);
nand U17927 (N_17927,N_14957,N_14366);
nor U17928 (N_17928,N_14620,N_15278);
nor U17929 (N_17929,N_15292,N_15768);
nand U17930 (N_17930,N_15890,N_14839);
nand U17931 (N_17931,N_15108,N_14810);
or U17932 (N_17932,N_14228,N_14183);
or U17933 (N_17933,N_14657,N_14787);
nand U17934 (N_17934,N_15256,N_15373);
nor U17935 (N_17935,N_14914,N_15915);
or U17936 (N_17936,N_15858,N_15397);
nor U17937 (N_17937,N_15814,N_14451);
or U17938 (N_17938,N_14013,N_15053);
or U17939 (N_17939,N_14722,N_15510);
nand U17940 (N_17940,N_14352,N_14215);
or U17941 (N_17941,N_14489,N_14737);
or U17942 (N_17942,N_15132,N_15570);
xor U17943 (N_17943,N_15434,N_15042);
and U17944 (N_17944,N_15823,N_15078);
and U17945 (N_17945,N_14498,N_14488);
or U17946 (N_17946,N_15900,N_14241);
nor U17947 (N_17947,N_14763,N_14917);
nor U17948 (N_17948,N_14119,N_15677);
and U17949 (N_17949,N_14890,N_15877);
nor U17950 (N_17950,N_14907,N_15769);
nor U17951 (N_17951,N_15623,N_14108);
and U17952 (N_17952,N_15505,N_14338);
nand U17953 (N_17953,N_15182,N_15014);
and U17954 (N_17954,N_15219,N_15913);
and U17955 (N_17955,N_15273,N_15487);
nor U17956 (N_17956,N_15954,N_14779);
nor U17957 (N_17957,N_14671,N_15755);
nand U17958 (N_17958,N_14806,N_15985);
or U17959 (N_17959,N_14235,N_15533);
nor U17960 (N_17960,N_15401,N_14889);
and U17961 (N_17961,N_14826,N_15643);
xor U17962 (N_17962,N_14525,N_15218);
or U17963 (N_17963,N_14547,N_14191);
nand U17964 (N_17964,N_15508,N_15667);
nor U17965 (N_17965,N_15716,N_14815);
nand U17966 (N_17966,N_15096,N_15447);
and U17967 (N_17967,N_15956,N_14633);
nand U17968 (N_17968,N_14350,N_14130);
and U17969 (N_17969,N_15727,N_15502);
nor U17970 (N_17970,N_15549,N_14882);
nand U17971 (N_17971,N_15782,N_15759);
nor U17972 (N_17972,N_15535,N_15158);
nor U17973 (N_17973,N_14430,N_14545);
and U17974 (N_17974,N_14519,N_14332);
nand U17975 (N_17975,N_14079,N_15084);
nand U17976 (N_17976,N_14096,N_14502);
and U17977 (N_17977,N_15757,N_15646);
nand U17978 (N_17978,N_15902,N_14952);
nand U17979 (N_17979,N_14185,N_15747);
nand U17980 (N_17980,N_14824,N_15904);
or U17981 (N_17981,N_14608,N_15397);
and U17982 (N_17982,N_14274,N_14746);
or U17983 (N_17983,N_14325,N_15364);
and U17984 (N_17984,N_15641,N_15730);
nor U17985 (N_17985,N_14285,N_15531);
nand U17986 (N_17986,N_14636,N_15468);
and U17987 (N_17987,N_15031,N_15605);
or U17988 (N_17988,N_14099,N_14028);
nand U17989 (N_17989,N_14862,N_15351);
or U17990 (N_17990,N_14460,N_15470);
or U17991 (N_17991,N_15795,N_14551);
nor U17992 (N_17992,N_14063,N_15737);
nand U17993 (N_17993,N_15138,N_15077);
nor U17994 (N_17994,N_15344,N_14337);
nand U17995 (N_17995,N_15197,N_15709);
nor U17996 (N_17996,N_14743,N_14134);
or U17997 (N_17997,N_15078,N_15931);
or U17998 (N_17998,N_15856,N_15438);
nor U17999 (N_17999,N_15368,N_14959);
and U18000 (N_18000,N_17483,N_16165);
or U18001 (N_18001,N_16463,N_17232);
or U18002 (N_18002,N_17616,N_16903);
and U18003 (N_18003,N_17996,N_16789);
and U18004 (N_18004,N_17693,N_16772);
nand U18005 (N_18005,N_17205,N_16769);
and U18006 (N_18006,N_16971,N_16107);
nand U18007 (N_18007,N_17136,N_17311);
and U18008 (N_18008,N_16965,N_17757);
or U18009 (N_18009,N_17192,N_17864);
nand U18010 (N_18010,N_16521,N_16699);
xor U18011 (N_18011,N_17357,N_16090);
or U18012 (N_18012,N_17097,N_16986);
nand U18013 (N_18013,N_16342,N_16371);
or U18014 (N_18014,N_17404,N_16786);
nand U18015 (N_18015,N_16201,N_17953);
nor U18016 (N_18016,N_16730,N_16678);
or U18017 (N_18017,N_16008,N_17037);
and U18018 (N_18018,N_16207,N_16992);
or U18019 (N_18019,N_17204,N_16263);
nor U18020 (N_18020,N_16141,N_17689);
nor U18021 (N_18021,N_17094,N_16654);
nand U18022 (N_18022,N_17303,N_16924);
nand U18023 (N_18023,N_17180,N_17459);
nand U18024 (N_18024,N_16102,N_16227);
nor U18025 (N_18025,N_16630,N_16778);
nor U18026 (N_18026,N_17776,N_17096);
nand U18027 (N_18027,N_17806,N_17251);
and U18028 (N_18028,N_16639,N_17805);
and U18029 (N_18029,N_17383,N_17932);
or U18030 (N_18030,N_17329,N_16100);
nor U18031 (N_18031,N_16856,N_16776);
or U18032 (N_18032,N_17914,N_16602);
nand U18033 (N_18033,N_17351,N_16503);
xor U18034 (N_18034,N_16363,N_16477);
or U18035 (N_18035,N_17601,N_17712);
nor U18036 (N_18036,N_17590,N_16328);
nor U18037 (N_18037,N_17596,N_17868);
xor U18038 (N_18038,N_16331,N_16407);
or U18039 (N_18039,N_16397,N_16016);
nor U18040 (N_18040,N_17397,N_17252);
nand U18041 (N_18041,N_17895,N_17777);
nand U18042 (N_18042,N_16012,N_17988);
nor U18043 (N_18043,N_17721,N_17407);
nand U18044 (N_18044,N_16246,N_17659);
xnor U18045 (N_18045,N_17774,N_17390);
nor U18046 (N_18046,N_17955,N_16905);
nand U18047 (N_18047,N_17962,N_16105);
nand U18048 (N_18048,N_16711,N_17950);
or U18049 (N_18049,N_16533,N_16709);
or U18050 (N_18050,N_16714,N_16514);
nand U18051 (N_18051,N_17733,N_17993);
nand U18052 (N_18052,N_16039,N_16023);
or U18053 (N_18053,N_16115,N_17385);
and U18054 (N_18054,N_17235,N_17754);
or U18055 (N_18055,N_17644,N_16546);
or U18056 (N_18056,N_16914,N_17770);
nand U18057 (N_18057,N_17358,N_16918);
or U18058 (N_18058,N_17120,N_16750);
nor U18059 (N_18059,N_17954,N_16351);
or U18060 (N_18060,N_16579,N_16308);
nor U18061 (N_18061,N_16266,N_17620);
nor U18062 (N_18062,N_16401,N_17403);
nor U18063 (N_18063,N_17038,N_17840);
xor U18064 (N_18064,N_16731,N_17849);
and U18065 (N_18065,N_16700,N_17700);
nand U18066 (N_18066,N_16632,N_17579);
or U18067 (N_18067,N_16673,N_17449);
nor U18068 (N_18068,N_16078,N_16495);
nand U18069 (N_18069,N_17133,N_17692);
and U18070 (N_18070,N_16135,N_16239);
nand U18071 (N_18071,N_16287,N_16046);
and U18072 (N_18072,N_16823,N_17285);
or U18073 (N_18073,N_16961,N_16468);
or U18074 (N_18074,N_16457,N_17345);
and U18075 (N_18075,N_17441,N_16313);
nand U18076 (N_18076,N_16524,N_16493);
nand U18077 (N_18077,N_17049,N_17350);
nand U18078 (N_18078,N_16688,N_16480);
nand U18079 (N_18079,N_16808,N_17947);
and U18080 (N_18080,N_16164,N_17181);
nor U18081 (N_18081,N_17978,N_16913);
nand U18082 (N_18082,N_16575,N_17123);
nor U18083 (N_18083,N_16230,N_16572);
and U18084 (N_18084,N_16253,N_17377);
and U18085 (N_18085,N_17142,N_17826);
and U18086 (N_18086,N_17023,N_17608);
nand U18087 (N_18087,N_16676,N_16446);
nand U18088 (N_18088,N_16416,N_17876);
or U18089 (N_18089,N_16071,N_16220);
xor U18090 (N_18090,N_17663,N_17881);
nand U18091 (N_18091,N_17786,N_17543);
nand U18092 (N_18092,N_16968,N_16073);
nor U18093 (N_18093,N_17905,N_16215);
and U18094 (N_18094,N_16228,N_17160);
nand U18095 (N_18095,N_16174,N_16364);
nand U18096 (N_18096,N_16947,N_16015);
nand U18097 (N_18097,N_17773,N_17986);
nor U18098 (N_18098,N_17005,N_16561);
nand U18099 (N_18099,N_16854,N_16837);
or U18100 (N_18100,N_16086,N_17018);
or U18101 (N_18101,N_17839,N_16002);
or U18102 (N_18102,N_16460,N_17353);
or U18103 (N_18103,N_17413,N_17201);
xnor U18104 (N_18104,N_17316,N_16643);
or U18105 (N_18105,N_16264,N_16221);
or U18106 (N_18106,N_16832,N_16896);
xor U18107 (N_18107,N_17735,N_16798);
and U18108 (N_18108,N_16384,N_17995);
nor U18109 (N_18109,N_16329,N_16439);
and U18110 (N_18110,N_16562,N_16319);
nand U18111 (N_18111,N_17150,N_16010);
nor U18112 (N_18112,N_16285,N_16345);
or U18113 (N_18113,N_16093,N_17869);
xor U18114 (N_18114,N_16998,N_16325);
and U18115 (N_18115,N_17083,N_16171);
or U18116 (N_18116,N_17804,N_16564);
nand U18117 (N_18117,N_16193,N_16558);
nor U18118 (N_18118,N_17918,N_17071);
nor U18119 (N_18119,N_17172,N_16894);
or U18120 (N_18120,N_16578,N_16565);
and U18121 (N_18121,N_16208,N_17922);
nor U18122 (N_18122,N_16871,N_17571);
xnor U18123 (N_18123,N_17450,N_16611);
or U18124 (N_18124,N_16391,N_17730);
or U18125 (N_18125,N_17535,N_16752);
and U18126 (N_18126,N_16747,N_16534);
and U18127 (N_18127,N_17743,N_17639);
nand U18128 (N_18128,N_16199,N_17425);
nor U18129 (N_18129,N_16055,N_17338);
and U18130 (N_18130,N_17623,N_16790);
or U18131 (N_18131,N_16252,N_17082);
nand U18132 (N_18132,N_17705,N_17269);
and U18133 (N_18133,N_16846,N_17737);
nand U18134 (N_18134,N_16210,N_17820);
nor U18135 (N_18135,N_16890,N_17877);
and U18136 (N_18136,N_17313,N_17809);
or U18137 (N_18137,N_16383,N_17759);
and U18138 (N_18138,N_16153,N_17222);
or U18139 (N_18139,N_17362,N_16906);
and U18140 (N_18140,N_17501,N_16693);
or U18141 (N_18141,N_16559,N_17344);
nor U18142 (N_18142,N_17432,N_17707);
and U18143 (N_18143,N_17346,N_16919);
nor U18144 (N_18144,N_17304,N_17716);
nand U18145 (N_18145,N_17655,N_17174);
or U18146 (N_18146,N_16825,N_17164);
and U18147 (N_18147,N_17395,N_16029);
nor U18148 (N_18148,N_17831,N_16161);
and U18149 (N_18149,N_17283,N_17044);
nor U18150 (N_18150,N_17463,N_16792);
or U18151 (N_18151,N_16387,N_17498);
or U18152 (N_18152,N_16075,N_16447);
and U18153 (N_18153,N_16249,N_16347);
nor U18154 (N_18154,N_17966,N_17112);
or U18155 (N_18155,N_16712,N_17682);
and U18156 (N_18156,N_17155,N_17267);
or U18157 (N_18157,N_16819,N_16054);
and U18158 (N_18158,N_16062,N_16355);
and U18159 (N_18159,N_16694,N_16038);
nor U18160 (N_18160,N_16425,N_16036);
or U18161 (N_18161,N_16405,N_16257);
nor U18162 (N_18162,N_17504,N_17074);
and U18163 (N_18163,N_17446,N_17633);
nand U18164 (N_18164,N_16501,N_17324);
or U18165 (N_18165,N_16788,N_17141);
or U18166 (N_18166,N_17190,N_16321);
nand U18167 (N_18167,N_17366,N_17177);
or U18168 (N_18168,N_16516,N_16589);
or U18169 (N_18169,N_16779,N_16410);
or U18170 (N_18170,N_16560,N_16755);
nand U18171 (N_18171,N_16007,N_17423);
and U18172 (N_18172,N_16224,N_17593);
nand U18173 (N_18173,N_17704,N_17884);
nand U18174 (N_18174,N_17054,N_16354);
nor U18175 (N_18175,N_17720,N_17581);
and U18176 (N_18176,N_16125,N_16352);
xor U18177 (N_18177,N_17233,N_17878);
nand U18178 (N_18178,N_16991,N_17008);
nor U18179 (N_18179,N_16323,N_16889);
nor U18180 (N_18180,N_16830,N_16626);
nand U18181 (N_18181,N_16796,N_17926);
nand U18182 (N_18182,N_17781,N_17144);
xor U18183 (N_18183,N_17855,N_17032);
and U18184 (N_18184,N_16852,N_17104);
nor U18185 (N_18185,N_17551,N_16486);
and U18186 (N_18186,N_17166,N_16618);
xnor U18187 (N_18187,N_17455,N_17400);
and U18188 (N_18188,N_16622,N_17179);
and U18189 (N_18189,N_16022,N_16908);
and U18190 (N_18190,N_17974,N_17456);
nand U18191 (N_18191,N_16256,N_17768);
or U18192 (N_18192,N_16528,N_17277);
nand U18193 (N_18193,N_17440,N_16196);
and U18194 (N_18194,N_17125,N_16953);
or U18195 (N_18195,N_17280,N_16955);
nor U18196 (N_18196,N_16743,N_17788);
nand U18197 (N_18197,N_17959,N_17453);
and U18198 (N_18198,N_16584,N_16537);
and U18199 (N_18199,N_17135,N_17131);
and U18200 (N_18200,N_16982,N_16301);
and U18201 (N_18201,N_17508,N_17028);
and U18202 (N_18202,N_17430,N_16030);
nand U18203 (N_18203,N_17818,N_16720);
nand U18204 (N_18204,N_16721,N_16137);
or U18205 (N_18205,N_16651,N_16428);
nand U18206 (N_18206,N_16344,N_17860);
xnor U18207 (N_18207,N_16979,N_17187);
nand U18208 (N_18208,N_16981,N_17365);
nor U18209 (N_18209,N_16116,N_16163);
nor U18210 (N_18210,N_17584,N_16198);
or U18211 (N_18211,N_16686,N_16223);
or U18212 (N_18212,N_17520,N_16214);
and U18213 (N_18213,N_16422,N_17673);
and U18214 (N_18214,N_17750,N_17376);
nor U18215 (N_18215,N_16318,N_17796);
nor U18216 (N_18216,N_17184,N_17019);
nor U18217 (N_18217,N_17761,N_16204);
and U18218 (N_18218,N_17823,N_16745);
and U18219 (N_18219,N_17065,N_17600);
xor U18220 (N_18220,N_16722,N_17696);
nor U18221 (N_18221,N_16431,N_17281);
nand U18222 (N_18222,N_17474,N_16236);
and U18223 (N_18223,N_16304,N_17002);
nand U18224 (N_18224,N_16276,N_17732);
and U18225 (N_18225,N_17972,N_16631);
and U18226 (N_18226,N_17087,N_17416);
xor U18227 (N_18227,N_16567,N_16727);
nand U18228 (N_18228,N_17225,N_16060);
or U18229 (N_18229,N_17115,N_17359);
and U18230 (N_18230,N_16254,N_16286);
and U18231 (N_18231,N_16202,N_16094);
nor U18232 (N_18232,N_16737,N_17848);
or U18233 (N_18233,N_17319,N_17265);
nor U18234 (N_18234,N_17744,N_17489);
and U18235 (N_18235,N_17957,N_16520);
or U18236 (N_18236,N_17722,N_16195);
or U18237 (N_18237,N_17837,N_17368);
nor U18238 (N_18238,N_16741,N_17838);
nor U18239 (N_18239,N_16928,N_16705);
or U18240 (N_18240,N_17827,N_16096);
nand U18241 (N_18241,N_17891,N_17654);
and U18242 (N_18242,N_16290,N_17226);
nand U18243 (N_18243,N_16880,N_17529);
nand U18244 (N_18244,N_16716,N_17154);
nor U18245 (N_18245,N_16515,N_16603);
or U18246 (N_18246,N_16884,N_17863);
nand U18247 (N_18247,N_17098,N_17921);
nand U18248 (N_18248,N_16988,N_17470);
and U18249 (N_18249,N_17106,N_17794);
nor U18250 (N_18250,N_17219,N_16898);
nand U18251 (N_18251,N_17011,N_17143);
nand U18252 (N_18252,N_17845,N_17084);
nor U18253 (N_18253,N_17152,N_17515);
or U18254 (N_18254,N_17814,N_16203);
nor U18255 (N_18255,N_16244,N_17363);
nand U18256 (N_18256,N_17749,N_16629);
and U18257 (N_18257,N_16556,N_17477);
nor U18258 (N_18258,N_16628,N_16269);
and U18259 (N_18259,N_17045,N_17553);
or U18260 (N_18260,N_17020,N_17917);
or U18261 (N_18261,N_17024,N_17661);
nor U18262 (N_18262,N_17641,N_17215);
and U18263 (N_18263,N_17414,N_16018);
nor U18264 (N_18264,N_16103,N_16152);
nand U18265 (N_18265,N_16554,N_16118);
nand U18266 (N_18266,N_17386,N_16912);
or U18267 (N_18267,N_16280,N_16855);
nor U18268 (N_18268,N_17672,N_17719);
or U18269 (N_18269,N_17830,N_17853);
nand U18270 (N_18270,N_16718,N_16014);
and U18271 (N_18271,N_17657,N_17651);
nand U18272 (N_18272,N_17635,N_16307);
nand U18273 (N_18273,N_16858,N_17724);
and U18274 (N_18274,N_16975,N_16582);
nand U18275 (N_18275,N_17667,N_16300);
or U18276 (N_18276,N_16985,N_17238);
or U18277 (N_18277,N_17236,N_17521);
nor U18278 (N_18278,N_16272,N_17979);
nor U18279 (N_18279,N_16485,N_17828);
nor U18280 (N_18280,N_17492,N_17116);
nand U18281 (N_18281,N_17412,N_17307);
or U18282 (N_18282,N_16156,N_17524);
nand U18283 (N_18283,N_17454,N_17287);
nor U18284 (N_18284,N_17481,N_17075);
nor U18285 (N_18285,N_16150,N_17890);
and U18286 (N_18286,N_16188,N_17250);
and U18287 (N_18287,N_16027,N_16540);
nor U18288 (N_18288,N_17726,N_16803);
xor U18289 (N_18289,N_16978,N_17711);
and U18290 (N_18290,N_16162,N_17572);
xnor U18291 (N_18291,N_17512,N_17419);
and U18292 (N_18292,N_17186,N_16935);
or U18293 (N_18293,N_16824,N_17217);
or U18294 (N_18294,N_17852,N_16158);
and U18295 (N_18295,N_16609,N_16845);
nand U18296 (N_18296,N_16343,N_17069);
nor U18297 (N_18297,N_17901,N_16114);
and U18298 (N_18298,N_16166,N_16084);
xnor U18299 (N_18299,N_16419,N_17882);
nor U18300 (N_18300,N_17025,N_17478);
nor U18301 (N_18301,N_16146,N_17218);
and U18302 (N_18302,N_16186,N_16034);
or U18303 (N_18303,N_17077,N_16931);
and U18304 (N_18304,N_17113,N_16719);
nor U18305 (N_18305,N_16691,N_16672);
and U18306 (N_18306,N_17471,N_16512);
or U18307 (N_18307,N_16109,N_17613);
or U18308 (N_18308,N_17885,N_16375);
or U18309 (N_18309,N_16314,N_17452);
nor U18310 (N_18310,N_17829,N_17398);
or U18311 (N_18311,N_17740,N_16145);
nand U18312 (N_18312,N_17485,N_16240);
nand U18313 (N_18313,N_16795,N_17710);
nand U18314 (N_18314,N_16664,N_17899);
or U18315 (N_18315,N_17771,N_16996);
or U18316 (N_18316,N_16513,N_17022);
nand U18317 (N_18317,N_16461,N_17325);
nor U18318 (N_18318,N_16108,N_17337);
nor U18319 (N_18319,N_17968,N_16088);
nand U18320 (N_18320,N_16888,N_16066);
and U18321 (N_18321,N_16592,N_16069);
and U18322 (N_18322,N_17348,N_17634);
xnor U18323 (N_18323,N_16764,N_17631);
or U18324 (N_18324,N_17132,N_17162);
nand U18325 (N_18325,N_17628,N_17944);
nor U18326 (N_18326,N_17394,N_17632);
or U18327 (N_18327,N_17246,N_16357);
nor U18328 (N_18328,N_17956,N_17706);
nand U18329 (N_18329,N_17393,N_17637);
nor U18330 (N_18330,N_16878,N_16827);
or U18331 (N_18331,N_16759,N_16491);
nor U18332 (N_18332,N_17668,N_16518);
or U18333 (N_18333,N_17486,N_17896);
and U18334 (N_18334,N_16360,N_16641);
and U18335 (N_18335,N_16531,N_17057);
nand U18336 (N_18336,N_17843,N_16294);
or U18337 (N_18337,N_17658,N_17662);
or U18338 (N_18338,N_17102,N_16708);
or U18339 (N_18339,N_16011,N_16599);
or U18340 (N_18340,N_16510,N_17148);
or U18341 (N_18341,N_16543,N_17111);
nor U18342 (N_18342,N_17292,N_17118);
or U18343 (N_18343,N_16509,N_17514);
nor U18344 (N_18344,N_16092,N_16448);
or U18345 (N_18345,N_17598,N_17650);
nor U18346 (N_18346,N_17437,N_17785);
or U18347 (N_18347,N_17643,N_17167);
or U18348 (N_18348,N_17985,N_17417);
and U18349 (N_18349,N_16939,N_17681);
or U18350 (N_18350,N_17370,N_17427);
nor U18351 (N_18351,N_16068,N_17889);
nor U18352 (N_18352,N_16650,N_17952);
or U18353 (N_18353,N_16095,N_17124);
and U18354 (N_18354,N_16455,N_17945);
or U18355 (N_18355,N_17467,N_17434);
or U18356 (N_18356,N_16870,N_16762);
and U18357 (N_18357,N_16175,N_17775);
and U18358 (N_18358,N_16051,N_17791);
and U18359 (N_18359,N_16653,N_17942);
nor U18360 (N_18360,N_16526,N_16800);
nand U18361 (N_18361,N_16774,N_17612);
nand U18362 (N_18362,N_17062,N_17745);
and U18363 (N_18363,N_16972,N_17936);
nand U18364 (N_18364,N_16283,N_16710);
or U18365 (N_18365,N_17444,N_17159);
nand U18366 (N_18366,N_17989,N_16459);
or U18367 (N_18367,N_17193,N_17462);
xnor U18368 (N_18368,N_16427,N_16079);
nor U18369 (N_18369,N_16123,N_16306);
or U18370 (N_18370,N_16184,N_17381);
and U18371 (N_18371,N_16751,N_16452);
or U18372 (N_18372,N_16942,N_16047);
nand U18373 (N_18373,N_16121,N_17169);
or U18374 (N_18374,N_16392,N_17870);
nand U18375 (N_18375,N_17765,N_17356);
and U18376 (N_18376,N_16035,N_16793);
and U18377 (N_18377,N_17725,N_17058);
nor U18378 (N_18378,N_16771,N_16989);
or U18379 (N_18379,N_17731,N_17779);
nor U18380 (N_18380,N_16633,N_16385);
nor U18381 (N_18381,N_17971,N_16365);
or U18382 (N_18382,N_17802,N_16019);
nand U18383 (N_18383,N_16684,N_17259);
nor U18384 (N_18384,N_17085,N_17861);
and U18385 (N_18385,N_17999,N_17274);
or U18386 (N_18386,N_16061,N_17461);
or U18387 (N_18387,N_16568,N_16615);
and U18388 (N_18388,N_17421,N_17026);
and U18389 (N_18389,N_16332,N_17374);
and U18390 (N_18390,N_17448,N_16675);
nand U18391 (N_18391,N_16733,N_17599);
and U18392 (N_18392,N_16857,N_16267);
or U18393 (N_18393,N_16013,N_17886);
or U18394 (N_18394,N_17566,N_16566);
nor U18395 (N_18395,N_17076,N_16056);
nand U18396 (N_18396,N_16541,N_17624);
or U18397 (N_18397,N_17089,N_17927);
or U18398 (N_18398,N_16973,N_16966);
and U18399 (N_18399,N_17875,N_16140);
and U18400 (N_18400,N_16320,N_16951);
or U18401 (N_18401,N_16235,N_17286);
or U18402 (N_18402,N_16368,N_17582);
and U18403 (N_18403,N_17698,N_16867);
and U18404 (N_18404,N_17549,N_16143);
nand U18405 (N_18405,N_17306,N_17300);
and U18406 (N_18406,N_16634,N_17264);
nand U18407 (N_18407,N_17602,N_16963);
nand U18408 (N_18408,N_16736,N_17016);
or U18409 (N_18409,N_16232,N_17327);
nor U18410 (N_18410,N_16456,N_16479);
nor U18411 (N_18411,N_16433,N_16671);
or U18412 (N_18412,N_16481,N_17742);
or U18413 (N_18413,N_16934,N_16261);
and U18414 (N_18414,N_16372,N_17161);
or U18415 (N_18415,N_16806,N_17975);
or U18416 (N_18416,N_16802,N_17607);
and U18417 (N_18417,N_16941,N_17301);
nor U18418 (N_18418,N_16729,N_16563);
and U18419 (N_18419,N_16926,N_17604);
or U18420 (N_18420,N_16277,N_17816);
nor U18421 (N_18421,N_17790,N_17756);
nand U18422 (N_18422,N_16209,N_16883);
nand U18423 (N_18423,N_16804,N_16995);
and U18424 (N_18424,N_17556,N_17795);
or U18425 (N_18425,N_16732,N_17940);
nor U18426 (N_18426,N_17029,N_16770);
and U18427 (N_18427,N_16658,N_17064);
nand U18428 (N_18428,N_17906,N_17552);
nand U18429 (N_18429,N_16065,N_16801);
nor U18430 (N_18430,N_17925,N_17223);
nand U18431 (N_18431,N_16500,N_17982);
nand U18432 (N_18432,N_17239,N_17800);
or U18433 (N_18433,N_16117,N_17276);
or U18434 (N_18434,N_17920,N_17782);
nand U18435 (N_18435,N_17762,N_16190);
and U18436 (N_18436,N_17929,N_16504);
nand U18437 (N_18437,N_16176,N_16127);
nor U18438 (N_18438,N_16453,N_16134);
and U18439 (N_18439,N_16271,N_17561);
nand U18440 (N_18440,N_16369,N_16021);
nor U18441 (N_18441,N_16050,N_17221);
nor U18442 (N_18442,N_16777,N_16902);
and U18443 (N_18443,N_17568,N_17475);
xnor U18444 (N_18444,N_16251,N_16668);
and U18445 (N_18445,N_17090,N_16585);
or U18446 (N_18446,N_17092,N_16378);
or U18447 (N_18447,N_16595,N_16701);
nor U18448 (N_18448,N_17380,N_17697);
nand U18449 (N_18449,N_16938,N_17151);
nor U18450 (N_18450,N_16259,N_17392);
nand U18451 (N_18451,N_16324,N_17355);
nand U18452 (N_18452,N_16445,N_16726);
or U18453 (N_18453,N_17734,N_16810);
or U18454 (N_18454,N_17488,N_16687);
or U18455 (N_18455,N_16958,N_16960);
nor U18456 (N_18456,N_17544,N_16768);
or U18457 (N_18457,N_17290,N_16980);
nand U18458 (N_18458,N_16130,N_16396);
nand U18459 (N_18459,N_17422,N_17997);
nand U18460 (N_18460,N_16311,N_17318);
or U18461 (N_18461,N_16645,N_16106);
nand U18462 (N_18462,N_16648,N_17396);
nor U18463 (N_18463,N_17606,N_16849);
or U18464 (N_18464,N_16882,N_16042);
nor U18465 (N_18465,N_17206,N_16723);
or U18466 (N_18466,N_16398,N_16218);
nand U18467 (N_18467,N_17931,N_17426);
or U18468 (N_18468,N_16948,N_17751);
nor U18469 (N_18469,N_17963,N_16703);
or U18470 (N_18470,N_17207,N_17589);
nand U18471 (N_18471,N_17034,N_17900);
and U18472 (N_18472,N_17811,N_17652);
and U18473 (N_18473,N_16949,N_17322);
and U18474 (N_18474,N_16349,N_17200);
nand U18475 (N_18475,N_17007,N_16893);
and U18476 (N_18476,N_17545,N_17114);
and U18477 (N_18477,N_17924,N_17237);
or U18478 (N_18478,N_17170,N_16172);
and U18479 (N_18479,N_17898,N_17801);
or U18480 (N_18480,N_16909,N_16532);
and U18481 (N_18481,N_17249,N_16403);
or U18482 (N_18482,N_17846,N_17465);
nor U18483 (N_18483,N_17302,N_17214);
and U18484 (N_18484,N_16783,N_16379);
nor U18485 (N_18485,N_16222,N_17014);
nor U18486 (N_18486,N_17506,N_17850);
nor U18487 (N_18487,N_17040,N_17676);
nor U18488 (N_18488,N_17729,N_17061);
or U18489 (N_18489,N_16576,N_17121);
nand U18490 (N_18490,N_17946,N_16284);
xor U18491 (N_18491,N_17268,N_16661);
or U18492 (N_18492,N_17323,N_16922);
xnor U18493 (N_18493,N_17298,N_16399);
and U18494 (N_18494,N_16338,N_17517);
and U18495 (N_18495,N_17594,N_17451);
nand U18496 (N_18496,N_17656,N_17564);
nor U18497 (N_18497,N_17728,N_16586);
or U18498 (N_18498,N_17531,N_17562);
or U18499 (N_18499,N_17767,N_16873);
and U18500 (N_18500,N_16037,N_17059);
and U18501 (N_18501,N_17039,N_16682);
or U18502 (N_18502,N_17766,N_17004);
nor U18503 (N_18503,N_17973,N_17110);
or U18504 (N_18504,N_16205,N_17783);
nand U18505 (N_18505,N_17163,N_17541);
nor U18506 (N_18506,N_16570,N_16757);
and U18507 (N_18507,N_17565,N_16738);
and U18508 (N_18508,N_16895,N_17149);
or U18509 (N_18509,N_16929,N_17715);
xnor U18510 (N_18510,N_16482,N_17364);
nor U18511 (N_18511,N_16892,N_17798);
and U18512 (N_18512,N_17983,N_16498);
and U18513 (N_18513,N_16813,N_17717);
or U18514 (N_18514,N_16519,N_17856);
or U18515 (N_18515,N_16613,N_16739);
or U18516 (N_18516,N_16600,N_17723);
or U18517 (N_18517,N_16962,N_16217);
and U18518 (N_18518,N_17070,N_17095);
and U18519 (N_18519,N_17000,N_16659);
or U18520 (N_18520,N_17006,N_16082);
and U18521 (N_18521,N_17342,N_16119);
nor U18522 (N_18522,N_17145,N_16597);
nor U18523 (N_18523,N_17406,N_16900);
or U18524 (N_18524,N_16869,N_16466);
or U18525 (N_18525,N_16728,N_17969);
and U18526 (N_18526,N_16706,N_17964);
nand U18527 (N_18527,N_17405,N_16367);
xnor U18528 (N_18528,N_17284,N_16590);
or U18529 (N_18529,N_17778,N_17042);
and U18530 (N_18530,N_16197,N_16098);
nand U18531 (N_18531,N_16921,N_17052);
and U18532 (N_18532,N_16473,N_17031);
or U18533 (N_18533,N_17701,N_16418);
nor U18534 (N_18534,N_16635,N_16970);
and U18535 (N_18535,N_16767,N_17763);
and U18536 (N_18536,N_16059,N_16506);
nor U18537 (N_18537,N_17428,N_17408);
or U18538 (N_18538,N_17862,N_16907);
nor U18539 (N_18539,N_16866,N_16758);
or U18540 (N_18540,N_16799,N_16402);
or U18541 (N_18541,N_16812,N_17185);
nand U18542 (N_18542,N_16848,N_16083);
nand U18543 (N_18543,N_17464,N_16154);
or U18544 (N_18544,N_17685,N_17188);
and U18545 (N_18545,N_17516,N_17139);
nand U18546 (N_18546,N_17326,N_17799);
and U18547 (N_18547,N_16434,N_16627);
nor U18548 (N_18548,N_16499,N_17888);
nand U18549 (N_18549,N_16474,N_17665);
nor U18550 (N_18550,N_17278,N_17919);
and U18551 (N_18551,N_17310,N_17242);
and U18552 (N_18552,N_17088,N_16829);
nor U18553 (N_18553,N_17067,N_16395);
and U18554 (N_18554,N_17048,N_17537);
nand U18555 (N_18555,N_16886,N_17105);
nand U18556 (N_18556,N_17339,N_16225);
and U18557 (N_18557,N_17738,N_17248);
and U18558 (N_18558,N_17540,N_16464);
and U18559 (N_18559,N_17894,N_16167);
nand U18560 (N_18560,N_16424,N_16112);
xor U18561 (N_18561,N_17867,N_16111);
and U18562 (N_18562,N_16358,N_17138);
and U18563 (N_18563,N_16977,N_16122);
or U18564 (N_18564,N_17960,N_17548);
and U18565 (N_18565,N_16679,N_17699);
nand U18566 (N_18566,N_17157,N_17709);
nor U18567 (N_18567,N_17690,N_17072);
nand U18568 (N_18568,N_16860,N_16614);
and U18569 (N_18569,N_16696,N_16185);
and U18570 (N_18570,N_17780,N_16927);
or U18571 (N_18571,N_17680,N_17758);
and U18572 (N_18572,N_17227,N_17760);
nand U18573 (N_18573,N_16621,N_17937);
nor U18574 (N_18574,N_17234,N_17509);
or U18575 (N_18575,N_17401,N_17107);
and U18576 (N_18576,N_17609,N_16219);
or U18577 (N_18577,N_17938,N_17748);
nand U18578 (N_18578,N_16189,N_17288);
nand U18579 (N_18579,N_16760,N_17499);
nor U18580 (N_18580,N_17727,N_17066);
or U18581 (N_18581,N_16393,N_17640);
and U18582 (N_18582,N_17610,N_17147);
or U18583 (N_18583,N_17216,N_17534);
and U18584 (N_18584,N_17271,N_16326);
xor U18585 (N_18585,N_17542,N_17511);
nor U18586 (N_18586,N_16472,N_17203);
nand U18587 (N_18587,N_17472,N_16872);
and U18588 (N_18588,N_16275,N_16089);
and U18589 (N_18589,N_17294,N_16454);
nor U18590 (N_18590,N_17354,N_16356);
and U18591 (N_18591,N_17684,N_17500);
nand U18592 (N_18592,N_17315,N_16292);
and U18593 (N_18593,N_16763,N_17495);
and U18594 (N_18594,N_17041,N_16087);
xnor U18595 (N_18595,N_17493,N_17714);
nor U18596 (N_18596,N_16032,N_16840);
or U18597 (N_18597,N_16754,N_16406);
nand U18598 (N_18598,N_16408,N_16946);
and U18599 (N_18599,N_16265,N_17646);
and U18600 (N_18600,N_16147,N_17879);
nor U18601 (N_18601,N_17411,N_17081);
nand U18602 (N_18602,N_16028,N_16707);
or U18603 (N_18603,N_16959,N_16610);
nor U18604 (N_18604,N_16553,N_16020);
nand U18605 (N_18605,N_17984,N_17415);
nand U18606 (N_18606,N_17261,N_17772);
nor U18607 (N_18607,N_17078,N_16303);
nand U18608 (N_18608,N_17279,N_17904);
nor U18609 (N_18609,N_17844,N_17605);
nor U18610 (N_18610,N_16901,N_17539);
nand U18611 (N_18611,N_16637,N_16862);
nor U18612 (N_18612,N_17442,N_17334);
nand U18613 (N_18613,N_17109,N_16148);
or U18614 (N_18614,N_17576,N_16580);
nand U18615 (N_18615,N_17675,N_17447);
nand U18616 (N_18616,N_17491,N_16875);
nor U18617 (N_18617,N_16327,N_17245);
nand U18618 (N_18618,N_16692,N_17951);
or U18619 (N_18619,N_17108,N_17841);
xnor U18620 (N_18620,N_17260,N_16822);
nor U18621 (N_18621,N_16557,N_17907);
nor U18622 (N_18622,N_16990,N_16785);
nor U18623 (N_18623,N_16389,N_16262);
nor U18624 (N_18624,N_17764,N_16291);
nor U18625 (N_18625,N_16381,N_17532);
or U18626 (N_18626,N_17948,N_17079);
or U18627 (N_18627,N_16954,N_16245);
nand U18628 (N_18628,N_17570,N_16891);
or U18629 (N_18629,N_16400,N_16449);
nand U18630 (N_18630,N_17998,N_17526);
nor U18631 (N_18631,N_16517,N_16191);
or U18632 (N_18632,N_17664,N_17484);
or U18633 (N_18633,N_17258,N_16539);
nand U18634 (N_18634,N_17547,N_16604);
nand U18635 (N_18635,N_16660,N_17817);
xor U18636 (N_18636,N_16296,N_16309);
or U18637 (N_18637,N_16655,N_16415);
or U18638 (N_18638,N_17976,N_16072);
or U18639 (N_18639,N_17916,N_17769);
nor U18640 (N_18640,N_16450,N_16511);
xor U18641 (N_18641,N_16766,N_17636);
or U18642 (N_18642,N_16471,N_16438);
xnor U18643 (N_18643,N_16807,N_17273);
nand U18644 (N_18644,N_17228,N_17595);
and U18645 (N_18645,N_17912,N_16877);
nand U18646 (N_18646,N_17436,N_16006);
and U18647 (N_18647,N_17202,N_17934);
nor U18648 (N_18648,N_16226,N_17010);
nor U18649 (N_18649,N_16282,N_16669);
and U18650 (N_18650,N_16350,N_16835);
and U18651 (N_18651,N_17880,N_16508);
and U18652 (N_18652,N_16530,N_16003);
nor U18653 (N_18653,N_16470,N_16674);
nor U18654 (N_18654,N_17457,N_16194);
nand U18655 (N_18655,N_17130,N_16746);
nand U18656 (N_18656,N_17443,N_16248);
or U18657 (N_18657,N_16335,N_16724);
nand U18658 (N_18658,N_17373,N_16206);
or U18659 (N_18659,N_17126,N_17068);
nor U18660 (N_18660,N_16289,N_16478);
and U18661 (N_18661,N_17178,N_16250);
or U18662 (N_18662,N_16952,N_16836);
nor U18663 (N_18663,N_16295,N_16945);
nand U18664 (N_18664,N_16552,N_16182);
nor U18665 (N_18665,N_17991,N_16697);
nor U18666 (N_18666,N_17789,N_17569);
or U18667 (N_18667,N_16067,N_17580);
or U18668 (N_18668,N_17482,N_17574);
nor U18669 (N_18669,N_17736,N_16734);
and U18670 (N_18670,N_16091,N_17911);
and U18671 (N_18671,N_17103,N_17585);
and U18672 (N_18672,N_16017,N_16964);
nor U18673 (N_18673,N_16666,N_16993);
and U18674 (N_18674,N_16169,N_17100);
nor U18675 (N_18675,N_16128,N_16270);
and U18676 (N_18676,N_16348,N_16717);
nand U18677 (N_18677,N_17479,N_16744);
or U18678 (N_18678,N_16784,N_16523);
or U18679 (N_18679,N_17653,N_16200);
nor U18680 (N_18680,N_16110,N_17210);
and U18681 (N_18681,N_17803,N_16753);
nand U18682 (N_18682,N_17558,N_16412);
nor U18683 (N_18683,N_17627,N_17755);
nand U18684 (N_18684,N_17686,N_17387);
nor U18685 (N_18685,N_16281,N_16237);
nand U18686 (N_18686,N_17429,N_16588);
xor U18687 (N_18687,N_16390,N_16587);
nor U18688 (N_18688,N_17171,N_16178);
nor U18689 (N_18689,N_17272,N_17001);
nor U18690 (N_18690,N_16861,N_17211);
nand U18691 (N_18691,N_17175,N_16937);
nand U18692 (N_18692,N_17043,N_17784);
nor U18693 (N_18693,N_16879,N_17035);
or U18694 (N_18694,N_17647,N_16525);
and U18695 (N_18695,N_17189,N_17713);
nand U18696 (N_18696,N_17528,N_17629);
nor U18697 (N_18697,N_17630,N_17433);
nor U18698 (N_18698,N_16081,N_17893);
or U18699 (N_18699,N_17523,N_16333);
or U18700 (N_18700,N_16815,N_16336);
xor U18701 (N_18701,N_16341,N_17053);
nor U18702 (N_18702,N_17967,N_16058);
or U18703 (N_18703,N_17332,N_17649);
and U18704 (N_18704,N_17367,N_16155);
or U18705 (N_18705,N_17928,N_16238);
nor U18706 (N_18706,N_16386,N_17091);
and U18707 (N_18707,N_16984,N_17687);
nor U18708 (N_18708,N_17017,N_16843);
or U18709 (N_18709,N_17469,N_16569);
or U18710 (N_18710,N_17859,N_17930);
and U18711 (N_18711,N_16917,N_16780);
nor U18712 (N_18712,N_17213,N_17546);
nand U18713 (N_18713,N_17923,N_16430);
and U18714 (N_18714,N_16487,N_16187);
nand U18715 (N_18715,N_16004,N_16548);
nor U18716 (N_18716,N_16009,N_17525);
nor U18717 (N_18717,N_16976,N_17458);
nand U18718 (N_18718,N_16640,N_16505);
nor U18719 (N_18719,N_17573,N_17263);
or U18720 (N_18720,N_17379,N_16126);
nand U18721 (N_18721,N_16120,N_16652);
xnor U18722 (N_18722,N_16380,N_16173);
or U18723 (N_18723,N_17939,N_17317);
nor U18724 (N_18724,N_16999,N_16443);
nor U18725 (N_18725,N_16550,N_16623);
xor U18726 (N_18726,N_16538,N_16944);
or U18727 (N_18727,N_17257,N_16484);
or U18728 (N_18728,N_16279,N_16192);
or U18729 (N_18729,N_17117,N_17312);
nand U18730 (N_18730,N_17009,N_16596);
or U18731 (N_18731,N_17497,N_17669);
or U18732 (N_18732,N_16834,N_16683);
or U18733 (N_18733,N_17195,N_16317);
nand U18734 (N_18734,N_16581,N_16841);
nor U18735 (N_18735,N_17490,N_17873);
nor U18736 (N_18736,N_17378,N_17987);
nor U18737 (N_18737,N_16142,N_17012);
nor U18738 (N_18738,N_17460,N_16334);
and U18739 (N_18739,N_16298,N_16969);
nor U18740 (N_18740,N_17321,N_17480);
or U18741 (N_18741,N_17063,N_17295);
nand U18742 (N_18742,N_17197,N_16492);
nand U18743 (N_18743,N_17625,N_16000);
nand U18744 (N_18744,N_17243,N_16657);
and U18745 (N_18745,N_16496,N_16070);
nor U18746 (N_18746,N_16956,N_16033);
nor U18747 (N_18747,N_16085,N_17244);
xor U18748 (N_18748,N_16647,N_16665);
nor U18749 (N_18749,N_17813,N_17518);
nand U18750 (N_18750,N_17741,N_16045);
nor U18751 (N_18751,N_16159,N_17372);
xnor U18752 (N_18752,N_16483,N_16216);
or U18753 (N_18753,N_17129,N_16646);
and U18754 (N_18754,N_17671,N_17949);
nor U18755 (N_18755,N_17638,N_16620);
nand U18756 (N_18756,N_17275,N_16920);
or U18757 (N_18757,N_16177,N_17262);
or U18758 (N_18758,N_16782,N_16583);
and U18759 (N_18759,N_17619,N_16781);
and U18760 (N_18760,N_17648,N_17753);
nand U18761 (N_18761,N_16451,N_17854);
and U18762 (N_18762,N_16702,N_17013);
nand U18763 (N_18763,N_17897,N_17341);
or U18764 (N_18764,N_17122,N_17563);
nor U18765 (N_18765,N_16409,N_17533);
nand U18766 (N_18766,N_17821,N_17309);
nand U18767 (N_18767,N_17617,N_16136);
nor U18768 (N_18768,N_16211,N_17858);
nor U18769 (N_18769,N_17583,N_17424);
nor U18770 (N_18770,N_17176,N_16361);
and U18771 (N_18771,N_16974,N_17165);
nand U18772 (N_18772,N_16535,N_17747);
nor U18773 (N_18773,N_17746,N_17941);
or U18774 (N_18774,N_16322,N_16288);
nor U18775 (N_18775,N_17902,N_16619);
nand U18776 (N_18776,N_17834,N_17153);
xor U18777 (N_18777,N_17883,N_17851);
xor U18778 (N_18778,N_16432,N_17787);
nand U18779 (N_18779,N_16598,N_16157);
nand U18780 (N_18780,N_17670,N_17328);
nand U18781 (N_18781,N_17320,N_17708);
nand U18782 (N_18782,N_17146,N_16099);
or U18783 (N_18783,N_16315,N_17822);
and U18784 (N_18784,N_17382,N_16049);
xor U18785 (N_18785,N_17502,N_17196);
nand U18786 (N_18786,N_16436,N_16041);
nor U18787 (N_18787,N_17618,N_16131);
nand U18788 (N_18788,N_16612,N_16574);
nor U18789 (N_18789,N_16469,N_17158);
or U18790 (N_18790,N_17981,N_16293);
or U18791 (N_18791,N_17892,N_16868);
nand U18792 (N_18792,N_17340,N_16353);
nor U18793 (N_18793,N_16359,N_16420);
and U18794 (N_18794,N_16213,N_17369);
or U18795 (N_18795,N_17055,N_17702);
nor U18796 (N_18796,N_16551,N_16820);
nand U18797 (N_18797,N_17718,N_17420);
nor U18798 (N_18798,N_17505,N_17033);
or U18799 (N_18799,N_17073,N_16404);
or U18800 (N_18800,N_17496,N_17874);
nand U18801 (N_18801,N_17527,N_16897);
nor U18802 (N_18802,N_16695,N_16475);
nor U18803 (N_18803,N_16234,N_17270);
nand U18804 (N_18804,N_17961,N_16444);
and U18805 (N_18805,N_17229,N_17409);
and U18806 (N_18806,N_17812,N_16899);
nor U18807 (N_18807,N_17127,N_16715);
nand U18808 (N_18808,N_16268,N_17445);
nor U18809 (N_18809,N_16005,N_16967);
or U18810 (N_18810,N_16689,N_17586);
nor U18811 (N_18811,N_17468,N_17810);
or U18812 (N_18812,N_16911,N_17674);
xnor U18813 (N_18813,N_17691,N_16053);
or U18814 (N_18814,N_17833,N_16278);
or U18815 (N_18815,N_16555,N_17550);
nor U18816 (N_18816,N_17913,N_16441);
and U18817 (N_18817,N_17857,N_16179);
nand U18818 (N_18818,N_17388,N_16104);
nand U18819 (N_18819,N_16077,N_17797);
and U18820 (N_18820,N_17473,N_16340);
nand U18821 (N_18821,N_16876,N_17435);
and U18822 (N_18822,N_17808,N_17555);
and U18823 (N_18823,N_16231,N_16851);
nand U18824 (N_18824,N_16242,N_16864);
nor U18825 (N_18825,N_16465,N_16681);
nor U18826 (N_18826,N_16542,N_17476);
and U18827 (N_18827,N_16816,N_16950);
nor U18828 (N_18828,N_17970,N_16742);
xor U18829 (N_18829,N_16670,N_16791);
and U18830 (N_18830,N_16940,N_17815);
or U18831 (N_18831,N_16685,N_17093);
or U18832 (N_18832,N_16310,N_17752);
or U18833 (N_18833,N_17677,N_17330);
nor U18834 (N_18834,N_16624,N_16168);
nand U18835 (N_18835,N_17438,N_17099);
and U18836 (N_18836,N_16302,N_16644);
nand U18837 (N_18837,N_17503,N_17695);
nand U18838 (N_18838,N_16435,N_17331);
or U18839 (N_18839,N_17194,N_16132);
or U18840 (N_18840,N_17291,N_16594);
nand U18841 (N_18841,N_17134,N_16987);
nor U18842 (N_18842,N_16821,N_16442);
nor U18843 (N_18843,N_16212,N_16773);
nor U18844 (N_18844,N_17519,N_17577);
nand U18845 (N_18845,N_16713,N_17101);
xnor U18846 (N_18846,N_16994,N_17824);
and U18847 (N_18847,N_16787,N_17567);
nor U18848 (N_18848,N_16522,N_16031);
xnor U18849 (N_18849,N_17626,N_17538);
and U18850 (N_18850,N_17992,N_17137);
nand U18851 (N_18851,N_16489,N_16337);
and U18852 (N_18852,N_16040,N_16616);
and U18853 (N_18853,N_16043,N_17299);
nand U18854 (N_18854,N_17047,N_17015);
and U18855 (N_18855,N_16181,N_17915);
and U18856 (N_18856,N_17908,N_17297);
or U18857 (N_18857,N_16887,N_16374);
or U18858 (N_18858,N_17021,N_16488);
and U18859 (N_18859,N_16057,N_17256);
nor U18860 (N_18860,N_16025,N_16885);
or U18861 (N_18861,N_17903,N_17391);
nand U18862 (N_18862,N_16113,N_16608);
or U18863 (N_18863,N_16847,N_17255);
or U18864 (N_18864,N_17418,N_16811);
or U18865 (N_18865,N_16052,N_16260);
nor U18866 (N_18866,N_16458,N_17399);
or U18867 (N_18867,N_16421,N_17513);
or U18868 (N_18868,N_16859,N_16930);
nand U18869 (N_18869,N_16074,N_17847);
and U18870 (N_18870,N_16133,N_17615);
nor U18871 (N_18871,N_17183,N_16339);
and U18872 (N_18872,N_17156,N_16698);
and U18873 (N_18873,N_16101,N_16607);
nand U18874 (N_18874,N_17835,N_16642);
and U18875 (N_18875,N_16440,N_17943);
or U18876 (N_18876,N_16794,N_16916);
nor U18877 (N_18877,N_17030,N_17683);
nor U18878 (N_18878,N_16170,N_17254);
or U18879 (N_18879,N_16026,N_17439);
nor U18880 (N_18880,N_16063,N_17208);
or U18881 (N_18881,N_16756,N_16923);
nor U18882 (N_18882,N_17603,N_17140);
nor U18883 (N_18883,N_16316,N_16299);
or U18884 (N_18884,N_16274,N_17352);
and U18885 (N_18885,N_16662,N_17086);
or U18886 (N_18886,N_17990,N_16573);
nand U18887 (N_18887,N_17592,N_17360);
or U18888 (N_18888,N_16549,N_17224);
nand U18889 (N_18889,N_16048,N_16388);
nand U18890 (N_18890,N_17253,N_16775);
nand U18891 (N_18891,N_17371,N_16865);
and U18892 (N_18892,N_17793,N_16863);
nand U18893 (N_18893,N_16625,N_17314);
and U18894 (N_18894,N_16838,N_16833);
and U18895 (N_18895,N_16366,N_16411);
nor U18896 (N_18896,N_16601,N_16502);
and U18897 (N_18897,N_17522,N_16817);
and U18898 (N_18898,N_16467,N_16797);
and U18899 (N_18899,N_17575,N_16160);
and U18900 (N_18900,N_16814,N_16839);
nor U18901 (N_18901,N_16748,N_16476);
and U18902 (N_18902,N_17494,N_16761);
nor U18903 (N_18903,N_17293,N_16139);
and U18904 (N_18904,N_17872,N_17910);
nand U18905 (N_18905,N_16229,N_16529);
or U18906 (N_18906,N_17343,N_16571);
nor U18907 (N_18907,N_17182,N_16933);
or U18908 (N_18908,N_17557,N_17554);
and U18909 (N_18909,N_16677,N_16129);
or U18910 (N_18910,N_16983,N_16394);
or U18911 (N_18911,N_16180,N_16636);
nor U18912 (N_18912,N_16080,N_17825);
and U18913 (N_18913,N_16765,N_16124);
nand U18914 (N_18914,N_16044,N_17703);
or U18915 (N_18915,N_17559,N_16957);
or U18916 (N_18916,N_17933,N_16377);
or U18917 (N_18917,N_16423,N_16490);
nand U18918 (N_18918,N_17887,N_17560);
xnor U18919 (N_18919,N_17240,N_16138);
or U18920 (N_18920,N_16547,N_16233);
or U18921 (N_18921,N_16638,N_16881);
nand U18922 (N_18922,N_16437,N_17199);
nor U18923 (N_18923,N_16429,N_16577);
or U18924 (N_18924,N_16842,N_16462);
xnor U18925 (N_18925,N_17694,N_16667);
nand U18926 (N_18926,N_17660,N_16617);
and U18927 (N_18927,N_16904,N_16915);
nand U18928 (N_18928,N_16704,N_17173);
and U18929 (N_18929,N_16874,N_17994);
and U18930 (N_18930,N_17621,N_17909);
or U18931 (N_18931,N_17410,N_17591);
nand U18932 (N_18932,N_16606,N_17588);
nor U18933 (N_18933,N_17347,N_17168);
nor U18934 (N_18934,N_17361,N_16183);
and U18935 (N_18935,N_17614,N_16312);
and U18936 (N_18936,N_17220,N_16809);
nand U18937 (N_18937,N_16426,N_16656);
nor U18938 (N_18938,N_16151,N_17935);
nand U18939 (N_18939,N_17209,N_17212);
nor U18940 (N_18940,N_17128,N_17375);
nor U18941 (N_18941,N_16943,N_16831);
nor U18942 (N_18942,N_17871,N_17308);
and U18943 (N_18943,N_17384,N_17688);
nand U18944 (N_18944,N_17333,N_17530);
nor U18945 (N_18945,N_16097,N_17431);
or U18946 (N_18946,N_16725,N_16024);
or U18947 (N_18947,N_17027,N_17060);
nor U18948 (N_18948,N_17739,N_16382);
nor U18949 (N_18949,N_16243,N_16910);
or U18950 (N_18950,N_16805,N_16376);
nor U18951 (N_18951,N_16828,N_16076);
nor U18952 (N_18952,N_16273,N_17050);
and U18953 (N_18953,N_17296,N_17578);
nand U18954 (N_18954,N_17866,N_16740);
xnor U18955 (N_18955,N_16373,N_17510);
nand U18956 (N_18956,N_16258,N_17487);
and U18957 (N_18957,N_17230,N_17807);
or U18958 (N_18958,N_17282,N_17977);
nand U18959 (N_18959,N_17402,N_16247);
nand U18960 (N_18960,N_16370,N_16735);
nor U18961 (N_18961,N_17965,N_16001);
or U18962 (N_18962,N_17679,N_16536);
nor U18963 (N_18963,N_17056,N_17642);
nor U18964 (N_18964,N_16853,N_17036);
nor U18965 (N_18965,N_16663,N_17645);
and U18966 (N_18966,N_16149,N_17231);
nor U18967 (N_18967,N_17191,N_16826);
xor U18968 (N_18968,N_17335,N_16527);
nor U18969 (N_18969,N_17119,N_17305);
or U18970 (N_18970,N_17842,N_17611);
nand U18971 (N_18971,N_17980,N_16144);
nor U18972 (N_18972,N_17466,N_17080);
nand U18973 (N_18973,N_17266,N_17241);
nor U18974 (N_18974,N_16593,N_17597);
and U18975 (N_18975,N_16591,N_16497);
and U18976 (N_18976,N_16346,N_17958);
nor U18977 (N_18977,N_16690,N_16305);
nand U18978 (N_18978,N_17336,N_16818);
and U18979 (N_18979,N_16997,N_17247);
nor U18980 (N_18980,N_16545,N_16850);
or U18981 (N_18981,N_17198,N_16749);
and U18982 (N_18982,N_17507,N_17536);
nor U18983 (N_18983,N_17003,N_17836);
nor U18984 (N_18984,N_16241,N_17832);
nor U18985 (N_18985,N_17587,N_16362);
nand U18986 (N_18986,N_17349,N_17792);
nor U18987 (N_18987,N_17678,N_17051);
or U18988 (N_18988,N_16936,N_16932);
nor U18989 (N_18989,N_16330,N_16414);
or U18990 (N_18990,N_16413,N_17389);
nor U18991 (N_18991,N_16507,N_17666);
nand U18992 (N_18992,N_17046,N_16297);
and U18993 (N_18993,N_16255,N_16544);
nand U18994 (N_18994,N_16064,N_16605);
or U18995 (N_18995,N_17865,N_17622);
or U18996 (N_18996,N_16494,N_16680);
nor U18997 (N_18997,N_16925,N_16844);
nand U18998 (N_18998,N_17819,N_16417);
nand U18999 (N_18999,N_17289,N_16649);
nand U19000 (N_19000,N_17592,N_16131);
nor U19001 (N_19001,N_17874,N_16210);
or U19002 (N_19002,N_17401,N_17399);
xor U19003 (N_19003,N_16941,N_16277);
nor U19004 (N_19004,N_16653,N_17876);
and U19005 (N_19005,N_17622,N_16396);
and U19006 (N_19006,N_16077,N_16421);
nor U19007 (N_19007,N_17271,N_16600);
and U19008 (N_19008,N_17864,N_16250);
and U19009 (N_19009,N_16335,N_17595);
nand U19010 (N_19010,N_16237,N_17469);
nand U19011 (N_19011,N_17608,N_16068);
and U19012 (N_19012,N_16472,N_16517);
nor U19013 (N_19013,N_17357,N_17760);
or U19014 (N_19014,N_16528,N_16347);
or U19015 (N_19015,N_17578,N_17935);
or U19016 (N_19016,N_17601,N_17239);
nor U19017 (N_19017,N_17198,N_17543);
nand U19018 (N_19018,N_17917,N_17895);
nor U19019 (N_19019,N_17369,N_16621);
xnor U19020 (N_19020,N_16551,N_16204);
and U19021 (N_19021,N_17884,N_17448);
and U19022 (N_19022,N_17423,N_17595);
and U19023 (N_19023,N_16136,N_16897);
and U19024 (N_19024,N_16212,N_16975);
nand U19025 (N_19025,N_16696,N_16698);
nor U19026 (N_19026,N_16425,N_16277);
nor U19027 (N_19027,N_17870,N_17917);
nand U19028 (N_19028,N_16401,N_17330);
or U19029 (N_19029,N_16256,N_16429);
nand U19030 (N_19030,N_17994,N_16802);
nand U19031 (N_19031,N_16053,N_16524);
and U19032 (N_19032,N_16482,N_17396);
and U19033 (N_19033,N_17705,N_17873);
nand U19034 (N_19034,N_16038,N_17086);
or U19035 (N_19035,N_16212,N_17862);
nor U19036 (N_19036,N_17857,N_16828);
or U19037 (N_19037,N_16830,N_17467);
xnor U19038 (N_19038,N_16846,N_17926);
and U19039 (N_19039,N_16720,N_17899);
xor U19040 (N_19040,N_16215,N_16798);
nor U19041 (N_19041,N_16105,N_17549);
and U19042 (N_19042,N_16454,N_16558);
or U19043 (N_19043,N_16972,N_16621);
nand U19044 (N_19044,N_17542,N_16773);
nor U19045 (N_19045,N_16750,N_16538);
nand U19046 (N_19046,N_17650,N_16135);
and U19047 (N_19047,N_16610,N_16186);
and U19048 (N_19048,N_17155,N_17320);
nand U19049 (N_19049,N_16433,N_17013);
nand U19050 (N_19050,N_16906,N_16310);
nand U19051 (N_19051,N_16976,N_17264);
nor U19052 (N_19052,N_17998,N_17406);
nand U19053 (N_19053,N_16812,N_17871);
or U19054 (N_19054,N_17839,N_17494);
nand U19055 (N_19055,N_17233,N_16265);
or U19056 (N_19056,N_17719,N_17882);
or U19057 (N_19057,N_16729,N_17485);
nor U19058 (N_19058,N_17276,N_16485);
nand U19059 (N_19059,N_17998,N_17784);
or U19060 (N_19060,N_16358,N_17558);
or U19061 (N_19061,N_16901,N_16535);
nand U19062 (N_19062,N_17446,N_17032);
nor U19063 (N_19063,N_17433,N_16828);
and U19064 (N_19064,N_16024,N_16171);
nand U19065 (N_19065,N_17897,N_16444);
or U19066 (N_19066,N_16002,N_17710);
nor U19067 (N_19067,N_17095,N_16745);
and U19068 (N_19068,N_17575,N_17622);
or U19069 (N_19069,N_17143,N_16057);
nor U19070 (N_19070,N_17196,N_16778);
nor U19071 (N_19071,N_17964,N_16171);
nor U19072 (N_19072,N_16070,N_17568);
and U19073 (N_19073,N_16766,N_17446);
or U19074 (N_19074,N_17191,N_16205);
nand U19075 (N_19075,N_17195,N_17093);
nand U19076 (N_19076,N_16656,N_17561);
and U19077 (N_19077,N_16869,N_16548);
nand U19078 (N_19078,N_16813,N_16612);
nor U19079 (N_19079,N_16188,N_17822);
or U19080 (N_19080,N_16773,N_16942);
or U19081 (N_19081,N_16130,N_16051);
nor U19082 (N_19082,N_17359,N_16132);
or U19083 (N_19083,N_17990,N_16129);
nor U19084 (N_19084,N_16468,N_16770);
and U19085 (N_19085,N_16242,N_17335);
or U19086 (N_19086,N_16929,N_16482);
nand U19087 (N_19087,N_17525,N_17993);
or U19088 (N_19088,N_17914,N_16616);
nor U19089 (N_19089,N_16769,N_17472);
nand U19090 (N_19090,N_16818,N_17250);
xor U19091 (N_19091,N_17677,N_16867);
and U19092 (N_19092,N_17077,N_16113);
nor U19093 (N_19093,N_16762,N_16230);
or U19094 (N_19094,N_17418,N_17962);
nand U19095 (N_19095,N_17693,N_16109);
nor U19096 (N_19096,N_16348,N_17451);
or U19097 (N_19097,N_16224,N_17106);
and U19098 (N_19098,N_16639,N_17691);
nand U19099 (N_19099,N_17681,N_16331);
and U19100 (N_19100,N_16444,N_17274);
nor U19101 (N_19101,N_17803,N_16436);
nand U19102 (N_19102,N_17617,N_17742);
nor U19103 (N_19103,N_17337,N_16255);
nor U19104 (N_19104,N_16597,N_16098);
or U19105 (N_19105,N_17489,N_16414);
and U19106 (N_19106,N_16587,N_17608);
nor U19107 (N_19107,N_17353,N_17035);
nor U19108 (N_19108,N_17562,N_17327);
or U19109 (N_19109,N_16831,N_16095);
nor U19110 (N_19110,N_16434,N_16125);
nor U19111 (N_19111,N_17896,N_16744);
or U19112 (N_19112,N_16117,N_17237);
nor U19113 (N_19113,N_17429,N_16035);
nor U19114 (N_19114,N_16871,N_16412);
or U19115 (N_19115,N_17744,N_16301);
or U19116 (N_19116,N_17758,N_17335);
nor U19117 (N_19117,N_16729,N_17804);
and U19118 (N_19118,N_17487,N_16988);
or U19119 (N_19119,N_16103,N_17355);
or U19120 (N_19120,N_17942,N_17978);
nor U19121 (N_19121,N_17144,N_17356);
xnor U19122 (N_19122,N_17324,N_17168);
or U19123 (N_19123,N_16485,N_16652);
or U19124 (N_19124,N_16437,N_17985);
nand U19125 (N_19125,N_17395,N_17541);
nand U19126 (N_19126,N_17772,N_16742);
nor U19127 (N_19127,N_17899,N_16612);
nand U19128 (N_19128,N_16883,N_17146);
nor U19129 (N_19129,N_16028,N_16638);
and U19130 (N_19130,N_16583,N_16509);
nor U19131 (N_19131,N_16225,N_16941);
and U19132 (N_19132,N_16574,N_16491);
nor U19133 (N_19133,N_17863,N_16372);
nor U19134 (N_19134,N_16202,N_17438);
nand U19135 (N_19135,N_17379,N_17508);
nor U19136 (N_19136,N_16722,N_16505);
nand U19137 (N_19137,N_17619,N_17869);
nor U19138 (N_19138,N_17780,N_17525);
and U19139 (N_19139,N_17066,N_17855);
nand U19140 (N_19140,N_16356,N_16179);
and U19141 (N_19141,N_17425,N_17367);
or U19142 (N_19142,N_17017,N_16205);
nor U19143 (N_19143,N_17954,N_16582);
or U19144 (N_19144,N_16853,N_16322);
xnor U19145 (N_19145,N_17837,N_16682);
nand U19146 (N_19146,N_16805,N_16773);
nand U19147 (N_19147,N_16072,N_17797);
nand U19148 (N_19148,N_17893,N_16906);
and U19149 (N_19149,N_17367,N_16106);
and U19150 (N_19150,N_16462,N_17092);
or U19151 (N_19151,N_17090,N_17261);
nor U19152 (N_19152,N_16582,N_16399);
nor U19153 (N_19153,N_17119,N_17001);
nor U19154 (N_19154,N_16119,N_17982);
or U19155 (N_19155,N_16173,N_17448);
or U19156 (N_19156,N_16334,N_16231);
or U19157 (N_19157,N_16127,N_17144);
and U19158 (N_19158,N_16258,N_16067);
nor U19159 (N_19159,N_16642,N_17229);
and U19160 (N_19160,N_16264,N_16010);
xor U19161 (N_19161,N_16845,N_16191);
xor U19162 (N_19162,N_16919,N_17017);
and U19163 (N_19163,N_16018,N_16674);
and U19164 (N_19164,N_17756,N_16458);
or U19165 (N_19165,N_16782,N_16067);
nor U19166 (N_19166,N_16701,N_16444);
or U19167 (N_19167,N_16632,N_17626);
or U19168 (N_19168,N_16017,N_16864);
nor U19169 (N_19169,N_16662,N_16369);
and U19170 (N_19170,N_16905,N_17526);
nand U19171 (N_19171,N_16294,N_16405);
or U19172 (N_19172,N_16188,N_17083);
or U19173 (N_19173,N_16955,N_16125);
or U19174 (N_19174,N_16353,N_17688);
or U19175 (N_19175,N_16302,N_16087);
and U19176 (N_19176,N_16710,N_17835);
or U19177 (N_19177,N_17329,N_16221);
or U19178 (N_19178,N_16862,N_17449);
nand U19179 (N_19179,N_17184,N_16373);
or U19180 (N_19180,N_17882,N_16165);
nor U19181 (N_19181,N_17950,N_17204);
xor U19182 (N_19182,N_17954,N_17190);
nand U19183 (N_19183,N_16221,N_17973);
and U19184 (N_19184,N_16663,N_17396);
and U19185 (N_19185,N_16308,N_16327);
nand U19186 (N_19186,N_16914,N_16606);
or U19187 (N_19187,N_16987,N_17058);
and U19188 (N_19188,N_17543,N_16016);
and U19189 (N_19189,N_16104,N_17005);
or U19190 (N_19190,N_16064,N_16320);
nand U19191 (N_19191,N_17749,N_16075);
nor U19192 (N_19192,N_16682,N_17881);
nand U19193 (N_19193,N_16301,N_17340);
and U19194 (N_19194,N_16178,N_17272);
nand U19195 (N_19195,N_17376,N_16278);
and U19196 (N_19196,N_16161,N_17198);
nor U19197 (N_19197,N_17670,N_17816);
and U19198 (N_19198,N_16033,N_16423);
xnor U19199 (N_19199,N_16225,N_16042);
nor U19200 (N_19200,N_17126,N_17880);
nor U19201 (N_19201,N_16023,N_17700);
nand U19202 (N_19202,N_16015,N_16170);
nor U19203 (N_19203,N_16475,N_16409);
and U19204 (N_19204,N_17658,N_16040);
or U19205 (N_19205,N_17424,N_16409);
xor U19206 (N_19206,N_16507,N_17092);
nor U19207 (N_19207,N_16038,N_17061);
and U19208 (N_19208,N_17216,N_17300);
and U19209 (N_19209,N_16265,N_16413);
nand U19210 (N_19210,N_16937,N_16522);
and U19211 (N_19211,N_17810,N_16457);
or U19212 (N_19212,N_17138,N_16566);
nand U19213 (N_19213,N_16382,N_16756);
and U19214 (N_19214,N_17524,N_16755);
or U19215 (N_19215,N_16441,N_16728);
or U19216 (N_19216,N_16378,N_16797);
and U19217 (N_19217,N_16196,N_16309);
and U19218 (N_19218,N_16783,N_16073);
and U19219 (N_19219,N_16238,N_17010);
nand U19220 (N_19220,N_17548,N_16844);
nor U19221 (N_19221,N_16341,N_16318);
nor U19222 (N_19222,N_17392,N_17264);
and U19223 (N_19223,N_17923,N_16096);
and U19224 (N_19224,N_17768,N_17642);
nor U19225 (N_19225,N_17699,N_17139);
nor U19226 (N_19226,N_17748,N_17023);
and U19227 (N_19227,N_17148,N_16868);
or U19228 (N_19228,N_17467,N_16579);
xor U19229 (N_19229,N_16227,N_16546);
and U19230 (N_19230,N_17916,N_17444);
or U19231 (N_19231,N_16059,N_17714);
or U19232 (N_19232,N_17292,N_16985);
xnor U19233 (N_19233,N_17903,N_16958);
and U19234 (N_19234,N_17810,N_16577);
nand U19235 (N_19235,N_16737,N_16224);
nand U19236 (N_19236,N_16923,N_17632);
and U19237 (N_19237,N_16986,N_16648);
nand U19238 (N_19238,N_17559,N_16007);
nand U19239 (N_19239,N_16951,N_16959);
or U19240 (N_19240,N_17593,N_17741);
nand U19241 (N_19241,N_16766,N_17445);
nor U19242 (N_19242,N_16562,N_17935);
and U19243 (N_19243,N_17739,N_17220);
nor U19244 (N_19244,N_17201,N_16468);
and U19245 (N_19245,N_16651,N_17794);
or U19246 (N_19246,N_17873,N_17001);
nor U19247 (N_19247,N_17749,N_16523);
nor U19248 (N_19248,N_16819,N_16021);
nor U19249 (N_19249,N_17913,N_16895);
and U19250 (N_19250,N_16995,N_17724);
or U19251 (N_19251,N_17446,N_17989);
and U19252 (N_19252,N_16918,N_17662);
nor U19253 (N_19253,N_16063,N_16657);
nor U19254 (N_19254,N_17392,N_17810);
nand U19255 (N_19255,N_16404,N_17593);
or U19256 (N_19256,N_16306,N_17838);
nand U19257 (N_19257,N_17645,N_16645);
or U19258 (N_19258,N_16228,N_16103);
nand U19259 (N_19259,N_17048,N_16241);
and U19260 (N_19260,N_17425,N_16588);
and U19261 (N_19261,N_16562,N_16459);
nor U19262 (N_19262,N_17231,N_16879);
nand U19263 (N_19263,N_16428,N_16983);
and U19264 (N_19264,N_17539,N_16707);
or U19265 (N_19265,N_17602,N_16909);
or U19266 (N_19266,N_16479,N_17605);
nor U19267 (N_19267,N_17764,N_17928);
or U19268 (N_19268,N_16030,N_16117);
nor U19269 (N_19269,N_17049,N_16367);
nand U19270 (N_19270,N_16139,N_16219);
or U19271 (N_19271,N_16804,N_16661);
or U19272 (N_19272,N_16149,N_16922);
nand U19273 (N_19273,N_17558,N_16469);
nor U19274 (N_19274,N_16896,N_17300);
nor U19275 (N_19275,N_16436,N_16312);
nand U19276 (N_19276,N_17070,N_17158);
and U19277 (N_19277,N_17072,N_17316);
nor U19278 (N_19278,N_17437,N_17532);
and U19279 (N_19279,N_16134,N_17617);
and U19280 (N_19280,N_17770,N_16647);
nand U19281 (N_19281,N_16769,N_16002);
nand U19282 (N_19282,N_17394,N_16420);
xor U19283 (N_19283,N_17396,N_17807);
nand U19284 (N_19284,N_16891,N_17354);
and U19285 (N_19285,N_17768,N_16608);
or U19286 (N_19286,N_16375,N_17842);
nor U19287 (N_19287,N_16084,N_17359);
and U19288 (N_19288,N_17012,N_17222);
nand U19289 (N_19289,N_16389,N_17091);
nand U19290 (N_19290,N_16538,N_17143);
nor U19291 (N_19291,N_16078,N_17194);
or U19292 (N_19292,N_16307,N_17750);
and U19293 (N_19293,N_17677,N_17196);
and U19294 (N_19294,N_16743,N_16046);
nand U19295 (N_19295,N_17866,N_16973);
nor U19296 (N_19296,N_17847,N_17992);
nand U19297 (N_19297,N_17015,N_17981);
and U19298 (N_19298,N_17283,N_17833);
and U19299 (N_19299,N_16197,N_17396);
nand U19300 (N_19300,N_16831,N_16726);
or U19301 (N_19301,N_16070,N_17497);
nand U19302 (N_19302,N_17567,N_16237);
and U19303 (N_19303,N_17020,N_17661);
nor U19304 (N_19304,N_16343,N_16865);
nor U19305 (N_19305,N_17777,N_16678);
or U19306 (N_19306,N_17613,N_16312);
nand U19307 (N_19307,N_16879,N_16435);
and U19308 (N_19308,N_16622,N_16747);
and U19309 (N_19309,N_16637,N_16595);
xor U19310 (N_19310,N_16444,N_17921);
or U19311 (N_19311,N_16445,N_17952);
xor U19312 (N_19312,N_16052,N_16627);
nor U19313 (N_19313,N_16756,N_17810);
nor U19314 (N_19314,N_16346,N_17295);
nand U19315 (N_19315,N_17935,N_16757);
or U19316 (N_19316,N_16683,N_17922);
and U19317 (N_19317,N_17401,N_17064);
nand U19318 (N_19318,N_17714,N_17810);
and U19319 (N_19319,N_16626,N_17728);
or U19320 (N_19320,N_17608,N_17203);
or U19321 (N_19321,N_16928,N_17176);
or U19322 (N_19322,N_17920,N_17648);
and U19323 (N_19323,N_16805,N_17172);
and U19324 (N_19324,N_17802,N_16510);
nor U19325 (N_19325,N_17603,N_17730);
nand U19326 (N_19326,N_17978,N_17354);
or U19327 (N_19327,N_16457,N_16417);
nand U19328 (N_19328,N_17638,N_16025);
nand U19329 (N_19329,N_17283,N_17503);
nand U19330 (N_19330,N_16569,N_17938);
or U19331 (N_19331,N_16108,N_17946);
nor U19332 (N_19332,N_17265,N_17358);
nand U19333 (N_19333,N_16697,N_17209);
nand U19334 (N_19334,N_17713,N_17136);
or U19335 (N_19335,N_17359,N_17375);
and U19336 (N_19336,N_17253,N_17966);
nor U19337 (N_19337,N_17853,N_17318);
nor U19338 (N_19338,N_16256,N_16258);
or U19339 (N_19339,N_16542,N_17691);
or U19340 (N_19340,N_16396,N_17858);
nand U19341 (N_19341,N_16889,N_16920);
nor U19342 (N_19342,N_17649,N_17253);
or U19343 (N_19343,N_17599,N_16402);
or U19344 (N_19344,N_16101,N_16601);
nand U19345 (N_19345,N_17845,N_17480);
nor U19346 (N_19346,N_17710,N_17401);
nor U19347 (N_19347,N_16791,N_17975);
or U19348 (N_19348,N_16172,N_17477);
nor U19349 (N_19349,N_17490,N_17790);
and U19350 (N_19350,N_16612,N_17784);
nor U19351 (N_19351,N_17604,N_17565);
nor U19352 (N_19352,N_16022,N_16013);
and U19353 (N_19353,N_16977,N_17119);
or U19354 (N_19354,N_16774,N_16751);
nand U19355 (N_19355,N_17508,N_17446);
nor U19356 (N_19356,N_17921,N_16513);
and U19357 (N_19357,N_16727,N_16191);
nand U19358 (N_19358,N_16701,N_17279);
or U19359 (N_19359,N_17439,N_16340);
and U19360 (N_19360,N_17015,N_16459);
or U19361 (N_19361,N_17760,N_16450);
nor U19362 (N_19362,N_16936,N_17897);
nor U19363 (N_19363,N_17105,N_16558);
or U19364 (N_19364,N_17020,N_16517);
nand U19365 (N_19365,N_17213,N_17349);
nand U19366 (N_19366,N_16702,N_17196);
or U19367 (N_19367,N_17827,N_17221);
nand U19368 (N_19368,N_17680,N_17906);
or U19369 (N_19369,N_16597,N_17108);
or U19370 (N_19370,N_16087,N_17329);
and U19371 (N_19371,N_17051,N_17184);
and U19372 (N_19372,N_17471,N_17713);
and U19373 (N_19373,N_17687,N_17078);
or U19374 (N_19374,N_16120,N_16012);
and U19375 (N_19375,N_16578,N_16631);
nor U19376 (N_19376,N_16869,N_16459);
or U19377 (N_19377,N_16298,N_16400);
nor U19378 (N_19378,N_16221,N_16857);
and U19379 (N_19379,N_17521,N_16984);
nand U19380 (N_19380,N_16906,N_16626);
or U19381 (N_19381,N_16508,N_17094);
nor U19382 (N_19382,N_16032,N_17932);
nand U19383 (N_19383,N_16804,N_16173);
nor U19384 (N_19384,N_16702,N_16112);
nand U19385 (N_19385,N_17369,N_17837);
and U19386 (N_19386,N_17370,N_17567);
nand U19387 (N_19387,N_16897,N_16661);
nor U19388 (N_19388,N_17587,N_17144);
or U19389 (N_19389,N_16606,N_17218);
nor U19390 (N_19390,N_16829,N_16975);
nand U19391 (N_19391,N_16214,N_16491);
or U19392 (N_19392,N_17212,N_17901);
and U19393 (N_19393,N_16646,N_16960);
and U19394 (N_19394,N_16818,N_16535);
or U19395 (N_19395,N_17242,N_17206);
xor U19396 (N_19396,N_16552,N_16339);
nor U19397 (N_19397,N_16829,N_17355);
nor U19398 (N_19398,N_17171,N_16494);
or U19399 (N_19399,N_17640,N_17463);
or U19400 (N_19400,N_17277,N_17561);
or U19401 (N_19401,N_16267,N_16925);
and U19402 (N_19402,N_17916,N_17248);
or U19403 (N_19403,N_17963,N_16042);
and U19404 (N_19404,N_16081,N_17765);
and U19405 (N_19405,N_17015,N_17754);
nand U19406 (N_19406,N_17703,N_16835);
nand U19407 (N_19407,N_17501,N_16417);
nor U19408 (N_19408,N_17700,N_16071);
and U19409 (N_19409,N_16233,N_17366);
nand U19410 (N_19410,N_17646,N_16577);
and U19411 (N_19411,N_17047,N_16062);
nand U19412 (N_19412,N_17225,N_16943);
nor U19413 (N_19413,N_17636,N_16297);
nand U19414 (N_19414,N_16168,N_17934);
or U19415 (N_19415,N_16835,N_17465);
nor U19416 (N_19416,N_17047,N_16105);
and U19417 (N_19417,N_17933,N_17135);
nor U19418 (N_19418,N_16954,N_17539);
and U19419 (N_19419,N_17517,N_16361);
nand U19420 (N_19420,N_16424,N_16936);
nand U19421 (N_19421,N_17867,N_16073);
or U19422 (N_19422,N_16767,N_16173);
xnor U19423 (N_19423,N_17606,N_17992);
nand U19424 (N_19424,N_17791,N_16793);
or U19425 (N_19425,N_16315,N_17155);
or U19426 (N_19426,N_17510,N_16656);
and U19427 (N_19427,N_16439,N_17895);
and U19428 (N_19428,N_17605,N_17791);
nor U19429 (N_19429,N_17458,N_16653);
nand U19430 (N_19430,N_16244,N_17703);
nand U19431 (N_19431,N_17765,N_16767);
nand U19432 (N_19432,N_16345,N_16406);
or U19433 (N_19433,N_16026,N_16628);
nand U19434 (N_19434,N_16187,N_17978);
nand U19435 (N_19435,N_16616,N_16172);
nor U19436 (N_19436,N_16280,N_16247);
and U19437 (N_19437,N_16649,N_17046);
and U19438 (N_19438,N_17204,N_16303);
and U19439 (N_19439,N_16810,N_17574);
nand U19440 (N_19440,N_16204,N_17858);
nand U19441 (N_19441,N_16235,N_16883);
and U19442 (N_19442,N_16293,N_16184);
or U19443 (N_19443,N_17854,N_16102);
or U19444 (N_19444,N_16708,N_17636);
or U19445 (N_19445,N_16466,N_17536);
or U19446 (N_19446,N_17718,N_17793);
nand U19447 (N_19447,N_17901,N_17561);
nand U19448 (N_19448,N_17810,N_16970);
xor U19449 (N_19449,N_17452,N_16953);
and U19450 (N_19450,N_17783,N_16620);
or U19451 (N_19451,N_17960,N_16367);
and U19452 (N_19452,N_17975,N_16691);
and U19453 (N_19453,N_17503,N_17811);
or U19454 (N_19454,N_17925,N_17972);
or U19455 (N_19455,N_16660,N_17729);
and U19456 (N_19456,N_17586,N_16519);
or U19457 (N_19457,N_16794,N_17955);
nor U19458 (N_19458,N_16698,N_17327);
or U19459 (N_19459,N_17046,N_16088);
nor U19460 (N_19460,N_16426,N_16813);
nor U19461 (N_19461,N_16155,N_16361);
nor U19462 (N_19462,N_17228,N_17141);
xnor U19463 (N_19463,N_17321,N_17487);
nand U19464 (N_19464,N_17030,N_17532);
xnor U19465 (N_19465,N_16461,N_17503);
and U19466 (N_19466,N_16415,N_16614);
and U19467 (N_19467,N_17158,N_16521);
nor U19468 (N_19468,N_16353,N_17085);
nand U19469 (N_19469,N_17260,N_16757);
nor U19470 (N_19470,N_16482,N_17320);
nand U19471 (N_19471,N_17396,N_16486);
nand U19472 (N_19472,N_16059,N_16752);
nand U19473 (N_19473,N_17714,N_17225);
nand U19474 (N_19474,N_16440,N_17408);
nor U19475 (N_19475,N_16406,N_16396);
or U19476 (N_19476,N_16672,N_16154);
nand U19477 (N_19477,N_16199,N_16725);
and U19478 (N_19478,N_16819,N_16459);
nor U19479 (N_19479,N_17984,N_16828);
nor U19480 (N_19480,N_16661,N_16201);
nor U19481 (N_19481,N_16517,N_17998);
nand U19482 (N_19482,N_16287,N_16701);
or U19483 (N_19483,N_16506,N_17675);
nor U19484 (N_19484,N_17849,N_16559);
and U19485 (N_19485,N_17793,N_17451);
or U19486 (N_19486,N_17300,N_17372);
or U19487 (N_19487,N_17148,N_16402);
or U19488 (N_19488,N_17518,N_16420);
or U19489 (N_19489,N_16057,N_17739);
nand U19490 (N_19490,N_16637,N_17543);
and U19491 (N_19491,N_17007,N_17944);
nor U19492 (N_19492,N_17031,N_16465);
nand U19493 (N_19493,N_17065,N_16902);
and U19494 (N_19494,N_16648,N_17033);
nor U19495 (N_19495,N_16187,N_16702);
and U19496 (N_19496,N_17111,N_17196);
or U19497 (N_19497,N_16503,N_17612);
or U19498 (N_19498,N_17768,N_16984);
nand U19499 (N_19499,N_17073,N_16494);
nor U19500 (N_19500,N_17745,N_17677);
and U19501 (N_19501,N_17206,N_17760);
nand U19502 (N_19502,N_17029,N_17442);
nor U19503 (N_19503,N_16632,N_17231);
or U19504 (N_19504,N_16129,N_17819);
or U19505 (N_19505,N_17272,N_17706);
nor U19506 (N_19506,N_16511,N_16980);
nand U19507 (N_19507,N_16566,N_17183);
and U19508 (N_19508,N_16151,N_17193);
or U19509 (N_19509,N_16009,N_17016);
and U19510 (N_19510,N_17311,N_17293);
nand U19511 (N_19511,N_17077,N_17946);
nor U19512 (N_19512,N_16196,N_17436);
nor U19513 (N_19513,N_17141,N_17836);
and U19514 (N_19514,N_16486,N_16368);
and U19515 (N_19515,N_17201,N_17949);
or U19516 (N_19516,N_16991,N_17238);
and U19517 (N_19517,N_17747,N_16818);
nor U19518 (N_19518,N_17868,N_17664);
nor U19519 (N_19519,N_16462,N_17965);
nand U19520 (N_19520,N_16555,N_16829);
nor U19521 (N_19521,N_17854,N_16570);
nand U19522 (N_19522,N_16107,N_17264);
and U19523 (N_19523,N_17537,N_17639);
or U19524 (N_19524,N_16709,N_17336);
or U19525 (N_19525,N_16628,N_16018);
and U19526 (N_19526,N_16355,N_17582);
nor U19527 (N_19527,N_16312,N_17778);
and U19528 (N_19528,N_16831,N_16548);
nand U19529 (N_19529,N_17027,N_17834);
nand U19530 (N_19530,N_17493,N_16224);
or U19531 (N_19531,N_17480,N_16875);
and U19532 (N_19532,N_16060,N_17792);
nand U19533 (N_19533,N_16171,N_17874);
nor U19534 (N_19534,N_16624,N_17927);
and U19535 (N_19535,N_17882,N_17720);
or U19536 (N_19536,N_16750,N_16957);
nor U19537 (N_19537,N_16254,N_17230);
nor U19538 (N_19538,N_16360,N_16052);
nor U19539 (N_19539,N_16633,N_17323);
nor U19540 (N_19540,N_16228,N_16564);
xor U19541 (N_19541,N_16921,N_17063);
nand U19542 (N_19542,N_16305,N_17885);
nand U19543 (N_19543,N_17785,N_17468);
and U19544 (N_19544,N_17263,N_16577);
nor U19545 (N_19545,N_17315,N_16412);
or U19546 (N_19546,N_16124,N_16250);
nor U19547 (N_19547,N_17190,N_16133);
and U19548 (N_19548,N_17718,N_17989);
or U19549 (N_19549,N_17949,N_17126);
xnor U19550 (N_19550,N_16487,N_17968);
nand U19551 (N_19551,N_16245,N_17709);
or U19552 (N_19552,N_17359,N_17851);
nand U19553 (N_19553,N_16603,N_17129);
nand U19554 (N_19554,N_16731,N_17622);
or U19555 (N_19555,N_16428,N_16366);
or U19556 (N_19556,N_16708,N_16099);
nor U19557 (N_19557,N_17527,N_17782);
nand U19558 (N_19558,N_17667,N_16319);
nand U19559 (N_19559,N_16458,N_16077);
or U19560 (N_19560,N_16606,N_16177);
nand U19561 (N_19561,N_17349,N_17702);
nand U19562 (N_19562,N_17433,N_17175);
and U19563 (N_19563,N_16143,N_16943);
xnor U19564 (N_19564,N_16551,N_16946);
and U19565 (N_19565,N_17348,N_17105);
nor U19566 (N_19566,N_17032,N_16909);
or U19567 (N_19567,N_17618,N_16939);
xor U19568 (N_19568,N_17232,N_16317);
nand U19569 (N_19569,N_17991,N_16537);
and U19570 (N_19570,N_17100,N_17415);
and U19571 (N_19571,N_16890,N_16932);
nor U19572 (N_19572,N_16737,N_17601);
nor U19573 (N_19573,N_16453,N_17324);
nor U19574 (N_19574,N_16220,N_16826);
nand U19575 (N_19575,N_17261,N_16346);
or U19576 (N_19576,N_16294,N_16295);
nand U19577 (N_19577,N_17412,N_16895);
nor U19578 (N_19578,N_16645,N_17626);
nand U19579 (N_19579,N_17380,N_16636);
nor U19580 (N_19580,N_17096,N_17237);
nor U19581 (N_19581,N_17241,N_16305);
and U19582 (N_19582,N_17729,N_17570);
nor U19583 (N_19583,N_16215,N_16145);
or U19584 (N_19584,N_16859,N_17578);
or U19585 (N_19585,N_17103,N_16234);
or U19586 (N_19586,N_17734,N_17518);
nor U19587 (N_19587,N_16811,N_17603);
and U19588 (N_19588,N_17177,N_16046);
or U19589 (N_19589,N_17588,N_17266);
nor U19590 (N_19590,N_17851,N_16152);
nor U19591 (N_19591,N_17005,N_17151);
and U19592 (N_19592,N_17209,N_17359);
or U19593 (N_19593,N_17039,N_17673);
or U19594 (N_19594,N_17504,N_16885);
or U19595 (N_19595,N_16033,N_16624);
or U19596 (N_19596,N_16135,N_16462);
nor U19597 (N_19597,N_16205,N_16741);
and U19598 (N_19598,N_17195,N_17916);
nor U19599 (N_19599,N_16901,N_16109);
and U19600 (N_19600,N_17235,N_16734);
nand U19601 (N_19601,N_16427,N_16756);
nand U19602 (N_19602,N_16947,N_17700);
xor U19603 (N_19603,N_17521,N_16450);
nor U19604 (N_19604,N_17950,N_17498);
or U19605 (N_19605,N_17068,N_16420);
or U19606 (N_19606,N_17160,N_17646);
nand U19607 (N_19607,N_17057,N_17766);
nand U19608 (N_19608,N_16487,N_17140);
or U19609 (N_19609,N_16364,N_16412);
and U19610 (N_19610,N_16800,N_16275);
nor U19611 (N_19611,N_16232,N_16167);
nor U19612 (N_19612,N_16432,N_17124);
nor U19613 (N_19613,N_17929,N_16431);
and U19614 (N_19614,N_16045,N_17701);
nand U19615 (N_19615,N_16203,N_17058);
nand U19616 (N_19616,N_16302,N_17467);
nand U19617 (N_19617,N_16708,N_17398);
nor U19618 (N_19618,N_17605,N_16760);
nor U19619 (N_19619,N_17159,N_16714);
nor U19620 (N_19620,N_17346,N_16343);
nand U19621 (N_19621,N_16660,N_17245);
and U19622 (N_19622,N_16089,N_17558);
and U19623 (N_19623,N_16501,N_16658);
nand U19624 (N_19624,N_16804,N_17631);
nand U19625 (N_19625,N_16147,N_17569);
nor U19626 (N_19626,N_16801,N_17688);
or U19627 (N_19627,N_17371,N_16068);
nand U19628 (N_19628,N_16036,N_16488);
nor U19629 (N_19629,N_16621,N_17400);
nand U19630 (N_19630,N_16476,N_17078);
or U19631 (N_19631,N_16718,N_16137);
nand U19632 (N_19632,N_16372,N_16853);
nor U19633 (N_19633,N_16139,N_17147);
nor U19634 (N_19634,N_16880,N_17378);
nand U19635 (N_19635,N_17553,N_16244);
or U19636 (N_19636,N_17251,N_17759);
nand U19637 (N_19637,N_16300,N_16099);
and U19638 (N_19638,N_17844,N_16123);
nand U19639 (N_19639,N_17600,N_16438);
and U19640 (N_19640,N_16922,N_17432);
nor U19641 (N_19641,N_16543,N_17063);
and U19642 (N_19642,N_17489,N_16136);
nor U19643 (N_19643,N_17960,N_17427);
and U19644 (N_19644,N_17072,N_16532);
nor U19645 (N_19645,N_16237,N_17684);
nor U19646 (N_19646,N_16037,N_17901);
nor U19647 (N_19647,N_16771,N_17733);
nor U19648 (N_19648,N_17860,N_16625);
or U19649 (N_19649,N_17564,N_17049);
nor U19650 (N_19650,N_17906,N_17255);
or U19651 (N_19651,N_16392,N_17692);
or U19652 (N_19652,N_17893,N_17465);
xnor U19653 (N_19653,N_17604,N_17166);
and U19654 (N_19654,N_17536,N_16973);
or U19655 (N_19655,N_16646,N_16893);
xor U19656 (N_19656,N_17896,N_16407);
and U19657 (N_19657,N_16012,N_16085);
and U19658 (N_19658,N_16067,N_16539);
and U19659 (N_19659,N_16691,N_17228);
xor U19660 (N_19660,N_17394,N_17204);
xor U19661 (N_19661,N_17619,N_16191);
or U19662 (N_19662,N_16101,N_17321);
nor U19663 (N_19663,N_16129,N_16295);
nor U19664 (N_19664,N_16503,N_17934);
or U19665 (N_19665,N_16628,N_16280);
or U19666 (N_19666,N_17103,N_17574);
nand U19667 (N_19667,N_16294,N_16223);
nor U19668 (N_19668,N_17093,N_17771);
and U19669 (N_19669,N_17155,N_17704);
and U19670 (N_19670,N_17751,N_17085);
xnor U19671 (N_19671,N_17177,N_16177);
nor U19672 (N_19672,N_17215,N_16148);
and U19673 (N_19673,N_16284,N_17951);
nor U19674 (N_19674,N_16455,N_16817);
nor U19675 (N_19675,N_17222,N_17139);
nand U19676 (N_19676,N_17408,N_16525);
nor U19677 (N_19677,N_16379,N_17598);
and U19678 (N_19678,N_17721,N_17729);
nor U19679 (N_19679,N_16728,N_16835);
and U19680 (N_19680,N_17085,N_17040);
and U19681 (N_19681,N_17033,N_16098);
xor U19682 (N_19682,N_16723,N_17964);
nor U19683 (N_19683,N_17559,N_16687);
nand U19684 (N_19684,N_17200,N_16097);
nand U19685 (N_19685,N_17175,N_16032);
nor U19686 (N_19686,N_17571,N_16961);
and U19687 (N_19687,N_17139,N_17560);
or U19688 (N_19688,N_17331,N_17100);
and U19689 (N_19689,N_16978,N_17744);
and U19690 (N_19690,N_17373,N_17118);
nor U19691 (N_19691,N_17519,N_16972);
and U19692 (N_19692,N_16856,N_16308);
or U19693 (N_19693,N_16821,N_16366);
and U19694 (N_19694,N_17190,N_17551);
and U19695 (N_19695,N_16177,N_17432);
nand U19696 (N_19696,N_16904,N_17459);
or U19697 (N_19697,N_16119,N_16035);
and U19698 (N_19698,N_16126,N_16683);
and U19699 (N_19699,N_17815,N_17072);
and U19700 (N_19700,N_16015,N_16369);
nor U19701 (N_19701,N_16239,N_17406);
nor U19702 (N_19702,N_17427,N_17510);
nor U19703 (N_19703,N_16180,N_16644);
nor U19704 (N_19704,N_16949,N_17465);
or U19705 (N_19705,N_16714,N_16414);
and U19706 (N_19706,N_17515,N_16970);
nor U19707 (N_19707,N_16476,N_17736);
nor U19708 (N_19708,N_17614,N_17814);
and U19709 (N_19709,N_16408,N_17521);
and U19710 (N_19710,N_17110,N_16807);
or U19711 (N_19711,N_17826,N_17306);
and U19712 (N_19712,N_16875,N_17994);
and U19713 (N_19713,N_16185,N_16985);
or U19714 (N_19714,N_17814,N_17711);
and U19715 (N_19715,N_17326,N_17771);
or U19716 (N_19716,N_17333,N_16808);
nand U19717 (N_19717,N_16634,N_17140);
nor U19718 (N_19718,N_17915,N_17095);
and U19719 (N_19719,N_16774,N_17873);
or U19720 (N_19720,N_16593,N_17271);
nor U19721 (N_19721,N_17264,N_16707);
nor U19722 (N_19722,N_17842,N_16457);
or U19723 (N_19723,N_17314,N_16048);
and U19724 (N_19724,N_17718,N_17026);
nor U19725 (N_19725,N_17318,N_17198);
nand U19726 (N_19726,N_16147,N_17299);
or U19727 (N_19727,N_17549,N_16746);
or U19728 (N_19728,N_17706,N_17299);
nand U19729 (N_19729,N_17249,N_17453);
nor U19730 (N_19730,N_17080,N_16022);
nand U19731 (N_19731,N_16298,N_16615);
nand U19732 (N_19732,N_16852,N_17909);
or U19733 (N_19733,N_17825,N_17583);
and U19734 (N_19734,N_16218,N_17179);
nor U19735 (N_19735,N_16566,N_16338);
and U19736 (N_19736,N_17782,N_17247);
and U19737 (N_19737,N_17580,N_16324);
and U19738 (N_19738,N_16189,N_17621);
or U19739 (N_19739,N_16506,N_17249);
and U19740 (N_19740,N_17365,N_16122);
and U19741 (N_19741,N_16493,N_16636);
nand U19742 (N_19742,N_17782,N_17394);
or U19743 (N_19743,N_17445,N_17795);
xor U19744 (N_19744,N_16744,N_17222);
and U19745 (N_19745,N_16572,N_17002);
and U19746 (N_19746,N_17437,N_16054);
or U19747 (N_19747,N_17447,N_16978);
or U19748 (N_19748,N_16290,N_17461);
xnor U19749 (N_19749,N_16847,N_17547);
and U19750 (N_19750,N_16464,N_17770);
or U19751 (N_19751,N_17631,N_16719);
nand U19752 (N_19752,N_16186,N_17532);
and U19753 (N_19753,N_16552,N_16018);
or U19754 (N_19754,N_17322,N_17628);
nor U19755 (N_19755,N_17685,N_17012);
or U19756 (N_19756,N_17626,N_17094);
or U19757 (N_19757,N_16665,N_17546);
nand U19758 (N_19758,N_17996,N_16063);
nor U19759 (N_19759,N_17115,N_17497);
nand U19760 (N_19760,N_16969,N_17430);
nor U19761 (N_19761,N_16742,N_17811);
nand U19762 (N_19762,N_16954,N_16932);
nand U19763 (N_19763,N_17910,N_17008);
and U19764 (N_19764,N_17654,N_17365);
and U19765 (N_19765,N_17791,N_16987);
or U19766 (N_19766,N_16791,N_16478);
and U19767 (N_19767,N_17757,N_16944);
and U19768 (N_19768,N_17647,N_16198);
and U19769 (N_19769,N_17583,N_17161);
nor U19770 (N_19770,N_16349,N_17897);
or U19771 (N_19771,N_16887,N_17370);
and U19772 (N_19772,N_16555,N_17048);
nor U19773 (N_19773,N_16452,N_17094);
and U19774 (N_19774,N_16394,N_17841);
nor U19775 (N_19775,N_17497,N_17913);
xnor U19776 (N_19776,N_16425,N_17273);
or U19777 (N_19777,N_16304,N_17464);
nor U19778 (N_19778,N_17489,N_17525);
nor U19779 (N_19779,N_17550,N_17790);
nand U19780 (N_19780,N_16773,N_16153);
or U19781 (N_19781,N_16115,N_17854);
nand U19782 (N_19782,N_17960,N_17578);
nor U19783 (N_19783,N_16324,N_16306);
or U19784 (N_19784,N_16184,N_16427);
nand U19785 (N_19785,N_16465,N_17924);
nand U19786 (N_19786,N_17045,N_16557);
nor U19787 (N_19787,N_16485,N_17934);
nor U19788 (N_19788,N_16335,N_16925);
and U19789 (N_19789,N_17456,N_16249);
or U19790 (N_19790,N_16279,N_17129);
and U19791 (N_19791,N_16342,N_17902);
nor U19792 (N_19792,N_16346,N_16132);
nand U19793 (N_19793,N_16585,N_17800);
nand U19794 (N_19794,N_17497,N_17108);
nor U19795 (N_19795,N_17253,N_17220);
and U19796 (N_19796,N_17488,N_16759);
nor U19797 (N_19797,N_16958,N_17424);
and U19798 (N_19798,N_17403,N_16275);
and U19799 (N_19799,N_17795,N_17477);
and U19800 (N_19800,N_17580,N_16487);
nand U19801 (N_19801,N_16167,N_16870);
nor U19802 (N_19802,N_17177,N_17501);
and U19803 (N_19803,N_17767,N_16060);
nand U19804 (N_19804,N_16102,N_17646);
and U19805 (N_19805,N_16561,N_17275);
and U19806 (N_19806,N_17786,N_17106);
and U19807 (N_19807,N_17727,N_16796);
nand U19808 (N_19808,N_16780,N_16595);
nand U19809 (N_19809,N_16819,N_17295);
xor U19810 (N_19810,N_17297,N_17728);
nor U19811 (N_19811,N_16371,N_17864);
and U19812 (N_19812,N_16192,N_17458);
or U19813 (N_19813,N_17851,N_17841);
nand U19814 (N_19814,N_16063,N_16478);
or U19815 (N_19815,N_16917,N_16544);
nor U19816 (N_19816,N_16384,N_16747);
and U19817 (N_19817,N_16320,N_17892);
and U19818 (N_19818,N_16000,N_16921);
and U19819 (N_19819,N_16202,N_17445);
and U19820 (N_19820,N_16666,N_16003);
nor U19821 (N_19821,N_17706,N_17949);
or U19822 (N_19822,N_16563,N_16875);
and U19823 (N_19823,N_16164,N_17281);
and U19824 (N_19824,N_17063,N_17298);
nor U19825 (N_19825,N_16254,N_16414);
and U19826 (N_19826,N_17967,N_16862);
nand U19827 (N_19827,N_17423,N_17686);
nand U19828 (N_19828,N_16680,N_16996);
nand U19829 (N_19829,N_16357,N_16996);
or U19830 (N_19830,N_17074,N_17397);
or U19831 (N_19831,N_17563,N_16042);
and U19832 (N_19832,N_17894,N_16779);
nand U19833 (N_19833,N_17071,N_16417);
and U19834 (N_19834,N_16399,N_17600);
nand U19835 (N_19835,N_17845,N_17240);
or U19836 (N_19836,N_16505,N_16178);
nand U19837 (N_19837,N_16898,N_16496);
and U19838 (N_19838,N_16451,N_16226);
and U19839 (N_19839,N_16770,N_17945);
nor U19840 (N_19840,N_16619,N_17004);
nand U19841 (N_19841,N_17273,N_16268);
nor U19842 (N_19842,N_17777,N_16143);
and U19843 (N_19843,N_16610,N_16571);
nor U19844 (N_19844,N_16049,N_16024);
nand U19845 (N_19845,N_17299,N_16106);
or U19846 (N_19846,N_16538,N_16351);
or U19847 (N_19847,N_16762,N_16136);
and U19848 (N_19848,N_16620,N_17750);
nand U19849 (N_19849,N_17147,N_16137);
nand U19850 (N_19850,N_16783,N_17344);
nand U19851 (N_19851,N_16698,N_17986);
or U19852 (N_19852,N_16551,N_16809);
or U19853 (N_19853,N_16217,N_17835);
or U19854 (N_19854,N_17140,N_17904);
or U19855 (N_19855,N_17045,N_17655);
nor U19856 (N_19856,N_16485,N_16197);
nand U19857 (N_19857,N_16965,N_17712);
and U19858 (N_19858,N_17493,N_16642);
or U19859 (N_19859,N_16310,N_16903);
and U19860 (N_19860,N_16332,N_17050);
nand U19861 (N_19861,N_16832,N_17896);
and U19862 (N_19862,N_16089,N_16187);
nand U19863 (N_19863,N_17218,N_16811);
nand U19864 (N_19864,N_16881,N_16092);
and U19865 (N_19865,N_16509,N_16326);
nor U19866 (N_19866,N_16404,N_17808);
and U19867 (N_19867,N_16303,N_17569);
nor U19868 (N_19868,N_16255,N_16246);
nor U19869 (N_19869,N_16277,N_17486);
nor U19870 (N_19870,N_17684,N_16440);
or U19871 (N_19871,N_16047,N_16567);
nor U19872 (N_19872,N_16918,N_16304);
nand U19873 (N_19873,N_16156,N_16248);
or U19874 (N_19874,N_17762,N_17469);
nor U19875 (N_19875,N_16879,N_17157);
nor U19876 (N_19876,N_16373,N_17677);
or U19877 (N_19877,N_16613,N_16576);
nor U19878 (N_19878,N_17935,N_16599);
nand U19879 (N_19879,N_17603,N_16319);
nor U19880 (N_19880,N_17808,N_16121);
nor U19881 (N_19881,N_16011,N_17146);
nand U19882 (N_19882,N_16425,N_16272);
nor U19883 (N_19883,N_16810,N_17938);
and U19884 (N_19884,N_16827,N_17369);
or U19885 (N_19885,N_17199,N_17767);
and U19886 (N_19886,N_16067,N_17955);
or U19887 (N_19887,N_17710,N_17747);
and U19888 (N_19888,N_17069,N_16745);
nand U19889 (N_19889,N_17144,N_17520);
or U19890 (N_19890,N_16887,N_17513);
or U19891 (N_19891,N_16880,N_17724);
nor U19892 (N_19892,N_16866,N_16267);
and U19893 (N_19893,N_16367,N_16190);
and U19894 (N_19894,N_17811,N_16229);
nand U19895 (N_19895,N_17118,N_16151);
or U19896 (N_19896,N_17461,N_17416);
and U19897 (N_19897,N_17014,N_16920);
nand U19898 (N_19898,N_16629,N_17494);
and U19899 (N_19899,N_17665,N_16553);
or U19900 (N_19900,N_17503,N_16951);
or U19901 (N_19901,N_17179,N_17814);
and U19902 (N_19902,N_17844,N_16828);
and U19903 (N_19903,N_16606,N_16690);
or U19904 (N_19904,N_17515,N_17917);
nor U19905 (N_19905,N_17842,N_17027);
nor U19906 (N_19906,N_16711,N_16553);
nor U19907 (N_19907,N_16341,N_16428);
and U19908 (N_19908,N_16201,N_17625);
and U19909 (N_19909,N_16236,N_16620);
xor U19910 (N_19910,N_16508,N_17136);
nand U19911 (N_19911,N_16157,N_16123);
and U19912 (N_19912,N_16611,N_16223);
nor U19913 (N_19913,N_17076,N_16670);
nor U19914 (N_19914,N_16261,N_17225);
or U19915 (N_19915,N_17503,N_16445);
and U19916 (N_19916,N_16415,N_17284);
nor U19917 (N_19917,N_16282,N_16072);
and U19918 (N_19918,N_16119,N_17392);
and U19919 (N_19919,N_16373,N_16914);
nor U19920 (N_19920,N_16351,N_17457);
nor U19921 (N_19921,N_16199,N_16853);
xnor U19922 (N_19922,N_16542,N_16132);
nand U19923 (N_19923,N_16896,N_16022);
nand U19924 (N_19924,N_16385,N_16149);
and U19925 (N_19925,N_17154,N_17909);
and U19926 (N_19926,N_17576,N_17722);
or U19927 (N_19927,N_17336,N_17106);
nand U19928 (N_19928,N_16033,N_17959);
nor U19929 (N_19929,N_16050,N_16068);
or U19930 (N_19930,N_17048,N_17144);
nor U19931 (N_19931,N_16667,N_16404);
or U19932 (N_19932,N_17823,N_16185);
or U19933 (N_19933,N_16727,N_17422);
or U19934 (N_19934,N_17022,N_17394);
nand U19935 (N_19935,N_16517,N_17070);
or U19936 (N_19936,N_16597,N_16076);
or U19937 (N_19937,N_16516,N_16277);
or U19938 (N_19938,N_16129,N_16493);
nand U19939 (N_19939,N_17791,N_17297);
and U19940 (N_19940,N_17360,N_16299);
and U19941 (N_19941,N_16408,N_17442);
xnor U19942 (N_19942,N_16839,N_16251);
nor U19943 (N_19943,N_17680,N_16943);
xor U19944 (N_19944,N_17130,N_17312);
nor U19945 (N_19945,N_17860,N_16446);
or U19946 (N_19946,N_17101,N_16567);
and U19947 (N_19947,N_16104,N_17167);
or U19948 (N_19948,N_16865,N_16857);
and U19949 (N_19949,N_16291,N_16881);
nor U19950 (N_19950,N_17160,N_17622);
or U19951 (N_19951,N_16548,N_17796);
and U19952 (N_19952,N_16798,N_17993);
nor U19953 (N_19953,N_17021,N_17333);
or U19954 (N_19954,N_17544,N_17602);
and U19955 (N_19955,N_17554,N_17977);
nor U19956 (N_19956,N_16045,N_17615);
nand U19957 (N_19957,N_17905,N_16784);
or U19958 (N_19958,N_16356,N_17877);
and U19959 (N_19959,N_16842,N_16152);
and U19960 (N_19960,N_17152,N_17793);
and U19961 (N_19961,N_16692,N_16684);
and U19962 (N_19962,N_16044,N_17669);
nand U19963 (N_19963,N_16222,N_17603);
and U19964 (N_19964,N_17183,N_17481);
or U19965 (N_19965,N_16140,N_17454);
nand U19966 (N_19966,N_16840,N_17730);
nor U19967 (N_19967,N_16887,N_17865);
nand U19968 (N_19968,N_17601,N_17854);
and U19969 (N_19969,N_17856,N_16242);
nand U19970 (N_19970,N_17943,N_17707);
or U19971 (N_19971,N_16459,N_16506);
nor U19972 (N_19972,N_16288,N_17274);
or U19973 (N_19973,N_17078,N_16389);
and U19974 (N_19974,N_16111,N_16247);
and U19975 (N_19975,N_17961,N_16264);
nand U19976 (N_19976,N_16495,N_17534);
or U19977 (N_19977,N_16365,N_16724);
nor U19978 (N_19978,N_17891,N_17339);
and U19979 (N_19979,N_17213,N_17068);
nor U19980 (N_19980,N_16503,N_16732);
and U19981 (N_19981,N_16873,N_16792);
or U19982 (N_19982,N_17195,N_16584);
nor U19983 (N_19983,N_16827,N_17343);
xor U19984 (N_19984,N_17645,N_17618);
nor U19985 (N_19985,N_17559,N_16953);
and U19986 (N_19986,N_17126,N_17792);
and U19987 (N_19987,N_16978,N_16630);
or U19988 (N_19988,N_16948,N_17587);
and U19989 (N_19989,N_16149,N_17820);
and U19990 (N_19990,N_17623,N_17065);
or U19991 (N_19991,N_16861,N_17515);
nor U19992 (N_19992,N_16860,N_17292);
and U19993 (N_19993,N_16634,N_17900);
or U19994 (N_19994,N_17842,N_16322);
or U19995 (N_19995,N_16043,N_16637);
nor U19996 (N_19996,N_16864,N_16612);
nand U19997 (N_19997,N_16771,N_16494);
or U19998 (N_19998,N_17066,N_16295);
nand U19999 (N_19999,N_17767,N_16389);
or U20000 (N_20000,N_19508,N_18684);
nand U20001 (N_20001,N_19161,N_19384);
or U20002 (N_20002,N_18665,N_18342);
nand U20003 (N_20003,N_18709,N_19077);
nand U20004 (N_20004,N_19179,N_18820);
nand U20005 (N_20005,N_18654,N_18178);
and U20006 (N_20006,N_18591,N_19403);
or U20007 (N_20007,N_19738,N_19210);
nor U20008 (N_20008,N_19919,N_18574);
and U20009 (N_20009,N_19338,N_18440);
nand U20010 (N_20010,N_18797,N_18495);
nand U20011 (N_20011,N_18229,N_19168);
or U20012 (N_20012,N_19498,N_19901);
nor U20013 (N_20013,N_19306,N_19702);
and U20014 (N_20014,N_19676,N_18103);
or U20015 (N_20015,N_18263,N_18607);
nand U20016 (N_20016,N_19626,N_18421);
or U20017 (N_20017,N_19223,N_18755);
or U20018 (N_20018,N_18208,N_19039);
or U20019 (N_20019,N_18959,N_19294);
nor U20020 (N_20020,N_19700,N_18774);
nand U20021 (N_20021,N_18882,N_19360);
xnor U20022 (N_20022,N_19097,N_19862);
nand U20023 (N_20023,N_19092,N_18622);
and U20024 (N_20024,N_18157,N_18334);
or U20025 (N_20025,N_19453,N_19318);
nor U20026 (N_20026,N_19510,N_19892);
nand U20027 (N_20027,N_18643,N_19049);
nor U20028 (N_20028,N_19851,N_18624);
or U20029 (N_20029,N_18687,N_19749);
nand U20030 (N_20030,N_18058,N_18854);
or U20031 (N_20031,N_19379,N_19973);
nand U20032 (N_20032,N_19727,N_18722);
nor U20033 (N_20033,N_19116,N_19916);
or U20034 (N_20034,N_19833,N_18748);
nor U20035 (N_20035,N_19088,N_18353);
nor U20036 (N_20036,N_19733,N_19528);
and U20037 (N_20037,N_18780,N_18679);
nand U20038 (N_20038,N_19705,N_19600);
or U20039 (N_20039,N_19767,N_19606);
nor U20040 (N_20040,N_19982,N_19840);
and U20041 (N_20041,N_19504,N_19740);
nor U20042 (N_20042,N_18620,N_19531);
or U20043 (N_20043,N_18473,N_18932);
nor U20044 (N_20044,N_19643,N_18828);
nor U20045 (N_20045,N_19741,N_18521);
nand U20046 (N_20046,N_18673,N_19932);
and U20047 (N_20047,N_18575,N_18518);
and U20048 (N_20048,N_19425,N_18723);
nor U20049 (N_20049,N_18137,N_18787);
or U20050 (N_20050,N_18918,N_19664);
nand U20051 (N_20051,N_19923,N_18803);
and U20052 (N_20052,N_18243,N_18339);
or U20053 (N_20053,N_18579,N_18319);
or U20054 (N_20054,N_18773,N_18795);
or U20055 (N_20055,N_19542,N_19291);
nor U20056 (N_20056,N_19969,N_18556);
or U20057 (N_20057,N_19458,N_18347);
or U20058 (N_20058,N_19133,N_18459);
nor U20059 (N_20059,N_18156,N_19823);
nor U20060 (N_20060,N_18540,N_19794);
or U20061 (N_20061,N_19480,N_19226);
nand U20062 (N_20062,N_19908,N_18593);
nand U20063 (N_20063,N_18976,N_19656);
and U20064 (N_20064,N_18983,N_18354);
nand U20065 (N_20065,N_19243,N_19264);
nor U20066 (N_20066,N_19107,N_18850);
and U20067 (N_20067,N_18202,N_18782);
nor U20068 (N_20068,N_18439,N_18890);
nand U20069 (N_20069,N_19361,N_18859);
or U20070 (N_20070,N_18199,N_18311);
and U20071 (N_20071,N_19772,N_18572);
or U20072 (N_20072,N_18701,N_18292);
nor U20073 (N_20073,N_19314,N_18594);
nor U20074 (N_20074,N_18635,N_18921);
or U20075 (N_20075,N_19565,N_19960);
or U20076 (N_20076,N_18857,N_18125);
or U20077 (N_20077,N_18499,N_19156);
nand U20078 (N_20078,N_19597,N_19878);
nor U20079 (N_20079,N_19102,N_19050);
or U20080 (N_20080,N_19985,N_19699);
or U20081 (N_20081,N_19225,N_18251);
nor U20082 (N_20082,N_18945,N_18379);
or U20083 (N_20083,N_19138,N_19165);
nand U20084 (N_20084,N_19274,N_19736);
and U20085 (N_20085,N_19959,N_19414);
and U20086 (N_20086,N_19559,N_18564);
nor U20087 (N_20087,N_19266,N_18588);
nand U20088 (N_20088,N_19351,N_18852);
nand U20089 (N_20089,N_19972,N_19182);
nor U20090 (N_20090,N_18650,N_18645);
or U20091 (N_20091,N_18470,N_19764);
and U20092 (N_20092,N_18066,N_18532);
and U20093 (N_20093,N_19158,N_19713);
nand U20094 (N_20094,N_18724,N_19680);
nor U20095 (N_20095,N_18326,N_19350);
and U20096 (N_20096,N_19029,N_18966);
nor U20097 (N_20097,N_18249,N_18336);
nor U20098 (N_20098,N_18169,N_18605);
and U20099 (N_20099,N_19711,N_18906);
and U20100 (N_20100,N_18506,N_19826);
or U20101 (N_20101,N_18592,N_19634);
or U20102 (N_20102,N_18908,N_18068);
and U20103 (N_20103,N_19560,N_19006);
or U20104 (N_20104,N_18919,N_18894);
and U20105 (N_20105,N_18410,N_18798);
nor U20106 (N_20106,N_18985,N_19513);
or U20107 (N_20107,N_19961,N_18734);
nor U20108 (N_20108,N_19954,N_18286);
nand U20109 (N_20109,N_19881,N_19455);
or U20110 (N_20110,N_18443,N_19089);
and U20111 (N_20111,N_19906,N_18660);
and U20112 (N_20112,N_18167,N_18562);
and U20113 (N_20113,N_19691,N_18267);
nand U20114 (N_20114,N_18806,N_18550);
nand U20115 (N_20115,N_19001,N_18314);
or U20116 (N_20116,N_19305,N_18427);
nand U20117 (N_20117,N_18638,N_18955);
or U20118 (N_20118,N_18519,N_18329);
nand U20119 (N_20119,N_18967,N_18998);
nor U20120 (N_20120,N_19048,N_19582);
nor U20121 (N_20121,N_18931,N_19682);
and U20122 (N_20122,N_18255,N_19693);
nor U20123 (N_20123,N_19619,N_18851);
or U20124 (N_20124,N_18747,N_18370);
or U20125 (N_20125,N_18390,N_18002);
or U20126 (N_20126,N_19992,N_18920);
and U20127 (N_20127,N_18980,N_18538);
xor U20128 (N_20128,N_18714,N_19020);
nor U20129 (N_20129,N_18301,N_18581);
nand U20130 (N_20130,N_18365,N_18358);
and U20131 (N_20131,N_19614,N_18783);
nor U20132 (N_20132,N_18460,N_18726);
or U20133 (N_20133,N_18106,N_18653);
nand U20134 (N_20134,N_18116,N_19363);
and U20135 (N_20135,N_18646,N_19777);
and U20136 (N_20136,N_18796,N_18320);
nor U20137 (N_20137,N_19476,N_18674);
and U20138 (N_20138,N_19256,N_18247);
or U20139 (N_20139,N_19041,N_18328);
and U20140 (N_20140,N_18299,N_19548);
nor U20141 (N_20141,N_18601,N_19339);
or U20142 (N_20142,N_18055,N_18992);
xor U20143 (N_20143,N_19530,N_18359);
and U20144 (N_20144,N_18203,N_19889);
nand U20145 (N_20145,N_19164,N_19971);
and U20146 (N_20146,N_19714,N_18697);
nor U20147 (N_20147,N_19364,N_18119);
nor U20148 (N_20148,N_18455,N_19445);
or U20149 (N_20149,N_19808,N_19975);
and U20150 (N_20150,N_18631,N_19467);
or U20151 (N_20151,N_19150,N_18128);
and U20152 (N_20152,N_18600,N_19538);
nand U20153 (N_20153,N_18212,N_18907);
nor U20154 (N_20154,N_19573,N_18392);
nor U20155 (N_20155,N_18472,N_18129);
and U20156 (N_20156,N_19842,N_18482);
nor U20157 (N_20157,N_19821,N_18713);
nand U20158 (N_20158,N_18911,N_18010);
nand U20159 (N_20159,N_19278,N_19797);
and U20160 (N_20160,N_19353,N_19724);
nor U20161 (N_20161,N_19601,N_19920);
or U20162 (N_20162,N_19781,N_18727);
or U20163 (N_20163,N_19084,N_18578);
or U20164 (N_20164,N_18205,N_18887);
and U20165 (N_20165,N_18544,N_18996);
nand U20166 (N_20166,N_18414,N_18166);
nor U20167 (N_20167,N_18929,N_18045);
nand U20168 (N_20168,N_19488,N_19236);
xnor U20169 (N_20169,N_18096,N_19146);
nand U20170 (N_20170,N_19240,N_19307);
and U20171 (N_20171,N_18982,N_18159);
nand U20172 (N_20172,N_18809,N_18260);
or U20173 (N_20173,N_18695,N_18073);
and U20174 (N_20174,N_18424,N_18355);
nor U20175 (N_20175,N_18056,N_19320);
or U20176 (N_20176,N_18386,N_18312);
and U20177 (N_20177,N_18017,N_18345);
nor U20178 (N_20178,N_19847,N_19782);
nand U20179 (N_20179,N_19864,N_19454);
or U20180 (N_20180,N_18102,N_18559);
nand U20181 (N_20181,N_18133,N_19227);
and U20182 (N_20182,N_19887,N_19061);
nor U20183 (N_20183,N_19543,N_18207);
nand U20184 (N_20184,N_18975,N_18739);
nand U20185 (N_20185,N_19673,N_18321);
and U20186 (N_20186,N_19469,N_18287);
or U20187 (N_20187,N_19378,N_18019);
nor U20188 (N_20188,N_19856,N_18836);
nor U20189 (N_20189,N_19417,N_18171);
nand U20190 (N_20190,N_18016,N_18174);
nand U20191 (N_20191,N_19261,N_18905);
nand U20192 (N_20192,N_19106,N_18496);
and U20193 (N_20193,N_18323,N_18131);
nor U20194 (N_20194,N_18953,N_19845);
nor U20195 (N_20195,N_18930,N_19463);
nor U20196 (N_20196,N_18669,N_18222);
or U20197 (N_20197,N_19428,N_18230);
and U20198 (N_20198,N_19792,N_19407);
and U20199 (N_20199,N_18121,N_19905);
and U20200 (N_20200,N_19046,N_18337);
or U20201 (N_20201,N_19745,N_18737);
and U20202 (N_20202,N_18611,N_18493);
and U20203 (N_20203,N_18134,N_19003);
or U20204 (N_20204,N_19562,N_19316);
nor U20205 (N_20205,N_19737,N_19841);
and U20206 (N_20206,N_19649,N_18030);
nor U20207 (N_20207,N_19547,N_19372);
nand U20208 (N_20208,N_18541,N_18510);
nor U20209 (N_20209,N_19686,N_19780);
nor U20210 (N_20210,N_18901,N_18457);
or U20211 (N_20211,N_19169,N_18252);
nand U20212 (N_20212,N_18954,N_19790);
and U20213 (N_20213,N_19394,N_18257);
or U20214 (N_20214,N_19366,N_19410);
and U20215 (N_20215,N_18123,N_19071);
nand U20216 (N_20216,N_19057,N_18762);
nor U20217 (N_20217,N_19712,N_18395);
or U20218 (N_20218,N_18240,N_19219);
nand U20219 (N_20219,N_19062,N_19857);
nor U20220 (N_20220,N_18034,N_18662);
and U20221 (N_20221,N_19073,N_19578);
or U20222 (N_20222,N_18098,N_19625);
nor U20223 (N_20223,N_19994,N_19086);
nor U20224 (N_20224,N_18136,N_19516);
nor U20225 (N_20225,N_19398,N_18808);
nor U20226 (N_20226,N_19861,N_18608);
and U20227 (N_20227,N_19438,N_18740);
or U20228 (N_20228,N_18776,N_18076);
and U20229 (N_20229,N_18213,N_19167);
nand U20230 (N_20230,N_18446,N_19060);
xnor U20231 (N_20231,N_19501,N_18602);
or U20232 (N_20232,N_18476,N_19154);
or U20233 (N_20233,N_19949,N_19837);
or U20234 (N_20234,N_19239,N_19276);
and U20235 (N_20235,N_19789,N_19687);
and U20236 (N_20236,N_18704,N_18143);
nand U20237 (N_20237,N_18441,N_19915);
nor U20238 (N_20238,N_19104,N_19660);
or U20239 (N_20239,N_18168,N_19828);
or U20240 (N_20240,N_18069,N_18027);
nor U20241 (N_20241,N_18743,N_19868);
nor U20242 (N_20242,N_18228,N_19388);
nor U20243 (N_20243,N_18616,N_19209);
nand U20244 (N_20244,N_18420,N_18313);
or U20245 (N_20245,N_19776,N_18490);
or U20246 (N_20246,N_19279,N_18138);
or U20247 (N_20247,N_18132,N_19173);
or U20248 (N_20248,N_18672,N_18369);
xor U20249 (N_20249,N_18682,N_18969);
nand U20250 (N_20250,N_19635,N_18663);
nor U20251 (N_20251,N_19936,N_19218);
and U20252 (N_20252,N_18481,N_19392);
xor U20253 (N_20253,N_19963,N_18511);
or U20254 (N_20254,N_18094,N_19537);
and U20255 (N_20255,N_18938,N_19103);
nor U20256 (N_20256,N_18195,N_18124);
and U20257 (N_20257,N_18527,N_18348);
and U20258 (N_20258,N_19967,N_19824);
or U20259 (N_20259,N_19918,N_18742);
or U20260 (N_20260,N_19630,N_19938);
nand U20261 (N_20261,N_19254,N_19836);
and U20262 (N_20262,N_19462,N_18553);
nor U20263 (N_20263,N_18135,N_18080);
nor U20264 (N_20264,N_18707,N_18877);
nor U20265 (N_20265,N_18396,N_18373);
nor U20266 (N_20266,N_18839,N_19008);
nand U20267 (N_20267,N_18934,N_19328);
nor U20268 (N_20268,N_19147,N_18351);
or U20269 (N_20269,N_18758,N_18084);
nor U20270 (N_20270,N_18560,N_19252);
and U20271 (N_20271,N_19611,N_18915);
nand U20272 (N_20272,N_19275,N_19436);
nor U20273 (N_20273,N_19246,N_19390);
nor U20274 (N_20274,N_18467,N_19335);
nand U20275 (N_20275,N_19739,N_18289);
or U20276 (N_20276,N_19087,N_19134);
nor U20277 (N_20277,N_19928,N_18997);
and U20278 (N_20278,N_18895,N_19897);
nand U20279 (N_20279,N_19669,N_19819);
nor U20280 (N_20280,N_18035,N_18264);
and U20281 (N_20281,N_18083,N_19137);
or U20282 (N_20282,N_18706,N_18528);
or U20283 (N_20283,N_19387,N_18403);
and U20284 (N_20284,N_18087,N_18215);
xnor U20285 (N_20285,N_19369,N_18829);
nand U20286 (N_20286,N_18306,N_19203);
or U20287 (N_20287,N_19082,N_18659);
nor U20288 (N_20288,N_18075,N_19984);
nor U20289 (N_20289,N_19610,N_19659);
and U20290 (N_20290,N_19675,N_18625);
nor U20291 (N_20291,N_18122,N_19486);
and U20292 (N_20292,N_19078,N_18352);
and U20293 (N_20293,N_19094,N_18817);
nand U20294 (N_20294,N_18064,N_18361);
nor U20295 (N_20295,N_18793,N_18120);
or U20296 (N_20296,N_19309,N_19948);
nor U20297 (N_20297,N_19592,N_19429);
nor U20298 (N_20298,N_19290,N_18177);
nor U20299 (N_20299,N_18023,N_18309);
nor U20300 (N_20300,N_18233,N_18590);
nor U20301 (N_20301,N_19603,N_19449);
nand U20302 (N_20302,N_18449,N_19470);
and U20303 (N_20303,N_18430,N_19709);
or U20304 (N_20304,N_18061,N_19802);
and U20305 (N_20305,N_18914,N_18629);
nand U20306 (N_20306,N_19051,N_19189);
nor U20307 (N_20307,N_18547,N_18007);
and U20308 (N_20308,N_19602,N_18194);
and U20309 (N_20309,N_18686,N_18760);
and U20310 (N_20310,N_19213,N_19632);
nand U20311 (N_20311,N_19523,N_18474);
and U20312 (N_20312,N_18847,N_19838);
nor U20313 (N_20313,N_18183,N_19262);
or U20314 (N_20314,N_18147,N_19993);
nor U20315 (N_20315,N_19551,N_19882);
nand U20316 (N_20316,N_18595,N_18318);
nor U20317 (N_20317,N_18520,N_18656);
or U20318 (N_20318,N_18478,N_18814);
nand U20319 (N_20319,N_19858,N_18118);
and U20320 (N_20320,N_18811,N_19645);
and U20321 (N_20321,N_18943,N_18881);
nor U20322 (N_20322,N_18282,N_18442);
and U20323 (N_20323,N_19299,N_19520);
nor U20324 (N_20324,N_18718,N_19304);
or U20325 (N_20325,N_19204,N_19295);
and U20326 (N_20326,N_18006,N_19518);
and U20327 (N_20327,N_18717,N_19452);
nand U20328 (N_20328,N_18418,N_19701);
or U20329 (N_20329,N_19337,N_18970);
nor U20330 (N_20330,N_19230,N_18861);
and U20331 (N_20331,N_19759,N_19689);
and U20332 (N_20332,N_18070,N_18021);
or U20333 (N_20333,N_18285,N_19970);
and U20334 (N_20334,N_18567,N_18041);
and U20335 (N_20335,N_19242,N_19177);
and U20336 (N_20336,N_18197,N_18204);
nor U20337 (N_20337,N_19143,N_18962);
nand U20338 (N_20338,N_19024,N_19464);
nand U20339 (N_20339,N_19980,N_18603);
nor U20340 (N_20340,N_18805,N_18150);
nor U20341 (N_20341,N_18071,N_18031);
or U20342 (N_20342,N_19093,N_19101);
and U20343 (N_20343,N_18261,N_18632);
or U20344 (N_20344,N_18305,N_19058);
or U20345 (N_20345,N_19260,N_18275);
and U20346 (N_20346,N_18028,N_18503);
nor U20347 (N_20347,N_19883,N_19342);
nand U20348 (N_20348,N_18813,N_18926);
or U20349 (N_20349,N_19529,N_18639);
nor U20350 (N_20350,N_19332,N_19770);
xnor U20351 (N_20351,N_19067,N_19572);
nand U20352 (N_20352,N_19633,N_18381);
nand U20353 (N_20353,N_18524,N_18617);
or U20354 (N_20354,N_19485,N_19743);
and U20355 (N_20355,N_19575,N_19413);
nand U20356 (N_20356,N_19427,N_19070);
nor U20357 (N_20357,N_19144,N_19323);
or U20358 (N_20358,N_18164,N_18163);
and U20359 (N_20359,N_19622,N_18343);
xnor U20360 (N_20360,N_18063,N_19271);
and U20361 (N_20361,N_18079,N_19217);
or U20362 (N_20362,N_18377,N_19566);
nor U20363 (N_20363,N_19004,N_18480);
nand U20364 (N_20364,N_18586,N_18840);
nand U20365 (N_20365,N_18763,N_18526);
xor U20366 (N_20366,N_18827,N_18040);
or U20367 (N_20367,N_19953,N_19742);
or U20368 (N_20368,N_19331,N_18271);
and U20369 (N_20369,N_19871,N_18698);
nand U20370 (N_20370,N_18580,N_19207);
nor U20371 (N_20371,N_19251,N_18715);
and U20372 (N_20372,N_19253,N_18870);
nand U20373 (N_20373,N_19435,N_18383);
nand U20374 (N_20374,N_19406,N_19846);
or U20375 (N_20375,N_18784,N_18298);
nand U20376 (N_20376,N_19411,N_18775);
nor U20377 (N_20377,N_18568,N_19991);
nor U20378 (N_20378,N_19118,N_19382);
and U20379 (N_20379,N_18552,N_18004);
or U20380 (N_20380,N_18615,N_18081);
nand U20381 (N_20381,N_18426,N_18692);
or U20382 (N_20382,N_18729,N_19431);
nor U20383 (N_20383,N_18049,N_19465);
or U20384 (N_20384,N_18022,N_18224);
or U20385 (N_20385,N_18502,N_19657);
nor U20386 (N_20386,N_18876,N_19157);
and U20387 (N_20387,N_19214,N_19031);
nand U20388 (N_20388,N_18752,N_18823);
nor U20389 (N_20389,N_19312,N_19809);
nor U20390 (N_20390,N_19939,N_19719);
nor U20391 (N_20391,N_19695,N_19870);
and U20392 (N_20392,N_18380,N_18332);
or U20393 (N_20393,N_19012,N_19886);
and U20394 (N_20394,N_19748,N_18963);
nand U20395 (N_20395,N_19865,N_19995);
and U20396 (N_20396,N_18325,N_19663);
and U20397 (N_20397,N_19640,N_18826);
and U20398 (N_20398,N_18099,N_19065);
nor U20399 (N_20399,N_18751,N_19224);
xnor U20400 (N_20400,N_18879,N_18254);
nor U20401 (N_20401,N_18330,N_19460);
nor U20402 (N_20402,N_18710,N_18529);
or U20403 (N_20403,N_19926,N_19755);
and U20404 (N_20404,N_19422,N_19440);
nand U20405 (N_20405,N_19302,N_18657);
and U20406 (N_20406,N_18072,N_19609);
nor U20407 (N_20407,N_18621,N_18464);
nor U20408 (N_20408,N_18111,N_19481);
nand U20409 (N_20409,N_19176,N_18487);
nand U20410 (N_20410,N_18533,N_18767);
nand U20411 (N_20411,N_18346,N_18530);
nand U20412 (N_20412,N_19913,N_19141);
nand U20413 (N_20413,N_19018,N_19268);
and U20414 (N_20414,N_18265,N_19549);
nand U20415 (N_20415,N_19015,N_18765);
or U20416 (N_20416,N_18219,N_19424);
and U20417 (N_20417,N_19025,N_18274);
and U20418 (N_20418,N_19720,N_18766);
and U20419 (N_20419,N_19800,N_18191);
nor U20420 (N_20420,N_18018,N_18180);
or U20421 (N_20421,N_19190,N_19880);
nand U20422 (N_20422,N_19175,N_18917);
and U20423 (N_20423,N_19681,N_18262);
xor U20424 (N_20424,N_19310,N_19943);
or U20425 (N_20425,N_18154,N_18618);
nand U20426 (N_20426,N_18725,N_18676);
nand U20427 (N_20427,N_18946,N_19345);
nor U20428 (N_20428,N_18733,N_18489);
nand U20429 (N_20429,N_19968,N_19126);
and U20430 (N_20430,N_18471,N_18768);
and U20431 (N_20431,N_19491,N_18720);
nor U20432 (N_20432,N_19801,N_19839);
and U20433 (N_20433,N_19115,N_18977);
or U20434 (N_20434,N_19957,N_19385);
nor U20435 (N_20435,N_18192,N_18226);
nand U20436 (N_20436,N_19618,N_18873);
nand U20437 (N_20437,N_19329,N_18317);
nor U20438 (N_20438,N_18090,N_19376);
nand U20439 (N_20439,N_19222,N_19571);
xnor U20440 (N_20440,N_19456,N_19248);
and U20441 (N_20441,N_19763,N_18754);
nand U20442 (N_20442,N_18477,N_18500);
nor U20443 (N_20443,N_19399,N_19546);
nor U20444 (N_20444,N_19433,N_18892);
nand U20445 (N_20445,N_19421,N_18566);
nand U20446 (N_20446,N_18104,N_19912);
nand U20447 (N_20447,N_18296,N_18961);
and U20448 (N_20448,N_19193,N_19958);
nor U20449 (N_20449,N_19757,N_19567);
nand U20450 (N_20450,N_19874,N_19232);
and U20451 (N_20451,N_19344,N_18689);
nor U20452 (N_20452,N_19080,N_19552);
nor U20453 (N_20453,N_19479,N_18843);
nor U20454 (N_20454,N_18450,N_19021);
and U20455 (N_20455,N_18721,N_19921);
or U20456 (N_20456,N_18649,N_19723);
nor U20457 (N_20457,N_19945,N_19375);
nand U20458 (N_20458,N_18188,N_19033);
and U20459 (N_20459,N_19053,N_18509);
or U20460 (N_20460,N_19888,N_19277);
nor U20461 (N_20461,N_18385,N_19721);
and U20462 (N_20462,N_19055,N_19670);
and U20463 (N_20463,N_19293,N_19202);
and U20464 (N_20464,N_18290,N_18612);
nand U20465 (N_20465,N_18910,N_19550);
or U20466 (N_20466,N_19125,N_18050);
or U20467 (N_20467,N_18790,N_18273);
and U20468 (N_20468,N_18468,N_18461);
xor U20469 (N_20469,N_19844,N_18761);
nand U20470 (N_20470,N_18548,N_19245);
nand U20471 (N_20471,N_19482,N_18042);
nand U20472 (N_20472,N_18181,N_18641);
or U20473 (N_20473,N_18062,N_19617);
and U20474 (N_20474,N_19056,N_19775);
nand U20475 (N_20475,N_18279,N_19408);
and U20476 (N_20476,N_18973,N_18270);
and U20477 (N_20477,N_18824,N_18732);
and U20478 (N_20478,N_19326,N_18026);
nand U20479 (N_20479,N_19574,N_18344);
nand U20480 (N_20480,N_19322,N_19666);
nand U20481 (N_20481,N_19181,N_19979);
or U20482 (N_20482,N_19383,N_19221);
and U20483 (N_20483,N_19624,N_19389);
nor U20484 (N_20484,N_18384,N_18788);
and U20485 (N_20485,N_19629,N_19473);
nand U20486 (N_20486,N_19330,N_19272);
or U20487 (N_20487,N_18438,N_19244);
nand U20488 (N_20488,N_18756,N_19358);
nand U20489 (N_20489,N_18869,N_19052);
or U20490 (N_20490,N_19589,N_19876);
nand U20491 (N_20491,N_19352,N_19752);
nand U20492 (N_20492,N_19521,N_18140);
or U20493 (N_20493,N_18451,N_18853);
nor U20494 (N_20494,N_18234,N_18677);
nand U20495 (N_20495,N_18001,N_18277);
nand U20496 (N_20496,N_18652,N_18184);
or U20497 (N_20497,N_18903,N_18845);
nand U20498 (N_20498,N_19698,N_18272);
xor U20499 (N_20499,N_19075,N_18880);
and U20500 (N_20500,N_19955,N_19929);
or U20501 (N_20501,N_19966,N_19186);
or U20502 (N_20502,N_18949,N_19990);
and U20503 (N_20503,N_18206,N_19798);
and U20504 (N_20504,N_19220,N_19668);
nand U20505 (N_20505,N_19494,N_19027);
or U20506 (N_20506,N_18902,N_19365);
and U20507 (N_20507,N_18736,N_19621);
and U20508 (N_20508,N_19771,N_18927);
and U20509 (N_20509,N_18097,N_18878);
and U20510 (N_20510,N_18712,N_19877);
nand U20511 (N_20511,N_18735,N_18968);
and U20512 (N_20512,N_19750,N_19799);
and U20513 (N_20513,N_19806,N_18400);
and U20514 (N_20514,N_18419,N_19072);
or U20515 (N_20515,N_18448,N_18816);
nor U20516 (N_20516,N_18047,N_19784);
nor U20517 (N_20517,N_19340,N_18582);
or U20518 (N_20518,N_19758,N_18413);
nand U20519 (N_20519,N_19639,N_18161);
nor U20520 (N_20520,N_18619,N_18680);
and U20521 (N_20521,N_19296,N_18990);
nand U20522 (N_20522,N_19989,N_18144);
or U20523 (N_20523,N_19869,N_18838);
nor U20524 (N_20524,N_19710,N_19348);
or U20525 (N_20525,N_19933,N_18340);
nand U20526 (N_20526,N_18916,N_19153);
or U20527 (N_20527,N_18974,N_18779);
or U20528 (N_20528,N_18866,N_18214);
nand U20529 (N_20529,N_19661,N_19527);
and U20530 (N_20530,N_18812,N_19769);
and U20531 (N_20531,N_19581,N_19987);
nor U20532 (N_20532,N_18065,N_19519);
xor U20533 (N_20533,N_19450,N_19437);
and U20534 (N_20534,N_18492,N_18871);
nor U20535 (N_20535,N_19211,N_19849);
nor U20536 (N_20536,N_19627,N_18505);
nand U20537 (N_20537,N_18232,N_19641);
nor U20538 (N_20538,N_19499,N_19514);
and U20539 (N_20539,N_18863,N_19047);
or U20540 (N_20540,N_18683,N_18523);
nand U20541 (N_20541,N_18000,N_19674);
and U20542 (N_20542,N_19947,N_19568);
nor U20543 (N_20543,N_18221,N_19558);
and U20544 (N_20544,N_19356,N_19884);
or U20545 (N_20545,N_19650,N_18694);
nand U20546 (N_20546,N_19079,N_19091);
nor U20547 (N_20547,N_18944,N_18988);
xnor U20548 (N_20548,N_19950,N_19259);
nor U20549 (N_20549,N_19124,N_19315);
nor U20550 (N_20550,N_19483,N_18415);
and U20551 (N_20551,N_19718,N_19145);
and U20552 (N_20552,N_19303,N_18210);
nand U20553 (N_20553,N_18807,N_18165);
nand U20554 (N_20554,N_18280,N_19812);
or U20555 (N_20555,N_18539,N_19678);
and U20556 (N_20556,N_19159,N_18658);
nor U20557 (N_20557,N_18598,N_18833);
nor U20558 (N_20558,N_18405,N_18092);
and U20559 (N_20559,N_19956,N_19255);
and U20560 (N_20560,N_19238,N_18584);
xor U20561 (N_20561,N_19178,N_19343);
nand U20562 (N_20562,N_18534,N_18514);
nor U20563 (N_20563,N_18454,N_18597);
nand U20564 (N_20564,N_18117,N_19317);
nand U20565 (N_20565,N_19234,N_18036);
and U20566 (N_20566,N_19119,N_19005);
and U20567 (N_20567,N_19997,N_18151);
and U20568 (N_20568,N_19000,N_19935);
and U20569 (N_20569,N_18542,N_19099);
or U20570 (N_20570,N_19911,N_19298);
or U20571 (N_20571,N_18770,N_19988);
nand U20572 (N_20572,N_19768,N_19325);
nor U20573 (N_20573,N_19615,N_18393);
nand U20574 (N_20574,N_18360,N_19019);
nand U20575 (N_20575,N_19667,N_19142);
nand U20576 (N_20576,N_19152,N_18925);
nand U20577 (N_20577,N_18746,N_19130);
or U20578 (N_20578,N_19623,N_19579);
nand U20579 (N_20579,N_19492,N_19263);
or U20580 (N_20580,N_18469,N_19250);
nor U20581 (N_20581,N_18085,N_19612);
nand U20582 (N_20582,N_19570,N_18404);
nor U20583 (N_20583,N_19907,N_19747);
nor U20584 (N_20584,N_18268,N_19292);
nor U20585 (N_20585,N_19732,N_18231);
nor U20586 (N_20586,N_19135,N_19914);
or U20587 (N_20587,N_18670,N_18302);
xor U20588 (N_20588,N_19396,N_19395);
nor U20589 (N_20589,N_18308,N_19194);
nand U20590 (N_20590,N_19022,N_18115);
nor U20591 (N_20591,N_18948,N_18749);
nor U20592 (N_20592,N_19442,N_18648);
nand U20593 (N_20593,N_18924,N_19814);
and U20594 (N_20594,N_19493,N_18284);
nor U20595 (N_20595,N_18623,N_18753);
nor U20596 (N_20596,N_18173,N_19148);
or U20597 (N_20597,N_18741,N_19962);
nor U20598 (N_20598,N_18909,N_18668);
or U20599 (N_20599,N_18630,N_18052);
or U20600 (N_20600,N_19409,N_18978);
and U20601 (N_20601,N_19564,N_18333);
and U20602 (N_20602,N_19620,N_18227);
or U20603 (N_20603,N_19321,N_18951);
nand U20604 (N_20604,N_18037,N_19810);
nor U20605 (N_20605,N_19829,N_18561);
nand U20606 (N_20606,N_18860,N_19439);
nor U20607 (N_20607,N_18862,N_19557);
nand U20608 (N_20608,N_18357,N_19269);
nor U20609 (N_20609,N_19998,N_19704);
nand U20610 (N_20610,N_19201,N_18664);
or U20611 (N_20611,N_19397,N_18485);
and U20612 (N_20612,N_19490,N_19553);
nor U20613 (N_20613,N_18310,N_19977);
or U20614 (N_20614,N_18757,N_18434);
nand U20615 (N_20615,N_18609,N_18417);
and U20616 (N_20616,N_18371,N_19703);
nand U20617 (N_20617,N_19444,N_18494);
nand U20618 (N_20618,N_18048,N_18259);
nor U20619 (N_20619,N_19308,N_18486);
nand U20620 (N_20620,N_18488,N_19655);
or U20621 (N_20621,N_19893,N_19140);
nand U20622 (N_20622,N_19605,N_18610);
and U20623 (N_20623,N_19942,N_18834);
or U20624 (N_20624,N_18190,N_18238);
or U20625 (N_20625,N_18504,N_18889);
and U20626 (N_20626,N_19081,N_19347);
and U20627 (N_20627,N_19083,N_18573);
nand U20628 (N_20628,N_18211,N_18537);
and U20629 (N_20629,N_18196,N_19690);
nor U20630 (N_20630,N_18952,N_18835);
or U20631 (N_20631,N_18789,N_18912);
or U20632 (N_20632,N_18844,N_19854);
nand U20633 (N_20633,N_18012,N_18335);
and U20634 (N_20634,N_18936,N_19672);
and U20635 (N_20635,N_19765,N_19859);
and U20636 (N_20636,N_19028,N_18475);
or U20637 (N_20637,N_18220,N_18113);
or U20638 (N_20638,N_18614,N_19517);
nor U20639 (N_20639,N_18549,N_18126);
nand U20640 (N_20640,N_19853,N_19813);
and U20641 (N_20641,N_19283,N_18432);
or U20642 (N_20642,N_19035,N_18571);
or U20643 (N_20643,N_19554,N_19286);
nor U20644 (N_20644,N_18209,N_19030);
nor U20645 (N_20645,N_19746,N_19412);
nor U20646 (N_20646,N_19662,N_19063);
nand U20647 (N_20647,N_18039,N_19287);
and U20648 (N_20648,N_18950,N_19525);
nand U20649 (N_20649,N_19927,N_18885);
or U20650 (N_20650,N_18433,N_19002);
or U20651 (N_20651,N_19852,N_19696);
nor U20652 (N_20652,N_18435,N_18057);
nor U20653 (N_20653,N_18922,N_19405);
nand U20654 (N_20654,N_19368,N_18792);
nor U20655 (N_20655,N_18005,N_18557);
nand U20656 (N_20656,N_18447,N_18785);
nor U20657 (N_20657,N_18256,N_18246);
or U20658 (N_20658,N_19754,N_18942);
or U20659 (N_20659,N_19362,N_18719);
nand U20660 (N_20660,N_18398,N_18107);
and U20661 (N_20661,N_18730,N_18110);
or U20662 (N_20662,N_18394,N_18244);
nand U20663 (N_20663,N_18367,N_18531);
nor U20664 (N_20664,N_18986,N_19477);
or U20665 (N_20665,N_19500,N_18008);
and U20666 (N_20666,N_18425,N_19779);
or U20667 (N_20667,N_19401,N_19653);
or U20668 (N_20668,N_18239,N_18685);
or U20669 (N_20669,N_19420,N_18728);
or U20670 (N_20670,N_19951,N_19580);
or U20671 (N_20671,N_19590,N_19237);
or U20672 (N_20672,N_19725,N_18316);
and U20673 (N_20673,N_18778,N_18013);
nor U20674 (N_20674,N_18160,N_19367);
nand U20675 (N_20675,N_19381,N_18744);
nor U20676 (N_20676,N_18388,N_18060);
or U20677 (N_20677,N_19180,N_18456);
or U20678 (N_20678,N_19900,N_19536);
nand U20679 (N_20679,N_18981,N_18416);
and U20680 (N_20680,N_18281,N_18362);
or U20681 (N_20681,N_19386,N_19679);
or U20682 (N_20682,N_19791,N_19684);
nand U20683 (N_20683,N_18038,N_18200);
nand U20684 (N_20684,N_19830,N_18216);
nand U20685 (N_20685,N_18577,N_19860);
nand U20686 (N_20686,N_19334,N_18904);
nor U20687 (N_20687,N_18772,N_18888);
nand U20688 (N_20688,N_18444,N_19016);
or U20689 (N_20689,N_19834,N_19235);
and U20690 (N_20690,N_19873,N_19478);
or U20691 (N_20691,N_18029,N_18536);
and U20692 (N_20692,N_18148,N_18971);
or U20693 (N_20693,N_18453,N_18821);
nor U20694 (N_20694,N_18248,N_18613);
and U20695 (N_20695,N_18170,N_18563);
and U20696 (N_20696,N_19503,N_18044);
and U20697 (N_20697,N_19818,N_18738);
nand U20698 (N_20698,N_18899,N_18015);
nand U20699 (N_20699,N_18516,N_19122);
or U20700 (N_20700,N_19965,N_18422);
and U20701 (N_20701,N_19585,N_19446);
nand U20702 (N_20702,N_19895,N_19647);
nand U20703 (N_20703,N_18837,N_19297);
or U20704 (N_20704,N_18984,N_19354);
and U20705 (N_20705,N_19875,N_19132);
nand U20706 (N_20706,N_18497,N_19391);
or U20707 (N_20707,N_19170,N_19090);
nand U20708 (N_20708,N_18596,N_18666);
nand U20709 (N_20709,N_18253,N_19171);
or U20710 (N_20710,N_18086,N_18832);
and U20711 (N_20711,N_19373,N_19247);
and U20712 (N_20712,N_18024,N_18428);
or U20713 (N_20713,N_19595,N_18452);
or U20714 (N_20714,N_19113,N_18185);
nor U20715 (N_20715,N_19577,N_18640);
or U20716 (N_20716,N_19333,N_18667);
nor U20717 (N_20717,N_19996,N_18297);
nor U20718 (N_20718,N_19096,N_19722);
nand U20719 (N_20719,N_18269,N_18583);
or U20720 (N_20720,N_19760,N_18389);
nor U20721 (N_20721,N_18585,N_19569);
or U20722 (N_20722,N_18831,N_18958);
and U20723 (N_20723,N_18223,N_18341);
and U20724 (N_20724,N_19336,N_19532);
and U20725 (N_20725,N_18324,N_18399);
and U20726 (N_20726,N_19074,N_19288);
or U20727 (N_20727,N_18484,N_19637);
nand U20728 (N_20728,N_19734,N_18093);
nand U20729 (N_20729,N_18303,N_19042);
or U20730 (N_20730,N_19430,N_19502);
nor U20731 (N_20731,N_18046,N_19540);
nand U20732 (N_20732,N_19114,N_19496);
or U20733 (N_20733,N_19835,N_19162);
and U20734 (N_20734,N_18960,N_18589);
or U20735 (N_20735,N_18014,N_18412);
and U20736 (N_20736,N_19054,N_18815);
or U20737 (N_20737,N_19805,N_19359);
and U20738 (N_20738,N_19867,N_18198);
nor U20739 (N_20739,N_19495,N_18033);
and U20740 (N_20740,N_19017,N_18376);
or U20741 (N_20741,N_19187,N_19576);
nand U20742 (N_20742,N_18896,N_19762);
nand U20743 (N_20743,N_19692,N_19489);
or U20744 (N_20744,N_19198,N_19716);
nor U20745 (N_20745,N_18928,N_18700);
or U20746 (N_20746,N_19265,N_18569);
and U20747 (N_20747,N_18794,N_19526);
and U20748 (N_20748,N_18708,N_19432);
or U20749 (N_20749,N_19043,N_18777);
or U20750 (N_20750,N_19036,N_19556);
or U20751 (N_20751,N_18236,N_18508);
or U20752 (N_20752,N_18802,N_19280);
and U20753 (N_20753,N_19466,N_19726);
nand U20754 (N_20754,N_19026,N_18993);
nand U20755 (N_20755,N_19974,N_19459);
nor U20756 (N_20756,N_19085,N_18408);
or U20757 (N_20757,N_18781,N_19163);
or U20758 (N_20758,N_19793,N_19843);
and U20759 (N_20759,N_18462,N_19059);
and U20760 (N_20760,N_19646,N_18633);
and U20761 (N_20761,N_19380,N_18304);
nor U20762 (N_20762,N_18109,N_19591);
nand U20763 (N_20763,N_18112,N_19931);
or U20764 (N_20764,N_18307,N_18483);
xnor U20765 (N_20765,N_19037,N_18702);
nand U20766 (N_20766,N_19108,N_18956);
and U20767 (N_20767,N_18897,N_19934);
or U20768 (N_20768,N_18020,N_19850);
nand U20769 (N_20769,N_18923,N_19281);
or U20770 (N_20770,N_19426,N_19418);
and U20771 (N_20771,N_18387,N_19636);
and U20772 (N_20772,N_18804,N_18245);
nor U20773 (N_20773,N_19946,N_19563);
and U20774 (N_20774,N_19471,N_19820);
and U20775 (N_20775,N_18522,N_19848);
nor U20776 (N_20776,N_18693,N_18051);
or U20777 (N_20777,N_19642,N_19665);
or U20778 (N_20778,N_19327,N_19902);
nor U20779 (N_20779,N_18501,N_18716);
nand U20780 (N_20780,N_19594,N_19756);
or U20781 (N_20781,N_19289,N_18543);
or U20782 (N_20782,N_18525,N_19069);
or U20783 (N_20783,N_18822,N_18498);
nand U20784 (N_20784,N_19894,N_18515);
nand U20785 (N_20785,N_19964,N_18647);
nor U20786 (N_20786,N_19899,N_18995);
and U20787 (N_20787,N_18101,N_18940);
nor U20788 (N_20788,N_19735,N_19199);
and U20789 (N_20789,N_19109,N_19694);
nand U20790 (N_20790,N_19952,N_18266);
nor U20791 (N_20791,N_18913,N_19282);
nor U20792 (N_20792,N_18237,N_19257);
and U20793 (N_20793,N_19941,N_18587);
and U20794 (N_20794,N_19472,N_18883);
and U20795 (N_20795,N_18546,N_19910);
nand U20796 (N_20796,N_18009,N_18661);
and U20797 (N_20797,N_18074,N_18053);
nand U20798 (N_20798,N_18819,N_19457);
and U20799 (N_20799,N_18858,N_18149);
or U20800 (N_20800,N_19783,N_19111);
and U20801 (N_20801,N_18406,N_19708);
nand U20802 (N_20802,N_19596,N_18162);
or U20803 (N_20803,N_19541,N_18372);
nor U20804 (N_20804,N_19930,N_19697);
nand U20805 (N_20805,N_19011,N_18846);
nor U20806 (N_20806,N_19443,N_18375);
or U20807 (N_20807,N_19785,N_18856);
and U20808 (N_20808,N_19423,N_19944);
or U20809 (N_20809,N_18604,N_18759);
and U20810 (N_20810,N_19487,N_19009);
and U20811 (N_20811,N_18875,N_18235);
nor U20812 (N_20812,N_19583,N_18276);
nor U20813 (N_20813,N_18554,N_18145);
xnor U20814 (N_20814,N_18655,N_18551);
nand U20815 (N_20815,N_19166,N_19903);
xnor U20816 (N_20816,N_19123,N_18189);
and U20817 (N_20817,N_18691,N_18886);
and U20818 (N_20818,N_18999,N_19811);
nor U20819 (N_20819,N_19197,N_18368);
xor U20820 (N_20820,N_19925,N_18745);
nor U20821 (N_20821,N_19896,N_18091);
nor U20822 (N_20822,N_18187,N_18391);
or U20823 (N_20823,N_19355,N_19651);
nand U20824 (N_20824,N_18437,N_19184);
nor U20825 (N_20825,N_19715,N_18872);
xnor U20826 (N_20826,N_19370,N_19855);
nand U20827 (N_20827,N_19795,N_18114);
nor U20828 (N_20828,N_19683,N_19825);
nor U20829 (N_20829,N_18293,N_18077);
nand U20830 (N_20830,N_18513,N_18423);
nor U20831 (N_20831,N_19509,N_19909);
nor U20832 (N_20832,N_18139,N_19522);
and U20833 (N_20833,N_19098,N_19284);
or U20834 (N_20834,N_19613,N_19117);
or U20835 (N_20835,N_18898,N_18512);
or U20836 (N_20836,N_19511,N_18397);
nor U20837 (N_20837,N_18651,N_19761);
nand U20838 (N_20838,N_19598,N_19535);
and U20839 (N_20839,N_19986,N_18193);
or U20840 (N_20840,N_19616,N_19707);
or U20841 (N_20841,N_18458,N_19155);
nor U20842 (N_20842,N_19604,N_19717);
nor U20843 (N_20843,N_18671,N_18374);
or U20844 (N_20844,N_19095,N_18078);
and U20845 (N_20845,N_18225,N_19195);
or U20846 (N_20846,N_19505,N_19434);
nand U20847 (N_20847,N_18644,N_19796);
nand U20848 (N_20848,N_19484,N_18105);
nand U20849 (N_20849,N_19751,N_19817);
and U20850 (N_20850,N_19545,N_18576);
nand U20851 (N_20851,N_18402,N_18095);
or U20852 (N_20852,N_18218,N_19128);
nand U20853 (N_20853,N_18678,N_19273);
and U20854 (N_20854,N_19728,N_18283);
and U20855 (N_20855,N_18295,N_19822);
nor U20856 (N_20856,N_19898,N_19753);
and U20857 (N_20857,N_19608,N_19937);
nor U20858 (N_20858,N_19815,N_18407);
xnor U20859 (N_20859,N_19249,N_19652);
and U20860 (N_20860,N_19447,N_18900);
nor U20861 (N_20861,N_19121,N_18642);
nand U20862 (N_20862,N_19032,N_18947);
nand U20863 (N_20863,N_19688,N_19448);
nand U20864 (N_20864,N_18032,N_19402);
or U20865 (N_20865,N_19010,N_19112);
nor U20866 (N_20866,N_18711,N_19419);
or U20867 (N_20867,N_18848,N_18146);
or U20868 (N_20868,N_18565,N_19533);
nor U20869 (N_20869,N_19586,N_18278);
nand U20870 (N_20870,N_19507,N_19976);
nor U20871 (N_20871,N_18626,N_19648);
nor U20872 (N_20872,N_19729,N_19584);
nor U20873 (N_20873,N_19131,N_19638);
or U20874 (N_20874,N_18841,N_19192);
nor U20875 (N_20875,N_18941,N_19827);
or U20876 (N_20876,N_18186,N_19208);
nand U20877 (N_20877,N_18141,N_19216);
or U20878 (N_20878,N_19461,N_18935);
and U20879 (N_20879,N_19766,N_18555);
nor U20880 (N_20880,N_19231,N_18445);
nand U20881 (N_20881,N_19832,N_19206);
or U20882 (N_20882,N_18933,N_18327);
nand U20883 (N_20883,N_18786,N_19200);
nor U20884 (N_20884,N_19120,N_18545);
nand U20885 (N_20885,N_19940,N_19773);
nor U20886 (N_20886,N_18964,N_18991);
or U20887 (N_20887,N_18842,N_18356);
or U20888 (N_20888,N_19515,N_19300);
nand U20889 (N_20889,N_18382,N_18054);
nand U20890 (N_20890,N_18818,N_18688);
nor U20891 (N_20891,N_19539,N_18799);
nor U20892 (N_20892,N_19804,N_18867);
or U20893 (N_20893,N_18830,N_18891);
nand U20894 (N_20894,N_19671,N_19497);
nor U20895 (N_20895,N_19045,N_19196);
nand U20896 (N_20896,N_18957,N_19677);
nor U20897 (N_20897,N_18937,N_19524);
nor U20898 (N_20898,N_19346,N_19191);
or U20899 (N_20899,N_18176,N_18411);
and U20900 (N_20900,N_19778,N_18331);
nand U20901 (N_20901,N_19924,N_19544);
nor U20902 (N_20902,N_19706,N_19685);
or U20903 (N_20903,N_18874,N_19731);
nand U20904 (N_20904,N_19205,N_19270);
or U20905 (N_20905,N_19983,N_19730);
xnor U20906 (N_20906,N_18628,N_19066);
or U20907 (N_20907,N_19258,N_18466);
nand U20908 (N_20908,N_19371,N_18634);
nor U20909 (N_20909,N_18463,N_18965);
nand U20910 (N_20910,N_18067,N_19229);
xnor U20911 (N_20911,N_18972,N_19023);
and U20912 (N_20912,N_19807,N_19534);
nand U20913 (N_20913,N_19357,N_19891);
and U20914 (N_20914,N_19160,N_19474);
nor U20915 (N_20915,N_19416,N_19349);
nor U20916 (N_20916,N_18465,N_19890);
or U20917 (N_20917,N_18801,N_18599);
and U20918 (N_20918,N_18939,N_18175);
and U20919 (N_20919,N_19076,N_19599);
nand U20920 (N_20920,N_19561,N_18409);
xnor U20921 (N_20921,N_19587,N_19904);
nand U20922 (N_20922,N_19788,N_18172);
nor U20923 (N_20923,N_18769,N_18258);
and U20924 (N_20924,N_19593,N_18750);
and U20925 (N_20925,N_18696,N_19212);
nor U20926 (N_20926,N_19644,N_19404);
or U20927 (N_20927,N_18059,N_19885);
nand U20928 (N_20928,N_19872,N_19007);
nor U20929 (N_20929,N_19174,N_19922);
nand U20930 (N_20930,N_19100,N_18884);
nor U20931 (N_20931,N_19506,N_19831);
nand U20932 (N_20932,N_19233,N_18636);
nand U20933 (N_20933,N_18681,N_18507);
and U20934 (N_20934,N_18003,N_18810);
nand U20935 (N_20935,N_19978,N_18675);
or U20936 (N_20936,N_19786,N_19311);
or U20937 (N_20937,N_19313,N_18158);
nor U20938 (N_20938,N_19879,N_18865);
nor U20939 (N_20939,N_18089,N_19228);
nor U20940 (N_20940,N_19044,N_18893);
and U20941 (N_20941,N_18155,N_19400);
or U20942 (N_20942,N_19415,N_18690);
or U20943 (N_20943,N_18364,N_19628);
or U20944 (N_20944,N_18250,N_19324);
or U20945 (N_20945,N_19863,N_19188);
nor U20946 (N_20946,N_19468,N_18994);
or U20947 (N_20947,N_19744,N_18291);
nor U20948 (N_20948,N_18300,N_19014);
nor U20949 (N_20949,N_18825,N_18517);
and U20950 (N_20950,N_19377,N_19064);
and U20951 (N_20951,N_18429,N_18989);
or U20952 (N_20952,N_18349,N_18025);
nand U20953 (N_20953,N_18731,N_18142);
nor U20954 (N_20954,N_19301,N_18535);
nand U20955 (N_20955,N_18868,N_19149);
nor U20956 (N_20956,N_19774,N_18288);
or U20957 (N_20957,N_18637,N_19475);
nand U20958 (N_20958,N_18217,N_18849);
nor U20959 (N_20959,N_19183,N_19451);
or U20960 (N_20960,N_19285,N_18241);
or U20961 (N_20961,N_18366,N_19981);
and U20962 (N_20962,N_19816,N_19241);
nand U20963 (N_20963,N_19136,N_18322);
nand U20964 (N_20964,N_19319,N_19034);
nand U20965 (N_20965,N_18771,N_19607);
nor U20966 (N_20966,N_19866,N_18242);
and U20967 (N_20967,N_18791,N_18987);
or U20968 (N_20968,N_19105,N_18979);
nand U20969 (N_20969,N_18855,N_18182);
or U20970 (N_20970,N_19040,N_18436);
nand U20971 (N_20971,N_19787,N_18570);
and U20972 (N_20972,N_18108,N_18699);
nand U20973 (N_20973,N_18043,N_18294);
nor U20974 (N_20974,N_18864,N_18088);
nor U20975 (N_20975,N_19803,N_18011);
nand U20976 (N_20976,N_19267,N_18401);
nor U20977 (N_20977,N_19013,N_18491);
and U20978 (N_20978,N_18800,N_19068);
xor U20979 (N_20979,N_18703,N_18082);
nor U20980 (N_20980,N_18130,N_18201);
nand U20981 (N_20981,N_19658,N_19374);
nor U20982 (N_20982,N_18606,N_19038);
nand U20983 (N_20983,N_19172,N_18350);
or U20984 (N_20984,N_18338,N_18764);
or U20985 (N_20985,N_18127,N_18153);
or U20986 (N_20986,N_18378,N_19512);
nand U20987 (N_20987,N_19917,N_19588);
xnor U20988 (N_20988,N_18627,N_19215);
nor U20989 (N_20989,N_18315,N_18558);
nor U20990 (N_20990,N_18100,N_19999);
nor U20991 (N_20991,N_19110,N_18363);
nor U20992 (N_20992,N_18152,N_19654);
nor U20993 (N_20993,N_19393,N_19631);
nor U20994 (N_20994,N_19555,N_19341);
nor U20995 (N_20995,N_19129,N_18479);
or U20996 (N_20996,N_19151,N_18179);
or U20997 (N_20997,N_19441,N_18705);
and U20998 (N_20998,N_19139,N_19185);
nand U20999 (N_20999,N_18431,N_19127);
nand U21000 (N_21000,N_19212,N_19361);
and U21001 (N_21001,N_18937,N_18713);
or U21002 (N_21002,N_19051,N_19016);
or U21003 (N_21003,N_18132,N_19710);
xnor U21004 (N_21004,N_19719,N_18013);
nor U21005 (N_21005,N_19019,N_18005);
and U21006 (N_21006,N_19307,N_19105);
nor U21007 (N_21007,N_18224,N_19022);
nor U21008 (N_21008,N_19223,N_19404);
or U21009 (N_21009,N_18994,N_18163);
or U21010 (N_21010,N_18890,N_18882);
nand U21011 (N_21011,N_19113,N_19536);
xor U21012 (N_21012,N_18606,N_19843);
nand U21013 (N_21013,N_18883,N_18435);
or U21014 (N_21014,N_19283,N_18731);
and U21015 (N_21015,N_19107,N_19199);
and U21016 (N_21016,N_19315,N_19100);
nand U21017 (N_21017,N_19949,N_19341);
or U21018 (N_21018,N_19849,N_18182);
nor U21019 (N_21019,N_18792,N_18540);
and U21020 (N_21020,N_19737,N_19856);
and U21021 (N_21021,N_19488,N_18068);
nand U21022 (N_21022,N_18157,N_19822);
or U21023 (N_21023,N_19907,N_19031);
and U21024 (N_21024,N_18874,N_18158);
nor U21025 (N_21025,N_18733,N_19731);
nand U21026 (N_21026,N_18945,N_19305);
nand U21027 (N_21027,N_19819,N_18426);
nor U21028 (N_21028,N_18436,N_19022);
nand U21029 (N_21029,N_18341,N_19396);
and U21030 (N_21030,N_19445,N_19733);
nor U21031 (N_21031,N_19519,N_19461);
or U21032 (N_21032,N_18613,N_19290);
and U21033 (N_21033,N_19295,N_19047);
nand U21034 (N_21034,N_19671,N_18836);
nand U21035 (N_21035,N_19248,N_18647);
and U21036 (N_21036,N_18578,N_19362);
and U21037 (N_21037,N_18028,N_19988);
or U21038 (N_21038,N_18695,N_18834);
or U21039 (N_21039,N_19305,N_19470);
nand U21040 (N_21040,N_19862,N_19254);
nor U21041 (N_21041,N_18041,N_19477);
or U21042 (N_21042,N_19992,N_18016);
or U21043 (N_21043,N_19347,N_18298);
or U21044 (N_21044,N_19065,N_19534);
or U21045 (N_21045,N_18782,N_18490);
nor U21046 (N_21046,N_18943,N_19104);
nor U21047 (N_21047,N_19756,N_19531);
or U21048 (N_21048,N_19412,N_19724);
nor U21049 (N_21049,N_18219,N_19191);
or U21050 (N_21050,N_19019,N_18114);
nand U21051 (N_21051,N_18822,N_19964);
or U21052 (N_21052,N_19872,N_18170);
and U21053 (N_21053,N_18245,N_18199);
nand U21054 (N_21054,N_19697,N_18653);
nor U21055 (N_21055,N_19830,N_18900);
nand U21056 (N_21056,N_18956,N_18663);
and U21057 (N_21057,N_19651,N_19810);
or U21058 (N_21058,N_18946,N_19733);
nand U21059 (N_21059,N_19943,N_19908);
nand U21060 (N_21060,N_19219,N_19735);
or U21061 (N_21061,N_19007,N_19537);
or U21062 (N_21062,N_18831,N_18490);
or U21063 (N_21063,N_18041,N_19072);
nand U21064 (N_21064,N_18993,N_18816);
and U21065 (N_21065,N_19822,N_18992);
nand U21066 (N_21066,N_19350,N_18270);
and U21067 (N_21067,N_18434,N_18650);
nor U21068 (N_21068,N_19037,N_18777);
nand U21069 (N_21069,N_18254,N_19674);
and U21070 (N_21070,N_19480,N_19105);
or U21071 (N_21071,N_18333,N_19294);
nor U21072 (N_21072,N_18665,N_18151);
nor U21073 (N_21073,N_19826,N_18212);
nor U21074 (N_21074,N_19195,N_18188);
and U21075 (N_21075,N_18193,N_19322);
and U21076 (N_21076,N_19070,N_19105);
and U21077 (N_21077,N_19107,N_19348);
nor U21078 (N_21078,N_18135,N_18058);
or U21079 (N_21079,N_18568,N_19945);
and U21080 (N_21080,N_18177,N_18343);
nor U21081 (N_21081,N_19233,N_18583);
or U21082 (N_21082,N_19540,N_19521);
and U21083 (N_21083,N_18086,N_19254);
xnor U21084 (N_21084,N_18433,N_19683);
or U21085 (N_21085,N_18695,N_19323);
nand U21086 (N_21086,N_18447,N_19945);
nand U21087 (N_21087,N_18485,N_18873);
nand U21088 (N_21088,N_19381,N_19097);
and U21089 (N_21089,N_19089,N_18708);
or U21090 (N_21090,N_19267,N_19248);
nor U21091 (N_21091,N_19798,N_19376);
and U21092 (N_21092,N_19011,N_18433);
or U21093 (N_21093,N_18408,N_19556);
and U21094 (N_21094,N_19074,N_18948);
nor U21095 (N_21095,N_18706,N_18525);
and U21096 (N_21096,N_18922,N_19354);
and U21097 (N_21097,N_19701,N_18731);
or U21098 (N_21098,N_18815,N_19301);
and U21099 (N_21099,N_19624,N_18414);
nand U21100 (N_21100,N_18793,N_19614);
nand U21101 (N_21101,N_19804,N_18037);
or U21102 (N_21102,N_19216,N_18190);
nor U21103 (N_21103,N_19495,N_18336);
and U21104 (N_21104,N_19857,N_18542);
or U21105 (N_21105,N_18311,N_18927);
or U21106 (N_21106,N_19937,N_19561);
nand U21107 (N_21107,N_19793,N_19081);
nor U21108 (N_21108,N_19470,N_18085);
or U21109 (N_21109,N_18524,N_19539);
or U21110 (N_21110,N_19011,N_18600);
and U21111 (N_21111,N_19858,N_18935);
nand U21112 (N_21112,N_19366,N_19285);
nand U21113 (N_21113,N_18140,N_18057);
and U21114 (N_21114,N_18402,N_19164);
and U21115 (N_21115,N_18857,N_18482);
nor U21116 (N_21116,N_18560,N_19153);
nor U21117 (N_21117,N_18574,N_19153);
and U21118 (N_21118,N_18937,N_19707);
nor U21119 (N_21119,N_18802,N_18414);
nor U21120 (N_21120,N_19062,N_19414);
or U21121 (N_21121,N_18896,N_18351);
xnor U21122 (N_21122,N_18539,N_18198);
or U21123 (N_21123,N_18971,N_19849);
nor U21124 (N_21124,N_18627,N_18021);
or U21125 (N_21125,N_18075,N_19497);
or U21126 (N_21126,N_19060,N_18549);
and U21127 (N_21127,N_18701,N_18581);
and U21128 (N_21128,N_19798,N_19628);
nor U21129 (N_21129,N_19056,N_18111);
or U21130 (N_21130,N_18084,N_19737);
or U21131 (N_21131,N_19404,N_19959);
or U21132 (N_21132,N_18296,N_18967);
or U21133 (N_21133,N_19428,N_19061);
and U21134 (N_21134,N_19592,N_19016);
or U21135 (N_21135,N_18135,N_18392);
and U21136 (N_21136,N_19478,N_19355);
and U21137 (N_21137,N_19291,N_19686);
nand U21138 (N_21138,N_18826,N_18623);
or U21139 (N_21139,N_19368,N_18901);
nor U21140 (N_21140,N_19372,N_18034);
or U21141 (N_21141,N_19021,N_18392);
or U21142 (N_21142,N_18078,N_18457);
or U21143 (N_21143,N_18700,N_18818);
or U21144 (N_21144,N_19508,N_18935);
nand U21145 (N_21145,N_19576,N_19444);
nand U21146 (N_21146,N_19619,N_18471);
nand U21147 (N_21147,N_18625,N_18020);
and U21148 (N_21148,N_18969,N_19055);
nor U21149 (N_21149,N_18772,N_19100);
nand U21150 (N_21150,N_19628,N_19725);
and U21151 (N_21151,N_18159,N_18555);
and U21152 (N_21152,N_18548,N_19246);
and U21153 (N_21153,N_18893,N_19469);
and U21154 (N_21154,N_19550,N_18186);
nand U21155 (N_21155,N_18687,N_19030);
nor U21156 (N_21156,N_18500,N_18685);
nor U21157 (N_21157,N_18768,N_18423);
nand U21158 (N_21158,N_19725,N_19635);
nand U21159 (N_21159,N_19434,N_18264);
or U21160 (N_21160,N_18509,N_19736);
nor U21161 (N_21161,N_18241,N_18479);
and U21162 (N_21162,N_19672,N_19846);
nor U21163 (N_21163,N_19561,N_19770);
and U21164 (N_21164,N_18223,N_18729);
nor U21165 (N_21165,N_19729,N_19677);
nand U21166 (N_21166,N_18304,N_18273);
and U21167 (N_21167,N_18584,N_18513);
nand U21168 (N_21168,N_18591,N_18691);
nand U21169 (N_21169,N_19488,N_19585);
nor U21170 (N_21170,N_19967,N_18028);
and U21171 (N_21171,N_19567,N_18107);
or U21172 (N_21172,N_18948,N_18609);
or U21173 (N_21173,N_18779,N_18210);
or U21174 (N_21174,N_18600,N_19246);
or U21175 (N_21175,N_19544,N_19070);
nand U21176 (N_21176,N_19490,N_19216);
or U21177 (N_21177,N_18304,N_19355);
nor U21178 (N_21178,N_19562,N_18766);
or U21179 (N_21179,N_18966,N_19502);
and U21180 (N_21180,N_18970,N_18000);
or U21181 (N_21181,N_18146,N_18291);
or U21182 (N_21182,N_19595,N_19046);
nor U21183 (N_21183,N_18512,N_19485);
and U21184 (N_21184,N_19661,N_18892);
nand U21185 (N_21185,N_18835,N_19818);
or U21186 (N_21186,N_18945,N_19001);
nand U21187 (N_21187,N_18346,N_19099);
or U21188 (N_21188,N_19317,N_19471);
and U21189 (N_21189,N_18409,N_18117);
nor U21190 (N_21190,N_19841,N_18064);
and U21191 (N_21191,N_18179,N_19842);
and U21192 (N_21192,N_18362,N_19715);
and U21193 (N_21193,N_19263,N_19668);
and U21194 (N_21194,N_18918,N_18632);
or U21195 (N_21195,N_18080,N_19608);
and U21196 (N_21196,N_18228,N_19766);
and U21197 (N_21197,N_19231,N_18344);
nor U21198 (N_21198,N_19000,N_19140);
and U21199 (N_21199,N_18324,N_18474);
nor U21200 (N_21200,N_18119,N_18929);
nand U21201 (N_21201,N_19260,N_19815);
and U21202 (N_21202,N_18146,N_18004);
nor U21203 (N_21203,N_19671,N_18000);
nand U21204 (N_21204,N_18423,N_18704);
and U21205 (N_21205,N_19737,N_18436);
nand U21206 (N_21206,N_18231,N_18095);
nor U21207 (N_21207,N_18222,N_19149);
nor U21208 (N_21208,N_18616,N_18711);
nand U21209 (N_21209,N_18960,N_18426);
and U21210 (N_21210,N_18860,N_19259);
or U21211 (N_21211,N_18745,N_18078);
nor U21212 (N_21212,N_18220,N_19797);
nand U21213 (N_21213,N_19699,N_19022);
and U21214 (N_21214,N_19260,N_18254);
nand U21215 (N_21215,N_19408,N_19018);
nor U21216 (N_21216,N_18805,N_19606);
nand U21217 (N_21217,N_18417,N_19922);
xor U21218 (N_21218,N_19462,N_18225);
nor U21219 (N_21219,N_19637,N_18970);
or U21220 (N_21220,N_19045,N_19355);
nand U21221 (N_21221,N_19128,N_19104);
or U21222 (N_21222,N_18604,N_18693);
nand U21223 (N_21223,N_19490,N_19752);
nor U21224 (N_21224,N_19181,N_18077);
or U21225 (N_21225,N_18356,N_18733);
xor U21226 (N_21226,N_19099,N_19197);
nand U21227 (N_21227,N_18246,N_18543);
nand U21228 (N_21228,N_18352,N_18024);
nor U21229 (N_21229,N_18337,N_18842);
nand U21230 (N_21230,N_19167,N_18279);
nand U21231 (N_21231,N_18504,N_18274);
nand U21232 (N_21232,N_18315,N_18322);
or U21233 (N_21233,N_19676,N_19207);
nor U21234 (N_21234,N_18659,N_18133);
and U21235 (N_21235,N_18164,N_19471);
nand U21236 (N_21236,N_19310,N_18086);
or U21237 (N_21237,N_18501,N_19879);
nor U21238 (N_21238,N_18193,N_19657);
nand U21239 (N_21239,N_18307,N_19082);
and U21240 (N_21240,N_18663,N_18603);
nand U21241 (N_21241,N_19470,N_19769);
or U21242 (N_21242,N_18562,N_19076);
xor U21243 (N_21243,N_18455,N_19157);
nor U21244 (N_21244,N_18527,N_19650);
or U21245 (N_21245,N_19682,N_19157);
and U21246 (N_21246,N_18347,N_19690);
or U21247 (N_21247,N_19915,N_19133);
nand U21248 (N_21248,N_18073,N_19287);
or U21249 (N_21249,N_18477,N_19080);
nor U21250 (N_21250,N_18877,N_18835);
or U21251 (N_21251,N_19398,N_18449);
nand U21252 (N_21252,N_19914,N_18548);
and U21253 (N_21253,N_19941,N_18455);
or U21254 (N_21254,N_19583,N_19468);
nand U21255 (N_21255,N_19871,N_19850);
nor U21256 (N_21256,N_18747,N_18462);
nor U21257 (N_21257,N_19716,N_19986);
nor U21258 (N_21258,N_18897,N_19543);
nand U21259 (N_21259,N_19961,N_19669);
and U21260 (N_21260,N_19491,N_19081);
nand U21261 (N_21261,N_19554,N_19262);
nor U21262 (N_21262,N_18939,N_19868);
or U21263 (N_21263,N_19255,N_19680);
or U21264 (N_21264,N_19922,N_18497);
nand U21265 (N_21265,N_19603,N_18577);
and U21266 (N_21266,N_18448,N_18058);
and U21267 (N_21267,N_18193,N_18952);
nor U21268 (N_21268,N_18808,N_19553);
or U21269 (N_21269,N_18607,N_19046);
xor U21270 (N_21270,N_19642,N_18420);
nor U21271 (N_21271,N_18804,N_19799);
or U21272 (N_21272,N_18565,N_19723);
nand U21273 (N_21273,N_19130,N_19182);
nor U21274 (N_21274,N_18957,N_18943);
nand U21275 (N_21275,N_19999,N_18766);
nand U21276 (N_21276,N_19919,N_18173);
nor U21277 (N_21277,N_19125,N_18388);
nand U21278 (N_21278,N_18729,N_19588);
nand U21279 (N_21279,N_19080,N_19219);
nor U21280 (N_21280,N_18993,N_18216);
or U21281 (N_21281,N_19226,N_19476);
nor U21282 (N_21282,N_19153,N_18106);
and U21283 (N_21283,N_18240,N_18541);
nand U21284 (N_21284,N_19838,N_18908);
or U21285 (N_21285,N_18051,N_19081);
or U21286 (N_21286,N_19003,N_18566);
and U21287 (N_21287,N_19581,N_18976);
nand U21288 (N_21288,N_19824,N_18555);
nand U21289 (N_21289,N_19748,N_18088);
nor U21290 (N_21290,N_18776,N_18833);
nand U21291 (N_21291,N_19006,N_19426);
nor U21292 (N_21292,N_18402,N_18089);
or U21293 (N_21293,N_19167,N_19411);
nor U21294 (N_21294,N_19958,N_19894);
nor U21295 (N_21295,N_19125,N_19108);
and U21296 (N_21296,N_19635,N_19237);
or U21297 (N_21297,N_18129,N_19094);
nand U21298 (N_21298,N_18126,N_18873);
and U21299 (N_21299,N_18350,N_18743);
or U21300 (N_21300,N_19399,N_19715);
nor U21301 (N_21301,N_19282,N_18908);
and U21302 (N_21302,N_18622,N_18183);
nor U21303 (N_21303,N_19004,N_18025);
nand U21304 (N_21304,N_19372,N_19094);
nor U21305 (N_21305,N_18201,N_19717);
nand U21306 (N_21306,N_18857,N_18293);
nor U21307 (N_21307,N_18695,N_18120);
xor U21308 (N_21308,N_19538,N_19959);
nor U21309 (N_21309,N_19828,N_18372);
and U21310 (N_21310,N_19093,N_18820);
nor U21311 (N_21311,N_19636,N_19092);
nor U21312 (N_21312,N_19371,N_19663);
nand U21313 (N_21313,N_18350,N_18346);
or U21314 (N_21314,N_18708,N_19236);
or U21315 (N_21315,N_18512,N_18656);
xnor U21316 (N_21316,N_18693,N_19518);
nor U21317 (N_21317,N_18671,N_19501);
or U21318 (N_21318,N_19524,N_19451);
or U21319 (N_21319,N_18007,N_19970);
or U21320 (N_21320,N_18017,N_19401);
nor U21321 (N_21321,N_19123,N_18452);
nor U21322 (N_21322,N_19039,N_18770);
or U21323 (N_21323,N_18215,N_18154);
nor U21324 (N_21324,N_19089,N_18328);
or U21325 (N_21325,N_19752,N_18425);
and U21326 (N_21326,N_19491,N_19846);
nor U21327 (N_21327,N_19985,N_18790);
nor U21328 (N_21328,N_18696,N_19771);
xor U21329 (N_21329,N_19300,N_19989);
nor U21330 (N_21330,N_19232,N_18137);
and U21331 (N_21331,N_18649,N_19447);
nor U21332 (N_21332,N_19981,N_19740);
or U21333 (N_21333,N_19944,N_18988);
and U21334 (N_21334,N_18202,N_19722);
nand U21335 (N_21335,N_18799,N_19013);
nand U21336 (N_21336,N_18275,N_19694);
or U21337 (N_21337,N_19663,N_18951);
and U21338 (N_21338,N_18754,N_19286);
nand U21339 (N_21339,N_19237,N_18315);
or U21340 (N_21340,N_19735,N_18659);
nand U21341 (N_21341,N_19797,N_18639);
and U21342 (N_21342,N_19704,N_19430);
or U21343 (N_21343,N_18299,N_18291);
nor U21344 (N_21344,N_18815,N_19308);
nor U21345 (N_21345,N_19209,N_19071);
nor U21346 (N_21346,N_19918,N_19613);
nor U21347 (N_21347,N_19753,N_18987);
or U21348 (N_21348,N_19150,N_18706);
or U21349 (N_21349,N_19853,N_18695);
nor U21350 (N_21350,N_19026,N_18648);
nor U21351 (N_21351,N_19755,N_19090);
or U21352 (N_21352,N_19585,N_18885);
nor U21353 (N_21353,N_18743,N_19415);
and U21354 (N_21354,N_18054,N_19300);
nor U21355 (N_21355,N_19164,N_19104);
or U21356 (N_21356,N_19030,N_19492);
or U21357 (N_21357,N_19723,N_19342);
nand U21358 (N_21358,N_18351,N_19592);
nor U21359 (N_21359,N_19052,N_18852);
or U21360 (N_21360,N_18321,N_19059);
and U21361 (N_21361,N_19733,N_18502);
nand U21362 (N_21362,N_18493,N_19486);
and U21363 (N_21363,N_19681,N_18420);
xnor U21364 (N_21364,N_19244,N_18764);
nor U21365 (N_21365,N_19394,N_18752);
nor U21366 (N_21366,N_19663,N_18258);
or U21367 (N_21367,N_19409,N_18864);
nor U21368 (N_21368,N_19576,N_19262);
nand U21369 (N_21369,N_19610,N_19462);
or U21370 (N_21370,N_18384,N_18110);
nor U21371 (N_21371,N_18664,N_19169);
or U21372 (N_21372,N_18235,N_18574);
nor U21373 (N_21373,N_19728,N_19174);
or U21374 (N_21374,N_18952,N_19001);
and U21375 (N_21375,N_18517,N_19814);
nand U21376 (N_21376,N_18247,N_19675);
and U21377 (N_21377,N_18956,N_18086);
or U21378 (N_21378,N_18351,N_19075);
or U21379 (N_21379,N_18662,N_18367);
nand U21380 (N_21380,N_18581,N_18792);
nor U21381 (N_21381,N_18333,N_19711);
or U21382 (N_21382,N_19379,N_19181);
and U21383 (N_21383,N_18000,N_18509);
nand U21384 (N_21384,N_19573,N_19314);
and U21385 (N_21385,N_18547,N_18303);
nor U21386 (N_21386,N_19498,N_18617);
or U21387 (N_21387,N_19536,N_18240);
and U21388 (N_21388,N_19983,N_19305);
nand U21389 (N_21389,N_18400,N_19893);
and U21390 (N_21390,N_18735,N_19119);
nand U21391 (N_21391,N_18343,N_18985);
nor U21392 (N_21392,N_19428,N_18123);
or U21393 (N_21393,N_19564,N_18507);
nand U21394 (N_21394,N_19729,N_19825);
nor U21395 (N_21395,N_19076,N_18880);
and U21396 (N_21396,N_18031,N_18886);
nand U21397 (N_21397,N_19484,N_18390);
nor U21398 (N_21398,N_19167,N_18217);
or U21399 (N_21399,N_19330,N_18394);
or U21400 (N_21400,N_19846,N_19514);
or U21401 (N_21401,N_19799,N_18509);
nor U21402 (N_21402,N_19686,N_19317);
nand U21403 (N_21403,N_18919,N_19069);
or U21404 (N_21404,N_18334,N_18457);
nor U21405 (N_21405,N_19034,N_19968);
or U21406 (N_21406,N_18662,N_19327);
nand U21407 (N_21407,N_18342,N_18577);
nand U21408 (N_21408,N_19744,N_18265);
nor U21409 (N_21409,N_18480,N_19397);
nand U21410 (N_21410,N_19638,N_19166);
nor U21411 (N_21411,N_19139,N_18410);
nor U21412 (N_21412,N_18831,N_18222);
nor U21413 (N_21413,N_19809,N_19284);
or U21414 (N_21414,N_18907,N_18512);
and U21415 (N_21415,N_19368,N_18208);
and U21416 (N_21416,N_19680,N_18332);
nor U21417 (N_21417,N_19506,N_18109);
nand U21418 (N_21418,N_19052,N_19352);
and U21419 (N_21419,N_18902,N_18797);
and U21420 (N_21420,N_18133,N_18306);
nand U21421 (N_21421,N_19722,N_18378);
or U21422 (N_21422,N_18410,N_19499);
nor U21423 (N_21423,N_19550,N_19522);
or U21424 (N_21424,N_19007,N_19094);
nand U21425 (N_21425,N_19147,N_18842);
nand U21426 (N_21426,N_19961,N_18915);
nand U21427 (N_21427,N_19530,N_18479);
nand U21428 (N_21428,N_19850,N_18173);
nor U21429 (N_21429,N_18075,N_19930);
nand U21430 (N_21430,N_19876,N_19674);
nand U21431 (N_21431,N_18610,N_19529);
nor U21432 (N_21432,N_19973,N_19329);
and U21433 (N_21433,N_18865,N_18747);
and U21434 (N_21434,N_19022,N_18598);
or U21435 (N_21435,N_19006,N_19464);
and U21436 (N_21436,N_19432,N_18518);
nand U21437 (N_21437,N_18905,N_19683);
nand U21438 (N_21438,N_19454,N_19912);
nand U21439 (N_21439,N_19257,N_18328);
nand U21440 (N_21440,N_19210,N_19775);
or U21441 (N_21441,N_19807,N_19765);
and U21442 (N_21442,N_18309,N_19576);
nor U21443 (N_21443,N_18526,N_18450);
and U21444 (N_21444,N_19434,N_19678);
and U21445 (N_21445,N_18872,N_18370);
or U21446 (N_21446,N_18891,N_19535);
and U21447 (N_21447,N_18956,N_19183);
and U21448 (N_21448,N_19338,N_19388);
nand U21449 (N_21449,N_18033,N_18898);
and U21450 (N_21450,N_19507,N_19844);
nor U21451 (N_21451,N_18490,N_19660);
or U21452 (N_21452,N_19661,N_18840);
nand U21453 (N_21453,N_18281,N_18452);
and U21454 (N_21454,N_19062,N_19238);
or U21455 (N_21455,N_19083,N_19810);
nor U21456 (N_21456,N_19161,N_18837);
or U21457 (N_21457,N_19025,N_19820);
nand U21458 (N_21458,N_19603,N_19322);
nor U21459 (N_21459,N_18807,N_18263);
nand U21460 (N_21460,N_19349,N_19396);
nor U21461 (N_21461,N_19088,N_18214);
nand U21462 (N_21462,N_18481,N_19056);
nand U21463 (N_21463,N_19593,N_19524);
nor U21464 (N_21464,N_18665,N_18947);
or U21465 (N_21465,N_18354,N_19783);
nor U21466 (N_21466,N_18277,N_18749);
nand U21467 (N_21467,N_18629,N_18887);
nand U21468 (N_21468,N_19970,N_19288);
nand U21469 (N_21469,N_18571,N_19927);
nor U21470 (N_21470,N_18452,N_18999);
and U21471 (N_21471,N_18683,N_19800);
nor U21472 (N_21472,N_19835,N_19418);
and U21473 (N_21473,N_19342,N_18417);
or U21474 (N_21474,N_19705,N_18288);
nor U21475 (N_21475,N_19587,N_18232);
nand U21476 (N_21476,N_19610,N_19381);
nand U21477 (N_21477,N_18222,N_18570);
nand U21478 (N_21478,N_18564,N_18411);
and U21479 (N_21479,N_18291,N_19325);
nand U21480 (N_21480,N_19245,N_18761);
and U21481 (N_21481,N_19362,N_18183);
nand U21482 (N_21482,N_18374,N_19806);
nand U21483 (N_21483,N_18923,N_19884);
or U21484 (N_21484,N_19718,N_19333);
nand U21485 (N_21485,N_18604,N_19027);
and U21486 (N_21486,N_19788,N_19766);
and U21487 (N_21487,N_18509,N_19317);
or U21488 (N_21488,N_18244,N_19472);
or U21489 (N_21489,N_19316,N_18148);
and U21490 (N_21490,N_18497,N_18576);
nand U21491 (N_21491,N_19835,N_19872);
or U21492 (N_21492,N_18381,N_19818);
nor U21493 (N_21493,N_19977,N_19065);
nor U21494 (N_21494,N_19958,N_18932);
nor U21495 (N_21495,N_19860,N_19034);
nand U21496 (N_21496,N_19653,N_19587);
nor U21497 (N_21497,N_18426,N_18357);
or U21498 (N_21498,N_18881,N_18547);
or U21499 (N_21499,N_19406,N_18025);
nor U21500 (N_21500,N_19862,N_18823);
nor U21501 (N_21501,N_19372,N_19384);
or U21502 (N_21502,N_19643,N_19504);
nand U21503 (N_21503,N_18826,N_19600);
and U21504 (N_21504,N_19351,N_18094);
or U21505 (N_21505,N_18576,N_18031);
nor U21506 (N_21506,N_19149,N_19054);
or U21507 (N_21507,N_18412,N_18537);
nor U21508 (N_21508,N_19303,N_19445);
nand U21509 (N_21509,N_19147,N_19090);
nand U21510 (N_21510,N_18581,N_19228);
nor U21511 (N_21511,N_19722,N_18563);
or U21512 (N_21512,N_18054,N_19257);
or U21513 (N_21513,N_18814,N_18742);
nor U21514 (N_21514,N_19146,N_19631);
nor U21515 (N_21515,N_19233,N_18960);
xor U21516 (N_21516,N_18351,N_18331);
nor U21517 (N_21517,N_19257,N_18156);
nand U21518 (N_21518,N_18880,N_19711);
and U21519 (N_21519,N_19096,N_19959);
nor U21520 (N_21520,N_19886,N_19625);
or U21521 (N_21521,N_19640,N_19375);
and U21522 (N_21522,N_19270,N_18498);
and U21523 (N_21523,N_18227,N_19243);
and U21524 (N_21524,N_19740,N_19240);
or U21525 (N_21525,N_19252,N_18805);
or U21526 (N_21526,N_19857,N_19373);
nor U21527 (N_21527,N_18303,N_18187);
or U21528 (N_21528,N_18505,N_19558);
and U21529 (N_21529,N_18545,N_18729);
nor U21530 (N_21530,N_18613,N_19529);
nand U21531 (N_21531,N_18049,N_18878);
nor U21532 (N_21532,N_18615,N_19740);
nand U21533 (N_21533,N_18674,N_19652);
and U21534 (N_21534,N_18829,N_18739);
nand U21535 (N_21535,N_19446,N_19760);
nand U21536 (N_21536,N_19490,N_19260);
nand U21537 (N_21537,N_19544,N_19151);
and U21538 (N_21538,N_19086,N_18768);
or U21539 (N_21539,N_19064,N_19756);
or U21540 (N_21540,N_19245,N_19088);
nand U21541 (N_21541,N_19215,N_19467);
nand U21542 (N_21542,N_19126,N_18858);
and U21543 (N_21543,N_18678,N_19245);
or U21544 (N_21544,N_19832,N_19783);
and U21545 (N_21545,N_19323,N_18756);
or U21546 (N_21546,N_19783,N_19515);
nor U21547 (N_21547,N_18994,N_19401);
nor U21548 (N_21548,N_18818,N_18617);
nor U21549 (N_21549,N_19433,N_19181);
and U21550 (N_21550,N_18382,N_18614);
and U21551 (N_21551,N_18861,N_19358);
or U21552 (N_21552,N_19695,N_18844);
nand U21553 (N_21553,N_19356,N_19674);
nor U21554 (N_21554,N_18541,N_19903);
or U21555 (N_21555,N_18202,N_18132);
nand U21556 (N_21556,N_19277,N_19622);
nand U21557 (N_21557,N_19370,N_18530);
nand U21558 (N_21558,N_19815,N_18491);
nor U21559 (N_21559,N_19100,N_18408);
nand U21560 (N_21560,N_18477,N_19814);
or U21561 (N_21561,N_19961,N_18465);
or U21562 (N_21562,N_18156,N_19525);
and U21563 (N_21563,N_19107,N_18024);
nand U21564 (N_21564,N_19170,N_19753);
and U21565 (N_21565,N_19509,N_18236);
or U21566 (N_21566,N_19851,N_18873);
or U21567 (N_21567,N_18639,N_19737);
nor U21568 (N_21568,N_19862,N_19228);
nor U21569 (N_21569,N_19646,N_18367);
nor U21570 (N_21570,N_19737,N_19993);
or U21571 (N_21571,N_19441,N_19551);
and U21572 (N_21572,N_18824,N_18929);
or U21573 (N_21573,N_19051,N_18251);
and U21574 (N_21574,N_19837,N_18004);
xor U21575 (N_21575,N_19550,N_18323);
nand U21576 (N_21576,N_19449,N_18227);
nand U21577 (N_21577,N_19856,N_19878);
and U21578 (N_21578,N_18114,N_18627);
nor U21579 (N_21579,N_19897,N_19503);
and U21580 (N_21580,N_18366,N_19301);
nor U21581 (N_21581,N_18488,N_19395);
nand U21582 (N_21582,N_19795,N_18151);
nor U21583 (N_21583,N_19050,N_18399);
nor U21584 (N_21584,N_19457,N_19308);
or U21585 (N_21585,N_18317,N_18059);
and U21586 (N_21586,N_19689,N_18669);
nand U21587 (N_21587,N_19601,N_18443);
nand U21588 (N_21588,N_19690,N_19216);
nand U21589 (N_21589,N_18680,N_19613);
and U21590 (N_21590,N_18756,N_19821);
nor U21591 (N_21591,N_18607,N_18710);
or U21592 (N_21592,N_19017,N_18496);
nor U21593 (N_21593,N_18988,N_19477);
nand U21594 (N_21594,N_19931,N_18715);
and U21595 (N_21595,N_18165,N_18274);
and U21596 (N_21596,N_19211,N_18416);
or U21597 (N_21597,N_18627,N_18719);
or U21598 (N_21598,N_19755,N_18339);
nor U21599 (N_21599,N_18109,N_19880);
or U21600 (N_21600,N_18726,N_19284);
nor U21601 (N_21601,N_19240,N_18204);
and U21602 (N_21602,N_19730,N_18977);
nor U21603 (N_21603,N_19983,N_19582);
nor U21604 (N_21604,N_19744,N_18573);
xor U21605 (N_21605,N_19970,N_18135);
nand U21606 (N_21606,N_19376,N_18022);
nand U21607 (N_21607,N_19953,N_19093);
and U21608 (N_21608,N_19748,N_19161);
or U21609 (N_21609,N_19798,N_18393);
or U21610 (N_21610,N_18886,N_19077);
nand U21611 (N_21611,N_19728,N_19687);
nand U21612 (N_21612,N_19064,N_18489);
xor U21613 (N_21613,N_19054,N_19687);
and U21614 (N_21614,N_18163,N_18593);
nor U21615 (N_21615,N_18924,N_19033);
and U21616 (N_21616,N_19013,N_18210);
nor U21617 (N_21617,N_18619,N_18263);
nor U21618 (N_21618,N_18460,N_19080);
nor U21619 (N_21619,N_18677,N_19794);
nand U21620 (N_21620,N_19218,N_18516);
or U21621 (N_21621,N_18057,N_18391);
nor U21622 (N_21622,N_19065,N_19540);
nor U21623 (N_21623,N_18785,N_18602);
nand U21624 (N_21624,N_19401,N_19008);
nand U21625 (N_21625,N_18200,N_18868);
or U21626 (N_21626,N_18356,N_18785);
or U21627 (N_21627,N_18340,N_19217);
or U21628 (N_21628,N_19004,N_18135);
or U21629 (N_21629,N_18538,N_19638);
nand U21630 (N_21630,N_19400,N_18682);
xnor U21631 (N_21631,N_18336,N_18444);
and U21632 (N_21632,N_19063,N_18083);
nor U21633 (N_21633,N_19061,N_18146);
and U21634 (N_21634,N_18476,N_18796);
nor U21635 (N_21635,N_19068,N_19005);
xor U21636 (N_21636,N_18221,N_18133);
or U21637 (N_21637,N_18887,N_18041);
and U21638 (N_21638,N_18247,N_19689);
and U21639 (N_21639,N_18544,N_18749);
and U21640 (N_21640,N_18650,N_18196);
and U21641 (N_21641,N_18383,N_19436);
and U21642 (N_21642,N_19742,N_18990);
nor U21643 (N_21643,N_19032,N_18250);
or U21644 (N_21644,N_18160,N_19359);
and U21645 (N_21645,N_19445,N_18377);
nand U21646 (N_21646,N_19927,N_18257);
or U21647 (N_21647,N_18529,N_19781);
xnor U21648 (N_21648,N_18370,N_18121);
or U21649 (N_21649,N_18318,N_18938);
or U21650 (N_21650,N_18203,N_18679);
nand U21651 (N_21651,N_18312,N_18160);
and U21652 (N_21652,N_19869,N_19664);
and U21653 (N_21653,N_18121,N_18897);
or U21654 (N_21654,N_19628,N_19291);
nor U21655 (N_21655,N_19024,N_19214);
or U21656 (N_21656,N_19453,N_18194);
and U21657 (N_21657,N_19395,N_18586);
and U21658 (N_21658,N_19237,N_18291);
and U21659 (N_21659,N_18874,N_19478);
nand U21660 (N_21660,N_18149,N_19670);
nand U21661 (N_21661,N_18215,N_19532);
or U21662 (N_21662,N_18827,N_18731);
and U21663 (N_21663,N_18563,N_19422);
or U21664 (N_21664,N_19157,N_19696);
or U21665 (N_21665,N_18616,N_19720);
nor U21666 (N_21666,N_18760,N_19406);
nor U21667 (N_21667,N_18782,N_18632);
or U21668 (N_21668,N_19024,N_18758);
nand U21669 (N_21669,N_18040,N_19017);
xor U21670 (N_21670,N_18655,N_18591);
and U21671 (N_21671,N_19943,N_18573);
nor U21672 (N_21672,N_19291,N_19076);
nand U21673 (N_21673,N_19458,N_19987);
and U21674 (N_21674,N_19936,N_19340);
and U21675 (N_21675,N_18025,N_18684);
nand U21676 (N_21676,N_18985,N_19255);
nand U21677 (N_21677,N_19216,N_19796);
or U21678 (N_21678,N_18912,N_19464);
nand U21679 (N_21679,N_18332,N_18537);
nor U21680 (N_21680,N_19762,N_18318);
and U21681 (N_21681,N_19692,N_19011);
or U21682 (N_21682,N_19302,N_18038);
nor U21683 (N_21683,N_18858,N_18910);
nor U21684 (N_21684,N_19814,N_19109);
nand U21685 (N_21685,N_18841,N_18684);
and U21686 (N_21686,N_18701,N_18786);
nand U21687 (N_21687,N_18177,N_18923);
nor U21688 (N_21688,N_19790,N_19742);
nor U21689 (N_21689,N_19133,N_18378);
nor U21690 (N_21690,N_18732,N_18151);
nor U21691 (N_21691,N_19838,N_19411);
or U21692 (N_21692,N_18003,N_19924);
nor U21693 (N_21693,N_19293,N_19973);
nand U21694 (N_21694,N_19659,N_18788);
or U21695 (N_21695,N_18486,N_19139);
nor U21696 (N_21696,N_18104,N_19166);
nor U21697 (N_21697,N_18556,N_19367);
or U21698 (N_21698,N_19269,N_19964);
nand U21699 (N_21699,N_18570,N_18730);
nor U21700 (N_21700,N_18201,N_18273);
nand U21701 (N_21701,N_18375,N_19596);
nor U21702 (N_21702,N_18075,N_19063);
nand U21703 (N_21703,N_18672,N_18514);
nor U21704 (N_21704,N_18064,N_19423);
or U21705 (N_21705,N_18966,N_18442);
nand U21706 (N_21706,N_19061,N_19415);
nand U21707 (N_21707,N_18314,N_19784);
or U21708 (N_21708,N_18773,N_19181);
and U21709 (N_21709,N_18380,N_18610);
or U21710 (N_21710,N_18353,N_19507);
nand U21711 (N_21711,N_18657,N_19989);
or U21712 (N_21712,N_19394,N_18495);
or U21713 (N_21713,N_18067,N_18501);
and U21714 (N_21714,N_19156,N_19822);
nor U21715 (N_21715,N_18496,N_18589);
nand U21716 (N_21716,N_19949,N_18313);
nand U21717 (N_21717,N_19641,N_18274);
nand U21718 (N_21718,N_19243,N_19271);
and U21719 (N_21719,N_18333,N_18053);
or U21720 (N_21720,N_19954,N_19363);
or U21721 (N_21721,N_18069,N_18578);
or U21722 (N_21722,N_18416,N_18359);
and U21723 (N_21723,N_18856,N_19495);
nand U21724 (N_21724,N_18943,N_19276);
and U21725 (N_21725,N_19531,N_18636);
and U21726 (N_21726,N_18916,N_19331);
nand U21727 (N_21727,N_19191,N_18460);
nand U21728 (N_21728,N_18346,N_18779);
nand U21729 (N_21729,N_19817,N_19837);
and U21730 (N_21730,N_19718,N_18720);
nor U21731 (N_21731,N_18809,N_19958);
or U21732 (N_21732,N_19136,N_19750);
or U21733 (N_21733,N_18827,N_18263);
nor U21734 (N_21734,N_19591,N_18939);
nor U21735 (N_21735,N_19997,N_18377);
or U21736 (N_21736,N_18893,N_19334);
or U21737 (N_21737,N_18906,N_19260);
nand U21738 (N_21738,N_18287,N_19933);
nand U21739 (N_21739,N_18201,N_18776);
nor U21740 (N_21740,N_19071,N_19916);
or U21741 (N_21741,N_19396,N_19250);
and U21742 (N_21742,N_18226,N_19590);
nor U21743 (N_21743,N_19240,N_19752);
nand U21744 (N_21744,N_19450,N_18521);
or U21745 (N_21745,N_19611,N_18358);
nand U21746 (N_21746,N_18390,N_18101);
nand U21747 (N_21747,N_19260,N_19410);
or U21748 (N_21748,N_18950,N_19677);
nor U21749 (N_21749,N_18324,N_19525);
nor U21750 (N_21750,N_19764,N_18042);
nand U21751 (N_21751,N_18593,N_18504);
and U21752 (N_21752,N_19272,N_18122);
or U21753 (N_21753,N_19236,N_18087);
and U21754 (N_21754,N_19238,N_18741);
nor U21755 (N_21755,N_18821,N_19796);
and U21756 (N_21756,N_18959,N_19573);
or U21757 (N_21757,N_19287,N_19043);
nor U21758 (N_21758,N_18994,N_19768);
nor U21759 (N_21759,N_18525,N_18046);
nor U21760 (N_21760,N_19980,N_18711);
nor U21761 (N_21761,N_19896,N_19492);
and U21762 (N_21762,N_19308,N_18998);
and U21763 (N_21763,N_19159,N_18819);
xnor U21764 (N_21764,N_19885,N_18941);
nand U21765 (N_21765,N_19985,N_18577);
or U21766 (N_21766,N_19551,N_18822);
nand U21767 (N_21767,N_18173,N_19975);
and U21768 (N_21768,N_18281,N_18902);
or U21769 (N_21769,N_19808,N_18124);
nor U21770 (N_21770,N_19070,N_19509);
nor U21771 (N_21771,N_18713,N_18093);
and U21772 (N_21772,N_19782,N_19051);
nand U21773 (N_21773,N_19232,N_18366);
or U21774 (N_21774,N_19273,N_19053);
nand U21775 (N_21775,N_19601,N_19511);
and U21776 (N_21776,N_18391,N_18233);
nor U21777 (N_21777,N_18323,N_19549);
nand U21778 (N_21778,N_19786,N_18758);
and U21779 (N_21779,N_18521,N_18589);
or U21780 (N_21780,N_19552,N_19304);
or U21781 (N_21781,N_18113,N_18963);
or U21782 (N_21782,N_18045,N_18441);
or U21783 (N_21783,N_19257,N_19012);
and U21784 (N_21784,N_18361,N_18328);
or U21785 (N_21785,N_19983,N_19720);
and U21786 (N_21786,N_19105,N_18327);
or U21787 (N_21787,N_18705,N_18937);
or U21788 (N_21788,N_19572,N_18628);
nand U21789 (N_21789,N_19709,N_18184);
nor U21790 (N_21790,N_18986,N_19407);
or U21791 (N_21791,N_19165,N_19262);
nand U21792 (N_21792,N_18863,N_18816);
nor U21793 (N_21793,N_18484,N_19188);
nand U21794 (N_21794,N_19514,N_18865);
nand U21795 (N_21795,N_18952,N_19560);
nand U21796 (N_21796,N_19186,N_19911);
nand U21797 (N_21797,N_19166,N_19685);
and U21798 (N_21798,N_18128,N_18778);
and U21799 (N_21799,N_18872,N_19348);
nor U21800 (N_21800,N_18348,N_18119);
or U21801 (N_21801,N_19503,N_18717);
xnor U21802 (N_21802,N_19321,N_19821);
nand U21803 (N_21803,N_18455,N_18805);
and U21804 (N_21804,N_18274,N_19124);
and U21805 (N_21805,N_19382,N_19296);
or U21806 (N_21806,N_18314,N_19763);
nor U21807 (N_21807,N_18895,N_18928);
and U21808 (N_21808,N_18779,N_19304);
nor U21809 (N_21809,N_19802,N_19919);
nand U21810 (N_21810,N_18340,N_18307);
nor U21811 (N_21811,N_18469,N_18091);
nand U21812 (N_21812,N_19909,N_18490);
or U21813 (N_21813,N_18441,N_19430);
nor U21814 (N_21814,N_18932,N_19022);
nor U21815 (N_21815,N_19575,N_18125);
xnor U21816 (N_21816,N_19580,N_19076);
nand U21817 (N_21817,N_18984,N_19307);
nand U21818 (N_21818,N_19556,N_18646);
nand U21819 (N_21819,N_18381,N_18247);
or U21820 (N_21820,N_19444,N_18611);
or U21821 (N_21821,N_19394,N_18584);
nor U21822 (N_21822,N_18909,N_18871);
nand U21823 (N_21823,N_19695,N_19817);
or U21824 (N_21824,N_19359,N_18144);
or U21825 (N_21825,N_18707,N_18413);
nand U21826 (N_21826,N_18714,N_18726);
nor U21827 (N_21827,N_18643,N_18303);
and U21828 (N_21828,N_19115,N_18955);
nand U21829 (N_21829,N_19257,N_18539);
nor U21830 (N_21830,N_19703,N_18367);
xnor U21831 (N_21831,N_18449,N_18642);
and U21832 (N_21832,N_18855,N_18919);
nor U21833 (N_21833,N_19750,N_19278);
nand U21834 (N_21834,N_19181,N_19688);
nor U21835 (N_21835,N_18331,N_19745);
nand U21836 (N_21836,N_19127,N_18576);
nand U21837 (N_21837,N_19151,N_19671);
and U21838 (N_21838,N_19457,N_19769);
nor U21839 (N_21839,N_19151,N_19244);
and U21840 (N_21840,N_19239,N_19685);
nand U21841 (N_21841,N_18180,N_18803);
or U21842 (N_21842,N_19780,N_18160);
nand U21843 (N_21843,N_18226,N_19930);
xnor U21844 (N_21844,N_18249,N_19611);
and U21845 (N_21845,N_19583,N_18542);
and U21846 (N_21846,N_19972,N_18124);
and U21847 (N_21847,N_18626,N_19516);
nor U21848 (N_21848,N_18941,N_19477);
nand U21849 (N_21849,N_19712,N_18034);
nor U21850 (N_21850,N_18698,N_18745);
and U21851 (N_21851,N_18465,N_18801);
nand U21852 (N_21852,N_19208,N_18742);
nand U21853 (N_21853,N_18258,N_19810);
nand U21854 (N_21854,N_18730,N_19216);
or U21855 (N_21855,N_18352,N_19725);
or U21856 (N_21856,N_18394,N_18108);
xnor U21857 (N_21857,N_18854,N_19701);
and U21858 (N_21858,N_19422,N_19112);
nand U21859 (N_21859,N_19956,N_19112);
nand U21860 (N_21860,N_19123,N_19963);
nor U21861 (N_21861,N_19416,N_18385);
and U21862 (N_21862,N_18476,N_19881);
or U21863 (N_21863,N_18848,N_18662);
or U21864 (N_21864,N_18400,N_18928);
nand U21865 (N_21865,N_18642,N_19882);
nand U21866 (N_21866,N_18702,N_18726);
and U21867 (N_21867,N_18828,N_18929);
nor U21868 (N_21868,N_19581,N_18775);
nand U21869 (N_21869,N_19240,N_19128);
or U21870 (N_21870,N_19546,N_18773);
and U21871 (N_21871,N_19715,N_18576);
nor U21872 (N_21872,N_19979,N_18602);
nand U21873 (N_21873,N_19663,N_18237);
and U21874 (N_21874,N_18287,N_19890);
and U21875 (N_21875,N_19900,N_19160);
nand U21876 (N_21876,N_18692,N_18987);
and U21877 (N_21877,N_18174,N_18467);
and U21878 (N_21878,N_19490,N_19882);
and U21879 (N_21879,N_19098,N_19849);
nor U21880 (N_21880,N_19234,N_18968);
nand U21881 (N_21881,N_18174,N_18973);
or U21882 (N_21882,N_19102,N_19436);
and U21883 (N_21883,N_18487,N_19192);
or U21884 (N_21884,N_18110,N_18189);
nor U21885 (N_21885,N_19606,N_19680);
nor U21886 (N_21886,N_18234,N_19485);
or U21887 (N_21887,N_18583,N_18446);
and U21888 (N_21888,N_19183,N_18337);
or U21889 (N_21889,N_19333,N_18830);
nor U21890 (N_21890,N_19429,N_19692);
nor U21891 (N_21891,N_19089,N_19717);
nor U21892 (N_21892,N_18830,N_19262);
or U21893 (N_21893,N_18105,N_19595);
nor U21894 (N_21894,N_18428,N_18448);
or U21895 (N_21895,N_18610,N_18153);
nand U21896 (N_21896,N_18165,N_18438);
xor U21897 (N_21897,N_18208,N_19795);
and U21898 (N_21898,N_19293,N_19448);
or U21899 (N_21899,N_18838,N_19036);
and U21900 (N_21900,N_19074,N_18469);
or U21901 (N_21901,N_18961,N_18545);
nand U21902 (N_21902,N_19207,N_18056);
and U21903 (N_21903,N_19610,N_18770);
and U21904 (N_21904,N_18179,N_18727);
and U21905 (N_21905,N_19933,N_18553);
and U21906 (N_21906,N_19093,N_18231);
nand U21907 (N_21907,N_18438,N_18737);
and U21908 (N_21908,N_19866,N_18357);
and U21909 (N_21909,N_19485,N_18507);
or U21910 (N_21910,N_19994,N_18541);
or U21911 (N_21911,N_18957,N_19402);
or U21912 (N_21912,N_19078,N_18566);
nor U21913 (N_21913,N_19566,N_19288);
nor U21914 (N_21914,N_19306,N_18229);
and U21915 (N_21915,N_19978,N_18876);
and U21916 (N_21916,N_19878,N_18420);
nor U21917 (N_21917,N_18467,N_18800);
nor U21918 (N_21918,N_19402,N_18671);
nor U21919 (N_21919,N_19611,N_18746);
nor U21920 (N_21920,N_18701,N_18214);
or U21921 (N_21921,N_19374,N_18251);
nor U21922 (N_21922,N_19008,N_18144);
nand U21923 (N_21923,N_19772,N_18156);
nor U21924 (N_21924,N_18014,N_18967);
or U21925 (N_21925,N_18851,N_19812);
or U21926 (N_21926,N_19174,N_18963);
nand U21927 (N_21927,N_18567,N_18289);
nand U21928 (N_21928,N_18970,N_19840);
nor U21929 (N_21929,N_18232,N_18401);
nand U21930 (N_21930,N_19574,N_19596);
nor U21931 (N_21931,N_19888,N_18364);
and U21932 (N_21932,N_18277,N_19742);
nand U21933 (N_21933,N_18649,N_18964);
and U21934 (N_21934,N_19863,N_18353);
or U21935 (N_21935,N_18718,N_19514);
nand U21936 (N_21936,N_19109,N_19560);
and U21937 (N_21937,N_19336,N_18221);
and U21938 (N_21938,N_18645,N_18620);
nand U21939 (N_21939,N_18173,N_18715);
and U21940 (N_21940,N_19088,N_19959);
and U21941 (N_21941,N_18657,N_19926);
nor U21942 (N_21942,N_19160,N_18950);
or U21943 (N_21943,N_19663,N_18604);
and U21944 (N_21944,N_19980,N_19333);
nand U21945 (N_21945,N_18362,N_18084);
or U21946 (N_21946,N_19519,N_18832);
or U21947 (N_21947,N_19462,N_19538);
nor U21948 (N_21948,N_19632,N_18498);
or U21949 (N_21949,N_19800,N_19499);
nor U21950 (N_21950,N_18545,N_19118);
nand U21951 (N_21951,N_19087,N_18545);
and U21952 (N_21952,N_19452,N_19205);
nor U21953 (N_21953,N_19534,N_18093);
and U21954 (N_21954,N_18785,N_19618);
nor U21955 (N_21955,N_18861,N_18827);
nand U21956 (N_21956,N_19246,N_19637);
and U21957 (N_21957,N_19851,N_18522);
and U21958 (N_21958,N_18913,N_19080);
xor U21959 (N_21959,N_19645,N_19099);
nor U21960 (N_21960,N_19281,N_18079);
nand U21961 (N_21961,N_19862,N_18589);
nor U21962 (N_21962,N_18901,N_19738);
or U21963 (N_21963,N_18044,N_18429);
nor U21964 (N_21964,N_18951,N_18445);
nand U21965 (N_21965,N_19323,N_18833);
nor U21966 (N_21966,N_19407,N_19755);
or U21967 (N_21967,N_19110,N_19530);
or U21968 (N_21968,N_19905,N_19052);
nor U21969 (N_21969,N_19892,N_19571);
nor U21970 (N_21970,N_19283,N_19855);
and U21971 (N_21971,N_19490,N_18861);
or U21972 (N_21972,N_19061,N_19272);
and U21973 (N_21973,N_19297,N_19841);
or U21974 (N_21974,N_18206,N_19166);
or U21975 (N_21975,N_19639,N_19321);
or U21976 (N_21976,N_18576,N_19585);
nand U21977 (N_21977,N_18140,N_19015);
nand U21978 (N_21978,N_18456,N_19560);
and U21979 (N_21979,N_18923,N_18338);
and U21980 (N_21980,N_18798,N_18680);
nor U21981 (N_21981,N_18609,N_18816);
nand U21982 (N_21982,N_18507,N_19012);
nor U21983 (N_21983,N_18725,N_19486);
nor U21984 (N_21984,N_19971,N_19604);
nor U21985 (N_21985,N_18718,N_18394);
and U21986 (N_21986,N_18049,N_19524);
or U21987 (N_21987,N_18522,N_19635);
nand U21988 (N_21988,N_19622,N_18099);
or U21989 (N_21989,N_18772,N_18014);
or U21990 (N_21990,N_18732,N_19928);
and U21991 (N_21991,N_18762,N_19988);
nor U21992 (N_21992,N_18336,N_19932);
and U21993 (N_21993,N_18166,N_19052);
nand U21994 (N_21994,N_18961,N_18152);
nor U21995 (N_21995,N_18304,N_18481);
nand U21996 (N_21996,N_19903,N_19061);
and U21997 (N_21997,N_19190,N_18995);
nand U21998 (N_21998,N_19036,N_18029);
nor U21999 (N_21999,N_19411,N_19607);
and U22000 (N_22000,N_21449,N_20915);
and U22001 (N_22001,N_21058,N_20319);
nand U22002 (N_22002,N_21101,N_20320);
nand U22003 (N_22003,N_21456,N_21170);
nand U22004 (N_22004,N_20761,N_20057);
nand U22005 (N_22005,N_21592,N_21577);
nor U22006 (N_22006,N_20542,N_21053);
or U22007 (N_22007,N_20874,N_20700);
or U22008 (N_22008,N_20070,N_21714);
and U22009 (N_22009,N_21502,N_20271);
nand U22010 (N_22010,N_20224,N_20938);
nor U22011 (N_22011,N_20382,N_21032);
or U22012 (N_22012,N_20090,N_20635);
nor U22013 (N_22013,N_20163,N_21768);
or U22014 (N_22014,N_20696,N_20653);
nand U22015 (N_22015,N_20363,N_20211);
and U22016 (N_22016,N_21850,N_21154);
or U22017 (N_22017,N_20752,N_20334);
nor U22018 (N_22018,N_20647,N_21744);
or U22019 (N_22019,N_21568,N_20468);
or U22020 (N_22020,N_21481,N_21855);
nand U22021 (N_22021,N_20709,N_21969);
nor U22022 (N_22022,N_21068,N_21124);
nor U22023 (N_22023,N_21927,N_20917);
or U22024 (N_22024,N_21440,N_20694);
nand U22025 (N_22025,N_20766,N_20238);
nor U22026 (N_22026,N_20093,N_21394);
nand U22027 (N_22027,N_21408,N_20423);
nor U22028 (N_22028,N_20489,N_20681);
xnor U22029 (N_22029,N_20975,N_20632);
or U22030 (N_22030,N_21480,N_21924);
and U22031 (N_22031,N_21912,N_20512);
nand U22032 (N_22032,N_21105,N_21683);
nand U22033 (N_22033,N_21729,N_20415);
nand U22034 (N_22034,N_21153,N_20302);
or U22035 (N_22035,N_20809,N_20114);
nand U22036 (N_22036,N_21229,N_21828);
nor U22037 (N_22037,N_21358,N_21051);
nor U22038 (N_22038,N_21548,N_21305);
and U22039 (N_22039,N_20013,N_20569);
nand U22040 (N_22040,N_20943,N_21605);
or U22041 (N_22041,N_21657,N_21133);
nor U22042 (N_22042,N_20050,N_20607);
or U22043 (N_22043,N_21600,N_20649);
or U22044 (N_22044,N_21926,N_20048);
and U22045 (N_22045,N_21553,N_21342);
and U22046 (N_22046,N_21696,N_21922);
nor U22047 (N_22047,N_21249,N_21015);
and U22048 (N_22048,N_21146,N_21441);
nor U22049 (N_22049,N_20007,N_21970);
or U22050 (N_22050,N_20893,N_21399);
nor U22051 (N_22051,N_21289,N_20092);
nor U22052 (N_22052,N_20557,N_20472);
or U22053 (N_22053,N_21836,N_20811);
nor U22054 (N_22054,N_20872,N_21754);
and U22055 (N_22055,N_21737,N_20418);
nand U22056 (N_22056,N_21673,N_21264);
and U22057 (N_22057,N_20828,N_21861);
nand U22058 (N_22058,N_21222,N_20169);
nand U22059 (N_22059,N_21516,N_21911);
and U22060 (N_22060,N_21870,N_21198);
and U22061 (N_22061,N_20179,N_20417);
or U22062 (N_22062,N_21023,N_20031);
and U22063 (N_22063,N_20160,N_20503);
and U22064 (N_22064,N_20913,N_21766);
and U22065 (N_22065,N_21920,N_20802);
nand U22066 (N_22066,N_21556,N_20433);
and U22067 (N_22067,N_21174,N_21290);
or U22068 (N_22068,N_21138,N_21535);
and U22069 (N_22069,N_20675,N_21518);
nand U22070 (N_22070,N_21971,N_20735);
nand U22071 (N_22071,N_21776,N_20736);
nand U22072 (N_22072,N_20219,N_21994);
nor U22073 (N_22073,N_20466,N_21671);
nor U22074 (N_22074,N_20812,N_21040);
or U22075 (N_22075,N_20208,N_20740);
nand U22076 (N_22076,N_20150,N_20107);
and U22077 (N_22077,N_21808,N_20676);
nand U22078 (N_22078,N_21352,N_21595);
nor U22079 (N_22079,N_20973,N_20102);
nor U22080 (N_22080,N_20544,N_20704);
nand U22081 (N_22081,N_20990,N_21016);
nand U22082 (N_22082,N_20964,N_20556);
nor U22083 (N_22083,N_21250,N_21246);
or U22084 (N_22084,N_21803,N_20778);
nand U22085 (N_22085,N_20367,N_20309);
nand U22086 (N_22086,N_21944,N_20531);
nand U22087 (N_22087,N_20223,N_20911);
nand U22088 (N_22088,N_21769,N_21667);
nand U22089 (N_22089,N_21462,N_21231);
or U22090 (N_22090,N_21355,N_20288);
nor U22091 (N_22091,N_21946,N_21644);
nor U22092 (N_22092,N_20516,N_21243);
nand U22093 (N_22093,N_21259,N_20027);
nor U22094 (N_22094,N_20316,N_20996);
or U22095 (N_22095,N_20793,N_20524);
nand U22096 (N_22096,N_21067,N_20714);
nor U22097 (N_22097,N_20554,N_20899);
nor U22098 (N_22098,N_21093,N_21149);
nand U22099 (N_22099,N_21654,N_20762);
nor U22100 (N_22100,N_20508,N_20876);
nor U22101 (N_22101,N_20442,N_20966);
nand U22102 (N_22102,N_20739,N_21147);
or U22103 (N_22103,N_21063,N_20283);
or U22104 (N_22104,N_21160,N_20963);
nand U22105 (N_22105,N_21003,N_20342);
or U22106 (N_22106,N_20940,N_20948);
or U22107 (N_22107,N_20687,N_21585);
and U22108 (N_22108,N_21418,N_20592);
or U22109 (N_22109,N_20474,N_20161);
nor U22110 (N_22110,N_20565,N_21491);
and U22111 (N_22111,N_21430,N_20346);
or U22112 (N_22112,N_21205,N_20581);
nand U22113 (N_22113,N_20492,N_20419);
or U22114 (N_22114,N_20133,N_20780);
xnor U22115 (N_22115,N_20236,N_21638);
nand U22116 (N_22116,N_20923,N_21433);
nand U22117 (N_22117,N_21843,N_20343);
nand U22118 (N_22118,N_20144,N_21561);
or U22119 (N_22119,N_20509,N_21165);
nand U22120 (N_22120,N_20193,N_21761);
and U22121 (N_22121,N_20256,N_20378);
nand U22122 (N_22122,N_21790,N_21361);
nand U22123 (N_22123,N_21747,N_20551);
and U22124 (N_22124,N_21451,N_21965);
nor U22125 (N_22125,N_20059,N_21457);
or U22126 (N_22126,N_21262,N_21185);
or U22127 (N_22127,N_20462,N_21034);
nor U22128 (N_22128,N_21385,N_21723);
nor U22129 (N_22129,N_21557,N_21917);
nor U22130 (N_22130,N_21712,N_21791);
nand U22131 (N_22131,N_20716,N_20603);
and U22132 (N_22132,N_20167,N_20620);
nor U22133 (N_22133,N_21158,N_21931);
and U22134 (N_22134,N_21607,N_20255);
or U22135 (N_22135,N_20612,N_20803);
nand U22136 (N_22136,N_21802,N_20623);
xnor U22137 (N_22137,N_20072,N_20200);
or U22138 (N_22138,N_21442,N_21637);
and U22139 (N_22139,N_20715,N_20616);
nor U22140 (N_22140,N_21123,N_21646);
nor U22141 (N_22141,N_20190,N_21307);
nand U22142 (N_22142,N_20527,N_20413);
nand U22143 (N_22143,N_20885,N_20499);
and U22144 (N_22144,N_20820,N_20595);
or U22145 (N_22145,N_20396,N_20630);
nor U22146 (N_22146,N_21951,N_21704);
nor U22147 (N_22147,N_20648,N_20670);
or U22148 (N_22148,N_20350,N_21255);
nor U22149 (N_22149,N_21446,N_21860);
nand U22150 (N_22150,N_20074,N_20584);
nand U22151 (N_22151,N_20362,N_20373);
nor U22152 (N_22152,N_20639,N_20277);
nor U22153 (N_22153,N_20446,N_20753);
or U22154 (N_22154,N_20852,N_21191);
and U22155 (N_22155,N_21291,N_21363);
nor U22156 (N_22156,N_20685,N_21950);
nor U22157 (N_22157,N_21360,N_20301);
or U22158 (N_22158,N_20022,N_21252);
or U22159 (N_22159,N_20510,N_21833);
or U22160 (N_22160,N_21292,N_21398);
nor U22161 (N_22161,N_21847,N_20545);
or U22162 (N_22162,N_21787,N_21349);
and U22163 (N_22163,N_20184,N_21296);
nand U22164 (N_22164,N_20197,N_21283);
nor U22165 (N_22165,N_20808,N_21055);
or U22166 (N_22166,N_20579,N_21665);
or U22167 (N_22167,N_20826,N_20490);
nand U22168 (N_22168,N_21771,N_20819);
and U22169 (N_22169,N_21054,N_21672);
and U22170 (N_22170,N_20981,N_21166);
and U22171 (N_22171,N_21366,N_20352);
nand U22172 (N_22172,N_21497,N_21883);
and U22173 (N_22173,N_21207,N_21545);
or U22174 (N_22174,N_21905,N_20798);
nand U22175 (N_22175,N_20563,N_21656);
and U22176 (N_22176,N_21437,N_21489);
or U22177 (N_22177,N_20930,N_21524);
or U22178 (N_22178,N_20712,N_20533);
xor U22179 (N_22179,N_20786,N_20307);
or U22180 (N_22180,N_21942,N_20773);
or U22181 (N_22181,N_21006,N_21980);
nor U22182 (N_22182,N_20389,N_20065);
nand U22183 (N_22183,N_21984,N_20049);
and U22184 (N_22184,N_20707,N_21907);
nand U22185 (N_22185,N_20546,N_20958);
or U22186 (N_22186,N_21428,N_20486);
or U22187 (N_22187,N_20482,N_21267);
nor U22188 (N_22188,N_21303,N_20829);
xor U22189 (N_22189,N_21986,N_20548);
xor U22190 (N_22190,N_20896,N_21429);
nand U22191 (N_22191,N_21127,N_21632);
nor U22192 (N_22192,N_21902,N_21914);
or U22193 (N_22193,N_20513,N_21613);
nor U22194 (N_22194,N_20275,N_21730);
nor U22195 (N_22195,N_20241,N_21356);
and U22196 (N_22196,N_21580,N_20760);
nor U22197 (N_22197,N_20344,N_20252);
and U22198 (N_22198,N_20838,N_21265);
nor U22199 (N_22199,N_21111,N_21135);
nand U22200 (N_22200,N_21716,N_20892);
nand U22201 (N_22201,N_20705,N_20183);
and U22202 (N_22202,N_21075,N_21972);
and U22203 (N_22203,N_21631,N_21699);
or U22204 (N_22204,N_21121,N_21517);
and U22205 (N_22205,N_21287,N_20186);
nor U22206 (N_22206,N_20666,N_21778);
nor U22207 (N_22207,N_21472,N_21223);
nor U22208 (N_22208,N_21519,N_21968);
or U22209 (N_22209,N_20312,N_21558);
or U22210 (N_22210,N_21314,N_20856);
nand U22211 (N_22211,N_21417,N_20475);
nor U22212 (N_22212,N_20310,N_20105);
and U22213 (N_22213,N_20906,N_20608);
nor U22214 (N_22214,N_20759,N_21711);
nor U22215 (N_22215,N_21196,N_20424);
nand U22216 (N_22216,N_20745,N_20397);
nand U22217 (N_22217,N_20481,N_20925);
nor U22218 (N_22218,N_20390,N_21899);
or U22219 (N_22219,N_21080,N_20098);
and U22220 (N_22220,N_21735,N_21688);
and U22221 (N_22221,N_20552,N_20591);
or U22222 (N_22222,N_20176,N_21234);
and U22223 (N_22223,N_21027,N_20199);
nand U22224 (N_22224,N_21005,N_21373);
or U22225 (N_22225,N_21715,N_21537);
or U22226 (N_22226,N_20033,N_20043);
nand U22227 (N_22227,N_20667,N_21348);
and U22228 (N_22228,N_21751,N_21526);
and U22229 (N_22229,N_21167,N_21288);
or U22230 (N_22230,N_20689,N_20845);
and U22231 (N_22231,N_21831,N_21993);
and U22232 (N_22232,N_21285,N_21892);
xnor U22233 (N_22233,N_20116,N_20306);
or U22234 (N_22234,N_20011,N_20227);
or U22235 (N_22235,N_21318,N_20678);
nand U22236 (N_22236,N_20052,N_21693);
xor U22237 (N_22237,N_21470,N_20790);
nand U22238 (N_22238,N_21013,N_20698);
or U22239 (N_22239,N_20519,N_21043);
nand U22240 (N_22240,N_21010,N_21176);
nor U22241 (N_22241,N_20430,N_21109);
or U22242 (N_22242,N_20748,N_21425);
or U22243 (N_22243,N_20853,N_21713);
or U22244 (N_22244,N_21884,N_21890);
nand U22245 (N_22245,N_20476,N_20369);
nor U22246 (N_22246,N_20897,N_20380);
nor U22247 (N_22247,N_20154,N_21513);
or U22248 (N_22248,N_20789,N_21499);
or U22249 (N_22249,N_20422,N_20438);
nor U22250 (N_22250,N_20847,N_20865);
or U22251 (N_22251,N_21137,N_20129);
or U22252 (N_22252,N_21849,N_20171);
nand U22253 (N_22253,N_21376,N_20741);
and U22254 (N_22254,N_20890,N_21838);
nand U22255 (N_22255,N_21465,N_21066);
nor U22256 (N_22256,N_21204,N_20775);
or U22257 (N_22257,N_21733,N_21708);
or U22258 (N_22258,N_20047,N_20815);
or U22259 (N_22259,N_20604,N_20693);
nand U22260 (N_22260,N_20041,N_21095);
nor U22261 (N_22261,N_20625,N_21966);
nand U22262 (N_22262,N_20493,N_21896);
or U22263 (N_22263,N_20629,N_21028);
nand U22264 (N_22264,N_21757,N_21698);
or U22265 (N_22265,N_20155,N_21742);
or U22266 (N_22266,N_21615,N_20426);
nand U22267 (N_22267,N_21351,N_21159);
nor U22268 (N_22268,N_20843,N_20992);
and U22269 (N_22269,N_21507,N_21520);
nor U22270 (N_22270,N_20453,N_21772);
nand U22271 (N_22271,N_20795,N_20977);
and U22272 (N_22272,N_21322,N_20257);
nor U22273 (N_22273,N_21113,N_20995);
or U22274 (N_22274,N_21203,N_21251);
nand U22275 (N_22275,N_21202,N_21813);
nand U22276 (N_22276,N_21219,N_21484);
nor U22277 (N_22277,N_20756,N_20198);
and U22278 (N_22278,N_21045,N_20807);
nand U22279 (N_22279,N_20268,N_20650);
or U22280 (N_22280,N_20537,N_20526);
nand U22281 (N_22281,N_20934,N_20960);
and U22282 (N_22282,N_20248,N_20641);
and U22283 (N_22283,N_21738,N_20018);
or U22284 (N_22284,N_21498,N_20101);
and U22285 (N_22285,N_21000,N_21389);
nand U22286 (N_22286,N_21603,N_21897);
nor U22287 (N_22287,N_20103,N_20726);
nand U22288 (N_22288,N_21581,N_20921);
nor U22289 (N_22289,N_20229,N_20850);
nor U22290 (N_22290,N_20463,N_21452);
and U22291 (N_22291,N_20001,N_20274);
nand U22292 (N_22292,N_21315,N_20794);
or U22293 (N_22293,N_20174,N_21227);
and U22294 (N_22294,N_21586,N_20928);
nand U22295 (N_22295,N_20166,N_21037);
and U22296 (N_22296,N_20159,N_21724);
nor U22297 (N_22297,N_21867,N_20673);
and U22298 (N_22298,N_21019,N_21645);
nor U22299 (N_22299,N_21435,N_21622);
or U22300 (N_22300,N_21770,N_20622);
nor U22301 (N_22301,N_21625,N_20860);
and U22302 (N_22302,N_21989,N_20528);
nor U22303 (N_22303,N_20353,N_20734);
nand U22304 (N_22304,N_20431,N_20547);
nand U22305 (N_22305,N_20286,N_21280);
xor U22306 (N_22306,N_21588,N_21739);
or U22307 (N_22307,N_21854,N_20540);
and U22308 (N_22308,N_20918,N_21574);
nor U22309 (N_22309,N_21431,N_21172);
and U22310 (N_22310,N_20699,N_20656);
nand U22311 (N_22311,N_20495,N_20952);
and U22312 (N_22312,N_21848,N_21070);
nand U22313 (N_22313,N_21990,N_20723);
nor U22314 (N_22314,N_20691,N_21760);
nor U22315 (N_22315,N_20162,N_20273);
or U22316 (N_22316,N_20040,N_20030);
or U22317 (N_22317,N_21378,N_21210);
nor U22318 (N_22318,N_21793,N_21514);
and U22319 (N_22319,N_20068,N_21081);
nand U22320 (N_22320,N_21852,N_21740);
nor U22321 (N_22321,N_21627,N_20924);
and U22322 (N_22322,N_21268,N_21961);
and U22323 (N_22323,N_20083,N_20796);
or U22324 (N_22324,N_20158,N_21959);
nand U22325 (N_22325,N_21344,N_21295);
or U22326 (N_22326,N_21256,N_20521);
and U22327 (N_22327,N_20605,N_21521);
nand U22328 (N_22328,N_21404,N_20835);
nand U22329 (N_22329,N_20323,N_20504);
and U22330 (N_22330,N_20765,N_21500);
and U22331 (N_22331,N_20772,N_20347);
nor U22332 (N_22332,N_21445,N_21395);
nand U22333 (N_22333,N_20553,N_21226);
and U22334 (N_22334,N_20168,N_21036);
nand U22335 (N_22335,N_21741,N_20237);
or U22336 (N_22336,N_21543,N_20132);
nand U22337 (N_22337,N_21842,N_21078);
and U22338 (N_22338,N_21379,N_21141);
or U22339 (N_22339,N_20412,N_20370);
nor U22340 (N_22340,N_21411,N_21569);
nor U22341 (N_22341,N_20821,N_20903);
or U22342 (N_22342,N_20870,N_20842);
nor U22343 (N_22343,N_21746,N_21840);
or U22344 (N_22344,N_20392,N_21731);
nand U22345 (N_22345,N_21187,N_21490);
and U22346 (N_22346,N_21386,N_21835);
and U22347 (N_22347,N_20559,N_21313);
or U22348 (N_22348,N_21257,N_20135);
or U22349 (N_22349,N_20119,N_21416);
or U22350 (N_22350,N_20919,N_20834);
and U22351 (N_22351,N_21998,N_21666);
nand U22352 (N_22352,N_21059,N_21281);
nand U22353 (N_22353,N_21049,N_21390);
or U22354 (N_22354,N_20242,N_21181);
nand U22355 (N_22355,N_21820,N_21539);
nor U22356 (N_22356,N_20364,N_21018);
or U22357 (N_22357,N_21818,N_21812);
and U22358 (N_22358,N_21664,N_20388);
and U22359 (N_22359,N_20863,N_20233);
nor U22360 (N_22360,N_21039,N_21589);
or U22361 (N_22361,N_20062,N_20871);
or U22362 (N_22362,N_20231,N_20152);
nor U22363 (N_22363,N_21794,N_21183);
nand U22364 (N_22364,N_20038,N_21504);
nand U22365 (N_22365,N_20783,N_21471);
and U22366 (N_22366,N_20538,N_20970);
nor U22367 (N_22367,N_20861,N_20279);
xor U22368 (N_22368,N_21367,N_20566);
or U22369 (N_22369,N_21649,N_20217);
nand U22370 (N_22370,N_20638,N_21947);
nand U22371 (N_22371,N_21674,N_21727);
or U22372 (N_22372,N_20543,N_21286);
and U22373 (N_22373,N_20447,N_20465);
nand U22374 (N_22374,N_20912,N_20900);
and U22375 (N_22375,N_20170,N_20439);
nand U22376 (N_22376,N_20376,N_20567);
nand U22377 (N_22377,N_21169,N_20429);
or U22378 (N_22378,N_21057,N_21525);
and U22379 (N_22379,N_20145,N_21321);
nand U22380 (N_22380,N_20998,N_21097);
or U22381 (N_22381,N_20212,N_21108);
nor U22382 (N_22382,N_20849,N_21997);
or U22383 (N_22383,N_21652,N_21035);
nor U22384 (N_22384,N_20056,N_21178);
or U22385 (N_22385,N_20905,N_20297);
nand U22386 (N_22386,N_20572,N_21269);
and U22387 (N_22387,N_20987,N_20243);
nor U22388 (N_22388,N_21459,N_20069);
nor U22389 (N_22389,N_20218,N_20806);
nor U22390 (N_22390,N_20602,N_20728);
or U22391 (N_22391,N_20532,N_21962);
nand U22392 (N_22392,N_21635,N_20276);
nand U22393 (N_22393,N_20530,N_21422);
and U22394 (N_22394,N_21975,N_21916);
nor U22395 (N_22395,N_20258,N_21939);
or U22396 (N_22396,N_21530,N_21242);
nor U22397 (N_22397,N_21346,N_20822);
xor U22398 (N_22398,N_20866,N_20522);
nand U22399 (N_22399,N_21682,N_21128);
or U22400 (N_22400,N_21162,N_20079);
and U22401 (N_22401,N_20725,N_20485);
nand U22402 (N_22402,N_21485,N_21247);
and U22403 (N_22403,N_21677,N_21212);
and U22404 (N_22404,N_20665,N_21120);
nand U22405 (N_22405,N_20470,N_21365);
or U22406 (N_22406,N_21522,N_21371);
and U22407 (N_22407,N_20383,N_21312);
and U22408 (N_22408,N_21756,N_20937);
nand U22409 (N_22409,N_20201,N_21201);
nand U22410 (N_22410,N_21115,N_20505);
nand U22411 (N_22411,N_20999,N_20182);
and U22412 (N_22412,N_20187,N_20535);
nand U22413 (N_22413,N_21012,N_20619);
or U22414 (N_22414,N_21815,N_20613);
nor U22415 (N_22415,N_21042,N_20731);
nor U22416 (N_22416,N_21239,N_20409);
nand U22417 (N_22417,N_20387,N_20916);
nand U22418 (N_22418,N_21573,N_20456);
and U22419 (N_22419,N_21347,N_20427);
or U22420 (N_22420,N_20721,N_20002);
nand U22421 (N_22421,N_20980,N_20374);
and U22422 (N_22422,N_20391,N_21050);
nor U22423 (N_22423,N_20889,N_21308);
and U22424 (N_22424,N_20264,N_20029);
and U22425 (N_22425,N_21200,N_20529);
nor U22426 (N_22426,N_20690,N_21228);
or U22427 (N_22427,N_21743,N_21173);
and U22428 (N_22428,N_21628,N_21636);
nor U22429 (N_22429,N_20882,N_20895);
or U22430 (N_22430,N_21327,N_21370);
nor U22431 (N_22431,N_20240,N_21134);
nand U22432 (N_22432,N_20337,N_20609);
nand U22433 (N_22433,N_20359,N_20063);
or U22434 (N_22434,N_21354,N_20901);
nor U22435 (N_22435,N_20280,N_21544);
nor U22436 (N_22436,N_21114,N_21685);
nand U22437 (N_22437,N_21444,N_21350);
nor U22438 (N_22438,N_20914,N_21074);
and U22439 (N_22439,N_20770,N_20053);
and U22440 (N_22440,N_20886,N_20894);
and U22441 (N_22441,N_21374,N_20281);
and U22442 (N_22442,N_21478,N_21443);
and U22443 (N_22443,N_21782,N_21083);
nor U22444 (N_22444,N_21025,N_21310);
xor U22445 (N_22445,N_20356,N_21538);
or U22446 (N_22446,N_20205,N_21875);
nand U22447 (N_22447,N_20073,N_20210);
and U22448 (N_22448,N_20750,N_20411);
nand U22449 (N_22449,N_20645,N_21616);
or U22450 (N_22450,N_20146,N_21197);
or U22451 (N_22451,N_21619,N_20873);
and U22452 (N_22452,N_20814,N_21213);
nor U22453 (N_22453,N_20137,N_21206);
nor U22454 (N_22454,N_20452,N_20403);
nand U22455 (N_22455,N_21454,N_20910);
nor U22456 (N_22456,N_20005,N_20965);
or U22457 (N_22457,N_20058,N_21868);
nand U22458 (N_22458,N_20165,N_20654);
nor U22459 (N_22459,N_21785,N_21795);
nor U22460 (N_22460,N_21862,N_20066);
nor U22461 (N_22461,N_20192,N_21161);
or U22462 (N_22462,N_20425,N_20071);
or U22463 (N_22463,N_21909,N_20488);
nand U22464 (N_22464,N_20751,N_21476);
xnor U22465 (N_22465,N_20117,N_21345);
nor U22466 (N_22466,N_21650,N_21858);
nand U22467 (N_22467,N_21887,N_21218);
nor U22468 (N_22468,N_20875,N_20982);
nor U22469 (N_22469,N_20597,N_21447);
and U22470 (N_22470,N_21273,N_20988);
nand U22471 (N_22471,N_20076,N_20339);
and U22472 (N_22472,N_20864,N_21670);
or U22473 (N_22473,N_21921,N_21701);
or U22474 (N_22474,N_21807,N_21575);
nand U22475 (N_22475,N_21817,N_21869);
or U22476 (N_22476,N_21608,N_20724);
and U22477 (N_22477,N_20278,N_21987);
nor U22478 (N_22478,N_21152,N_21254);
nor U22479 (N_22479,N_21918,N_21913);
nand U22480 (N_22480,N_21925,N_20008);
or U22481 (N_22481,N_20046,N_21092);
or U22482 (N_22482,N_20743,N_21566);
nor U22483 (N_22483,N_20386,N_20846);
xor U22484 (N_22484,N_21572,N_20340);
or U22485 (N_22485,N_20404,N_20232);
nor U22486 (N_22486,N_20112,N_20644);
or U22487 (N_22487,N_20782,N_21208);
nor U22488 (N_22488,N_21427,N_20784);
nor U22489 (N_22489,N_20123,N_20124);
nand U22490 (N_22490,N_20614,N_21709);
nor U22491 (N_22491,N_20313,N_21046);
and U22492 (N_22492,N_21695,N_21957);
or U22493 (N_22493,N_21583,N_21224);
and U22494 (N_22494,N_20496,N_21872);
and U22495 (N_22495,N_20000,N_21689);
or U22496 (N_22496,N_20322,N_21678);
or U22497 (N_22497,N_21407,N_21309);
or U22498 (N_22498,N_21238,N_21482);
or U22499 (N_22499,N_20445,N_21311);
nor U22500 (N_22500,N_21935,N_21617);
nor U22501 (N_22501,N_21610,N_20448);
and U22502 (N_22502,N_20295,N_21258);
nand U22503 (N_22503,N_20020,N_20877);
and U22504 (N_22504,N_20483,N_21992);
and U22505 (N_22505,N_21819,N_20081);
nor U22506 (N_22506,N_21941,N_20298);
or U22507 (N_22507,N_21122,N_20148);
nor U22508 (N_22508,N_20536,N_21542);
or U22509 (N_22509,N_20269,N_21372);
and U22510 (N_22510,N_21274,N_21004);
nor U22511 (N_22511,N_20779,N_20574);
nand U22512 (N_22512,N_20832,N_21851);
nand U22513 (N_22513,N_20157,N_21294);
and U22514 (N_22514,N_20037,N_21387);
and U22515 (N_22515,N_21148,N_20111);
and U22516 (N_22516,N_21209,N_20984);
or U22517 (N_22517,N_20953,N_21936);
nand U22518 (N_22518,N_20078,N_20402);
or U22519 (N_22519,N_21827,N_21506);
nand U22520 (N_22520,N_21629,N_20345);
and U22521 (N_22521,N_21675,N_20075);
xor U22522 (N_22522,N_21823,N_21079);
or U22523 (N_22523,N_20147,N_21419);
and U22524 (N_22524,N_20333,N_21302);
nor U22525 (N_22525,N_21030,N_20140);
xor U22526 (N_22526,N_21624,N_21948);
and U22527 (N_22527,N_20096,N_21879);
nor U22528 (N_22528,N_20351,N_21216);
nor U22529 (N_22529,N_21895,N_21773);
nand U22530 (N_22530,N_21021,N_21136);
nor U22531 (N_22531,N_21719,N_20697);
nand U22532 (N_22532,N_21565,N_21455);
or U22533 (N_22533,N_21420,N_20325);
nor U22534 (N_22534,N_20511,N_21692);
nor U22535 (N_22535,N_21752,N_21151);
and U22536 (N_22536,N_21943,N_21973);
or U22537 (N_22537,N_21547,N_20799);
nor U22538 (N_22538,N_21659,N_20003);
or U22539 (N_22539,N_20944,N_20661);
and U22540 (N_22540,N_20664,N_20507);
nor U22541 (N_22541,N_21956,N_20769);
nand U22542 (N_22542,N_21690,N_20473);
nor U22543 (N_22543,N_20328,N_20213);
nor U22544 (N_22544,N_20080,N_20143);
nand U22545 (N_22545,N_21955,N_21026);
and U22546 (N_22546,N_21974,N_20599);
nand U22547 (N_22547,N_21103,N_21594);
or U22548 (N_22548,N_21272,N_20195);
and U22549 (N_22549,N_20267,N_20432);
or U22550 (N_22550,N_20589,N_20467);
or U22551 (N_22551,N_20330,N_20787);
or U22552 (N_22552,N_20859,N_20776);
and U22553 (N_22553,N_21089,N_20142);
nor U22554 (N_22554,N_20130,N_20881);
nor U22555 (N_22555,N_21100,N_21339);
or U22556 (N_22556,N_21319,N_21501);
nor U22557 (N_22557,N_21687,N_20457);
or U22558 (N_22558,N_20015,N_20416);
or U22559 (N_22559,N_21597,N_20055);
nor U22560 (N_22560,N_21653,N_20106);
or U22561 (N_22561,N_21235,N_20720);
and U22562 (N_22562,N_20290,N_20520);
or U22563 (N_22563,N_21156,N_20922);
and U22564 (N_22564,N_21402,N_20936);
nand U22565 (N_22565,N_20164,N_20573);
nor U22566 (N_22566,N_21523,N_21007);
or U22567 (N_22567,N_20019,N_20180);
nor U22568 (N_22568,N_20365,N_21621);
and U22569 (N_22569,N_21877,N_21033);
nor U22570 (N_22570,N_21903,N_20869);
or U22571 (N_22571,N_20021,N_21211);
nor U22572 (N_22572,N_20194,N_21816);
or U22573 (N_22573,N_20515,N_20539);
nand U22574 (N_22574,N_20810,N_21278);
nand U22575 (N_22575,N_21150,N_20974);
nor U22576 (N_22576,N_21634,N_20266);
or U22577 (N_22577,N_21087,N_20758);
nand U22578 (N_22578,N_21072,N_20746);
nor U22579 (N_22579,N_21091,N_21179);
and U22580 (N_22580,N_20642,N_20014);
nand U22581 (N_22581,N_20986,N_21486);
nor U22582 (N_22582,N_21978,N_21641);
nand U22583 (N_22583,N_21930,N_21382);
and U22584 (N_22584,N_21805,N_20099);
nor U22585 (N_22585,N_21806,N_20598);
nor U22586 (N_22586,N_21069,N_21932);
and U22587 (N_22587,N_20957,N_20851);
and U22588 (N_22588,N_21736,N_20477);
nand U22589 (N_22589,N_20110,N_20631);
nand U22590 (N_22590,N_20042,N_21192);
or U22591 (N_22591,N_20315,N_21056);
or U22592 (N_22592,N_20805,N_21604);
or U22593 (N_22593,N_20054,N_20713);
nand U22594 (N_22594,N_20800,N_20643);
and U22595 (N_22595,N_20458,N_20379);
or U22596 (N_22596,N_20023,N_20480);
nor U22597 (N_22597,N_21977,N_21810);
xnor U22598 (N_22598,N_21963,N_20304);
nor U22599 (N_22599,N_21403,N_21300);
nor U22600 (N_22600,N_20317,N_20366);
or U22601 (N_22601,N_21999,N_20601);
nand U22602 (N_22602,N_20484,N_21062);
nor U22603 (N_22603,N_20742,N_21044);
nor U22604 (N_22604,N_20109,N_21774);
nand U22605 (N_22605,N_21298,N_21383);
nand U22606 (N_22606,N_21052,N_20191);
or U22607 (N_22607,N_20972,N_21065);
and U22608 (N_22608,N_21560,N_21177);
or U22609 (N_22609,N_20259,N_20097);
or U22610 (N_22610,N_21126,N_21364);
or U22611 (N_22611,N_20051,N_21225);
nand U22612 (N_22612,N_20993,N_21106);
nor U22613 (N_22613,N_21316,N_21591);
and U22614 (N_22614,N_20253,N_20122);
or U22615 (N_22615,N_20077,N_20121);
nor U22616 (N_22616,N_21663,N_21882);
nand U22617 (N_22617,N_21047,N_21651);
and U22618 (N_22618,N_20247,N_21157);
and U22619 (N_22619,N_21144,N_21555);
nand U22620 (N_22620,N_21017,N_21564);
or U22621 (N_22621,N_21775,N_20064);
nand U22622 (N_22622,N_20891,N_21578);
or U22623 (N_22623,N_20491,N_21777);
or U22624 (N_22624,N_20420,N_20082);
nand U22625 (N_22625,N_20733,N_20153);
or U22626 (N_22626,N_20088,N_20655);
nor U22627 (N_22627,N_20585,N_21118);
nor U22628 (N_22628,N_21116,N_21786);
nor U22629 (N_22629,N_20904,N_20289);
or U22630 (N_22630,N_21643,N_21381);
nor U22631 (N_22631,N_21304,N_20296);
and U22632 (N_22632,N_21898,N_20932);
or U22633 (N_22633,N_20131,N_20825);
xor U22634 (N_22634,N_21864,N_21117);
and U22635 (N_22635,N_20497,N_21531);
and U22636 (N_22636,N_20270,N_20888);
and U22637 (N_22637,N_20621,N_21570);
nand U22638 (N_22638,N_21182,N_21853);
or U22639 (N_22639,N_21844,N_21995);
xor U22640 (N_22640,N_21184,N_20824);
and U22641 (N_22641,N_20868,N_21814);
nand U22642 (N_22642,N_20450,N_20931);
nor U22643 (N_22643,N_20469,N_21541);
xnor U22644 (N_22644,N_20061,N_21549);
nor U22645 (N_22645,N_20568,N_20087);
and U22646 (N_22646,N_21532,N_21085);
and U22647 (N_22647,N_20823,N_21496);
nor U22648 (N_22648,N_21333,N_20261);
xnor U22649 (N_22649,N_21276,N_21606);
or U22650 (N_22650,N_21002,N_20571);
or U22651 (N_22651,N_21090,N_20985);
nor U22652 (N_22652,N_20583,N_21391);
nand U22653 (N_22653,N_20857,N_21414);
and U22654 (N_22654,N_20950,N_21904);
or U22655 (N_22655,N_20300,N_21163);
nand U22656 (N_22656,N_20514,N_20220);
or U22657 (N_22657,N_20335,N_21846);
nand U22658 (N_22658,N_20032,N_21832);
and U22659 (N_22659,N_21473,N_21194);
nand U22660 (N_22660,N_20813,N_21323);
nand U22661 (N_22661,N_20178,N_20706);
nand U22662 (N_22662,N_21084,N_21540);
nand U22663 (N_22663,N_21796,N_20414);
or U22664 (N_22664,N_20405,N_21626);
nor U22665 (N_22665,N_21392,N_21559);
and U22666 (N_22666,N_20060,N_20215);
and U22667 (N_22667,N_20672,N_21188);
and U22668 (N_22668,N_20969,N_21421);
nor U22669 (N_22669,N_20978,N_20744);
and U22670 (N_22670,N_20935,N_20327);
and U22671 (N_22671,N_20549,N_20225);
or U22672 (N_22672,N_20506,N_21099);
nor U22673 (N_22673,N_20141,N_20606);
and U22674 (N_22674,N_21856,N_21086);
and U22675 (N_22675,N_21934,N_20265);
nand U22676 (N_22676,N_20209,N_21076);
and U22677 (N_22677,N_21684,N_21691);
nand U22678 (N_22678,N_21718,N_20303);
and U22679 (N_22679,N_20398,N_20671);
nand U22680 (N_22680,N_21789,N_20839);
and U22681 (N_22681,N_20501,N_21061);
nand U22682 (N_22682,N_20381,N_20207);
and U22683 (N_22683,N_21369,N_21885);
nor U22684 (N_22684,N_21112,N_20311);
nand U22685 (N_22685,N_20045,N_20577);
and U22686 (N_22686,N_20624,N_21767);
nor U22687 (N_22687,N_21438,N_21038);
nor U22688 (N_22688,N_20627,N_20637);
and U22689 (N_22689,N_21505,N_20177);
nand U22690 (N_22690,N_21906,N_21071);
xor U22691 (N_22691,N_21655,N_20156);
or U22692 (N_22692,N_20262,N_20768);
nor U22693 (N_22693,N_20994,N_20658);
and U22694 (N_22694,N_20785,N_21171);
nor U22695 (N_22695,N_20360,N_21784);
nor U22696 (N_22696,N_20626,N_21186);
nand U22697 (N_22697,N_21241,N_20586);
xnor U22698 (N_22698,N_20234,N_20593);
and U22699 (N_22699,N_20695,N_21306);
nand U22700 (N_22700,N_20848,N_20729);
and U22701 (N_22701,N_20833,N_21728);
or U22702 (N_22702,N_20118,N_21865);
and U22703 (N_22703,N_20855,N_20884);
nor U22704 (N_22704,N_20717,N_20206);
nor U22705 (N_22705,N_21140,N_20108);
nand U22706 (N_22706,N_21593,N_21073);
or U22707 (N_22707,N_21464,N_21668);
and U22708 (N_22708,N_20004,N_21263);
nand U22709 (N_22709,N_20732,N_20436);
xor U22710 (N_22710,N_21001,N_21357);
nand U22711 (N_22711,N_20084,N_21020);
or U22712 (N_22712,N_21230,N_20677);
or U22713 (N_22713,N_20594,N_21011);
and U22714 (N_22714,N_20669,N_21602);
nor U22715 (N_22715,N_20285,N_20039);
nand U22716 (N_22716,N_21536,N_21396);
and U22717 (N_22717,N_21797,N_21563);
or U22718 (N_22718,N_20272,N_21401);
or U22719 (N_22719,N_21270,N_21640);
and U22720 (N_22720,N_21788,N_20139);
xnor U22721 (N_22721,N_21494,N_21244);
or U22722 (N_22722,N_20010,N_21094);
or U22723 (N_22723,N_20471,N_20332);
nor U22724 (N_22724,N_21271,N_20518);
nand U22725 (N_22725,N_21991,N_20730);
nor U22726 (N_22726,N_20375,N_20771);
nand U22727 (N_22727,N_20686,N_20883);
or U22728 (N_22728,N_20500,N_21623);
or U22729 (N_22729,N_21804,N_21609);
nand U22730 (N_22730,N_20827,N_21064);
nor U22731 (N_22731,N_20326,N_21088);
and U22732 (N_22732,N_20578,N_20949);
and U22733 (N_22733,N_21686,N_21822);
nand U22734 (N_22734,N_20867,N_20434);
nand U22735 (N_22735,N_21240,N_20575);
and U22736 (N_22736,N_20927,N_21359);
and U22737 (N_22737,N_20781,N_20100);
nor U22738 (N_22738,N_20384,N_20091);
or U22739 (N_22739,N_21720,N_20588);
nand U22740 (N_22740,N_20909,N_21562);
xnor U22741 (N_22741,N_20104,N_20738);
nand U22742 (N_22742,N_20517,N_21880);
nand U22743 (N_22743,N_21145,N_20816);
or U22744 (N_22744,N_20149,N_20006);
nor U22745 (N_22745,N_20763,N_21722);
nand U22746 (N_22746,N_20245,N_21528);
and U22747 (N_22747,N_21131,N_21949);
and U22748 (N_22748,N_21981,N_20094);
nand U22749 (N_22749,N_21759,N_21405);
nor U22750 (N_22750,N_21669,N_21334);
or U22751 (N_22751,N_20555,N_20920);
nand U22752 (N_22752,N_20525,N_21590);
or U22753 (N_22753,N_21436,N_21923);
nor U22754 (N_22754,N_21060,N_20293);
nand U22755 (N_22755,N_21253,N_21878);
nor U22756 (N_22756,N_21460,N_20216);
nor U22757 (N_22757,N_20461,N_20902);
nor U22758 (N_22758,N_20034,N_20692);
nand U22759 (N_22759,N_21458,N_21825);
or U22760 (N_22760,N_20044,N_20951);
nor U22761 (N_22761,N_21612,N_21576);
nor U22762 (N_22762,N_20338,N_21180);
and U22763 (N_22763,N_21279,N_20459);
and U22764 (N_22764,N_20983,N_21964);
and U22765 (N_22765,N_20214,N_20017);
and U22766 (N_22766,N_20451,N_20134);
or U22767 (N_22767,N_20976,N_20228);
and U22768 (N_22768,N_20230,N_20354);
nor U22769 (N_22769,N_21900,N_20455);
or U22770 (N_22770,N_21393,N_21679);
nand U22771 (N_22771,N_21193,N_21753);
nor U22772 (N_22772,N_21077,N_21529);
or U22773 (N_22773,N_21550,N_21873);
nand U22774 (N_22774,N_21676,N_20946);
nor U22775 (N_22775,N_20336,N_21781);
or U22776 (N_22776,N_21233,N_21190);
nand U22777 (N_22777,N_21618,N_20067);
and U22778 (N_22778,N_20125,N_21412);
nor U22779 (N_22779,N_21330,N_21368);
or U22780 (N_22780,N_20837,N_21132);
or U22781 (N_22781,N_21960,N_21706);
xnor U22782 (N_22782,N_20804,N_21214);
or U22783 (N_22783,N_21337,N_20962);
or U22784 (N_22784,N_20498,N_20652);
nand U22785 (N_22785,N_21929,N_21658);
nand U22786 (N_22786,N_21220,N_20926);
and U22787 (N_22787,N_20400,N_21857);
or U22788 (N_22788,N_20942,N_20858);
nor U22789 (N_22789,N_21979,N_21792);
and U22790 (N_22790,N_21982,N_21726);
or U22791 (N_22791,N_21245,N_21765);
nand U22792 (N_22792,N_21515,N_20331);
nand U22793 (N_22793,N_21014,N_20659);
nor U22794 (N_22794,N_21596,N_20701);
or U22795 (N_22795,N_20879,N_20576);
nor U22796 (N_22796,N_21467,N_20749);
and U22797 (N_22797,N_21894,N_21217);
or U22798 (N_22798,N_21889,N_20341);
nand U22799 (N_22799,N_20523,N_20703);
or U22800 (N_22800,N_20175,N_20239);
or U22801 (N_22801,N_21426,N_20560);
or U22802 (N_22802,N_21915,N_21110);
nand U22803 (N_22803,N_20817,N_21189);
nor U22804 (N_22804,N_21567,N_21988);
nor U22805 (N_22805,N_20128,N_20862);
and U22806 (N_22806,N_21450,N_21758);
nor U22807 (N_22807,N_20126,N_21763);
and U22808 (N_22808,N_20136,N_21527);
nand U22809 (N_22809,N_20841,N_20600);
nor U22810 (N_22810,N_20929,N_21380);
and U22811 (N_22811,N_20836,N_20587);
nor U22812 (N_22812,N_20487,N_20089);
nor U22813 (N_22813,N_20688,N_20550);
and U22814 (N_22814,N_21483,N_20314);
nor U22815 (N_22815,N_21697,N_21362);
nor U22816 (N_22816,N_21409,N_20291);
nor U22817 (N_22817,N_21275,N_20222);
nor U22818 (N_22818,N_21953,N_21410);
or U22819 (N_22819,N_21700,N_20294);
and U22820 (N_22820,N_20646,N_20792);
or U22821 (N_22821,N_20737,N_20840);
nand U22822 (N_22822,N_20844,N_21142);
or U22823 (N_22823,N_20399,N_21461);
nor U22824 (N_22824,N_20189,N_21463);
and U22825 (N_22825,N_21983,N_20299);
nand U22826 (N_22826,N_20898,N_21508);
nor U22827 (N_22827,N_21694,N_21841);
nor U22828 (N_22828,N_21384,N_21910);
xor U22829 (N_22829,N_21824,N_20558);
or U22830 (N_22830,N_21863,N_20421);
nor U22831 (N_22831,N_20961,N_21725);
xor U22832 (N_22832,N_21248,N_20887);
nand U22833 (N_22833,N_20401,N_21809);
nand U22834 (N_22834,N_20203,N_21874);
and U22835 (N_22835,N_20657,N_21143);
nor U22836 (N_22836,N_21029,N_21579);
nor U22837 (N_22837,N_20454,N_20997);
and U22838 (N_22838,N_20959,N_20502);
or U22839 (N_22839,N_20138,N_21448);
and U22840 (N_22840,N_21707,N_21940);
or U22841 (N_22841,N_20757,N_20305);
and U22842 (N_22842,N_20711,N_21022);
or U22843 (N_22843,N_21282,N_21891);
nor U22844 (N_22844,N_20682,N_21749);
or U22845 (N_22845,N_21908,N_20660);
nand U22846 (N_22846,N_20410,N_21933);
and U22847 (N_22847,N_21780,N_21375);
and U22848 (N_22848,N_21888,N_20633);
or U22849 (N_22849,N_20797,N_20443);
nand U22850 (N_22850,N_21901,N_20036);
or U22851 (N_22851,N_20086,N_20127);
or U22852 (N_22852,N_20615,N_21830);
nor U22853 (N_22853,N_21199,N_20854);
or U22854 (N_22854,N_20611,N_21468);
nand U22855 (N_22855,N_21475,N_20610);
and U22856 (N_22856,N_21801,N_21512);
nor U22857 (N_22857,N_21236,N_20460);
and U22858 (N_22858,N_20395,N_21477);
nor U22859 (N_22859,N_21320,N_21967);
nand U22860 (N_22860,N_21284,N_20408);
and U22861 (N_22861,N_21434,N_20791);
or U22862 (N_22862,N_20818,N_20246);
and U22863 (N_22863,N_20181,N_21232);
nor U22864 (N_22864,N_21340,N_21871);
or U22865 (N_22865,N_21107,N_21976);
or U22866 (N_22866,N_21024,N_20250);
and U22867 (N_22867,N_20954,N_20634);
xor U22868 (N_22868,N_21620,N_21601);
nand U22869 (N_22869,N_20394,N_20235);
nand U22870 (N_22870,N_20651,N_21168);
and U22871 (N_22871,N_21928,N_21750);
nand U22872 (N_22872,N_21876,N_21783);
or U22873 (N_22873,N_20722,N_21299);
nor U22874 (N_22874,N_21552,N_20348);
nand U22875 (N_22875,N_21301,N_20085);
and U22876 (N_22876,N_21996,N_20968);
and U22877 (N_22877,N_21845,N_21493);
or U22878 (N_22878,N_21893,N_20016);
nand U22879 (N_22879,N_20878,N_20406);
and U22880 (N_22880,N_21764,N_21798);
and U22881 (N_22881,N_21377,N_20979);
nand U22882 (N_22882,N_21510,N_20441);
and U22883 (N_22883,N_20662,N_21938);
nor U22884 (N_22884,N_20009,N_21648);
or U22885 (N_22885,N_21985,N_20479);
or U22886 (N_22886,N_20989,N_21584);
or U22887 (N_22887,N_20908,N_20933);
or U22888 (N_22888,N_21479,N_20151);
nand U22889 (N_22889,N_21102,N_21125);
nand U22890 (N_22890,N_20095,N_21582);
nand U22891 (N_22891,N_21082,N_20324);
or U22892 (N_22892,N_20260,N_21551);
nor U22893 (N_22893,N_20284,N_21266);
and U22894 (N_22894,N_21661,N_20115);
and U22895 (N_22895,N_21487,N_21511);
nor U22896 (N_22896,N_20035,N_20357);
or U22897 (N_22897,N_21332,N_21702);
nand U22898 (N_22898,N_21647,N_20880);
nor U22899 (N_22899,N_21546,N_20718);
or U22900 (N_22900,N_20727,N_20582);
or U22901 (N_22901,N_20371,N_21119);
nor U22902 (N_22902,N_21329,N_20282);
nand U22903 (N_22903,N_21826,N_21633);
or U22904 (N_22904,N_20393,N_21474);
nand U22905 (N_22905,N_21954,N_20012);
nor U22906 (N_22906,N_20435,N_21415);
nor U22907 (N_22907,N_21424,N_21571);
or U22908 (N_22908,N_21453,N_21336);
or U22909 (N_22909,N_21732,N_20955);
or U22910 (N_22910,N_21705,N_20710);
nor U22911 (N_22911,N_20226,N_21139);
or U22912 (N_22912,N_21614,N_21839);
nor U22913 (N_22913,N_21413,N_20628);
or U22914 (N_22914,N_20120,N_20358);
or U22915 (N_22915,N_20907,N_20640);
nor U22916 (N_22916,N_21492,N_20534);
nor U22917 (N_22917,N_21662,N_20449);
nor U22918 (N_22918,N_21881,N_20372);
and U22919 (N_22919,N_21261,N_21945);
nand U22920 (N_22920,N_21821,N_20494);
nand U22921 (N_22921,N_21779,N_20777);
or U22922 (N_22922,N_20188,N_20967);
nor U22923 (N_22923,N_21829,N_21587);
or U22924 (N_22924,N_21104,N_21129);
or U22925 (N_22925,N_21745,N_20251);
and U22926 (N_22926,N_21554,N_20026);
or U22927 (N_22927,N_21293,N_20618);
and U22928 (N_22928,N_21755,N_21397);
nor U22929 (N_22929,N_21703,N_21533);
or U22930 (N_22930,N_20185,N_20478);
nand U22931 (N_22931,N_20385,N_20831);
nand U22932 (N_22932,N_21215,N_21098);
nor U22933 (N_22933,N_20674,N_21406);
nand U22934 (N_22934,N_21297,N_21096);
nand U22935 (N_22935,N_21660,N_20945);
and U22936 (N_22936,N_20747,N_20254);
nand U22937 (N_22937,N_20202,N_20596);
or U22938 (N_22938,N_20590,N_20349);
or U22939 (N_22939,N_20407,N_20580);
and U22940 (N_22940,N_20702,N_21837);
or U22941 (N_22941,N_21325,N_21680);
nand U22942 (N_22942,N_20113,N_21353);
nand U22943 (N_22943,N_21041,N_20318);
and U22944 (N_22944,N_21495,N_20755);
or U22945 (N_22945,N_20679,N_20368);
or U22946 (N_22946,N_21031,N_20428);
and U22947 (N_22947,N_21221,N_20764);
nand U22948 (N_22948,N_21630,N_20440);
nand U22949 (N_22949,N_20562,N_20683);
nand U22950 (N_22950,N_20561,N_21639);
or U22951 (N_22951,N_20774,N_20991);
and U22952 (N_22952,N_20767,N_20287);
and U22953 (N_22953,N_21423,N_21734);
and U22954 (N_22954,N_20464,N_21331);
nor U22955 (N_22955,N_21611,N_20941);
nand U22956 (N_22956,N_21598,N_20172);
and U22957 (N_22957,N_21195,N_20024);
nor U22958 (N_22958,N_20377,N_20939);
nor U22959 (N_22959,N_21009,N_20437);
nor U22960 (N_22960,N_20668,N_21717);
and U22961 (N_22961,N_20754,N_20355);
nor U22962 (N_22962,N_21317,N_21952);
or U22963 (N_22963,N_21237,N_20329);
nand U22964 (N_22964,N_20719,N_21710);
nand U22965 (N_22965,N_21048,N_20971);
nand U22966 (N_22966,N_20244,N_21335);
nand U22967 (N_22967,N_21130,N_21800);
or U22968 (N_22968,N_20564,N_21534);
nor U22969 (N_22969,N_21008,N_21338);
or U22970 (N_22970,N_20708,N_21834);
or U22971 (N_22971,N_20830,N_21642);
and U22972 (N_22972,N_20321,N_20221);
nor U22973 (N_22973,N_20541,N_21326);
nor U22974 (N_22974,N_20636,N_21341);
or U22975 (N_22975,N_20801,N_20263);
and U22976 (N_22976,N_21466,N_21509);
nand U22977 (N_22977,N_21164,N_20570);
and U22978 (N_22978,N_21400,N_21439);
nand U22979 (N_22979,N_21324,N_21469);
or U22980 (N_22980,N_21919,N_20663);
nor U22981 (N_22981,N_21388,N_20173);
nor U22982 (N_22982,N_21748,N_21155);
or U22983 (N_22983,N_21681,N_21811);
nor U22984 (N_22984,N_21277,N_21432);
nor U22985 (N_22985,N_20617,N_21799);
and U22986 (N_22986,N_20196,N_21260);
nor U22987 (N_22987,N_20684,N_20947);
nand U22988 (N_22988,N_21503,N_21328);
and U22989 (N_22989,N_21937,N_20444);
nand U22990 (N_22990,N_21599,N_20956);
or U22991 (N_22991,N_21488,N_21866);
nand U22992 (N_22992,N_20249,N_21175);
and U22993 (N_22993,N_20788,N_20028);
and U22994 (N_22994,N_20025,N_21859);
nor U22995 (N_22995,N_21762,N_21886);
xor U22996 (N_22996,N_20292,N_20680);
nor U22997 (N_22997,N_21343,N_20308);
nand U22998 (N_22998,N_21958,N_20361);
nand U22999 (N_22999,N_20204,N_21721);
and U23000 (N_23000,N_20371,N_21206);
or U23001 (N_23001,N_21114,N_21605);
nand U23002 (N_23002,N_21382,N_21919);
or U23003 (N_23003,N_20236,N_20783);
and U23004 (N_23004,N_20454,N_20942);
nor U23005 (N_23005,N_20762,N_21220);
or U23006 (N_23006,N_21860,N_21929);
xor U23007 (N_23007,N_20575,N_20564);
or U23008 (N_23008,N_21662,N_21106);
or U23009 (N_23009,N_21067,N_21063);
nor U23010 (N_23010,N_20561,N_21326);
and U23011 (N_23011,N_20662,N_20308);
xnor U23012 (N_23012,N_21965,N_21509);
nor U23013 (N_23013,N_21877,N_21921);
and U23014 (N_23014,N_21046,N_20506);
and U23015 (N_23015,N_21541,N_20718);
or U23016 (N_23016,N_20282,N_21919);
or U23017 (N_23017,N_21184,N_21358);
and U23018 (N_23018,N_21330,N_20556);
nand U23019 (N_23019,N_20770,N_21735);
or U23020 (N_23020,N_21416,N_21618);
nor U23021 (N_23021,N_20425,N_20195);
and U23022 (N_23022,N_20980,N_20399);
nor U23023 (N_23023,N_21568,N_20475);
and U23024 (N_23024,N_20702,N_20234);
nand U23025 (N_23025,N_20372,N_20374);
nor U23026 (N_23026,N_20829,N_20039);
nand U23027 (N_23027,N_20508,N_20643);
nand U23028 (N_23028,N_20058,N_20825);
nor U23029 (N_23029,N_20520,N_21396);
nand U23030 (N_23030,N_21419,N_20724);
or U23031 (N_23031,N_21627,N_21562);
or U23032 (N_23032,N_21771,N_21106);
or U23033 (N_23033,N_20567,N_20545);
nor U23034 (N_23034,N_20205,N_20756);
nor U23035 (N_23035,N_21791,N_21849);
nor U23036 (N_23036,N_20149,N_20815);
or U23037 (N_23037,N_21175,N_20610);
nand U23038 (N_23038,N_20783,N_20660);
nand U23039 (N_23039,N_21723,N_21352);
and U23040 (N_23040,N_20236,N_20354);
or U23041 (N_23041,N_21322,N_21583);
nand U23042 (N_23042,N_21884,N_20034);
and U23043 (N_23043,N_20661,N_20045);
nor U23044 (N_23044,N_20573,N_21947);
and U23045 (N_23045,N_21970,N_21381);
nand U23046 (N_23046,N_21245,N_21800);
nor U23047 (N_23047,N_21061,N_20608);
nand U23048 (N_23048,N_20404,N_20426);
and U23049 (N_23049,N_20983,N_20595);
or U23050 (N_23050,N_20678,N_20207);
and U23051 (N_23051,N_21553,N_21507);
nor U23052 (N_23052,N_21697,N_20938);
and U23053 (N_23053,N_21716,N_21528);
nand U23054 (N_23054,N_20577,N_21006);
nor U23055 (N_23055,N_20233,N_20028);
or U23056 (N_23056,N_20091,N_20082);
nor U23057 (N_23057,N_21925,N_20136);
nor U23058 (N_23058,N_20344,N_21050);
nand U23059 (N_23059,N_20437,N_20644);
nor U23060 (N_23060,N_21575,N_20927);
or U23061 (N_23061,N_20010,N_20263);
xor U23062 (N_23062,N_20604,N_21258);
nand U23063 (N_23063,N_21921,N_21177);
or U23064 (N_23064,N_21747,N_21410);
and U23065 (N_23065,N_21012,N_20411);
nand U23066 (N_23066,N_21185,N_20041);
or U23067 (N_23067,N_20295,N_20769);
and U23068 (N_23068,N_20641,N_20170);
nor U23069 (N_23069,N_21743,N_21807);
and U23070 (N_23070,N_21301,N_21011);
nor U23071 (N_23071,N_20445,N_21174);
and U23072 (N_23072,N_20172,N_20818);
or U23073 (N_23073,N_20024,N_20857);
or U23074 (N_23074,N_21368,N_20817);
or U23075 (N_23075,N_21410,N_20138);
nor U23076 (N_23076,N_20397,N_21535);
or U23077 (N_23077,N_20047,N_21827);
nor U23078 (N_23078,N_20538,N_20219);
or U23079 (N_23079,N_21114,N_20234);
and U23080 (N_23080,N_21241,N_20620);
nor U23081 (N_23081,N_20171,N_21491);
and U23082 (N_23082,N_21424,N_20020);
or U23083 (N_23083,N_20647,N_20952);
or U23084 (N_23084,N_20132,N_20592);
nor U23085 (N_23085,N_21065,N_21678);
nor U23086 (N_23086,N_21057,N_21887);
or U23087 (N_23087,N_21302,N_20768);
nand U23088 (N_23088,N_20521,N_21890);
and U23089 (N_23089,N_20599,N_21551);
or U23090 (N_23090,N_20848,N_21734);
or U23091 (N_23091,N_21158,N_21697);
or U23092 (N_23092,N_21031,N_21908);
or U23093 (N_23093,N_20470,N_21784);
or U23094 (N_23094,N_20407,N_21812);
and U23095 (N_23095,N_21052,N_20776);
nand U23096 (N_23096,N_20523,N_21604);
nand U23097 (N_23097,N_21442,N_20924);
and U23098 (N_23098,N_21032,N_20743);
nor U23099 (N_23099,N_20551,N_21326);
or U23100 (N_23100,N_21022,N_21485);
and U23101 (N_23101,N_21556,N_20642);
nor U23102 (N_23102,N_21473,N_20061);
and U23103 (N_23103,N_20241,N_20772);
and U23104 (N_23104,N_21993,N_20400);
nand U23105 (N_23105,N_20631,N_20421);
or U23106 (N_23106,N_21465,N_20504);
or U23107 (N_23107,N_20085,N_20927);
and U23108 (N_23108,N_21663,N_21134);
or U23109 (N_23109,N_20288,N_21841);
nand U23110 (N_23110,N_20493,N_21563);
nand U23111 (N_23111,N_21481,N_20519);
nand U23112 (N_23112,N_21864,N_21844);
or U23113 (N_23113,N_20065,N_21994);
nor U23114 (N_23114,N_21702,N_20871);
xnor U23115 (N_23115,N_20756,N_21644);
and U23116 (N_23116,N_20543,N_20054);
nand U23117 (N_23117,N_21333,N_20497);
or U23118 (N_23118,N_20078,N_20107);
and U23119 (N_23119,N_21167,N_21697);
or U23120 (N_23120,N_21622,N_20286);
or U23121 (N_23121,N_20179,N_20899);
nand U23122 (N_23122,N_20215,N_21917);
nor U23123 (N_23123,N_21619,N_20097);
and U23124 (N_23124,N_20012,N_20362);
or U23125 (N_23125,N_21520,N_20833);
and U23126 (N_23126,N_20339,N_20591);
and U23127 (N_23127,N_21102,N_20759);
nand U23128 (N_23128,N_21204,N_21510);
xnor U23129 (N_23129,N_20575,N_20489);
nor U23130 (N_23130,N_21225,N_20702);
nor U23131 (N_23131,N_20709,N_20538);
or U23132 (N_23132,N_21699,N_21532);
nor U23133 (N_23133,N_20173,N_21662);
nand U23134 (N_23134,N_20777,N_21203);
or U23135 (N_23135,N_20310,N_21384);
and U23136 (N_23136,N_21273,N_20024);
or U23137 (N_23137,N_20684,N_21983);
nor U23138 (N_23138,N_21565,N_21525);
nand U23139 (N_23139,N_20153,N_21712);
and U23140 (N_23140,N_21864,N_20251);
nand U23141 (N_23141,N_21742,N_20040);
nand U23142 (N_23142,N_21716,N_20591);
and U23143 (N_23143,N_20625,N_21864);
and U23144 (N_23144,N_20752,N_20807);
or U23145 (N_23145,N_21016,N_21895);
and U23146 (N_23146,N_20346,N_21888);
and U23147 (N_23147,N_21042,N_20789);
or U23148 (N_23148,N_20825,N_21569);
or U23149 (N_23149,N_21939,N_20388);
xnor U23150 (N_23150,N_21566,N_21094);
nand U23151 (N_23151,N_20961,N_21559);
nor U23152 (N_23152,N_21134,N_20196);
or U23153 (N_23153,N_20597,N_20391);
nand U23154 (N_23154,N_21587,N_21302);
nor U23155 (N_23155,N_21140,N_21822);
or U23156 (N_23156,N_20638,N_21432);
xor U23157 (N_23157,N_20590,N_20250);
or U23158 (N_23158,N_21380,N_21993);
nor U23159 (N_23159,N_20599,N_21031);
nand U23160 (N_23160,N_21017,N_21967);
nand U23161 (N_23161,N_20224,N_21471);
and U23162 (N_23162,N_20420,N_20075);
or U23163 (N_23163,N_20729,N_21637);
nor U23164 (N_23164,N_20116,N_21901);
or U23165 (N_23165,N_20653,N_20528);
nor U23166 (N_23166,N_21051,N_20604);
or U23167 (N_23167,N_20014,N_20083);
nand U23168 (N_23168,N_20523,N_20796);
xor U23169 (N_23169,N_21238,N_20583);
and U23170 (N_23170,N_20016,N_21640);
and U23171 (N_23171,N_21079,N_21572);
or U23172 (N_23172,N_21766,N_20624);
or U23173 (N_23173,N_20766,N_21403);
and U23174 (N_23174,N_20034,N_21084);
or U23175 (N_23175,N_20922,N_20389);
nand U23176 (N_23176,N_21985,N_20367);
or U23177 (N_23177,N_21327,N_20859);
and U23178 (N_23178,N_20248,N_20528);
nand U23179 (N_23179,N_21267,N_21341);
nand U23180 (N_23180,N_21803,N_20198);
nor U23181 (N_23181,N_20902,N_21561);
or U23182 (N_23182,N_20745,N_21682);
or U23183 (N_23183,N_20467,N_20708);
nand U23184 (N_23184,N_21675,N_20025);
nor U23185 (N_23185,N_20937,N_21864);
nand U23186 (N_23186,N_21914,N_20825);
and U23187 (N_23187,N_21865,N_20737);
nor U23188 (N_23188,N_21118,N_21317);
nor U23189 (N_23189,N_20774,N_20463);
nor U23190 (N_23190,N_20193,N_21134);
or U23191 (N_23191,N_21863,N_21498);
nand U23192 (N_23192,N_21927,N_21628);
nor U23193 (N_23193,N_20649,N_21352);
nand U23194 (N_23194,N_21636,N_20936);
or U23195 (N_23195,N_21321,N_21446);
and U23196 (N_23196,N_21960,N_21701);
and U23197 (N_23197,N_20287,N_21769);
or U23198 (N_23198,N_20523,N_20410);
or U23199 (N_23199,N_21465,N_20298);
xor U23200 (N_23200,N_20953,N_20503);
or U23201 (N_23201,N_21639,N_20551);
and U23202 (N_23202,N_20928,N_21511);
nor U23203 (N_23203,N_21891,N_21188);
nand U23204 (N_23204,N_21338,N_21040);
nand U23205 (N_23205,N_21594,N_21574);
nand U23206 (N_23206,N_20797,N_21760);
nand U23207 (N_23207,N_20957,N_21908);
and U23208 (N_23208,N_21063,N_20986);
and U23209 (N_23209,N_20622,N_21433);
nor U23210 (N_23210,N_20955,N_20403);
nand U23211 (N_23211,N_21804,N_20113);
and U23212 (N_23212,N_21219,N_21570);
xor U23213 (N_23213,N_20519,N_21594);
and U23214 (N_23214,N_21562,N_21536);
and U23215 (N_23215,N_20097,N_20629);
and U23216 (N_23216,N_21390,N_21723);
nor U23217 (N_23217,N_20729,N_21438);
or U23218 (N_23218,N_21933,N_20135);
or U23219 (N_23219,N_20629,N_21447);
and U23220 (N_23220,N_21338,N_20001);
or U23221 (N_23221,N_21864,N_20188);
and U23222 (N_23222,N_20188,N_21155);
nand U23223 (N_23223,N_21986,N_20775);
nand U23224 (N_23224,N_20706,N_20166);
nor U23225 (N_23225,N_20641,N_21725);
nand U23226 (N_23226,N_20330,N_21537);
or U23227 (N_23227,N_20294,N_21430);
or U23228 (N_23228,N_21359,N_21873);
or U23229 (N_23229,N_20495,N_20574);
nor U23230 (N_23230,N_21073,N_20489);
nor U23231 (N_23231,N_21954,N_21990);
and U23232 (N_23232,N_20003,N_21299);
and U23233 (N_23233,N_20376,N_21611);
nor U23234 (N_23234,N_21153,N_21284);
nor U23235 (N_23235,N_21295,N_21860);
and U23236 (N_23236,N_21939,N_21394);
nor U23237 (N_23237,N_21412,N_20891);
xor U23238 (N_23238,N_20170,N_20740);
and U23239 (N_23239,N_20882,N_21611);
or U23240 (N_23240,N_21011,N_20360);
nor U23241 (N_23241,N_21899,N_21970);
nand U23242 (N_23242,N_20437,N_21074);
and U23243 (N_23243,N_20522,N_21898);
nand U23244 (N_23244,N_21529,N_21501);
nor U23245 (N_23245,N_21049,N_21169);
or U23246 (N_23246,N_20367,N_20167);
nor U23247 (N_23247,N_21808,N_21611);
xor U23248 (N_23248,N_21640,N_21850);
or U23249 (N_23249,N_21647,N_21325);
and U23250 (N_23250,N_20339,N_21765);
nand U23251 (N_23251,N_20823,N_20425);
xnor U23252 (N_23252,N_21647,N_20035);
nor U23253 (N_23253,N_21138,N_21366);
xor U23254 (N_23254,N_20799,N_20802);
xor U23255 (N_23255,N_20876,N_21121);
or U23256 (N_23256,N_20457,N_20902);
nand U23257 (N_23257,N_21750,N_20402);
nand U23258 (N_23258,N_21104,N_20165);
nand U23259 (N_23259,N_20605,N_20214);
or U23260 (N_23260,N_21136,N_20604);
or U23261 (N_23261,N_20758,N_21948);
nand U23262 (N_23262,N_20549,N_21175);
and U23263 (N_23263,N_20780,N_21530);
nand U23264 (N_23264,N_21817,N_21067);
nor U23265 (N_23265,N_20442,N_20816);
or U23266 (N_23266,N_21434,N_20110);
nand U23267 (N_23267,N_21031,N_21473);
and U23268 (N_23268,N_21902,N_20087);
or U23269 (N_23269,N_21082,N_20224);
xnor U23270 (N_23270,N_21341,N_20892);
nor U23271 (N_23271,N_20461,N_21118);
or U23272 (N_23272,N_21546,N_20074);
nor U23273 (N_23273,N_21018,N_21564);
nor U23274 (N_23274,N_21517,N_20265);
or U23275 (N_23275,N_21746,N_20250);
nand U23276 (N_23276,N_20340,N_20764);
or U23277 (N_23277,N_21409,N_21825);
nor U23278 (N_23278,N_21202,N_21352);
or U23279 (N_23279,N_21264,N_21833);
and U23280 (N_23280,N_21618,N_20303);
nand U23281 (N_23281,N_20519,N_20115);
nor U23282 (N_23282,N_21798,N_20987);
xor U23283 (N_23283,N_20502,N_21647);
or U23284 (N_23284,N_20994,N_20630);
and U23285 (N_23285,N_20120,N_21160);
and U23286 (N_23286,N_21957,N_21791);
nor U23287 (N_23287,N_21033,N_21471);
or U23288 (N_23288,N_21773,N_20357);
xor U23289 (N_23289,N_20272,N_21615);
and U23290 (N_23290,N_21694,N_21145);
or U23291 (N_23291,N_20781,N_20924);
nor U23292 (N_23292,N_20065,N_21802);
nor U23293 (N_23293,N_21180,N_21958);
nand U23294 (N_23294,N_20740,N_20480);
and U23295 (N_23295,N_21413,N_20453);
nand U23296 (N_23296,N_21926,N_20586);
nor U23297 (N_23297,N_21817,N_20967);
xnor U23298 (N_23298,N_21632,N_21407);
and U23299 (N_23299,N_20278,N_21743);
nand U23300 (N_23300,N_20186,N_20571);
and U23301 (N_23301,N_20050,N_21436);
nand U23302 (N_23302,N_20762,N_20099);
or U23303 (N_23303,N_20668,N_20124);
and U23304 (N_23304,N_20836,N_20614);
and U23305 (N_23305,N_21443,N_21156);
nor U23306 (N_23306,N_21836,N_20937);
or U23307 (N_23307,N_21999,N_20086);
and U23308 (N_23308,N_20434,N_20971);
nor U23309 (N_23309,N_21688,N_21707);
nor U23310 (N_23310,N_20525,N_21430);
nand U23311 (N_23311,N_21648,N_20752);
and U23312 (N_23312,N_21506,N_20786);
nor U23313 (N_23313,N_20158,N_20815);
and U23314 (N_23314,N_20929,N_21589);
and U23315 (N_23315,N_20374,N_20359);
and U23316 (N_23316,N_21672,N_20218);
and U23317 (N_23317,N_21233,N_20507);
nand U23318 (N_23318,N_21831,N_20567);
and U23319 (N_23319,N_21404,N_21694);
or U23320 (N_23320,N_20522,N_20822);
nor U23321 (N_23321,N_21723,N_20673);
nor U23322 (N_23322,N_20675,N_21860);
xor U23323 (N_23323,N_20918,N_21911);
nor U23324 (N_23324,N_20235,N_20206);
nand U23325 (N_23325,N_20775,N_20330);
nor U23326 (N_23326,N_20678,N_21124);
nor U23327 (N_23327,N_21735,N_21886);
nand U23328 (N_23328,N_21378,N_20010);
nor U23329 (N_23329,N_21221,N_21239);
nand U23330 (N_23330,N_20938,N_21671);
and U23331 (N_23331,N_20992,N_20922);
or U23332 (N_23332,N_20269,N_21755);
or U23333 (N_23333,N_21864,N_21936);
or U23334 (N_23334,N_20466,N_21616);
or U23335 (N_23335,N_20932,N_21430);
nand U23336 (N_23336,N_20339,N_21524);
nand U23337 (N_23337,N_20685,N_20317);
xnor U23338 (N_23338,N_21896,N_21336);
nor U23339 (N_23339,N_21781,N_21992);
nor U23340 (N_23340,N_20212,N_21425);
and U23341 (N_23341,N_20942,N_21638);
or U23342 (N_23342,N_21553,N_21049);
or U23343 (N_23343,N_21722,N_20094);
nand U23344 (N_23344,N_21497,N_21945);
and U23345 (N_23345,N_21293,N_20559);
and U23346 (N_23346,N_20247,N_20738);
nand U23347 (N_23347,N_20080,N_21509);
and U23348 (N_23348,N_21304,N_20355);
and U23349 (N_23349,N_20997,N_20884);
or U23350 (N_23350,N_21365,N_21428);
nand U23351 (N_23351,N_21681,N_21390);
and U23352 (N_23352,N_20506,N_21630);
nand U23353 (N_23353,N_20229,N_21513);
nand U23354 (N_23354,N_20305,N_21609);
and U23355 (N_23355,N_21439,N_20907);
or U23356 (N_23356,N_21679,N_21714);
nor U23357 (N_23357,N_20381,N_21697);
or U23358 (N_23358,N_20754,N_21361);
nand U23359 (N_23359,N_20982,N_21418);
nor U23360 (N_23360,N_21535,N_20843);
and U23361 (N_23361,N_21318,N_20595);
or U23362 (N_23362,N_21778,N_20792);
nand U23363 (N_23363,N_21148,N_21241);
nand U23364 (N_23364,N_20392,N_20411);
nand U23365 (N_23365,N_20312,N_21746);
xnor U23366 (N_23366,N_21277,N_21065);
nand U23367 (N_23367,N_20786,N_20710);
nor U23368 (N_23368,N_21195,N_21200);
xor U23369 (N_23369,N_20381,N_20258);
nand U23370 (N_23370,N_21234,N_21001);
and U23371 (N_23371,N_20568,N_21578);
or U23372 (N_23372,N_21006,N_21005);
nand U23373 (N_23373,N_21140,N_21099);
or U23374 (N_23374,N_20702,N_20264);
and U23375 (N_23375,N_21599,N_20698);
nand U23376 (N_23376,N_21675,N_20861);
or U23377 (N_23377,N_20748,N_20835);
xor U23378 (N_23378,N_21974,N_20498);
nand U23379 (N_23379,N_20742,N_21307);
nor U23380 (N_23380,N_21807,N_21182);
xnor U23381 (N_23381,N_21962,N_20701);
or U23382 (N_23382,N_20902,N_20425);
nor U23383 (N_23383,N_20189,N_20539);
or U23384 (N_23384,N_21604,N_21701);
nor U23385 (N_23385,N_21084,N_20962);
and U23386 (N_23386,N_21661,N_20359);
nand U23387 (N_23387,N_21118,N_21811);
xor U23388 (N_23388,N_21302,N_20571);
nor U23389 (N_23389,N_20096,N_21661);
nand U23390 (N_23390,N_21199,N_20090);
and U23391 (N_23391,N_21206,N_21308);
nor U23392 (N_23392,N_21745,N_21775);
or U23393 (N_23393,N_21385,N_20899);
or U23394 (N_23394,N_21739,N_20000);
and U23395 (N_23395,N_20204,N_21476);
or U23396 (N_23396,N_21489,N_21531);
or U23397 (N_23397,N_20942,N_21757);
nand U23398 (N_23398,N_21641,N_21876);
and U23399 (N_23399,N_21040,N_21991);
nand U23400 (N_23400,N_20769,N_20153);
nor U23401 (N_23401,N_21882,N_20766);
and U23402 (N_23402,N_21679,N_20925);
or U23403 (N_23403,N_20472,N_21425);
nand U23404 (N_23404,N_20707,N_20266);
or U23405 (N_23405,N_21512,N_21655);
nor U23406 (N_23406,N_20438,N_20371);
nand U23407 (N_23407,N_20724,N_20131);
nand U23408 (N_23408,N_21798,N_21538);
nor U23409 (N_23409,N_21681,N_20077);
and U23410 (N_23410,N_20861,N_21428);
or U23411 (N_23411,N_20125,N_20613);
xor U23412 (N_23412,N_20241,N_21613);
and U23413 (N_23413,N_20669,N_21199);
nor U23414 (N_23414,N_21653,N_20530);
and U23415 (N_23415,N_21898,N_21492);
nor U23416 (N_23416,N_20513,N_20338);
or U23417 (N_23417,N_21564,N_21859);
or U23418 (N_23418,N_20967,N_21366);
nand U23419 (N_23419,N_21449,N_20096);
nand U23420 (N_23420,N_21811,N_20714);
or U23421 (N_23421,N_20454,N_20895);
or U23422 (N_23422,N_21661,N_21880);
nand U23423 (N_23423,N_20871,N_20033);
nor U23424 (N_23424,N_21484,N_20417);
and U23425 (N_23425,N_21055,N_21508);
and U23426 (N_23426,N_21207,N_20994);
or U23427 (N_23427,N_21568,N_21730);
or U23428 (N_23428,N_20500,N_21065);
or U23429 (N_23429,N_21868,N_20786);
nor U23430 (N_23430,N_21714,N_20351);
nor U23431 (N_23431,N_21923,N_21592);
or U23432 (N_23432,N_20542,N_20422);
nor U23433 (N_23433,N_20741,N_20666);
and U23434 (N_23434,N_21900,N_21950);
nor U23435 (N_23435,N_21462,N_20369);
nand U23436 (N_23436,N_20786,N_21639);
xnor U23437 (N_23437,N_21521,N_21026);
or U23438 (N_23438,N_21905,N_20220);
and U23439 (N_23439,N_21279,N_21698);
nor U23440 (N_23440,N_20721,N_21594);
and U23441 (N_23441,N_21779,N_20305);
nor U23442 (N_23442,N_20216,N_21743);
nand U23443 (N_23443,N_21720,N_20467);
or U23444 (N_23444,N_20241,N_20291);
and U23445 (N_23445,N_20742,N_21712);
nand U23446 (N_23446,N_20662,N_20011);
xnor U23447 (N_23447,N_21104,N_21314);
or U23448 (N_23448,N_21752,N_21791);
nor U23449 (N_23449,N_20513,N_21901);
or U23450 (N_23450,N_20072,N_20471);
xor U23451 (N_23451,N_20799,N_20178);
or U23452 (N_23452,N_21937,N_21983);
xnor U23453 (N_23453,N_20478,N_21544);
and U23454 (N_23454,N_21092,N_21579);
or U23455 (N_23455,N_21095,N_20951);
or U23456 (N_23456,N_20232,N_20348);
and U23457 (N_23457,N_20396,N_20443);
or U23458 (N_23458,N_20569,N_20697);
and U23459 (N_23459,N_21509,N_21967);
or U23460 (N_23460,N_21850,N_20539);
or U23461 (N_23461,N_21563,N_21700);
and U23462 (N_23462,N_21033,N_20634);
or U23463 (N_23463,N_21962,N_20246);
nand U23464 (N_23464,N_21982,N_20456);
xor U23465 (N_23465,N_21345,N_21508);
nand U23466 (N_23466,N_20826,N_21710);
nand U23467 (N_23467,N_21852,N_20330);
and U23468 (N_23468,N_20477,N_20093);
and U23469 (N_23469,N_20234,N_21957);
nand U23470 (N_23470,N_21827,N_21409);
nand U23471 (N_23471,N_20123,N_21349);
and U23472 (N_23472,N_21664,N_20224);
and U23473 (N_23473,N_21344,N_20698);
nor U23474 (N_23474,N_21095,N_21910);
or U23475 (N_23475,N_21349,N_21078);
or U23476 (N_23476,N_20415,N_21233);
nand U23477 (N_23477,N_21999,N_21862);
nand U23478 (N_23478,N_21199,N_21229);
and U23479 (N_23479,N_20264,N_21627);
or U23480 (N_23480,N_21333,N_21115);
and U23481 (N_23481,N_21926,N_21227);
nand U23482 (N_23482,N_20827,N_20767);
or U23483 (N_23483,N_20169,N_20286);
nand U23484 (N_23484,N_21812,N_21484);
or U23485 (N_23485,N_21786,N_21145);
nor U23486 (N_23486,N_21980,N_21208);
and U23487 (N_23487,N_21963,N_21194);
nor U23488 (N_23488,N_20267,N_21070);
nor U23489 (N_23489,N_21677,N_21421);
or U23490 (N_23490,N_21062,N_21020);
and U23491 (N_23491,N_20813,N_20871);
and U23492 (N_23492,N_20297,N_21274);
nand U23493 (N_23493,N_20068,N_20298);
nor U23494 (N_23494,N_20195,N_21769);
and U23495 (N_23495,N_21300,N_20699);
or U23496 (N_23496,N_20876,N_21583);
and U23497 (N_23497,N_20276,N_21328);
and U23498 (N_23498,N_20235,N_21340);
or U23499 (N_23499,N_20928,N_21515);
nand U23500 (N_23500,N_20980,N_21743);
nor U23501 (N_23501,N_21526,N_21517);
nor U23502 (N_23502,N_21081,N_20683);
and U23503 (N_23503,N_20352,N_20732);
or U23504 (N_23504,N_21253,N_21434);
nand U23505 (N_23505,N_21096,N_20312);
and U23506 (N_23506,N_21716,N_20896);
and U23507 (N_23507,N_21714,N_20275);
nor U23508 (N_23508,N_20829,N_21001);
or U23509 (N_23509,N_20860,N_21177);
and U23510 (N_23510,N_21744,N_21295);
and U23511 (N_23511,N_20810,N_20999);
nor U23512 (N_23512,N_21223,N_21350);
nor U23513 (N_23513,N_21551,N_21319);
nand U23514 (N_23514,N_20737,N_21538);
nand U23515 (N_23515,N_20048,N_21639);
nor U23516 (N_23516,N_20681,N_20727);
or U23517 (N_23517,N_20659,N_21045);
nand U23518 (N_23518,N_20659,N_20374);
nand U23519 (N_23519,N_21545,N_21046);
xor U23520 (N_23520,N_21828,N_20309);
nor U23521 (N_23521,N_20165,N_21727);
nor U23522 (N_23522,N_20995,N_20768);
nand U23523 (N_23523,N_21459,N_20608);
and U23524 (N_23524,N_20696,N_21794);
nand U23525 (N_23525,N_20349,N_21454);
and U23526 (N_23526,N_21391,N_21448);
or U23527 (N_23527,N_21750,N_21540);
or U23528 (N_23528,N_20682,N_21680);
and U23529 (N_23529,N_21308,N_20379);
and U23530 (N_23530,N_21986,N_20991);
nand U23531 (N_23531,N_21457,N_21209);
xor U23532 (N_23532,N_21434,N_20676);
nand U23533 (N_23533,N_20591,N_21122);
and U23534 (N_23534,N_21556,N_20690);
and U23535 (N_23535,N_21968,N_21480);
nor U23536 (N_23536,N_20527,N_20116);
and U23537 (N_23537,N_21003,N_21138);
nand U23538 (N_23538,N_20422,N_20097);
or U23539 (N_23539,N_20352,N_20033);
and U23540 (N_23540,N_20452,N_20749);
nand U23541 (N_23541,N_20485,N_21965);
and U23542 (N_23542,N_20554,N_20592);
or U23543 (N_23543,N_20701,N_20413);
nor U23544 (N_23544,N_20661,N_20425);
or U23545 (N_23545,N_20763,N_20727);
nand U23546 (N_23546,N_21455,N_21575);
and U23547 (N_23547,N_20698,N_20559);
nand U23548 (N_23548,N_21427,N_20681);
nor U23549 (N_23549,N_20093,N_21002);
xnor U23550 (N_23550,N_20580,N_20386);
nor U23551 (N_23551,N_21677,N_20116);
nand U23552 (N_23552,N_21811,N_20009);
or U23553 (N_23553,N_21644,N_21670);
and U23554 (N_23554,N_21058,N_21978);
or U23555 (N_23555,N_21025,N_20536);
nand U23556 (N_23556,N_20884,N_20910);
nor U23557 (N_23557,N_20210,N_21275);
nand U23558 (N_23558,N_20957,N_21353);
nand U23559 (N_23559,N_21893,N_20680);
or U23560 (N_23560,N_20083,N_21499);
nor U23561 (N_23561,N_21262,N_21371);
and U23562 (N_23562,N_20487,N_21489);
nand U23563 (N_23563,N_20739,N_21690);
and U23564 (N_23564,N_20993,N_20393);
and U23565 (N_23565,N_21776,N_20354);
nand U23566 (N_23566,N_21869,N_20984);
nor U23567 (N_23567,N_20372,N_20380);
xor U23568 (N_23568,N_21486,N_21176);
nand U23569 (N_23569,N_21037,N_20953);
xor U23570 (N_23570,N_21797,N_20111);
nor U23571 (N_23571,N_20254,N_21450);
or U23572 (N_23572,N_21874,N_21437);
or U23573 (N_23573,N_20159,N_21033);
and U23574 (N_23574,N_20187,N_20899);
nor U23575 (N_23575,N_21463,N_20542);
and U23576 (N_23576,N_21116,N_21241);
xnor U23577 (N_23577,N_21012,N_21757);
and U23578 (N_23578,N_21103,N_20801);
and U23579 (N_23579,N_21246,N_20760);
xor U23580 (N_23580,N_20831,N_21659);
and U23581 (N_23581,N_20467,N_20045);
nand U23582 (N_23582,N_20287,N_21997);
nor U23583 (N_23583,N_20434,N_20691);
or U23584 (N_23584,N_20707,N_20427);
and U23585 (N_23585,N_21893,N_21363);
nand U23586 (N_23586,N_20575,N_20015);
and U23587 (N_23587,N_21600,N_21886);
or U23588 (N_23588,N_20694,N_20529);
or U23589 (N_23589,N_20051,N_20575);
nand U23590 (N_23590,N_20188,N_21506);
xnor U23591 (N_23591,N_21053,N_20933);
nor U23592 (N_23592,N_20339,N_20528);
nand U23593 (N_23593,N_20814,N_20861);
nand U23594 (N_23594,N_20221,N_21089);
nand U23595 (N_23595,N_21546,N_21713);
nand U23596 (N_23596,N_21190,N_21077);
nor U23597 (N_23597,N_20870,N_20595);
or U23598 (N_23598,N_20901,N_20139);
nor U23599 (N_23599,N_20705,N_20533);
and U23600 (N_23600,N_20117,N_21745);
nor U23601 (N_23601,N_20207,N_20655);
nor U23602 (N_23602,N_21054,N_21398);
or U23603 (N_23603,N_21856,N_20072);
nor U23604 (N_23604,N_20389,N_20959);
and U23605 (N_23605,N_20843,N_21772);
nor U23606 (N_23606,N_21730,N_20479);
or U23607 (N_23607,N_20373,N_21085);
nor U23608 (N_23608,N_21956,N_20454);
and U23609 (N_23609,N_20312,N_20225);
and U23610 (N_23610,N_21125,N_20116);
nand U23611 (N_23611,N_21352,N_20753);
and U23612 (N_23612,N_21396,N_21711);
and U23613 (N_23613,N_21528,N_21784);
xor U23614 (N_23614,N_20285,N_20548);
nand U23615 (N_23615,N_20059,N_21084);
nand U23616 (N_23616,N_21486,N_20174);
nor U23617 (N_23617,N_21602,N_20414);
nor U23618 (N_23618,N_20883,N_20285);
or U23619 (N_23619,N_21766,N_21031);
nand U23620 (N_23620,N_21131,N_20713);
xnor U23621 (N_23621,N_20758,N_20291);
nand U23622 (N_23622,N_20642,N_21277);
nand U23623 (N_23623,N_21454,N_20357);
nand U23624 (N_23624,N_21237,N_20947);
nand U23625 (N_23625,N_20301,N_20356);
or U23626 (N_23626,N_20498,N_21010);
or U23627 (N_23627,N_21482,N_20037);
or U23628 (N_23628,N_20913,N_21685);
or U23629 (N_23629,N_20591,N_20763);
or U23630 (N_23630,N_20776,N_20091);
and U23631 (N_23631,N_20636,N_20902);
and U23632 (N_23632,N_21048,N_21277);
xnor U23633 (N_23633,N_20505,N_20234);
and U23634 (N_23634,N_20028,N_21025);
xor U23635 (N_23635,N_21299,N_20395);
or U23636 (N_23636,N_20931,N_21454);
nand U23637 (N_23637,N_21291,N_20987);
or U23638 (N_23638,N_20456,N_21651);
or U23639 (N_23639,N_20228,N_20595);
or U23640 (N_23640,N_21471,N_21053);
nand U23641 (N_23641,N_21679,N_20526);
nor U23642 (N_23642,N_21810,N_20849);
nand U23643 (N_23643,N_20359,N_20313);
or U23644 (N_23644,N_21666,N_20756);
nor U23645 (N_23645,N_20985,N_21564);
nor U23646 (N_23646,N_21210,N_21811);
or U23647 (N_23647,N_21199,N_20309);
or U23648 (N_23648,N_20781,N_21867);
nand U23649 (N_23649,N_21406,N_20086);
nor U23650 (N_23650,N_20200,N_21156);
or U23651 (N_23651,N_21987,N_21557);
xnor U23652 (N_23652,N_20353,N_20112);
nor U23653 (N_23653,N_20768,N_21801);
nor U23654 (N_23654,N_20662,N_21438);
or U23655 (N_23655,N_21608,N_21265);
nor U23656 (N_23656,N_21501,N_20394);
and U23657 (N_23657,N_21713,N_21952);
nor U23658 (N_23658,N_21721,N_21973);
and U23659 (N_23659,N_21214,N_20576);
and U23660 (N_23660,N_21315,N_20002);
nand U23661 (N_23661,N_20140,N_20937);
nor U23662 (N_23662,N_20095,N_20391);
nand U23663 (N_23663,N_21420,N_21184);
nor U23664 (N_23664,N_20952,N_21375);
nand U23665 (N_23665,N_20514,N_20673);
nand U23666 (N_23666,N_21317,N_20792);
and U23667 (N_23667,N_21927,N_20860);
nand U23668 (N_23668,N_20668,N_20155);
or U23669 (N_23669,N_20968,N_21515);
and U23670 (N_23670,N_20510,N_20982);
or U23671 (N_23671,N_20990,N_20263);
nor U23672 (N_23672,N_21110,N_20786);
nand U23673 (N_23673,N_21053,N_21016);
or U23674 (N_23674,N_20534,N_21733);
and U23675 (N_23675,N_21079,N_21321);
and U23676 (N_23676,N_21724,N_20878);
nor U23677 (N_23677,N_20053,N_21470);
and U23678 (N_23678,N_20797,N_21510);
and U23679 (N_23679,N_20482,N_20970);
and U23680 (N_23680,N_20032,N_21433);
and U23681 (N_23681,N_20817,N_21053);
nand U23682 (N_23682,N_20472,N_21912);
and U23683 (N_23683,N_20028,N_20967);
or U23684 (N_23684,N_20612,N_21062);
nand U23685 (N_23685,N_20403,N_21169);
or U23686 (N_23686,N_21180,N_21930);
or U23687 (N_23687,N_21455,N_21004);
xnor U23688 (N_23688,N_21370,N_20232);
and U23689 (N_23689,N_21355,N_21640);
and U23690 (N_23690,N_21047,N_20874);
and U23691 (N_23691,N_20235,N_21516);
and U23692 (N_23692,N_20033,N_21873);
and U23693 (N_23693,N_20598,N_21465);
or U23694 (N_23694,N_20793,N_20710);
nor U23695 (N_23695,N_21169,N_20482);
nor U23696 (N_23696,N_21524,N_21782);
or U23697 (N_23697,N_21065,N_21533);
or U23698 (N_23698,N_21931,N_20938);
and U23699 (N_23699,N_21544,N_21591);
or U23700 (N_23700,N_21634,N_21069);
nand U23701 (N_23701,N_21236,N_20879);
nor U23702 (N_23702,N_21974,N_20784);
nor U23703 (N_23703,N_20290,N_21787);
nand U23704 (N_23704,N_20086,N_21250);
nor U23705 (N_23705,N_20462,N_20701);
nand U23706 (N_23706,N_20184,N_20803);
or U23707 (N_23707,N_20638,N_21440);
and U23708 (N_23708,N_21164,N_21713);
or U23709 (N_23709,N_20202,N_20773);
nor U23710 (N_23710,N_20605,N_21524);
nand U23711 (N_23711,N_21175,N_20294);
or U23712 (N_23712,N_20932,N_20056);
or U23713 (N_23713,N_20463,N_20817);
or U23714 (N_23714,N_21970,N_21661);
and U23715 (N_23715,N_20288,N_20356);
nor U23716 (N_23716,N_20194,N_20918);
or U23717 (N_23717,N_20636,N_20848);
nor U23718 (N_23718,N_20227,N_21242);
and U23719 (N_23719,N_21264,N_20052);
or U23720 (N_23720,N_20469,N_20498);
and U23721 (N_23721,N_20062,N_21709);
or U23722 (N_23722,N_21228,N_20775);
nor U23723 (N_23723,N_20834,N_20442);
nor U23724 (N_23724,N_20132,N_20347);
and U23725 (N_23725,N_21519,N_20883);
or U23726 (N_23726,N_20861,N_20318);
nand U23727 (N_23727,N_20652,N_20092);
and U23728 (N_23728,N_21735,N_21506);
or U23729 (N_23729,N_20034,N_21352);
and U23730 (N_23730,N_20784,N_20113);
nand U23731 (N_23731,N_21161,N_21952);
nand U23732 (N_23732,N_21583,N_20283);
nand U23733 (N_23733,N_21351,N_20728);
and U23734 (N_23734,N_20116,N_21662);
and U23735 (N_23735,N_21754,N_21140);
or U23736 (N_23736,N_21461,N_20871);
and U23737 (N_23737,N_21635,N_21039);
nand U23738 (N_23738,N_20610,N_20194);
or U23739 (N_23739,N_20764,N_20091);
and U23740 (N_23740,N_20015,N_20574);
or U23741 (N_23741,N_21873,N_20385);
nor U23742 (N_23742,N_20311,N_21949);
nor U23743 (N_23743,N_21767,N_20581);
nand U23744 (N_23744,N_20119,N_20975);
and U23745 (N_23745,N_21246,N_21427);
or U23746 (N_23746,N_21424,N_21691);
and U23747 (N_23747,N_21425,N_21652);
and U23748 (N_23748,N_20683,N_20075);
nor U23749 (N_23749,N_20791,N_21101);
nor U23750 (N_23750,N_20036,N_20564);
or U23751 (N_23751,N_20201,N_20002);
or U23752 (N_23752,N_20256,N_21071);
nand U23753 (N_23753,N_21662,N_20457);
or U23754 (N_23754,N_20649,N_21372);
or U23755 (N_23755,N_20930,N_20072);
nor U23756 (N_23756,N_20363,N_20530);
nand U23757 (N_23757,N_20919,N_21983);
nand U23758 (N_23758,N_20441,N_20783);
or U23759 (N_23759,N_21589,N_20942);
or U23760 (N_23760,N_21711,N_20224);
nand U23761 (N_23761,N_21906,N_21217);
or U23762 (N_23762,N_21856,N_20384);
and U23763 (N_23763,N_20274,N_20518);
nor U23764 (N_23764,N_20454,N_20710);
and U23765 (N_23765,N_21623,N_21238);
and U23766 (N_23766,N_20484,N_21556);
and U23767 (N_23767,N_20063,N_21405);
nand U23768 (N_23768,N_21986,N_21836);
nand U23769 (N_23769,N_20390,N_21618);
nand U23770 (N_23770,N_21407,N_21328);
nor U23771 (N_23771,N_21099,N_20784);
or U23772 (N_23772,N_21630,N_21823);
nor U23773 (N_23773,N_21342,N_21989);
nor U23774 (N_23774,N_20191,N_20153);
nand U23775 (N_23775,N_20776,N_21963);
or U23776 (N_23776,N_20606,N_20907);
nor U23777 (N_23777,N_21294,N_21299);
and U23778 (N_23778,N_20750,N_20365);
and U23779 (N_23779,N_20556,N_20546);
nor U23780 (N_23780,N_20830,N_21536);
or U23781 (N_23781,N_21763,N_21281);
or U23782 (N_23782,N_20520,N_21752);
and U23783 (N_23783,N_20264,N_20522);
nand U23784 (N_23784,N_20274,N_21092);
or U23785 (N_23785,N_21785,N_20512);
nor U23786 (N_23786,N_21098,N_20500);
and U23787 (N_23787,N_20811,N_21839);
and U23788 (N_23788,N_20116,N_20951);
and U23789 (N_23789,N_21868,N_21395);
nand U23790 (N_23790,N_20050,N_21172);
and U23791 (N_23791,N_21116,N_21404);
nand U23792 (N_23792,N_21127,N_20305);
nor U23793 (N_23793,N_20322,N_21521);
and U23794 (N_23794,N_21416,N_20718);
or U23795 (N_23795,N_20038,N_20198);
and U23796 (N_23796,N_20699,N_21945);
or U23797 (N_23797,N_21772,N_21409);
and U23798 (N_23798,N_21730,N_21549);
or U23799 (N_23799,N_21701,N_21903);
or U23800 (N_23800,N_21739,N_20949);
xor U23801 (N_23801,N_21792,N_20954);
nand U23802 (N_23802,N_20394,N_20643);
nand U23803 (N_23803,N_21986,N_21351);
nor U23804 (N_23804,N_21511,N_21720);
xnor U23805 (N_23805,N_21959,N_20890);
nand U23806 (N_23806,N_21120,N_20434);
nor U23807 (N_23807,N_20401,N_21378);
nor U23808 (N_23808,N_21375,N_21654);
nand U23809 (N_23809,N_21239,N_20386);
or U23810 (N_23810,N_20553,N_21196);
or U23811 (N_23811,N_21104,N_20258);
nor U23812 (N_23812,N_20839,N_20311);
and U23813 (N_23813,N_20166,N_20096);
nand U23814 (N_23814,N_20828,N_20493);
and U23815 (N_23815,N_20359,N_20400);
or U23816 (N_23816,N_20732,N_20549);
or U23817 (N_23817,N_20998,N_20833);
and U23818 (N_23818,N_21832,N_21287);
or U23819 (N_23819,N_21240,N_21211);
xnor U23820 (N_23820,N_21838,N_20438);
nand U23821 (N_23821,N_21570,N_21812);
or U23822 (N_23822,N_20703,N_20330);
nand U23823 (N_23823,N_20556,N_20457);
nor U23824 (N_23824,N_21498,N_20312);
nor U23825 (N_23825,N_21258,N_21073);
and U23826 (N_23826,N_21571,N_21666);
or U23827 (N_23827,N_20547,N_21962);
or U23828 (N_23828,N_21155,N_20760);
and U23829 (N_23829,N_20572,N_21311);
nor U23830 (N_23830,N_21921,N_20841);
nand U23831 (N_23831,N_21099,N_20625);
nand U23832 (N_23832,N_20272,N_20843);
or U23833 (N_23833,N_21949,N_20017);
and U23834 (N_23834,N_20309,N_21439);
nand U23835 (N_23835,N_21770,N_21101);
and U23836 (N_23836,N_21208,N_20271);
and U23837 (N_23837,N_21444,N_21077);
nand U23838 (N_23838,N_20783,N_21601);
nor U23839 (N_23839,N_20731,N_21034);
nand U23840 (N_23840,N_21188,N_21806);
and U23841 (N_23841,N_20929,N_21330);
nor U23842 (N_23842,N_20709,N_20860);
nand U23843 (N_23843,N_21266,N_21989);
nand U23844 (N_23844,N_21099,N_21963);
nand U23845 (N_23845,N_20547,N_20976);
or U23846 (N_23846,N_20161,N_21181);
and U23847 (N_23847,N_21980,N_20181);
nor U23848 (N_23848,N_20744,N_20400);
nand U23849 (N_23849,N_21196,N_21644);
or U23850 (N_23850,N_21225,N_20271);
nor U23851 (N_23851,N_21951,N_21361);
or U23852 (N_23852,N_20142,N_20609);
nor U23853 (N_23853,N_21719,N_21335);
xnor U23854 (N_23854,N_20958,N_20630);
or U23855 (N_23855,N_21101,N_20756);
nor U23856 (N_23856,N_21076,N_20871);
or U23857 (N_23857,N_21429,N_21569);
and U23858 (N_23858,N_20123,N_20125);
or U23859 (N_23859,N_21608,N_20106);
nand U23860 (N_23860,N_21070,N_20493);
nand U23861 (N_23861,N_21444,N_20106);
nor U23862 (N_23862,N_21996,N_20843);
nand U23863 (N_23863,N_21797,N_21006);
and U23864 (N_23864,N_20405,N_20228);
nand U23865 (N_23865,N_20587,N_20928);
nand U23866 (N_23866,N_21130,N_21492);
or U23867 (N_23867,N_21923,N_20363);
and U23868 (N_23868,N_20619,N_20355);
nor U23869 (N_23869,N_21769,N_20103);
nand U23870 (N_23870,N_20104,N_21007);
and U23871 (N_23871,N_21043,N_21495);
xnor U23872 (N_23872,N_20711,N_20356);
and U23873 (N_23873,N_20198,N_21852);
nand U23874 (N_23874,N_21437,N_20111);
and U23875 (N_23875,N_20159,N_21565);
or U23876 (N_23876,N_21964,N_21940);
or U23877 (N_23877,N_20423,N_21044);
nor U23878 (N_23878,N_21010,N_20976);
xnor U23879 (N_23879,N_20848,N_20182);
and U23880 (N_23880,N_21534,N_20582);
nand U23881 (N_23881,N_20020,N_20460);
nor U23882 (N_23882,N_21644,N_21311);
nand U23883 (N_23883,N_21094,N_20004);
and U23884 (N_23884,N_21843,N_21072);
and U23885 (N_23885,N_21194,N_21185);
nor U23886 (N_23886,N_20069,N_21655);
and U23887 (N_23887,N_20660,N_21627);
and U23888 (N_23888,N_20341,N_20065);
nand U23889 (N_23889,N_20613,N_21252);
nand U23890 (N_23890,N_20107,N_21369);
nor U23891 (N_23891,N_21907,N_21704);
or U23892 (N_23892,N_21872,N_20898);
or U23893 (N_23893,N_20819,N_20503);
and U23894 (N_23894,N_20176,N_20264);
nand U23895 (N_23895,N_20037,N_21370);
and U23896 (N_23896,N_21227,N_21928);
nor U23897 (N_23897,N_21972,N_21119);
nand U23898 (N_23898,N_21940,N_21332);
or U23899 (N_23899,N_20155,N_21385);
nor U23900 (N_23900,N_20481,N_21318);
nor U23901 (N_23901,N_20022,N_20981);
nor U23902 (N_23902,N_20149,N_21769);
or U23903 (N_23903,N_20585,N_20959);
or U23904 (N_23904,N_20477,N_20472);
and U23905 (N_23905,N_20648,N_21161);
or U23906 (N_23906,N_21834,N_20261);
and U23907 (N_23907,N_21893,N_21297);
nor U23908 (N_23908,N_21908,N_20136);
nor U23909 (N_23909,N_21780,N_20236);
or U23910 (N_23910,N_21253,N_21470);
nor U23911 (N_23911,N_20706,N_21674);
nand U23912 (N_23912,N_20349,N_20863);
and U23913 (N_23913,N_20581,N_20035);
or U23914 (N_23914,N_21966,N_20052);
nor U23915 (N_23915,N_20878,N_21307);
nand U23916 (N_23916,N_20819,N_21056);
or U23917 (N_23917,N_21660,N_20693);
or U23918 (N_23918,N_21868,N_20759);
or U23919 (N_23919,N_21912,N_20661);
or U23920 (N_23920,N_20143,N_20349);
nor U23921 (N_23921,N_20916,N_21434);
and U23922 (N_23922,N_21854,N_21353);
or U23923 (N_23923,N_20220,N_21916);
or U23924 (N_23924,N_21691,N_21869);
or U23925 (N_23925,N_21435,N_20531);
nand U23926 (N_23926,N_21509,N_21814);
and U23927 (N_23927,N_20334,N_20740);
and U23928 (N_23928,N_21867,N_20808);
nor U23929 (N_23929,N_21655,N_20073);
nand U23930 (N_23930,N_21897,N_20419);
or U23931 (N_23931,N_21041,N_21914);
or U23932 (N_23932,N_21097,N_20113);
nand U23933 (N_23933,N_20857,N_21251);
nand U23934 (N_23934,N_20132,N_21588);
nand U23935 (N_23935,N_20294,N_20980);
nand U23936 (N_23936,N_21785,N_20878);
or U23937 (N_23937,N_20165,N_21028);
or U23938 (N_23938,N_21951,N_20031);
nand U23939 (N_23939,N_20851,N_21134);
or U23940 (N_23940,N_20753,N_20356);
nand U23941 (N_23941,N_20349,N_21742);
and U23942 (N_23942,N_21644,N_20684);
and U23943 (N_23943,N_21407,N_20545);
or U23944 (N_23944,N_20672,N_21890);
nor U23945 (N_23945,N_20275,N_21578);
or U23946 (N_23946,N_21845,N_20439);
nand U23947 (N_23947,N_21383,N_20620);
or U23948 (N_23948,N_20413,N_21057);
or U23949 (N_23949,N_20952,N_21331);
nand U23950 (N_23950,N_20265,N_21258);
and U23951 (N_23951,N_21246,N_21466);
nand U23952 (N_23952,N_20473,N_20419);
nand U23953 (N_23953,N_20246,N_21377);
or U23954 (N_23954,N_21685,N_21133);
and U23955 (N_23955,N_20671,N_21754);
and U23956 (N_23956,N_21510,N_20466);
nand U23957 (N_23957,N_21632,N_21854);
or U23958 (N_23958,N_21274,N_21426);
nor U23959 (N_23959,N_21218,N_20827);
nand U23960 (N_23960,N_20013,N_20688);
nor U23961 (N_23961,N_20511,N_21382);
xnor U23962 (N_23962,N_20172,N_21629);
and U23963 (N_23963,N_20645,N_20070);
nor U23964 (N_23964,N_20559,N_21649);
or U23965 (N_23965,N_20023,N_21194);
or U23966 (N_23966,N_21716,N_21680);
or U23967 (N_23967,N_20519,N_20029);
nor U23968 (N_23968,N_20669,N_21353);
and U23969 (N_23969,N_21830,N_21773);
nor U23970 (N_23970,N_21877,N_21567);
nor U23971 (N_23971,N_20245,N_20273);
or U23972 (N_23972,N_20912,N_21942);
nor U23973 (N_23973,N_20243,N_20307);
and U23974 (N_23974,N_21702,N_21461);
and U23975 (N_23975,N_20792,N_21664);
nand U23976 (N_23976,N_21962,N_21457);
nor U23977 (N_23977,N_21883,N_20340);
nor U23978 (N_23978,N_21881,N_21297);
or U23979 (N_23979,N_20030,N_21818);
nand U23980 (N_23980,N_21345,N_21480);
nor U23981 (N_23981,N_21209,N_21846);
nand U23982 (N_23982,N_20791,N_20139);
xor U23983 (N_23983,N_20339,N_20533);
nand U23984 (N_23984,N_20126,N_20645);
nor U23985 (N_23985,N_20840,N_21031);
nand U23986 (N_23986,N_20438,N_21102);
nor U23987 (N_23987,N_20886,N_21591);
and U23988 (N_23988,N_21430,N_20598);
and U23989 (N_23989,N_21242,N_20820);
nand U23990 (N_23990,N_20181,N_20312);
nor U23991 (N_23991,N_20106,N_20109);
and U23992 (N_23992,N_20747,N_20321);
and U23993 (N_23993,N_21193,N_20005);
and U23994 (N_23994,N_20668,N_21044);
or U23995 (N_23995,N_20073,N_21914);
nand U23996 (N_23996,N_21740,N_20685);
or U23997 (N_23997,N_20287,N_21681);
and U23998 (N_23998,N_20772,N_20801);
nand U23999 (N_23999,N_20134,N_20916);
or U24000 (N_24000,N_22513,N_23000);
nand U24001 (N_24001,N_23298,N_22465);
nor U24002 (N_24002,N_22499,N_23759);
or U24003 (N_24003,N_22474,N_22198);
nor U24004 (N_24004,N_22832,N_23895);
nor U24005 (N_24005,N_22150,N_23102);
and U24006 (N_24006,N_22429,N_22939);
and U24007 (N_24007,N_23055,N_22693);
nor U24008 (N_24008,N_23056,N_23530);
and U24009 (N_24009,N_23259,N_23945);
nor U24010 (N_24010,N_23890,N_22619);
nor U24011 (N_24011,N_22354,N_22196);
and U24012 (N_24012,N_23263,N_22719);
and U24013 (N_24013,N_22769,N_22563);
nor U24014 (N_24014,N_22866,N_22153);
nor U24015 (N_24015,N_22065,N_22730);
nand U24016 (N_24016,N_23333,N_22040);
nor U24017 (N_24017,N_22301,N_23558);
and U24018 (N_24018,N_23765,N_23423);
nand U24019 (N_24019,N_23038,N_22620);
xor U24020 (N_24020,N_22439,N_22736);
and U24021 (N_24021,N_22741,N_22917);
or U24022 (N_24022,N_22701,N_23585);
nor U24023 (N_24023,N_23215,N_23450);
nor U24024 (N_24024,N_22064,N_23911);
and U24025 (N_24025,N_22863,N_23819);
nand U24026 (N_24026,N_22371,N_22823);
or U24027 (N_24027,N_22096,N_22852);
nor U24028 (N_24028,N_23374,N_22283);
nand U24029 (N_24029,N_23609,N_22277);
nor U24030 (N_24030,N_23933,N_22697);
and U24031 (N_24031,N_23412,N_23972);
or U24032 (N_24032,N_22647,N_23288);
or U24033 (N_24033,N_22790,N_22530);
or U24034 (N_24034,N_23481,N_23318);
nor U24035 (N_24035,N_23902,N_23161);
or U24036 (N_24036,N_22882,N_23560);
or U24037 (N_24037,N_23218,N_23232);
nor U24038 (N_24038,N_23206,N_22038);
nor U24039 (N_24039,N_22255,N_22613);
or U24040 (N_24040,N_22779,N_22510);
or U24041 (N_24041,N_22893,N_22614);
or U24042 (N_24042,N_22341,N_22228);
and U24043 (N_24043,N_23705,N_23150);
or U24044 (N_24044,N_23135,N_22644);
and U24045 (N_24045,N_23873,N_23758);
or U24046 (N_24046,N_22567,N_22186);
nand U24047 (N_24047,N_22957,N_22658);
nand U24048 (N_24048,N_23036,N_22720);
and U24049 (N_24049,N_22526,N_22623);
and U24050 (N_24050,N_23269,N_22133);
and U24051 (N_24051,N_23906,N_22488);
or U24052 (N_24052,N_23790,N_23293);
nand U24053 (N_24053,N_23248,N_22905);
or U24054 (N_24054,N_22185,N_22080);
and U24055 (N_24055,N_22586,N_23787);
nor U24056 (N_24056,N_22290,N_22217);
nor U24057 (N_24057,N_22073,N_22551);
nand U24058 (N_24058,N_22809,N_22011);
nor U24059 (N_24059,N_22532,N_23305);
and U24060 (N_24060,N_22386,N_23573);
nor U24061 (N_24061,N_22345,N_23177);
or U24062 (N_24062,N_23769,N_22662);
nand U24063 (N_24063,N_23313,N_22523);
and U24064 (N_24064,N_23154,N_22868);
nand U24065 (N_24065,N_22580,N_23068);
xor U24066 (N_24066,N_22826,N_22943);
nor U24067 (N_24067,N_22028,N_23818);
nand U24068 (N_24068,N_22578,N_23181);
nand U24069 (N_24069,N_23006,N_23381);
nor U24070 (N_24070,N_22505,N_22980);
nand U24071 (N_24071,N_22140,N_23957);
or U24072 (N_24072,N_23777,N_22956);
nor U24073 (N_24073,N_23458,N_22267);
nand U24074 (N_24074,N_23625,N_22101);
nand U24075 (N_24075,N_22709,N_23871);
or U24076 (N_24076,N_23986,N_22740);
xor U24077 (N_24077,N_23223,N_22787);
or U24078 (N_24078,N_22684,N_23802);
nand U24079 (N_24079,N_23007,N_22460);
nand U24080 (N_24080,N_22397,N_22400);
nand U24081 (N_24081,N_22954,N_22773);
or U24082 (N_24082,N_23084,N_22655);
and U24083 (N_24083,N_23728,N_22804);
or U24084 (N_24084,N_22595,N_23196);
and U24085 (N_24085,N_23311,N_23165);
nor U24086 (N_24086,N_23315,N_23071);
nand U24087 (N_24087,N_22728,N_23265);
or U24088 (N_24088,N_22057,N_23783);
nand U24089 (N_24089,N_22334,N_22471);
nand U24090 (N_24090,N_23119,N_23193);
nand U24091 (N_24091,N_23785,N_23881);
and U24092 (N_24092,N_22287,N_22357);
nor U24093 (N_24093,N_22243,N_23060);
and U24094 (N_24094,N_23489,N_22405);
or U24095 (N_24095,N_23394,N_23058);
or U24096 (N_24096,N_23240,N_22733);
nand U24097 (N_24097,N_22162,N_22346);
nor U24098 (N_24098,N_23171,N_23516);
or U24099 (N_24099,N_23294,N_22169);
or U24100 (N_24100,N_23901,N_22884);
nor U24101 (N_24101,N_23525,N_23396);
nand U24102 (N_24102,N_23994,N_22172);
and U24103 (N_24103,N_22971,N_22187);
or U24104 (N_24104,N_22049,N_22092);
or U24105 (N_24105,N_23456,N_22381);
and U24106 (N_24106,N_22679,N_22835);
or U24107 (N_24107,N_22218,N_22326);
and U24108 (N_24108,N_22780,N_23428);
nor U24109 (N_24109,N_23740,N_23581);
nand U24110 (N_24110,N_22053,N_22200);
nand U24111 (N_24111,N_23051,N_22710);
nor U24112 (N_24112,N_23284,N_22144);
nand U24113 (N_24113,N_23047,N_23101);
nor U24114 (N_24114,N_23766,N_22543);
nand U24115 (N_24115,N_22293,N_22932);
nor U24116 (N_24116,N_23267,N_23100);
nor U24117 (N_24117,N_23488,N_23366);
nor U24118 (N_24118,N_22492,N_22820);
or U24119 (N_24119,N_23182,N_23649);
or U24120 (N_24120,N_22981,N_23549);
nor U24121 (N_24121,N_22180,N_23002);
nand U24122 (N_24122,N_22700,N_23106);
and U24123 (N_24123,N_22422,N_22575);
or U24124 (N_24124,N_22383,N_23761);
nand U24125 (N_24125,N_22136,N_23984);
and U24126 (N_24126,N_23667,N_22161);
or U24127 (N_24127,N_22621,N_23420);
nor U24128 (N_24128,N_23998,N_22858);
or U24129 (N_24129,N_22122,N_23245);
xnor U24130 (N_24130,N_23822,N_22408);
xnor U24131 (N_24131,N_23132,N_22359);
nand U24132 (N_24132,N_23561,N_23476);
and U24133 (N_24133,N_22128,N_22247);
or U24134 (N_24134,N_23629,N_23437);
or U24135 (N_24135,N_22164,N_22690);
nor U24136 (N_24136,N_22625,N_22753);
nand U24137 (N_24137,N_23997,N_23061);
and U24138 (N_24138,N_22432,N_23274);
and U24139 (N_24139,N_23500,N_23037);
nand U24140 (N_24140,N_23435,N_23121);
nor U24141 (N_24141,N_22507,N_23467);
or U24142 (N_24142,N_23341,N_23568);
xnor U24143 (N_24143,N_22076,N_22781);
or U24144 (N_24144,N_22275,N_22377);
or U24145 (N_24145,N_23534,N_23795);
and U24146 (N_24146,N_23138,N_23856);
nor U24147 (N_24147,N_22688,N_22888);
xor U24148 (N_24148,N_22969,N_23014);
and U24149 (N_24149,N_23421,N_23262);
nand U24150 (N_24150,N_22444,N_23666);
and U24151 (N_24151,N_22410,N_23065);
and U24152 (N_24152,N_22665,N_23433);
nand U24153 (N_24153,N_23029,N_22426);
xor U24154 (N_24154,N_22585,N_22480);
or U24155 (N_24155,N_22135,N_23637);
and U24156 (N_24156,N_23094,N_22175);
nor U24157 (N_24157,N_22178,N_22201);
or U24158 (N_24158,N_23916,N_23108);
or U24159 (N_24159,N_22236,N_22987);
nand U24160 (N_24160,N_23964,N_23466);
nor U24161 (N_24161,N_22843,N_22627);
nor U24162 (N_24162,N_22203,N_22145);
or U24163 (N_24163,N_23820,N_22651);
nor U24164 (N_24164,N_22152,N_22366);
nor U24165 (N_24165,N_23087,N_22114);
nand U24166 (N_24166,N_23079,N_23967);
nor U24167 (N_24167,N_22725,N_23180);
and U24168 (N_24168,N_23811,N_22123);
and U24169 (N_24169,N_23713,N_23979);
nand U24170 (N_24170,N_22495,N_23867);
nand U24171 (N_24171,N_22258,N_23331);
xnor U24172 (N_24172,N_22524,N_23021);
and U24173 (N_24173,N_23570,N_23010);
nor U24174 (N_24174,N_22265,N_23781);
or U24175 (N_24175,N_23879,N_22830);
and U24176 (N_24176,N_23271,N_23127);
and U24177 (N_24177,N_22276,N_23226);
or U24178 (N_24178,N_23515,N_22403);
and U24179 (N_24179,N_23589,N_23049);
and U24180 (N_24180,N_23490,N_22663);
nand U24181 (N_24181,N_23139,N_22516);
and U24182 (N_24182,N_23844,N_23813);
or U24183 (N_24183,N_23556,N_22167);
nand U24184 (N_24184,N_23767,N_23362);
nor U24185 (N_24185,N_22896,N_22810);
and U24186 (N_24186,N_23675,N_22353);
nor U24187 (N_24187,N_22482,N_23639);
nor U24188 (N_24188,N_23640,N_23375);
xnor U24189 (N_24189,N_23725,N_22702);
or U24190 (N_24190,N_22996,N_22494);
nand U24191 (N_24191,N_22682,N_22842);
and U24192 (N_24192,N_23185,N_23377);
nand U24193 (N_24193,N_23721,N_22925);
or U24194 (N_24194,N_23775,N_23214);
and U24195 (N_24195,N_23630,N_23949);
and U24196 (N_24196,N_23114,N_23706);
nor U24197 (N_24197,N_23338,N_23988);
and U24198 (N_24198,N_22840,N_22850);
or U24199 (N_24199,N_22085,N_22770);
and U24200 (N_24200,N_22999,N_23908);
and U24201 (N_24201,N_23339,N_23314);
nor U24202 (N_24202,N_23557,N_23920);
or U24203 (N_24203,N_23163,N_22238);
and U24204 (N_24204,N_22940,N_22250);
nor U24205 (N_24205,N_22531,N_23440);
or U24206 (N_24206,N_22522,N_23932);
and U24207 (N_24207,N_22583,N_22428);
and U24208 (N_24208,N_22929,N_22927);
nor U24209 (N_24209,N_23567,N_23553);
nor U24210 (N_24210,N_23363,N_23418);
nand U24211 (N_24211,N_23103,N_23368);
nor U24212 (N_24212,N_22572,N_23716);
and U24213 (N_24213,N_23528,N_22691);
or U24214 (N_24214,N_22489,N_23050);
or U24215 (N_24215,N_22681,N_23659);
nand U24216 (N_24216,N_23472,N_22105);
or U24217 (N_24217,N_23179,N_23442);
or U24218 (N_24218,N_23829,N_23275);
nand U24219 (N_24219,N_23173,N_22836);
or U24220 (N_24220,N_22311,N_22219);
nor U24221 (N_24221,N_23416,N_22883);
nor U24222 (N_24222,N_23438,N_23796);
nor U24223 (N_24223,N_22446,N_23823);
and U24224 (N_24224,N_23306,N_22194);
nand U24225 (N_24225,N_22376,N_22387);
and U24226 (N_24226,N_22078,N_23616);
and U24227 (N_24227,N_22562,N_23624);
nand U24228 (N_24228,N_22897,N_22796);
and U24229 (N_24229,N_23771,N_23631);
xnor U24230 (N_24230,N_23757,N_23976);
and U24231 (N_24231,N_22090,N_22212);
or U24232 (N_24232,N_23210,N_23146);
and U24233 (N_24233,N_23657,N_22802);
or U24234 (N_24234,N_22822,N_22284);
nor U24235 (N_24235,N_22760,N_22766);
nor U24236 (N_24236,N_22867,N_23504);
or U24237 (N_24237,N_23510,N_22019);
nand U24238 (N_24238,N_22642,N_22244);
or U24239 (N_24239,N_22632,N_22759);
nor U24240 (N_24240,N_23993,N_22292);
and U24241 (N_24241,N_23209,N_22479);
nand U24242 (N_24242,N_23544,N_23373);
nor U24243 (N_24243,N_23661,N_23251);
and U24244 (N_24244,N_22685,N_22870);
nor U24245 (N_24245,N_22329,N_22211);
nor U24246 (N_24246,N_23043,N_23016);
nor U24247 (N_24247,N_22549,N_23076);
nor U24248 (N_24248,N_22789,N_22829);
nand U24249 (N_24249,N_23794,N_23012);
and U24250 (N_24250,N_23239,N_22319);
nor U24251 (N_24251,N_22340,N_23940);
and U24252 (N_24252,N_22002,N_23548);
nor U24253 (N_24253,N_23198,N_23158);
nor U24254 (N_24254,N_23491,N_22001);
nand U24255 (N_24255,N_23144,N_22674);
or U24256 (N_24256,N_22747,N_23199);
and U24257 (N_24257,N_22317,N_22298);
and U24258 (N_24258,N_22856,N_23046);
and U24259 (N_24259,N_22536,N_22449);
nand U24260 (N_24260,N_23393,N_23460);
and U24261 (N_24261,N_22445,N_23332);
nor U24262 (N_24262,N_22242,N_23961);
nand U24263 (N_24263,N_22640,N_22389);
and U24264 (N_24264,N_22959,N_23833);
or U24265 (N_24265,N_23022,N_23941);
or U24266 (N_24266,N_22286,N_23749);
nand U24267 (N_24267,N_22483,N_22636);
and U24268 (N_24268,N_22812,N_23751);
nor U24269 (N_24269,N_23807,N_22699);
nor U24270 (N_24270,N_22738,N_23300);
nand U24271 (N_24271,N_23285,N_23449);
nand U24272 (N_24272,N_22608,N_22159);
and U24273 (N_24273,N_23635,N_22007);
nand U24274 (N_24274,N_23859,N_23505);
nand U24275 (N_24275,N_22052,N_23847);
and U24276 (N_24276,N_22241,N_23292);
and U24277 (N_24277,N_22908,N_22231);
nand U24278 (N_24278,N_23734,N_23598);
nand U24279 (N_24279,N_22107,N_22548);
or U24280 (N_24280,N_22800,N_23602);
or U24281 (N_24281,N_22020,N_22204);
and U24282 (N_24282,N_22245,N_22094);
and U24283 (N_24283,N_23768,N_23008);
or U24284 (N_24284,N_22361,N_23521);
or U24285 (N_24285,N_22768,N_23367);
or U24286 (N_24286,N_23782,N_23559);
xnor U24287 (N_24287,N_23980,N_23919);
nor U24288 (N_24288,N_22677,N_23444);
and U24289 (N_24289,N_23981,N_22666);
or U24290 (N_24290,N_22503,N_23398);
nor U24291 (N_24291,N_23664,N_23231);
nand U24292 (N_24292,N_22827,N_22390);
or U24293 (N_24293,N_22995,N_23115);
nor U24294 (N_24294,N_23962,N_23801);
or U24295 (N_24295,N_23638,N_23024);
and U24296 (N_24296,N_23914,N_23303);
xor U24297 (N_24297,N_23357,N_23863);
and U24298 (N_24298,N_22055,N_22617);
nor U24299 (N_24299,N_23612,N_23898);
nor U24300 (N_24300,N_23607,N_23434);
nor U24301 (N_24301,N_22861,N_23574);
nor U24302 (N_24302,N_22086,N_23647);
nand U24303 (N_24303,N_23089,N_22680);
nand U24304 (N_24304,N_22698,N_23027);
or U24305 (N_24305,N_23955,N_22072);
nand U24306 (N_24306,N_23344,N_23235);
or U24307 (N_24307,N_23918,N_23969);
or U24308 (N_24308,N_23028,N_22900);
nand U24309 (N_24309,N_22915,N_23774);
and U24310 (N_24310,N_23968,N_22638);
or U24311 (N_24311,N_22594,N_23673);
nand U24312 (N_24312,N_23539,N_22034);
and U24313 (N_24313,N_22000,N_23773);
nor U24314 (N_24314,N_22117,N_22997);
and U24315 (N_24315,N_22440,N_22914);
and U24316 (N_24316,N_22542,N_22425);
xor U24317 (N_24317,N_22259,N_22857);
nand U24318 (N_24318,N_23874,N_22875);
nor U24319 (N_24319,N_23526,N_22230);
and U24320 (N_24320,N_23860,N_23841);
and U24321 (N_24321,N_22312,N_23383);
nor U24322 (N_24322,N_22582,N_22365);
or U24323 (N_24323,N_22240,N_23464);
nand U24324 (N_24324,N_23569,N_22207);
or U24325 (N_24325,N_22629,N_23970);
and U24326 (N_24326,N_23883,N_23846);
and U24327 (N_24327,N_22552,N_22059);
or U24328 (N_24328,N_23854,N_22331);
and U24329 (N_24329,N_22024,N_23717);
and U24330 (N_24330,N_22831,N_22182);
nor U24331 (N_24331,N_23307,N_23861);
or U24332 (N_24332,N_22650,N_23959);
and U24333 (N_24333,N_23278,N_22137);
and U24334 (N_24334,N_23042,N_23302);
nor U24335 (N_24335,N_23066,N_22430);
or U24336 (N_24336,N_22036,N_22202);
or U24337 (N_24337,N_23772,N_22919);
nand U24338 (N_24338,N_22676,N_23776);
or U24339 (N_24339,N_23120,N_23457);
nor U24340 (N_24340,N_23475,N_23204);
xor U24341 (N_24341,N_23763,N_23935);
and U24342 (N_24342,N_23312,N_22058);
nor U24343 (N_24343,N_22579,N_22491);
nand U24344 (N_24344,N_23352,N_22824);
nor U24345 (N_24345,N_23893,N_22392);
or U24346 (N_24346,N_23878,N_22886);
and U24347 (N_24347,N_23360,N_22149);
nor U24348 (N_24348,N_22950,N_22782);
or U24349 (N_24349,N_22944,N_22795);
and U24350 (N_24350,N_22894,N_22328);
or U24351 (N_24351,N_23821,N_23628);
nor U24352 (N_24352,N_23054,N_23756);
and U24353 (N_24353,N_22902,N_23279);
nor U24354 (N_24354,N_23237,N_23222);
and U24355 (N_24355,N_23831,N_23334);
or U24356 (N_24356,N_23229,N_22414);
nor U24357 (N_24357,N_23364,N_22988);
or U24358 (N_24358,N_22731,N_22171);
nor U24359 (N_24359,N_22213,N_23839);
nor U24360 (N_24360,N_22717,N_23851);
and U24361 (N_24361,N_23128,N_23153);
or U24362 (N_24362,N_23205,N_22571);
and U24363 (N_24363,N_22904,N_22718);
nand U24364 (N_24364,N_22504,N_23952);
and U24365 (N_24365,N_23186,N_23018);
nor U24366 (N_24366,N_23454,N_23170);
nand U24367 (N_24367,N_23936,N_23216);
nand U24368 (N_24368,N_23620,N_23063);
or U24369 (N_24369,N_22553,N_22457);
nor U24370 (N_24370,N_23934,N_23172);
or U24371 (N_24371,N_23891,N_22139);
nand U24372 (N_24372,N_22555,N_23496);
nor U24373 (N_24373,N_22714,N_22689);
or U24374 (N_24374,N_22108,N_22515);
nor U24375 (N_24375,N_22890,N_22509);
and U24376 (N_24376,N_23401,N_23075);
nand U24377 (N_24377,N_22788,N_23169);
nand U24378 (N_24378,N_23720,N_22307);
and U24379 (N_24379,N_22871,N_22584);
or U24380 (N_24380,N_23155,N_22442);
and U24381 (N_24381,N_22846,N_22813);
or U24382 (N_24382,N_23411,N_23889);
or U24383 (N_24383,N_23611,N_23258);
nor U24384 (N_24384,N_22481,N_22336);
and U24385 (N_24385,N_23092,N_22558);
and U24386 (N_24386,N_22179,N_23129);
and U24387 (N_24387,N_23634,N_22556);
nor U24388 (N_24388,N_23403,N_23555);
nand U24389 (N_24389,N_23482,N_22746);
or U24390 (N_24390,N_23136,N_23862);
or U24391 (N_24391,N_22313,N_23359);
nand U24392 (N_24392,N_22734,N_22538);
nor U24393 (N_24393,N_23414,N_22616);
nor U24394 (N_24394,N_23184,N_22342);
xor U24395 (N_24395,N_23966,N_22132);
nand U24396 (N_24396,N_22909,N_23137);
nand U24397 (N_24397,N_23584,N_23701);
nand U24398 (N_24398,N_22082,N_23670);
and U24399 (N_24399,N_23563,N_23287);
nor U24400 (N_24400,N_22015,N_22272);
nor U24401 (N_24401,N_22756,N_23388);
nand U24402 (N_24402,N_22325,N_22966);
nand U24403 (N_24403,N_22839,N_23944);
xor U24404 (N_24404,N_22310,N_22239);
and U24405 (N_24405,N_22808,N_22044);
or U24406 (N_24406,N_23590,N_22156);
and U24407 (N_24407,N_22281,N_23806);
nand U24408 (N_24408,N_22401,N_22014);
nand U24409 (N_24409,N_22777,N_22569);
or U24410 (N_24410,N_23770,N_22023);
or U24411 (N_24411,N_23712,N_22976);
or U24412 (N_24412,N_22517,N_22093);
nor U24413 (N_24413,N_23384,N_22188);
or U24414 (N_24414,N_23200,N_22437);
nand U24415 (N_24415,N_23726,N_22407);
or U24416 (N_24416,N_23105,N_23126);
nand U24417 (N_24417,N_23365,N_23264);
nand U24418 (N_24418,N_23358,N_22295);
or U24419 (N_24419,N_22417,N_23619);
nand U24420 (N_24420,N_23755,N_23192);
nand U24421 (N_24421,N_22142,N_22931);
nand U24422 (N_24422,N_23330,N_22355);
or U24423 (N_24423,N_22633,N_23147);
xnor U24424 (N_24424,N_22865,N_22936);
or U24425 (N_24425,N_23636,N_22013);
or U24426 (N_24426,N_23737,N_23015);
or U24427 (N_24427,N_23912,N_22322);
or U24428 (N_24428,N_23211,N_22380);
nor U24429 (N_24429,N_23402,N_22912);
and U24430 (N_24430,N_22634,N_22948);
nand U24431 (N_24431,N_22262,N_23238);
nor U24432 (N_24432,N_23910,N_22043);
xor U24433 (N_24433,N_22089,N_23082);
nor U24434 (N_24434,N_22972,N_23729);
or U24435 (N_24435,N_23183,N_22296);
nor U24436 (N_24436,N_23395,N_23816);
or U24437 (N_24437,N_22887,N_22134);
nand U24438 (N_24438,N_22450,N_23840);
or U24439 (N_24439,N_23201,N_23099);
nor U24440 (N_24440,N_23814,N_23834);
nor U24441 (N_24441,N_22237,N_23680);
and U24442 (N_24442,N_22451,N_23578);
nand U24443 (N_24443,N_22889,N_22109);
or U24444 (N_24444,N_22994,N_22018);
and U24445 (N_24445,N_23234,N_22593);
nor U24446 (N_24446,N_22129,N_22084);
nand U24447 (N_24447,N_23989,N_23035);
and U24448 (N_24448,N_22022,N_23225);
and U24449 (N_24449,N_22339,N_23599);
nand U24450 (N_24450,N_23371,N_23546);
nor U24451 (N_24451,N_22723,N_22210);
nor U24452 (N_24452,N_23784,N_22416);
and U24453 (N_24453,N_22924,N_23188);
nor U24454 (N_24454,N_23658,N_23954);
or U24455 (N_24455,N_23124,N_22166);
nor U24456 (N_24456,N_23244,N_22192);
or U24457 (N_24457,N_22358,N_22111);
nor U24458 (N_24458,N_22257,N_23999);
and U24459 (N_24459,N_23978,N_22529);
nand U24460 (N_24460,N_23554,N_22039);
or U24461 (N_24461,N_23439,N_23415);
and U24462 (N_24462,N_22854,N_23571);
or U24463 (N_24463,N_23261,N_22163);
or U24464 (N_24464,N_22127,N_23744);
nand U24465 (N_24465,N_22233,N_22113);
or U24466 (N_24466,N_22844,N_22977);
nand U24467 (N_24467,N_22098,N_22251);
nor U24468 (N_24468,N_22799,N_22916);
nand U24469 (N_24469,N_23745,N_23922);
and U24470 (N_24470,N_22285,N_22027);
nor U24471 (N_24471,N_22138,N_23336);
or U24472 (N_24472,N_22268,N_23497);
nand U24473 (N_24473,N_22472,N_22657);
nand U24474 (N_24474,N_23309,N_23501);
xor U24475 (N_24475,N_22347,N_23270);
nor U24476 (N_24476,N_23436,N_23130);
nand U24477 (N_24477,N_22938,N_22630);
and U24478 (N_24478,N_23896,N_23797);
or U24479 (N_24479,N_23156,N_22845);
and U24480 (N_24480,N_22775,N_23943);
nor U24481 (N_24481,N_22304,N_22935);
xnor U24482 (N_24482,N_22892,N_23618);
and U24483 (N_24483,N_23764,N_22356);
and U24484 (N_24484,N_22853,N_23202);
and U24485 (N_24485,N_23122,N_22256);
nand U24486 (N_24486,N_23779,N_22876);
nor U24487 (N_24487,N_22466,N_22221);
nor U24488 (N_24488,N_23674,N_22683);
and U24489 (N_24489,N_22974,N_23702);
nor U24490 (N_24490,N_22302,N_22315);
nor U24491 (N_24491,N_22497,N_22631);
nor U24492 (N_24492,N_23842,N_22501);
or U24493 (N_24493,N_22891,N_22545);
nor U24494 (N_24494,N_22661,N_23946);
nand U24495 (N_24495,N_23353,N_22722);
xnor U24496 (N_24496,N_23026,N_22266);
nor U24497 (N_24497,N_22306,N_22415);
and U24498 (N_24498,N_22447,N_22771);
and U24499 (N_24499,N_22518,N_23885);
nand U24500 (N_24500,N_22124,N_22490);
nor U24501 (N_24501,N_23409,N_22335);
nand U24502 (N_24502,N_23899,N_23791);
nand U24503 (N_24503,N_22962,N_22565);
or U24504 (N_24504,N_22743,N_23707);
or U24505 (N_24505,N_22975,N_23480);
nand U24506 (N_24506,N_23512,N_23113);
nand U24507 (N_24507,N_22601,N_22807);
nor U24508 (N_24508,N_23662,N_22946);
nand U24509 (N_24509,N_22273,N_23809);
or U24510 (N_24510,N_22878,N_22157);
nor U24511 (N_24511,N_22656,N_22318);
nor U24512 (N_24512,N_23532,N_22798);
nand U24513 (N_24513,N_22933,N_23255);
and U24514 (N_24514,N_23652,N_23552);
and U24515 (N_24515,N_22112,N_23960);
nor U24516 (N_24516,N_23213,N_22745);
or U24517 (N_24517,N_23531,N_22654);
nor U24518 (N_24518,N_23579,N_22215);
nor U24519 (N_24519,N_22811,N_22581);
and U24520 (N_24520,N_22475,N_23681);
nor U24521 (N_24521,N_23875,N_22352);
and U24522 (N_24522,N_22083,N_23746);
or U24523 (N_24523,N_22269,N_23217);
nand U24524 (N_24524,N_22819,N_22305);
and U24525 (N_24525,N_22786,N_22821);
nor U24526 (N_24526,N_22847,N_23550);
and U24527 (N_24527,N_23346,N_22671);
nand U24528 (N_24528,N_22270,N_23738);
or U24529 (N_24529,N_22533,N_23040);
nand U24530 (N_24530,N_22794,N_23614);
or U24531 (N_24531,N_23174,N_22004);
or U24532 (N_24532,N_22227,N_22455);
or U24533 (N_24533,N_23276,N_22732);
nand U24534 (N_24534,N_22762,N_22404);
and U24535 (N_24535,N_22992,N_22667);
or U24536 (N_24536,N_23096,N_22729);
nor U24537 (N_24537,N_22297,N_23151);
nand U24538 (N_24538,N_22332,N_23167);
nor U24539 (N_24539,N_22784,N_22873);
or U24540 (N_24540,N_22079,N_23565);
nor U24541 (N_24541,N_22805,N_22051);
xnor U24542 (N_24542,N_23686,N_23289);
xnor U24543 (N_24543,N_22993,N_23533);
nand U24544 (N_24544,N_22859,N_22309);
nor U24545 (N_24545,N_23870,N_23088);
nor U24546 (N_24546,N_22487,N_22041);
or U24547 (N_24547,N_22983,N_22716);
and U24548 (N_24548,N_23097,N_23788);
and U24549 (N_24549,N_23965,N_23692);
xnor U24550 (N_24550,N_23626,N_22448);
and U24551 (N_24551,N_22104,N_23653);
and U24552 (N_24552,N_22607,N_23723);
nand U24553 (N_24553,N_22849,N_23538);
and U24554 (N_24554,N_23117,N_22061);
or U24555 (N_24555,N_23576,N_23310);
nor U24556 (N_24556,N_22222,N_23937);
nand U24557 (N_24557,N_22554,N_22727);
nand U24558 (N_24558,N_22115,N_22125);
nand U24559 (N_24559,N_22006,N_22314);
nand U24560 (N_24560,N_23321,N_23112);
or U24561 (N_24561,N_22409,N_23203);
nand U24562 (N_24562,N_22453,N_22622);
or U24563 (N_24563,N_23507,N_23280);
and U24564 (N_24564,N_23857,N_22514);
or U24565 (N_24565,N_23951,N_22512);
nand U24566 (N_24566,N_23741,N_23090);
nor U24567 (N_24567,N_22478,N_23724);
nand U24568 (N_24568,N_22063,N_22181);
nand U24569 (N_24569,N_23677,N_22960);
or U24570 (N_24570,N_23343,N_23350);
nand U24571 (N_24571,N_22208,N_22364);
nor U24572 (N_24572,N_22639,N_23266);
nand U24573 (N_24573,N_23408,N_23956);
nand U24574 (N_24574,N_23694,N_23017);
nand U24575 (N_24575,N_22791,N_23425);
nor U24576 (N_24576,N_22459,N_22712);
or U24577 (N_24577,N_22828,N_23727);
nand U24578 (N_24578,N_22561,N_22223);
nand U24579 (N_24579,N_22991,N_22848);
and U24580 (N_24580,N_23732,N_22197);
and U24581 (N_24581,N_22327,N_23236);
nor U24582 (N_24582,N_23925,N_23317);
nand U24583 (N_24583,N_23950,N_23067);
or U24584 (N_24584,N_23518,N_22921);
nand U24585 (N_24585,N_22042,N_22818);
nor U24586 (N_24586,N_23448,N_23683);
or U24587 (N_24587,N_23104,N_22303);
or U24588 (N_24588,N_22402,N_23260);
nor U24589 (N_24589,N_23019,N_22618);
nor U24590 (N_24590,N_23013,N_23592);
nand U24591 (N_24591,N_22978,N_22652);
and U24592 (N_24592,N_23987,N_23011);
and U24593 (N_24593,N_23044,N_22424);
and U24594 (N_24594,N_22032,N_23325);
or U24595 (N_24595,N_23308,N_22158);
nor U24596 (N_24596,N_23900,N_23514);
or U24597 (N_24597,N_22476,N_22559);
and U24598 (N_24598,N_23283,N_23977);
or U24599 (N_24599,N_23233,N_23864);
or U24600 (N_24600,N_23752,N_23324);
nand U24601 (N_24601,N_22168,N_23340);
or U24602 (N_24602,N_22901,N_22816);
or U24603 (N_24603,N_23277,N_22735);
and U24604 (N_24604,N_22570,N_23417);
nor U24605 (N_24605,N_22418,N_23939);
nor U24606 (N_24606,N_22232,N_23005);
and U24607 (N_24607,N_22350,N_23178);
nor U24608 (N_24608,N_23710,N_23868);
nand U24609 (N_24609,N_23928,N_23641);
and U24610 (N_24610,N_23335,N_22783);
nand U24611 (N_24611,N_22100,N_23676);
or U24612 (N_24612,N_23708,N_22419);
or U24613 (N_24613,N_23399,N_23973);
and U24614 (N_24614,N_22757,N_22374);
and U24615 (N_24615,N_22160,N_23572);
nand U24616 (N_24616,N_23651,N_23836);
and U24617 (N_24617,N_22420,N_22926);
nand U24618 (N_24618,N_22669,N_23345);
or U24619 (N_24619,N_22675,N_23250);
or U24620 (N_24620,N_22707,N_23004);
or U24621 (N_24621,N_22395,N_23164);
or U24622 (N_24622,N_23850,N_22220);
nor U24623 (N_24623,N_23424,N_22391);
nand U24624 (N_24624,N_23663,N_22984);
nor U24625 (N_24625,N_22838,N_22141);
nand U24626 (N_24626,N_22216,N_23110);
and U24627 (N_24627,N_23931,N_23524);
nand U24628 (N_24628,N_22349,N_23463);
and U24629 (N_24629,N_23975,N_23133);
or U24630 (N_24630,N_22527,N_22368);
nor U24631 (N_24631,N_22099,N_23134);
nand U24632 (N_24632,N_23689,N_23053);
nor U24633 (N_24633,N_22945,N_23429);
and U24634 (N_24634,N_23913,N_23838);
nor U24635 (N_24635,N_22263,N_22033);
nor U24636 (N_24636,N_23824,N_22970);
nor U24637 (N_24637,N_23443,N_23479);
and U24638 (N_24638,N_22715,N_22934);
nand U24639 (N_24639,N_22367,N_22234);
xnor U24640 (N_24640,N_23529,N_22300);
or U24641 (N_24641,N_23486,N_23654);
nor U24642 (N_24642,N_23580,N_23081);
nand U24643 (N_24643,N_23958,N_22748);
and U24644 (N_24644,N_22016,N_23672);
nor U24645 (N_24645,N_23595,N_23577);
or U24646 (N_24646,N_23921,N_22557);
and U24647 (N_24647,N_23601,N_23656);
or U24648 (N_24648,N_23039,N_22737);
nand U24649 (N_24649,N_23522,N_23608);
or U24650 (N_24650,N_22467,N_23074);
and U24651 (N_24651,N_22337,N_22120);
nor U24652 (N_24652,N_23915,N_23208);
nor U24653 (N_24653,N_23621,N_22443);
nor U24654 (N_24654,N_23326,N_22648);
nand U24655 (N_24655,N_23419,N_23080);
and U24656 (N_24656,N_22519,N_23669);
nand U24657 (N_24657,N_22772,N_23753);
xnor U24658 (N_24658,N_23062,N_22384);
nand U24659 (N_24659,N_23031,N_23385);
nor U24660 (N_24660,N_23286,N_22010);
and U24661 (N_24661,N_22922,N_23455);
and U24662 (N_24662,N_22612,N_23888);
and U24663 (N_24663,N_23886,N_23591);
nor U24664 (N_24664,N_23246,N_22047);
nor U24665 (N_24665,N_22056,N_23498);
and U24666 (N_24666,N_22037,N_23354);
nand U24667 (N_24667,N_22003,N_22911);
or U24668 (N_24668,N_22695,N_23907);
nor U24669 (N_24669,N_23495,N_22500);
and U24670 (N_24670,N_22989,N_23805);
or U24671 (N_24671,N_22421,N_22814);
and U24672 (N_24672,N_22463,N_23483);
and U24673 (N_24673,N_22229,N_22485);
nor U24674 (N_24674,N_23249,N_22592);
or U24675 (N_24675,N_22299,N_22797);
and U24676 (N_24676,N_23502,N_23897);
or U24677 (N_24677,N_22338,N_23316);
or U24678 (N_24678,N_23527,N_22199);
nand U24679 (N_24679,N_23992,N_22841);
nor U24680 (N_24680,N_22393,N_23033);
and U24681 (N_24681,N_22920,N_23095);
nand U24682 (N_24682,N_23668,N_23320);
or U24683 (N_24683,N_22708,N_22541);
nand U24684 (N_24684,N_23093,N_22323);
and U24685 (N_24685,N_22967,N_22473);
and U24686 (N_24686,N_23942,N_23537);
nand U24687 (N_24687,N_22986,N_23780);
nand U24688 (N_24688,N_22624,N_22330);
nor U24689 (N_24689,N_23827,N_22106);
nor U24690 (N_24690,N_23465,N_22825);
nand U24691 (N_24691,N_23826,N_22602);
nor U24692 (N_24692,N_22635,N_23461);
and U24693 (N_24693,N_22597,N_23032);
nand U24694 (N_24694,N_23003,N_23372);
nor U24695 (N_24695,N_23125,N_23142);
and U24696 (N_24696,N_22528,N_23623);
and U24697 (N_24697,N_22399,N_22628);
nor U24698 (N_24698,N_23722,N_23078);
and U24699 (N_24699,N_22641,N_22225);
nor U24700 (N_24700,N_23176,N_22869);
nor U24701 (N_24701,N_22362,N_22441);
and U24702 (N_24702,N_23508,N_22343);
and U24703 (N_24703,N_23253,N_23297);
or U24704 (N_24704,N_23351,N_23152);
or U24705 (N_24705,N_23149,N_22637);
nor U24706 (N_24706,N_22851,N_23610);
nand U24707 (N_24707,N_22253,N_23445);
and U24708 (N_24708,N_23869,N_22493);
nand U24709 (N_24709,N_22462,N_23830);
nor U24710 (N_24710,N_23877,N_22694);
nand U24711 (N_24711,N_22435,N_23410);
xnor U24712 (N_24712,N_23545,N_22062);
or U24713 (N_24713,N_23190,N_22070);
nor U24714 (N_24714,N_22792,N_22880);
or U24715 (N_24715,N_22095,N_22021);
and U24716 (N_24716,N_22653,N_23882);
or U24717 (N_24717,N_22646,N_23982);
nor U24718 (N_24718,N_23487,N_22110);
nor U24719 (N_24719,N_22692,N_22573);
and U24720 (N_24720,N_22705,N_22672);
and U24721 (N_24721,N_22382,N_22075);
nand U24722 (N_24722,N_22091,N_22235);
and U24723 (N_24723,N_22670,N_22952);
and U24724 (N_24724,N_22360,N_23441);
or U24725 (N_24725,N_23947,N_23690);
and U24726 (N_24726,N_23810,N_23693);
nor U24727 (N_24727,N_22603,N_23189);
and U24728 (N_24728,N_22568,N_22965);
and U24729 (N_24729,N_23743,N_23212);
nor U24730 (N_24730,N_22615,N_22664);
or U24731 (N_24731,N_22486,N_22009);
nor U24732 (N_24732,N_23123,N_22765);
xor U24733 (N_24733,N_23207,N_23034);
or U24734 (N_24734,N_23400,N_22899);
and U24735 (N_24735,N_23804,N_23930);
nand U24736 (N_24736,N_22577,N_22496);
nor U24737 (N_24737,N_22596,N_23519);
or U24738 (N_24738,N_23430,N_22279);
and U24739 (N_24739,N_23739,N_22961);
nor U24740 (N_24740,N_23903,N_23426);
nor U24741 (N_24741,N_22855,N_22379);
and U24742 (N_24742,N_22396,N_22165);
nor U24743 (N_24743,N_22434,N_22566);
nand U24744 (N_24744,N_23887,N_23687);
nor U24745 (N_24745,N_23845,N_23477);
and U24746 (N_24746,N_22289,N_23397);
or U24747 (N_24747,N_22763,N_22468);
nand U24748 (N_24748,N_22659,N_22029);
or U24749 (N_24749,N_23422,N_23597);
nand U24750 (N_24750,N_22193,N_23586);
nand U24751 (N_24751,N_22776,N_22316);
nand U24752 (N_24752,N_22755,N_23268);
or U24753 (N_24753,N_22508,N_23224);
nand U24754 (N_24754,N_23600,N_23905);
nor U24755 (N_24755,N_23923,N_22758);
or U24756 (N_24756,N_22862,N_22604);
or U24757 (N_24757,N_23835,N_22547);
nor U24758 (N_24758,N_23832,N_23665);
nand U24759 (N_24759,N_23220,N_22834);
and U24760 (N_24760,N_22333,N_22879);
nor U24761 (N_24761,N_23760,N_22031);
nor U24762 (N_24762,N_22546,N_22146);
or U24763 (N_24763,N_23471,N_22143);
or U24764 (N_24764,N_23349,N_23116);
nand U24765 (N_24765,N_23247,N_23131);
or U24766 (N_24766,N_23704,N_23855);
or U24767 (N_24767,N_22308,N_22540);
nand U24768 (N_24768,N_22173,N_23187);
or U24769 (N_24769,N_22274,N_22121);
or U24770 (N_24770,N_23175,N_23605);
or U24771 (N_24771,N_22060,N_22599);
nor U24772 (N_24772,N_22126,N_22588);
or U24773 (N_24773,N_22282,N_22248);
nand U24774 (N_24774,N_22726,N_23494);
nor U24775 (N_24775,N_23858,N_22195);
nor U24776 (N_24776,N_23347,N_23281);
or U24777 (N_24777,N_23162,N_22949);
or U24778 (N_24778,N_22154,N_22953);
and U24779 (N_24779,N_23513,N_23356);
nand U24780 (N_24780,N_22264,N_22436);
nand U24781 (N_24781,N_22910,N_23837);
or U24782 (N_24782,N_22294,N_22260);
nor U24783 (N_24783,N_23077,N_23413);
and U24784 (N_24784,N_22525,N_22958);
and U24785 (N_24785,N_23812,N_22833);
nand U24786 (N_24786,N_23160,N_22406);
nor U24787 (N_24787,N_22484,N_23322);
nor U24788 (N_24788,N_22793,N_23098);
nor U24789 (N_24789,N_22643,N_23143);
and U24790 (N_24790,N_22687,N_23748);
or U24791 (N_24791,N_22706,N_23355);
and U24792 (N_24792,N_23086,N_22937);
nand U24793 (N_24793,N_23370,N_23485);
nand U24794 (N_24794,N_22351,N_22686);
or U24795 (N_24795,N_22645,N_23715);
and U24796 (N_24796,N_23111,N_22456);
xnor U24797 (N_24797,N_23499,N_23319);
nand U24798 (N_24798,N_23617,N_22982);
and U24799 (N_24799,N_22906,N_22877);
nor U24800 (N_24800,N_23678,N_23378);
nand U24801 (N_24801,N_22458,N_23730);
nor U24802 (N_24802,N_23703,N_23478);
nand U24803 (N_24803,N_22767,N_22990);
nor U24804 (N_24804,N_23073,N_23736);
and U24805 (N_24805,N_23030,N_23904);
and U24806 (N_24806,N_23323,N_22177);
nor U24807 (N_24807,N_23361,N_22427);
or U24808 (N_24808,N_22750,N_23695);
and U24809 (N_24809,N_23750,N_22673);
nand U24810 (N_24810,N_23843,N_22363);
nand U24811 (N_24811,N_23219,N_22885);
or U24812 (N_24812,N_23273,N_22544);
and U24813 (N_24813,N_22148,N_22291);
or U24814 (N_24814,N_22097,N_22591);
nand U24815 (N_24815,N_22261,N_23786);
nor U24816 (N_24816,N_22469,N_23020);
nor U24817 (N_24817,N_22534,N_23825);
nand U24818 (N_24818,N_22801,N_23282);
xnor U24819 (N_24819,N_23052,N_22506);
nand U24820 (N_24820,N_22560,N_23853);
nand U24821 (N_24821,N_22249,N_22626);
or U24822 (N_24822,N_23996,N_23583);
and U24823 (N_24823,N_23141,N_23221);
nor U24824 (N_24824,N_23985,N_23547);
and U24825 (N_24825,N_22087,N_23242);
nand U24826 (N_24826,N_23733,N_23711);
and U24827 (N_24827,N_23872,N_22749);
and U24828 (N_24828,N_22170,N_22385);
nor U24829 (N_24829,N_22721,N_23971);
or U24830 (N_24830,N_23257,N_22046);
nand U24831 (N_24831,N_23194,N_22521);
or U24832 (N_24832,N_23803,N_23230);
and U24833 (N_24833,N_23064,N_23604);
and U24834 (N_24834,N_23195,N_22067);
nand U24835 (N_24835,N_22744,N_23511);
and U24836 (N_24836,N_22461,N_23543);
nand U24837 (N_24837,N_23747,N_23386);
nand U24838 (N_24838,N_23622,N_23650);
nand U24839 (N_24839,N_23698,N_22589);
and U24840 (N_24840,N_22898,N_22190);
nand U24841 (N_24841,N_22324,N_23328);
nor U24842 (N_24842,N_23995,N_22069);
or U24843 (N_24843,N_22184,N_22071);
or U24844 (N_24844,N_23575,N_22711);
and U24845 (N_24845,N_23072,N_22209);
or U24846 (N_24846,N_22035,N_22649);
nor U24847 (N_24847,N_23407,N_22742);
or U24848 (N_24848,N_22502,N_22806);
and U24849 (N_24849,N_23157,N_23252);
nor U24850 (N_24850,N_22176,N_22151);
nor U24851 (N_24851,N_23432,N_23390);
nand U24852 (N_24852,N_22537,N_23679);
and U24853 (N_24853,N_22288,N_22751);
nand U24854 (N_24854,N_23369,N_23542);
and U24855 (N_24855,N_22609,N_22520);
nor U24856 (N_24856,N_23892,N_23691);
and U24857 (N_24857,N_23938,N_23389);
nand U24858 (N_24858,N_23564,N_23168);
nor U24859 (N_24859,N_23817,N_23884);
or U24860 (N_24860,N_22088,N_22963);
and U24861 (N_24861,N_23948,N_23762);
and U24862 (N_24862,N_23789,N_23718);
and U24863 (N_24863,N_23057,N_22411);
nor U24864 (N_24864,N_22116,N_23387);
nand U24865 (N_24865,N_23243,N_22774);
nand U24866 (N_24866,N_23301,N_22373);
nand U24867 (N_24867,N_23427,N_23688);
or U24868 (N_24868,N_23593,N_23963);
nand U24869 (N_24869,N_22754,N_23974);
nor U24870 (N_24870,N_22923,N_22668);
or U24871 (N_24871,N_22918,N_22378);
nor U24872 (N_24872,N_22008,N_23808);
or U24873 (N_24873,N_23462,N_23025);
nand U24874 (N_24874,N_23468,N_23405);
nor U24875 (N_24875,N_22955,N_22907);
and U24876 (N_24876,N_23719,N_23391);
xnor U24877 (N_24877,N_22550,N_23517);
and U24878 (N_24878,N_22131,N_22077);
nand U24879 (N_24879,N_22930,N_23256);
and U24880 (N_24880,N_22068,N_23700);
nand U24881 (N_24881,N_23731,N_22803);
and U24882 (N_24882,N_22598,N_22713);
nand U24883 (N_24883,N_23492,N_22423);
and U24884 (N_24884,N_23228,N_23894);
or U24885 (N_24885,N_22511,N_23392);
nor U24886 (N_24886,N_22454,N_23509);
and U24887 (N_24887,N_23085,N_23459);
or U24888 (N_24888,N_23587,N_23337);
and U24889 (N_24889,N_23376,N_23699);
xnor U24890 (N_24890,N_23227,N_22913);
or U24891 (N_24891,N_22189,N_22815);
nor U24892 (N_24892,N_22066,N_23909);
nor U24893 (N_24893,N_23643,N_23566);
and U24894 (N_24894,N_22205,N_22752);
nand U24895 (N_24895,N_23197,N_23083);
and U24896 (N_24896,N_23642,N_23983);
nand U24897 (N_24897,N_23540,N_22174);
nand U24898 (N_24898,N_23241,N_22224);
nor U24899 (N_24899,N_23469,N_23926);
or U24900 (N_24900,N_23329,N_22005);
nand U24901 (N_24901,N_23990,N_23431);
and U24902 (N_24902,N_22412,N_23446);
and U24903 (N_24903,N_22660,N_23451);
nor U24904 (N_24904,N_22369,N_23633);
and U24905 (N_24905,N_23627,N_23917);
nor U24906 (N_24906,N_22895,N_22452);
nand U24907 (N_24907,N_22498,N_22872);
and U24908 (N_24908,N_23109,N_22470);
xor U24909 (N_24909,N_23107,N_22817);
xor U24910 (N_24910,N_23644,N_22985);
nand U24911 (N_24911,N_23535,N_23865);
nand U24912 (N_24912,N_23059,N_22119);
or U24913 (N_24913,N_22903,N_22464);
nor U24914 (N_24914,N_23406,N_22147);
or U24915 (N_24915,N_23536,N_23735);
nand U24916 (N_24916,N_23754,N_22252);
xnor U24917 (N_24917,N_23296,N_22081);
and U24918 (N_24918,N_22576,N_22600);
or U24919 (N_24919,N_22394,N_22045);
nand U24920 (N_24920,N_22764,N_22864);
and U24921 (N_24921,N_23924,N_22206);
and U24922 (N_24922,N_23140,N_23470);
and U24923 (N_24923,N_23596,N_23815);
nor U24924 (N_24924,N_23852,N_22012);
and U24925 (N_24925,N_22785,N_23474);
nor U24926 (N_24926,N_22761,N_22348);
nor U24927 (N_24927,N_23148,N_23551);
or U24928 (N_24928,N_23304,N_23453);
nor U24929 (N_24929,N_22979,N_23299);
or U24930 (N_24930,N_23380,N_22941);
and U24931 (N_24931,N_22130,N_23091);
nand U24932 (N_24932,N_23685,N_23473);
or U24933 (N_24933,N_23159,N_22928);
and U24934 (N_24934,N_23493,N_23696);
or U24935 (N_24935,N_22278,N_23348);
or U24936 (N_24936,N_22271,N_23001);
nor U24937 (N_24937,N_22610,N_23953);
and U24938 (N_24938,N_23828,N_23291);
or U24939 (N_24939,N_22191,N_23645);
and U24940 (N_24940,N_22696,N_22118);
nand U24941 (N_24941,N_22017,N_23045);
nor U24942 (N_24942,N_22246,N_23655);
nor U24943 (N_24943,N_22431,N_22320);
and U24944 (N_24944,N_22438,N_22433);
and U24945 (N_24945,N_22535,N_23646);
or U24946 (N_24946,N_22477,N_22388);
xnor U24947 (N_24947,N_23070,N_23848);
nor U24948 (N_24948,N_23876,N_23880);
or U24949 (N_24949,N_22964,N_23023);
or U24950 (N_24950,N_22778,N_22605);
nor U24951 (N_24951,N_23632,N_23382);
and U24952 (N_24952,N_22590,N_22103);
nand U24953 (N_24953,N_23606,N_22375);
and U24954 (N_24954,N_22611,N_23682);
and U24955 (N_24955,N_22539,N_23582);
nor U24956 (N_24956,N_23191,N_22951);
or U24957 (N_24957,N_23615,N_23798);
nor U24958 (N_24958,N_22678,N_22998);
nand U24959 (N_24959,N_22704,N_22214);
or U24960 (N_24960,N_23069,N_22947);
nand U24961 (N_24961,N_23118,N_22606);
nand U24962 (N_24962,N_22254,N_23849);
nor U24963 (N_24963,N_23048,N_23295);
nand U24964 (N_24964,N_23799,N_22102);
and U24965 (N_24965,N_23927,N_22155);
and U24966 (N_24966,N_22030,N_22587);
nor U24967 (N_24967,N_22942,N_22054);
and U24968 (N_24968,N_23613,N_22564);
nor U24969 (N_24969,N_23342,N_23648);
nor U24970 (N_24970,N_22074,N_23145);
nand U24971 (N_24971,N_22881,N_22574);
or U24972 (N_24972,N_22226,N_23562);
or U24973 (N_24973,N_23327,N_22874);
or U24974 (N_24974,N_22183,N_22344);
and U24975 (N_24975,N_23452,N_22973);
nand U24976 (N_24976,N_22860,N_23991);
and U24977 (N_24977,N_22050,N_22280);
and U24978 (N_24978,N_23588,N_23866);
and U24979 (N_24979,N_23009,N_23603);
or U24980 (N_24980,N_23447,N_22370);
and U24981 (N_24981,N_22321,N_23793);
or U24982 (N_24982,N_23484,N_23041);
and U24983 (N_24983,N_23671,N_22025);
nand U24984 (N_24984,N_23541,N_23660);
or U24985 (N_24985,N_23254,N_23709);
nand U24986 (N_24986,N_22724,N_23594);
nor U24987 (N_24987,N_23503,N_22413);
nand U24988 (N_24988,N_23404,N_23778);
or U24989 (N_24989,N_22026,N_23714);
or U24990 (N_24990,N_23800,N_23684);
or U24991 (N_24991,N_22398,N_23272);
nor U24992 (N_24992,N_23290,N_22968);
and U24993 (N_24993,N_22837,N_23742);
or U24994 (N_24994,N_23792,N_22048);
and U24995 (N_24995,N_23697,N_23506);
nand U24996 (N_24996,N_23166,N_23523);
or U24997 (N_24997,N_22739,N_22703);
xnor U24998 (N_24998,N_23929,N_23379);
nor U24999 (N_24999,N_23520,N_22372);
and U25000 (N_25000,N_23296,N_22407);
and U25001 (N_25001,N_22657,N_22279);
nor U25002 (N_25002,N_23126,N_23544);
and U25003 (N_25003,N_22109,N_22513);
or U25004 (N_25004,N_23353,N_22192);
nor U25005 (N_25005,N_23405,N_23060);
and U25006 (N_25006,N_23748,N_23485);
nand U25007 (N_25007,N_22609,N_23187);
or U25008 (N_25008,N_22444,N_22390);
nand U25009 (N_25009,N_23141,N_23436);
nand U25010 (N_25010,N_22122,N_22100);
and U25011 (N_25011,N_22507,N_22014);
or U25012 (N_25012,N_23829,N_23653);
nor U25013 (N_25013,N_23527,N_22061);
nand U25014 (N_25014,N_23595,N_23233);
and U25015 (N_25015,N_22093,N_22480);
nand U25016 (N_25016,N_22635,N_23681);
and U25017 (N_25017,N_23554,N_23933);
or U25018 (N_25018,N_23901,N_22335);
nor U25019 (N_25019,N_23638,N_22102);
and U25020 (N_25020,N_22194,N_23788);
and U25021 (N_25021,N_22982,N_22475);
nand U25022 (N_25022,N_23901,N_23584);
and U25023 (N_25023,N_23970,N_22100);
and U25024 (N_25024,N_23878,N_23517);
nor U25025 (N_25025,N_23466,N_22893);
and U25026 (N_25026,N_23525,N_23432);
or U25027 (N_25027,N_22878,N_22402);
nand U25028 (N_25028,N_23676,N_22781);
and U25029 (N_25029,N_23008,N_23266);
nand U25030 (N_25030,N_22641,N_22210);
and U25031 (N_25031,N_22015,N_22287);
nand U25032 (N_25032,N_22368,N_23636);
nor U25033 (N_25033,N_22720,N_22810);
nand U25034 (N_25034,N_23413,N_22220);
and U25035 (N_25035,N_23792,N_23543);
and U25036 (N_25036,N_23256,N_22207);
and U25037 (N_25037,N_22913,N_23424);
or U25038 (N_25038,N_23156,N_22823);
or U25039 (N_25039,N_22537,N_23918);
and U25040 (N_25040,N_23917,N_22776);
or U25041 (N_25041,N_22724,N_22690);
and U25042 (N_25042,N_23580,N_23949);
nor U25043 (N_25043,N_23888,N_23838);
xnor U25044 (N_25044,N_23270,N_22002);
nand U25045 (N_25045,N_23913,N_22813);
or U25046 (N_25046,N_22174,N_22424);
nor U25047 (N_25047,N_22097,N_23269);
xnor U25048 (N_25048,N_22515,N_22636);
and U25049 (N_25049,N_22129,N_22974);
and U25050 (N_25050,N_22527,N_22299);
and U25051 (N_25051,N_22674,N_23820);
nand U25052 (N_25052,N_23267,N_23477);
and U25053 (N_25053,N_23339,N_23398);
and U25054 (N_25054,N_22015,N_23174);
and U25055 (N_25055,N_23285,N_22257);
nor U25056 (N_25056,N_23414,N_23496);
or U25057 (N_25057,N_23559,N_23982);
nand U25058 (N_25058,N_23848,N_22759);
nor U25059 (N_25059,N_22559,N_23612);
or U25060 (N_25060,N_22480,N_22906);
nor U25061 (N_25061,N_23520,N_23536);
nor U25062 (N_25062,N_23857,N_22521);
or U25063 (N_25063,N_22651,N_22380);
nand U25064 (N_25064,N_22478,N_22097);
xor U25065 (N_25065,N_23257,N_23970);
or U25066 (N_25066,N_22716,N_23124);
and U25067 (N_25067,N_22647,N_23391);
or U25068 (N_25068,N_22388,N_22335);
nor U25069 (N_25069,N_23953,N_23793);
or U25070 (N_25070,N_23249,N_22188);
and U25071 (N_25071,N_23683,N_23769);
nand U25072 (N_25072,N_22747,N_22295);
and U25073 (N_25073,N_22804,N_23462);
nand U25074 (N_25074,N_23722,N_22472);
nor U25075 (N_25075,N_23620,N_22113);
and U25076 (N_25076,N_22928,N_22474);
and U25077 (N_25077,N_22776,N_22718);
nor U25078 (N_25078,N_22764,N_23811);
nand U25079 (N_25079,N_23431,N_23331);
nand U25080 (N_25080,N_22355,N_23354);
and U25081 (N_25081,N_23445,N_23750);
or U25082 (N_25082,N_22240,N_23098);
nand U25083 (N_25083,N_23601,N_22760);
or U25084 (N_25084,N_23489,N_22673);
or U25085 (N_25085,N_22689,N_22386);
and U25086 (N_25086,N_23703,N_23183);
and U25087 (N_25087,N_22111,N_23772);
and U25088 (N_25088,N_22570,N_23543);
nand U25089 (N_25089,N_23969,N_23449);
nand U25090 (N_25090,N_22767,N_23749);
nand U25091 (N_25091,N_22402,N_23842);
nand U25092 (N_25092,N_22702,N_23535);
and U25093 (N_25093,N_23193,N_23939);
nand U25094 (N_25094,N_22051,N_23447);
nor U25095 (N_25095,N_23036,N_23500);
and U25096 (N_25096,N_23577,N_22543);
nor U25097 (N_25097,N_22387,N_23302);
and U25098 (N_25098,N_23457,N_23827);
nor U25099 (N_25099,N_22083,N_22501);
nand U25100 (N_25100,N_22677,N_22938);
nand U25101 (N_25101,N_22675,N_22333);
or U25102 (N_25102,N_22893,N_22030);
or U25103 (N_25103,N_23596,N_22780);
or U25104 (N_25104,N_23027,N_22928);
or U25105 (N_25105,N_22119,N_23634);
or U25106 (N_25106,N_23140,N_23833);
nor U25107 (N_25107,N_22484,N_23272);
nand U25108 (N_25108,N_22915,N_23694);
or U25109 (N_25109,N_22680,N_22634);
nor U25110 (N_25110,N_22404,N_23054);
or U25111 (N_25111,N_23703,N_22829);
nand U25112 (N_25112,N_23510,N_23763);
nand U25113 (N_25113,N_22774,N_23376);
nor U25114 (N_25114,N_22010,N_22858);
or U25115 (N_25115,N_22558,N_22149);
nand U25116 (N_25116,N_22348,N_23282);
and U25117 (N_25117,N_22316,N_22893);
nand U25118 (N_25118,N_22314,N_23616);
nor U25119 (N_25119,N_23630,N_22737);
nor U25120 (N_25120,N_22057,N_22158);
and U25121 (N_25121,N_23953,N_22564);
xnor U25122 (N_25122,N_22565,N_22474);
nor U25123 (N_25123,N_22357,N_23616);
nand U25124 (N_25124,N_23781,N_22891);
nor U25125 (N_25125,N_23799,N_23773);
nand U25126 (N_25126,N_22974,N_23359);
nand U25127 (N_25127,N_23541,N_23525);
nand U25128 (N_25128,N_22670,N_23317);
or U25129 (N_25129,N_23101,N_23921);
nor U25130 (N_25130,N_23108,N_22697);
and U25131 (N_25131,N_23620,N_23869);
nand U25132 (N_25132,N_22288,N_23319);
and U25133 (N_25133,N_23320,N_22375);
and U25134 (N_25134,N_23435,N_22744);
nand U25135 (N_25135,N_23669,N_23471);
nor U25136 (N_25136,N_23593,N_22287);
nor U25137 (N_25137,N_23093,N_22817);
nand U25138 (N_25138,N_23740,N_22043);
nor U25139 (N_25139,N_23860,N_22626);
nand U25140 (N_25140,N_22023,N_23780);
nand U25141 (N_25141,N_22007,N_23898);
nor U25142 (N_25142,N_22428,N_22940);
nor U25143 (N_25143,N_22695,N_22336);
and U25144 (N_25144,N_22635,N_22830);
and U25145 (N_25145,N_22489,N_22816);
nand U25146 (N_25146,N_23703,N_23742);
nor U25147 (N_25147,N_23342,N_23980);
nand U25148 (N_25148,N_22416,N_23495);
or U25149 (N_25149,N_23752,N_23163);
or U25150 (N_25150,N_22227,N_22610);
nor U25151 (N_25151,N_22642,N_23343);
and U25152 (N_25152,N_23397,N_23412);
and U25153 (N_25153,N_22508,N_22912);
or U25154 (N_25154,N_23788,N_22138);
xnor U25155 (N_25155,N_23457,N_23760);
and U25156 (N_25156,N_23284,N_23861);
and U25157 (N_25157,N_23022,N_22311);
nand U25158 (N_25158,N_23849,N_23401);
nor U25159 (N_25159,N_22793,N_23285);
and U25160 (N_25160,N_23784,N_23672);
nand U25161 (N_25161,N_23248,N_22223);
nand U25162 (N_25162,N_23139,N_22700);
nand U25163 (N_25163,N_23980,N_22825);
nand U25164 (N_25164,N_22597,N_22007);
nor U25165 (N_25165,N_23653,N_23425);
or U25166 (N_25166,N_23901,N_23753);
and U25167 (N_25167,N_23765,N_22075);
xnor U25168 (N_25168,N_23506,N_22874);
nor U25169 (N_25169,N_23286,N_23208);
nor U25170 (N_25170,N_22390,N_23281);
nor U25171 (N_25171,N_23954,N_22215);
nor U25172 (N_25172,N_23083,N_22470);
nor U25173 (N_25173,N_22816,N_22108);
nor U25174 (N_25174,N_22021,N_23547);
nand U25175 (N_25175,N_22490,N_23464);
nor U25176 (N_25176,N_22699,N_22794);
nand U25177 (N_25177,N_22376,N_22313);
and U25178 (N_25178,N_22733,N_23059);
and U25179 (N_25179,N_22311,N_22941);
or U25180 (N_25180,N_23969,N_23790);
or U25181 (N_25181,N_22750,N_23602);
nand U25182 (N_25182,N_22617,N_22755);
and U25183 (N_25183,N_22293,N_22103);
nand U25184 (N_25184,N_22402,N_23428);
or U25185 (N_25185,N_22661,N_22114);
nand U25186 (N_25186,N_23707,N_23782);
or U25187 (N_25187,N_23833,N_23570);
and U25188 (N_25188,N_23231,N_23742);
and U25189 (N_25189,N_22358,N_22362);
nor U25190 (N_25190,N_22000,N_22552);
nor U25191 (N_25191,N_23568,N_22789);
nor U25192 (N_25192,N_23301,N_23967);
nand U25193 (N_25193,N_22144,N_22746);
nand U25194 (N_25194,N_22902,N_23567);
and U25195 (N_25195,N_23287,N_23819);
nor U25196 (N_25196,N_22538,N_22704);
or U25197 (N_25197,N_22786,N_22186);
nand U25198 (N_25198,N_23440,N_23412);
nand U25199 (N_25199,N_23593,N_22956);
nand U25200 (N_25200,N_22885,N_23984);
nand U25201 (N_25201,N_22985,N_23027);
nand U25202 (N_25202,N_23573,N_23133);
nand U25203 (N_25203,N_22176,N_23048);
nor U25204 (N_25204,N_22555,N_23075);
nor U25205 (N_25205,N_22896,N_23013);
nor U25206 (N_25206,N_22512,N_23336);
nor U25207 (N_25207,N_23016,N_23215);
or U25208 (N_25208,N_23256,N_22550);
and U25209 (N_25209,N_22042,N_22600);
and U25210 (N_25210,N_23340,N_23009);
and U25211 (N_25211,N_22703,N_22408);
nor U25212 (N_25212,N_23424,N_23482);
nand U25213 (N_25213,N_23539,N_22339);
or U25214 (N_25214,N_23831,N_23724);
and U25215 (N_25215,N_23286,N_23545);
nor U25216 (N_25216,N_22614,N_23444);
and U25217 (N_25217,N_22121,N_22685);
and U25218 (N_25218,N_22086,N_23866);
nor U25219 (N_25219,N_23225,N_22405);
nand U25220 (N_25220,N_22303,N_22469);
nand U25221 (N_25221,N_23584,N_22501);
and U25222 (N_25222,N_22136,N_22035);
xor U25223 (N_25223,N_23173,N_22988);
nand U25224 (N_25224,N_23436,N_23093);
and U25225 (N_25225,N_22007,N_23856);
or U25226 (N_25226,N_22556,N_22260);
nor U25227 (N_25227,N_22442,N_23807);
nand U25228 (N_25228,N_22650,N_22260);
nor U25229 (N_25229,N_23510,N_22314);
nand U25230 (N_25230,N_22510,N_23244);
nor U25231 (N_25231,N_22322,N_22031);
and U25232 (N_25232,N_22949,N_22219);
nand U25233 (N_25233,N_22048,N_22316);
or U25234 (N_25234,N_23117,N_22220);
and U25235 (N_25235,N_23475,N_23266);
or U25236 (N_25236,N_23197,N_22015);
and U25237 (N_25237,N_22996,N_23543);
nor U25238 (N_25238,N_22095,N_22875);
nor U25239 (N_25239,N_22248,N_23514);
or U25240 (N_25240,N_23352,N_22430);
and U25241 (N_25241,N_23171,N_22104);
or U25242 (N_25242,N_22742,N_23469);
nor U25243 (N_25243,N_23602,N_23179);
nor U25244 (N_25244,N_23899,N_23949);
or U25245 (N_25245,N_22198,N_23611);
xnor U25246 (N_25246,N_22899,N_22156);
nand U25247 (N_25247,N_22140,N_23806);
nand U25248 (N_25248,N_22031,N_22689);
or U25249 (N_25249,N_22237,N_22273);
nand U25250 (N_25250,N_22655,N_22046);
nor U25251 (N_25251,N_22070,N_23270);
nor U25252 (N_25252,N_22556,N_23405);
nor U25253 (N_25253,N_23815,N_23046);
or U25254 (N_25254,N_22578,N_23711);
xor U25255 (N_25255,N_22885,N_23803);
nand U25256 (N_25256,N_22323,N_22427);
nand U25257 (N_25257,N_23235,N_22296);
nor U25258 (N_25258,N_22509,N_23812);
nand U25259 (N_25259,N_23889,N_22414);
nor U25260 (N_25260,N_23898,N_23341);
or U25261 (N_25261,N_22077,N_23652);
nand U25262 (N_25262,N_22156,N_22578);
nor U25263 (N_25263,N_23779,N_22577);
nand U25264 (N_25264,N_22856,N_22585);
nand U25265 (N_25265,N_23298,N_22162);
xnor U25266 (N_25266,N_23675,N_22615);
nand U25267 (N_25267,N_23915,N_23927);
or U25268 (N_25268,N_23860,N_22153);
or U25269 (N_25269,N_23087,N_23734);
nor U25270 (N_25270,N_22114,N_23718);
or U25271 (N_25271,N_22895,N_22033);
nor U25272 (N_25272,N_23856,N_23714);
and U25273 (N_25273,N_22402,N_23832);
or U25274 (N_25274,N_22231,N_22415);
nand U25275 (N_25275,N_22643,N_22733);
and U25276 (N_25276,N_22176,N_23819);
nor U25277 (N_25277,N_23238,N_23914);
nand U25278 (N_25278,N_23225,N_22224);
and U25279 (N_25279,N_22850,N_23339);
or U25280 (N_25280,N_22365,N_22094);
and U25281 (N_25281,N_22510,N_22647);
nand U25282 (N_25282,N_23165,N_22254);
and U25283 (N_25283,N_22489,N_23180);
nand U25284 (N_25284,N_22414,N_23572);
or U25285 (N_25285,N_23739,N_22484);
nand U25286 (N_25286,N_22025,N_23181);
or U25287 (N_25287,N_22697,N_23200);
nand U25288 (N_25288,N_23087,N_23003);
and U25289 (N_25289,N_22620,N_22303);
nor U25290 (N_25290,N_23149,N_23846);
nor U25291 (N_25291,N_22686,N_23611);
nand U25292 (N_25292,N_23343,N_22667);
nor U25293 (N_25293,N_22284,N_23316);
nand U25294 (N_25294,N_22353,N_23153);
or U25295 (N_25295,N_23805,N_23172);
or U25296 (N_25296,N_23097,N_22228);
and U25297 (N_25297,N_23822,N_22013);
or U25298 (N_25298,N_23453,N_23322);
nor U25299 (N_25299,N_23243,N_23440);
nor U25300 (N_25300,N_22919,N_23920);
and U25301 (N_25301,N_22768,N_22415);
and U25302 (N_25302,N_23731,N_23847);
or U25303 (N_25303,N_23328,N_22486);
and U25304 (N_25304,N_23564,N_22582);
nand U25305 (N_25305,N_22621,N_23761);
nand U25306 (N_25306,N_23004,N_22031);
and U25307 (N_25307,N_22594,N_23536);
and U25308 (N_25308,N_23111,N_23942);
nand U25309 (N_25309,N_22588,N_23494);
or U25310 (N_25310,N_22789,N_22684);
and U25311 (N_25311,N_23504,N_22882);
nand U25312 (N_25312,N_23777,N_23829);
nor U25313 (N_25313,N_22926,N_22537);
and U25314 (N_25314,N_23698,N_23653);
and U25315 (N_25315,N_23358,N_23014);
and U25316 (N_25316,N_22117,N_23734);
nand U25317 (N_25317,N_23274,N_22196);
nand U25318 (N_25318,N_23226,N_22070);
nor U25319 (N_25319,N_23875,N_23138);
and U25320 (N_25320,N_23255,N_22157);
nand U25321 (N_25321,N_23511,N_23746);
nor U25322 (N_25322,N_22385,N_23580);
nor U25323 (N_25323,N_22516,N_23080);
nor U25324 (N_25324,N_22268,N_23377);
nor U25325 (N_25325,N_23344,N_22158);
nand U25326 (N_25326,N_23155,N_23204);
or U25327 (N_25327,N_23426,N_23042);
nand U25328 (N_25328,N_23660,N_22794);
and U25329 (N_25329,N_22744,N_22810);
nor U25330 (N_25330,N_23170,N_22840);
nand U25331 (N_25331,N_23827,N_22520);
nand U25332 (N_25332,N_23210,N_23966);
and U25333 (N_25333,N_22200,N_22132);
nand U25334 (N_25334,N_23704,N_22782);
or U25335 (N_25335,N_23820,N_23172);
nor U25336 (N_25336,N_22567,N_22745);
nor U25337 (N_25337,N_23414,N_23556);
nor U25338 (N_25338,N_23885,N_22860);
nor U25339 (N_25339,N_23245,N_22723);
nand U25340 (N_25340,N_22148,N_23479);
nand U25341 (N_25341,N_23874,N_22399);
or U25342 (N_25342,N_23035,N_23794);
or U25343 (N_25343,N_23105,N_22718);
and U25344 (N_25344,N_22157,N_22779);
or U25345 (N_25345,N_22189,N_22586);
or U25346 (N_25346,N_23909,N_22987);
nor U25347 (N_25347,N_22018,N_23606);
nor U25348 (N_25348,N_22812,N_22638);
nor U25349 (N_25349,N_23625,N_22689);
nand U25350 (N_25350,N_23342,N_23197);
and U25351 (N_25351,N_22628,N_23129);
nand U25352 (N_25352,N_23376,N_23544);
nor U25353 (N_25353,N_23534,N_23707);
and U25354 (N_25354,N_23088,N_22446);
nand U25355 (N_25355,N_22702,N_23573);
or U25356 (N_25356,N_22500,N_22084);
nor U25357 (N_25357,N_22564,N_22919);
nand U25358 (N_25358,N_22285,N_23229);
and U25359 (N_25359,N_23759,N_22962);
and U25360 (N_25360,N_22685,N_22034);
or U25361 (N_25361,N_22810,N_22206);
and U25362 (N_25362,N_23813,N_23105);
nand U25363 (N_25363,N_23757,N_22196);
nand U25364 (N_25364,N_22495,N_23715);
nor U25365 (N_25365,N_22077,N_23266);
nor U25366 (N_25366,N_23045,N_22672);
nand U25367 (N_25367,N_23477,N_23103);
and U25368 (N_25368,N_23083,N_23245);
nor U25369 (N_25369,N_22657,N_23886);
nor U25370 (N_25370,N_23736,N_22121);
and U25371 (N_25371,N_23634,N_23346);
nand U25372 (N_25372,N_23609,N_23113);
nor U25373 (N_25373,N_23146,N_22765);
nand U25374 (N_25374,N_23534,N_23097);
nor U25375 (N_25375,N_22362,N_23015);
or U25376 (N_25376,N_22986,N_23349);
and U25377 (N_25377,N_22576,N_23360);
or U25378 (N_25378,N_22856,N_23903);
and U25379 (N_25379,N_23325,N_22332);
or U25380 (N_25380,N_22790,N_23291);
or U25381 (N_25381,N_23354,N_23107);
and U25382 (N_25382,N_23680,N_23725);
nor U25383 (N_25383,N_23398,N_23358);
and U25384 (N_25384,N_22642,N_22079);
and U25385 (N_25385,N_23174,N_22124);
xor U25386 (N_25386,N_22248,N_22701);
or U25387 (N_25387,N_23355,N_22524);
nand U25388 (N_25388,N_22872,N_22367);
nor U25389 (N_25389,N_23329,N_23840);
nand U25390 (N_25390,N_22529,N_22629);
and U25391 (N_25391,N_23321,N_22369);
or U25392 (N_25392,N_23899,N_23415);
nand U25393 (N_25393,N_22048,N_22918);
nand U25394 (N_25394,N_22408,N_22780);
nand U25395 (N_25395,N_23223,N_22159);
or U25396 (N_25396,N_23763,N_22830);
and U25397 (N_25397,N_23677,N_22750);
and U25398 (N_25398,N_22958,N_22487);
or U25399 (N_25399,N_23116,N_22594);
nor U25400 (N_25400,N_22167,N_22298);
or U25401 (N_25401,N_22867,N_23994);
and U25402 (N_25402,N_22110,N_23505);
and U25403 (N_25403,N_22521,N_23261);
nand U25404 (N_25404,N_22011,N_22377);
and U25405 (N_25405,N_23115,N_23714);
nand U25406 (N_25406,N_23858,N_22387);
and U25407 (N_25407,N_22145,N_22609);
nand U25408 (N_25408,N_22928,N_22124);
nor U25409 (N_25409,N_22694,N_23250);
nor U25410 (N_25410,N_22753,N_22214);
nand U25411 (N_25411,N_22010,N_22106);
nand U25412 (N_25412,N_23725,N_22981);
and U25413 (N_25413,N_23017,N_22228);
nor U25414 (N_25414,N_22631,N_23020);
or U25415 (N_25415,N_22536,N_23751);
or U25416 (N_25416,N_23958,N_23223);
nor U25417 (N_25417,N_23260,N_23592);
or U25418 (N_25418,N_22774,N_22787);
nor U25419 (N_25419,N_23968,N_23941);
nand U25420 (N_25420,N_22527,N_22646);
or U25421 (N_25421,N_22783,N_23539);
nand U25422 (N_25422,N_22984,N_23744);
nor U25423 (N_25423,N_23599,N_23156);
nand U25424 (N_25424,N_23329,N_22701);
and U25425 (N_25425,N_23983,N_23107);
and U25426 (N_25426,N_23161,N_22803);
or U25427 (N_25427,N_23718,N_22982);
or U25428 (N_25428,N_23971,N_23176);
or U25429 (N_25429,N_22811,N_22903);
or U25430 (N_25430,N_23021,N_22295);
and U25431 (N_25431,N_22539,N_23780);
or U25432 (N_25432,N_23434,N_23524);
nand U25433 (N_25433,N_23636,N_23252);
nand U25434 (N_25434,N_22108,N_22923);
nand U25435 (N_25435,N_23650,N_22468);
or U25436 (N_25436,N_22291,N_22804);
nand U25437 (N_25437,N_22893,N_23789);
nor U25438 (N_25438,N_23077,N_23393);
or U25439 (N_25439,N_22392,N_22586);
nor U25440 (N_25440,N_23393,N_22696);
or U25441 (N_25441,N_22841,N_23743);
and U25442 (N_25442,N_22912,N_22306);
or U25443 (N_25443,N_23128,N_23004);
nand U25444 (N_25444,N_23842,N_22588);
or U25445 (N_25445,N_23925,N_22879);
or U25446 (N_25446,N_22066,N_22576);
xnor U25447 (N_25447,N_22649,N_23739);
nand U25448 (N_25448,N_23514,N_22531);
nor U25449 (N_25449,N_22466,N_22108);
or U25450 (N_25450,N_23871,N_22915);
nor U25451 (N_25451,N_22234,N_22893);
nor U25452 (N_25452,N_23882,N_23418);
nand U25453 (N_25453,N_23526,N_23341);
nand U25454 (N_25454,N_22311,N_23412);
or U25455 (N_25455,N_23044,N_23765);
or U25456 (N_25456,N_22502,N_22647);
or U25457 (N_25457,N_23260,N_23496);
and U25458 (N_25458,N_22003,N_23584);
and U25459 (N_25459,N_22939,N_23467);
or U25460 (N_25460,N_23889,N_23261);
nor U25461 (N_25461,N_22061,N_23427);
nor U25462 (N_25462,N_22394,N_23054);
or U25463 (N_25463,N_22996,N_22867);
nor U25464 (N_25464,N_22741,N_22596);
xor U25465 (N_25465,N_22887,N_22301);
or U25466 (N_25466,N_22121,N_22705);
or U25467 (N_25467,N_22690,N_23276);
nor U25468 (N_25468,N_23040,N_23637);
and U25469 (N_25469,N_23029,N_22436);
nand U25470 (N_25470,N_22916,N_22673);
and U25471 (N_25471,N_23234,N_23200);
nand U25472 (N_25472,N_22804,N_22571);
nand U25473 (N_25473,N_22988,N_22918);
nand U25474 (N_25474,N_23465,N_23201);
nand U25475 (N_25475,N_23602,N_23724);
nor U25476 (N_25476,N_23308,N_23788);
nor U25477 (N_25477,N_22562,N_23405);
or U25478 (N_25478,N_22015,N_22683);
nor U25479 (N_25479,N_23077,N_22340);
nor U25480 (N_25480,N_22691,N_23840);
and U25481 (N_25481,N_22512,N_23661);
nand U25482 (N_25482,N_22169,N_23766);
and U25483 (N_25483,N_23091,N_22626);
or U25484 (N_25484,N_22291,N_22553);
or U25485 (N_25485,N_23475,N_23650);
nand U25486 (N_25486,N_22461,N_22973);
nor U25487 (N_25487,N_22354,N_23421);
and U25488 (N_25488,N_23906,N_23400);
nand U25489 (N_25489,N_23542,N_23286);
nor U25490 (N_25490,N_23771,N_23479);
nand U25491 (N_25491,N_23692,N_23543);
and U25492 (N_25492,N_23929,N_23651);
nand U25493 (N_25493,N_23512,N_22246);
or U25494 (N_25494,N_23649,N_22065);
nand U25495 (N_25495,N_22537,N_23960);
nor U25496 (N_25496,N_22074,N_23638);
nor U25497 (N_25497,N_23976,N_23633);
or U25498 (N_25498,N_22211,N_22102);
nor U25499 (N_25499,N_23750,N_22084);
or U25500 (N_25500,N_22965,N_22112);
nor U25501 (N_25501,N_22582,N_23750);
or U25502 (N_25502,N_22872,N_23472);
or U25503 (N_25503,N_22236,N_23850);
or U25504 (N_25504,N_23003,N_22635);
nor U25505 (N_25505,N_23149,N_22553);
or U25506 (N_25506,N_23694,N_23205);
nor U25507 (N_25507,N_22921,N_22895);
or U25508 (N_25508,N_22219,N_22881);
and U25509 (N_25509,N_23777,N_22448);
or U25510 (N_25510,N_23612,N_22929);
nor U25511 (N_25511,N_23372,N_23593);
or U25512 (N_25512,N_23305,N_22524);
nor U25513 (N_25513,N_23870,N_22861);
nand U25514 (N_25514,N_23804,N_23703);
or U25515 (N_25515,N_22755,N_23039);
nor U25516 (N_25516,N_22064,N_22900);
nand U25517 (N_25517,N_23496,N_22628);
nor U25518 (N_25518,N_23478,N_22417);
nor U25519 (N_25519,N_22357,N_22994);
and U25520 (N_25520,N_22159,N_22361);
nor U25521 (N_25521,N_23936,N_23593);
or U25522 (N_25522,N_23682,N_23918);
nand U25523 (N_25523,N_22683,N_23497);
nand U25524 (N_25524,N_22847,N_23599);
nor U25525 (N_25525,N_23665,N_22085);
nand U25526 (N_25526,N_23929,N_23532);
and U25527 (N_25527,N_22825,N_22719);
and U25528 (N_25528,N_22621,N_22372);
and U25529 (N_25529,N_22913,N_23582);
nand U25530 (N_25530,N_23406,N_22390);
nor U25531 (N_25531,N_22554,N_23009);
nor U25532 (N_25532,N_22698,N_23460);
or U25533 (N_25533,N_22663,N_22971);
or U25534 (N_25534,N_22864,N_22204);
or U25535 (N_25535,N_22923,N_23108);
or U25536 (N_25536,N_22530,N_23074);
or U25537 (N_25537,N_22786,N_23368);
nand U25538 (N_25538,N_23577,N_22970);
xnor U25539 (N_25539,N_22795,N_23080);
and U25540 (N_25540,N_23306,N_22154);
or U25541 (N_25541,N_22369,N_23030);
and U25542 (N_25542,N_23149,N_22421);
or U25543 (N_25543,N_22163,N_23946);
or U25544 (N_25544,N_22094,N_22678);
nor U25545 (N_25545,N_23971,N_23522);
nand U25546 (N_25546,N_23486,N_22219);
or U25547 (N_25547,N_22756,N_23411);
nand U25548 (N_25548,N_22573,N_23432);
nor U25549 (N_25549,N_22609,N_23155);
and U25550 (N_25550,N_23220,N_23059);
nor U25551 (N_25551,N_23932,N_22890);
or U25552 (N_25552,N_23003,N_22575);
or U25553 (N_25553,N_23757,N_22356);
xor U25554 (N_25554,N_23388,N_22627);
nor U25555 (N_25555,N_22013,N_23770);
nand U25556 (N_25556,N_22789,N_22943);
nand U25557 (N_25557,N_22836,N_22820);
and U25558 (N_25558,N_22437,N_22067);
nor U25559 (N_25559,N_23695,N_23218);
and U25560 (N_25560,N_22453,N_22241);
or U25561 (N_25561,N_22017,N_23672);
and U25562 (N_25562,N_22714,N_23802);
nor U25563 (N_25563,N_22634,N_23974);
nor U25564 (N_25564,N_22980,N_23703);
nand U25565 (N_25565,N_23455,N_23791);
or U25566 (N_25566,N_23636,N_23524);
nand U25567 (N_25567,N_23687,N_22219);
nand U25568 (N_25568,N_23340,N_23151);
and U25569 (N_25569,N_22631,N_23126);
nand U25570 (N_25570,N_22981,N_22900);
nor U25571 (N_25571,N_22353,N_22163);
or U25572 (N_25572,N_22870,N_23236);
and U25573 (N_25573,N_22499,N_22066);
and U25574 (N_25574,N_22088,N_23082);
nor U25575 (N_25575,N_22250,N_23502);
or U25576 (N_25576,N_23085,N_22400);
and U25577 (N_25577,N_22381,N_22384);
nand U25578 (N_25578,N_22062,N_23808);
nor U25579 (N_25579,N_23603,N_22076);
or U25580 (N_25580,N_23733,N_23992);
nor U25581 (N_25581,N_23721,N_22715);
nand U25582 (N_25582,N_23220,N_23331);
or U25583 (N_25583,N_22170,N_22158);
and U25584 (N_25584,N_23636,N_23881);
nor U25585 (N_25585,N_23101,N_23522);
nand U25586 (N_25586,N_22781,N_23349);
nor U25587 (N_25587,N_23420,N_23751);
nor U25588 (N_25588,N_23715,N_23021);
nand U25589 (N_25589,N_23515,N_22437);
nand U25590 (N_25590,N_22916,N_22419);
and U25591 (N_25591,N_22363,N_22044);
nand U25592 (N_25592,N_22855,N_23769);
or U25593 (N_25593,N_23176,N_22453);
or U25594 (N_25594,N_23159,N_23629);
nor U25595 (N_25595,N_23213,N_22114);
and U25596 (N_25596,N_22304,N_22835);
xnor U25597 (N_25597,N_23706,N_22170);
nor U25598 (N_25598,N_23132,N_23014);
nand U25599 (N_25599,N_23076,N_22479);
and U25600 (N_25600,N_22908,N_22265);
nand U25601 (N_25601,N_23393,N_22275);
xor U25602 (N_25602,N_23361,N_22171);
and U25603 (N_25603,N_23480,N_22105);
nand U25604 (N_25604,N_22512,N_23511);
nor U25605 (N_25605,N_23907,N_23732);
or U25606 (N_25606,N_22985,N_23577);
or U25607 (N_25607,N_22991,N_22736);
nand U25608 (N_25608,N_23203,N_22348);
or U25609 (N_25609,N_22262,N_22488);
and U25610 (N_25610,N_23500,N_22835);
or U25611 (N_25611,N_22007,N_22537);
nand U25612 (N_25612,N_22907,N_23674);
xnor U25613 (N_25613,N_23809,N_23245);
and U25614 (N_25614,N_22805,N_22860);
nand U25615 (N_25615,N_22221,N_22639);
and U25616 (N_25616,N_22673,N_23859);
or U25617 (N_25617,N_23771,N_23491);
nor U25618 (N_25618,N_23732,N_23917);
nand U25619 (N_25619,N_22135,N_22998);
or U25620 (N_25620,N_22998,N_22515);
xor U25621 (N_25621,N_22047,N_23115);
nor U25622 (N_25622,N_23672,N_22257);
or U25623 (N_25623,N_22273,N_22488);
nand U25624 (N_25624,N_22809,N_23481);
nor U25625 (N_25625,N_22146,N_23809);
or U25626 (N_25626,N_22539,N_22433);
and U25627 (N_25627,N_22479,N_23111);
nand U25628 (N_25628,N_23861,N_23243);
or U25629 (N_25629,N_22060,N_22274);
and U25630 (N_25630,N_22842,N_22634);
or U25631 (N_25631,N_23637,N_23216);
nand U25632 (N_25632,N_23337,N_23935);
and U25633 (N_25633,N_23681,N_22593);
nor U25634 (N_25634,N_23207,N_23950);
nor U25635 (N_25635,N_23738,N_23235);
or U25636 (N_25636,N_23301,N_23446);
nand U25637 (N_25637,N_23687,N_22808);
nand U25638 (N_25638,N_22695,N_23940);
or U25639 (N_25639,N_23885,N_22804);
xor U25640 (N_25640,N_22108,N_22538);
or U25641 (N_25641,N_23038,N_22829);
and U25642 (N_25642,N_22910,N_23510);
or U25643 (N_25643,N_22997,N_22071);
nand U25644 (N_25644,N_22343,N_22901);
or U25645 (N_25645,N_22239,N_22992);
or U25646 (N_25646,N_23976,N_22616);
or U25647 (N_25647,N_23018,N_22868);
nand U25648 (N_25648,N_22080,N_23533);
nor U25649 (N_25649,N_23207,N_22431);
or U25650 (N_25650,N_23273,N_23457);
and U25651 (N_25651,N_23064,N_23789);
nor U25652 (N_25652,N_23234,N_23982);
or U25653 (N_25653,N_22305,N_23711);
nor U25654 (N_25654,N_22704,N_23752);
nor U25655 (N_25655,N_23744,N_22260);
or U25656 (N_25656,N_23792,N_23931);
or U25657 (N_25657,N_22691,N_23456);
xnor U25658 (N_25658,N_23025,N_22697);
or U25659 (N_25659,N_22220,N_22182);
nand U25660 (N_25660,N_22149,N_22530);
nor U25661 (N_25661,N_22319,N_22118);
or U25662 (N_25662,N_23311,N_23922);
and U25663 (N_25663,N_23006,N_23641);
nor U25664 (N_25664,N_22765,N_23157);
nor U25665 (N_25665,N_22807,N_23330);
or U25666 (N_25666,N_22123,N_22055);
and U25667 (N_25667,N_22900,N_22018);
xor U25668 (N_25668,N_22967,N_23463);
or U25669 (N_25669,N_22018,N_22523);
or U25670 (N_25670,N_22694,N_23803);
nand U25671 (N_25671,N_23464,N_23101);
nand U25672 (N_25672,N_23967,N_23065);
and U25673 (N_25673,N_22102,N_23743);
or U25674 (N_25674,N_23460,N_23506);
nor U25675 (N_25675,N_23207,N_22009);
or U25676 (N_25676,N_22935,N_23823);
and U25677 (N_25677,N_22880,N_23808);
and U25678 (N_25678,N_23370,N_23125);
or U25679 (N_25679,N_22256,N_23683);
and U25680 (N_25680,N_22724,N_23301);
and U25681 (N_25681,N_23417,N_22731);
nand U25682 (N_25682,N_22214,N_23969);
and U25683 (N_25683,N_23570,N_23124);
nand U25684 (N_25684,N_23242,N_22003);
nand U25685 (N_25685,N_23432,N_23217);
nand U25686 (N_25686,N_23681,N_23133);
or U25687 (N_25687,N_23907,N_22392);
or U25688 (N_25688,N_22676,N_23798);
nand U25689 (N_25689,N_23648,N_22016);
and U25690 (N_25690,N_22674,N_22172);
nand U25691 (N_25691,N_23323,N_22878);
nand U25692 (N_25692,N_23066,N_23956);
or U25693 (N_25693,N_23255,N_22990);
nand U25694 (N_25694,N_23406,N_22007);
and U25695 (N_25695,N_23123,N_22729);
nor U25696 (N_25696,N_22176,N_23575);
nor U25697 (N_25697,N_23260,N_23896);
and U25698 (N_25698,N_23509,N_22027);
and U25699 (N_25699,N_22967,N_23219);
nor U25700 (N_25700,N_22802,N_23280);
or U25701 (N_25701,N_22216,N_22143);
and U25702 (N_25702,N_23133,N_22266);
nand U25703 (N_25703,N_22596,N_22248);
nor U25704 (N_25704,N_22234,N_23091);
or U25705 (N_25705,N_22093,N_23338);
nor U25706 (N_25706,N_22186,N_22930);
and U25707 (N_25707,N_22563,N_22577);
nand U25708 (N_25708,N_23274,N_23868);
or U25709 (N_25709,N_22625,N_22265);
or U25710 (N_25710,N_23888,N_22831);
or U25711 (N_25711,N_22786,N_23151);
nor U25712 (N_25712,N_22941,N_22747);
and U25713 (N_25713,N_23206,N_23795);
and U25714 (N_25714,N_23478,N_22661);
nor U25715 (N_25715,N_22932,N_23321);
and U25716 (N_25716,N_23695,N_22173);
nand U25717 (N_25717,N_23841,N_22950);
and U25718 (N_25718,N_23557,N_23430);
or U25719 (N_25719,N_23885,N_22840);
nand U25720 (N_25720,N_22582,N_22866);
xnor U25721 (N_25721,N_23001,N_23374);
nor U25722 (N_25722,N_23304,N_23109);
nor U25723 (N_25723,N_22859,N_22538);
or U25724 (N_25724,N_22334,N_23398);
nand U25725 (N_25725,N_22909,N_23181);
nor U25726 (N_25726,N_22489,N_23206);
or U25727 (N_25727,N_22592,N_23064);
and U25728 (N_25728,N_23501,N_23193);
nor U25729 (N_25729,N_23101,N_23630);
nor U25730 (N_25730,N_22675,N_23798);
nand U25731 (N_25731,N_23482,N_22851);
or U25732 (N_25732,N_22987,N_23380);
or U25733 (N_25733,N_22542,N_23646);
and U25734 (N_25734,N_22539,N_23649);
or U25735 (N_25735,N_22149,N_23460);
or U25736 (N_25736,N_23133,N_22021);
and U25737 (N_25737,N_22485,N_22830);
nand U25738 (N_25738,N_23355,N_22662);
nand U25739 (N_25739,N_23854,N_22904);
or U25740 (N_25740,N_22503,N_22188);
nand U25741 (N_25741,N_22165,N_22241);
or U25742 (N_25742,N_22661,N_22555);
and U25743 (N_25743,N_23464,N_22459);
nand U25744 (N_25744,N_22406,N_22060);
nand U25745 (N_25745,N_23226,N_22786);
nand U25746 (N_25746,N_23469,N_23782);
and U25747 (N_25747,N_22546,N_22736);
nor U25748 (N_25748,N_23947,N_22215);
nor U25749 (N_25749,N_23695,N_22955);
nand U25750 (N_25750,N_23683,N_23583);
nor U25751 (N_25751,N_22986,N_22167);
or U25752 (N_25752,N_23391,N_23754);
and U25753 (N_25753,N_23623,N_22635);
nand U25754 (N_25754,N_23057,N_23272);
and U25755 (N_25755,N_23014,N_22298);
or U25756 (N_25756,N_22379,N_22928);
nor U25757 (N_25757,N_23256,N_23892);
and U25758 (N_25758,N_22592,N_22203);
and U25759 (N_25759,N_22369,N_23822);
nand U25760 (N_25760,N_22474,N_23580);
xor U25761 (N_25761,N_22329,N_22539);
or U25762 (N_25762,N_23412,N_23825);
and U25763 (N_25763,N_23740,N_23632);
or U25764 (N_25764,N_22599,N_22320);
and U25765 (N_25765,N_23683,N_22759);
or U25766 (N_25766,N_23182,N_23596);
nor U25767 (N_25767,N_23677,N_22628);
nor U25768 (N_25768,N_22051,N_22171);
or U25769 (N_25769,N_23948,N_23314);
and U25770 (N_25770,N_22575,N_23816);
or U25771 (N_25771,N_22936,N_23845);
xor U25772 (N_25772,N_23859,N_23403);
xor U25773 (N_25773,N_23523,N_23952);
nor U25774 (N_25774,N_23002,N_22717);
nor U25775 (N_25775,N_23800,N_22554);
nand U25776 (N_25776,N_22849,N_23539);
nand U25777 (N_25777,N_22807,N_22525);
nand U25778 (N_25778,N_23756,N_23450);
nand U25779 (N_25779,N_22955,N_23317);
and U25780 (N_25780,N_23298,N_22056);
nor U25781 (N_25781,N_22672,N_23518);
nand U25782 (N_25782,N_22617,N_23850);
nor U25783 (N_25783,N_22528,N_22098);
nand U25784 (N_25784,N_23562,N_23319);
nand U25785 (N_25785,N_23802,N_23344);
or U25786 (N_25786,N_22262,N_23256);
nor U25787 (N_25787,N_22089,N_23603);
nand U25788 (N_25788,N_23880,N_22206);
nand U25789 (N_25789,N_22303,N_23096);
and U25790 (N_25790,N_22920,N_22414);
nor U25791 (N_25791,N_22435,N_22704);
and U25792 (N_25792,N_22303,N_23624);
or U25793 (N_25793,N_23255,N_22866);
nor U25794 (N_25794,N_22010,N_23600);
nor U25795 (N_25795,N_22818,N_23224);
or U25796 (N_25796,N_23537,N_22799);
nand U25797 (N_25797,N_23286,N_22394);
nand U25798 (N_25798,N_22589,N_22671);
and U25799 (N_25799,N_23591,N_22443);
or U25800 (N_25800,N_23694,N_23952);
and U25801 (N_25801,N_22335,N_23391);
or U25802 (N_25802,N_22479,N_22918);
xnor U25803 (N_25803,N_22372,N_23144);
nand U25804 (N_25804,N_22590,N_23538);
xor U25805 (N_25805,N_23691,N_22137);
nor U25806 (N_25806,N_22313,N_22094);
nand U25807 (N_25807,N_22251,N_23985);
nand U25808 (N_25808,N_22513,N_22533);
nand U25809 (N_25809,N_22546,N_22816);
nand U25810 (N_25810,N_22127,N_22121);
nor U25811 (N_25811,N_23019,N_22874);
nand U25812 (N_25812,N_23281,N_22363);
or U25813 (N_25813,N_22977,N_23844);
nand U25814 (N_25814,N_23417,N_23323);
nand U25815 (N_25815,N_22844,N_23254);
and U25816 (N_25816,N_22678,N_23157);
nor U25817 (N_25817,N_22076,N_22816);
nor U25818 (N_25818,N_23179,N_23937);
nand U25819 (N_25819,N_22524,N_23287);
and U25820 (N_25820,N_23431,N_23744);
nor U25821 (N_25821,N_23107,N_23825);
or U25822 (N_25822,N_23545,N_23384);
nor U25823 (N_25823,N_22578,N_23846);
nor U25824 (N_25824,N_23466,N_23080);
nor U25825 (N_25825,N_22923,N_22645);
xnor U25826 (N_25826,N_23762,N_23562);
and U25827 (N_25827,N_22069,N_23198);
nor U25828 (N_25828,N_23699,N_23985);
and U25829 (N_25829,N_23308,N_22138);
nand U25830 (N_25830,N_22213,N_22804);
or U25831 (N_25831,N_22284,N_23501);
or U25832 (N_25832,N_23843,N_23998);
xnor U25833 (N_25833,N_23843,N_23159);
and U25834 (N_25834,N_22080,N_22186);
and U25835 (N_25835,N_23289,N_23827);
nor U25836 (N_25836,N_23001,N_23788);
nand U25837 (N_25837,N_22103,N_23751);
nand U25838 (N_25838,N_23626,N_23610);
and U25839 (N_25839,N_23523,N_22872);
or U25840 (N_25840,N_22682,N_23251);
or U25841 (N_25841,N_22509,N_22820);
nand U25842 (N_25842,N_22591,N_22651);
nand U25843 (N_25843,N_23379,N_23468);
nor U25844 (N_25844,N_22463,N_23328);
nand U25845 (N_25845,N_23064,N_22025);
nand U25846 (N_25846,N_22203,N_23510);
nand U25847 (N_25847,N_23141,N_23373);
nor U25848 (N_25848,N_23460,N_23607);
and U25849 (N_25849,N_22501,N_22474);
nor U25850 (N_25850,N_23665,N_23655);
nand U25851 (N_25851,N_22402,N_22884);
and U25852 (N_25852,N_22325,N_22633);
nor U25853 (N_25853,N_23754,N_23839);
nand U25854 (N_25854,N_23110,N_23387);
or U25855 (N_25855,N_22472,N_22492);
nor U25856 (N_25856,N_22601,N_23416);
or U25857 (N_25857,N_22343,N_23439);
nor U25858 (N_25858,N_23413,N_22507);
or U25859 (N_25859,N_22868,N_22813);
nor U25860 (N_25860,N_22565,N_22178);
nand U25861 (N_25861,N_22905,N_23261);
nand U25862 (N_25862,N_23553,N_22146);
nand U25863 (N_25863,N_22995,N_22069);
nand U25864 (N_25864,N_23155,N_22286);
and U25865 (N_25865,N_22695,N_22215);
or U25866 (N_25866,N_23000,N_22915);
nand U25867 (N_25867,N_22770,N_22211);
and U25868 (N_25868,N_22120,N_22354);
nand U25869 (N_25869,N_23697,N_23609);
nor U25870 (N_25870,N_22277,N_23102);
nand U25871 (N_25871,N_23099,N_22199);
and U25872 (N_25872,N_23747,N_23284);
nand U25873 (N_25873,N_23311,N_22113);
or U25874 (N_25874,N_22344,N_22732);
or U25875 (N_25875,N_22367,N_23728);
nand U25876 (N_25876,N_23452,N_22770);
nor U25877 (N_25877,N_23725,N_23094);
and U25878 (N_25878,N_22115,N_23266);
nand U25879 (N_25879,N_22200,N_23196);
nor U25880 (N_25880,N_23170,N_22806);
or U25881 (N_25881,N_23082,N_22236);
nor U25882 (N_25882,N_22315,N_22517);
xor U25883 (N_25883,N_23912,N_23289);
nand U25884 (N_25884,N_23339,N_22423);
nand U25885 (N_25885,N_23156,N_23113);
and U25886 (N_25886,N_22913,N_23001);
nand U25887 (N_25887,N_23150,N_23638);
and U25888 (N_25888,N_22853,N_22178);
or U25889 (N_25889,N_22987,N_23557);
or U25890 (N_25890,N_23436,N_22633);
nand U25891 (N_25891,N_23782,N_23520);
or U25892 (N_25892,N_22872,N_22913);
and U25893 (N_25893,N_23725,N_22425);
and U25894 (N_25894,N_23428,N_23016);
nand U25895 (N_25895,N_22546,N_23875);
or U25896 (N_25896,N_22959,N_22899);
and U25897 (N_25897,N_22261,N_23711);
and U25898 (N_25898,N_23448,N_23280);
nand U25899 (N_25899,N_22785,N_23368);
nor U25900 (N_25900,N_23838,N_23319);
nand U25901 (N_25901,N_23371,N_22402);
or U25902 (N_25902,N_22093,N_22389);
and U25903 (N_25903,N_22209,N_23931);
or U25904 (N_25904,N_22918,N_23956);
nand U25905 (N_25905,N_23796,N_23125);
or U25906 (N_25906,N_23443,N_22094);
or U25907 (N_25907,N_23973,N_23188);
nand U25908 (N_25908,N_23300,N_23802);
and U25909 (N_25909,N_23418,N_23981);
or U25910 (N_25910,N_23282,N_23959);
nand U25911 (N_25911,N_23086,N_22442);
or U25912 (N_25912,N_22933,N_22854);
nand U25913 (N_25913,N_22120,N_22985);
and U25914 (N_25914,N_23129,N_22116);
and U25915 (N_25915,N_22622,N_23517);
or U25916 (N_25916,N_23045,N_23584);
and U25917 (N_25917,N_22798,N_22652);
nor U25918 (N_25918,N_23710,N_22404);
nor U25919 (N_25919,N_23691,N_22232);
and U25920 (N_25920,N_23326,N_22682);
nor U25921 (N_25921,N_22269,N_23235);
nand U25922 (N_25922,N_23795,N_23183);
or U25923 (N_25923,N_23075,N_22568);
nor U25924 (N_25924,N_23091,N_22584);
nand U25925 (N_25925,N_23106,N_23956);
nand U25926 (N_25926,N_23007,N_22354);
nand U25927 (N_25927,N_22524,N_22126);
nand U25928 (N_25928,N_22969,N_22580);
nand U25929 (N_25929,N_22401,N_22104);
nor U25930 (N_25930,N_22947,N_22086);
nand U25931 (N_25931,N_22813,N_23095);
nand U25932 (N_25932,N_22925,N_22011);
or U25933 (N_25933,N_23263,N_23120);
nand U25934 (N_25934,N_22105,N_23151);
or U25935 (N_25935,N_22706,N_23985);
nand U25936 (N_25936,N_23336,N_22357);
nand U25937 (N_25937,N_23901,N_22215);
or U25938 (N_25938,N_23184,N_22566);
nor U25939 (N_25939,N_22829,N_23718);
nand U25940 (N_25940,N_23729,N_23559);
and U25941 (N_25941,N_23012,N_23551);
or U25942 (N_25942,N_22713,N_22694);
or U25943 (N_25943,N_23303,N_23922);
or U25944 (N_25944,N_23600,N_23058);
or U25945 (N_25945,N_23123,N_22300);
or U25946 (N_25946,N_22870,N_22618);
and U25947 (N_25947,N_23441,N_23445);
xnor U25948 (N_25948,N_22524,N_22208);
nor U25949 (N_25949,N_23918,N_23292);
or U25950 (N_25950,N_22473,N_23161);
and U25951 (N_25951,N_23048,N_23092);
nand U25952 (N_25952,N_23762,N_23026);
and U25953 (N_25953,N_23424,N_22801);
or U25954 (N_25954,N_23018,N_22895);
and U25955 (N_25955,N_23108,N_23580);
nand U25956 (N_25956,N_22566,N_22974);
nand U25957 (N_25957,N_22638,N_22484);
or U25958 (N_25958,N_23257,N_23236);
and U25959 (N_25959,N_22927,N_22157);
nor U25960 (N_25960,N_23207,N_22751);
or U25961 (N_25961,N_22774,N_22034);
nor U25962 (N_25962,N_23835,N_22627);
and U25963 (N_25963,N_23921,N_23670);
nand U25964 (N_25964,N_22448,N_23253);
nand U25965 (N_25965,N_22992,N_22378);
nand U25966 (N_25966,N_22688,N_22150);
nand U25967 (N_25967,N_22436,N_22729);
and U25968 (N_25968,N_22965,N_23057);
and U25969 (N_25969,N_22558,N_22545);
nand U25970 (N_25970,N_22758,N_22573);
and U25971 (N_25971,N_23367,N_22704);
or U25972 (N_25972,N_23006,N_23692);
nand U25973 (N_25973,N_22918,N_22023);
xor U25974 (N_25974,N_23234,N_22790);
or U25975 (N_25975,N_23050,N_22959);
nand U25976 (N_25976,N_22740,N_23391);
nand U25977 (N_25977,N_23305,N_22890);
nor U25978 (N_25978,N_22435,N_23467);
and U25979 (N_25979,N_23428,N_22544);
and U25980 (N_25980,N_23388,N_22295);
or U25981 (N_25981,N_23074,N_22902);
or U25982 (N_25982,N_23314,N_22273);
nand U25983 (N_25983,N_23321,N_22416);
nor U25984 (N_25984,N_23058,N_23342);
and U25985 (N_25985,N_22859,N_23777);
nor U25986 (N_25986,N_22359,N_22751);
and U25987 (N_25987,N_22234,N_23253);
or U25988 (N_25988,N_23547,N_22126);
nand U25989 (N_25989,N_22704,N_23402);
nor U25990 (N_25990,N_22715,N_23584);
or U25991 (N_25991,N_22421,N_23548);
nor U25992 (N_25992,N_22120,N_22121);
and U25993 (N_25993,N_23935,N_23405);
nor U25994 (N_25994,N_23146,N_22405);
nand U25995 (N_25995,N_23274,N_23294);
nor U25996 (N_25996,N_22994,N_22808);
nor U25997 (N_25997,N_23301,N_23728);
nor U25998 (N_25998,N_22666,N_22613);
and U25999 (N_25999,N_22782,N_22872);
or U26000 (N_26000,N_24267,N_25263);
or U26001 (N_26001,N_25148,N_24700);
and U26002 (N_26002,N_25428,N_24086);
xnor U26003 (N_26003,N_24957,N_24364);
nand U26004 (N_26004,N_24632,N_25438);
nand U26005 (N_26005,N_24475,N_24803);
nor U26006 (N_26006,N_24900,N_25118);
nand U26007 (N_26007,N_25312,N_24822);
nor U26008 (N_26008,N_24864,N_25711);
nor U26009 (N_26009,N_24600,N_25480);
nand U26010 (N_26010,N_25752,N_24356);
nor U26011 (N_26011,N_24482,N_25835);
nand U26012 (N_26012,N_24402,N_24946);
and U26013 (N_26013,N_24150,N_25491);
and U26014 (N_26014,N_24184,N_25522);
nor U26015 (N_26015,N_24341,N_25067);
or U26016 (N_26016,N_25115,N_24065);
nand U26017 (N_26017,N_25797,N_24607);
nand U26018 (N_26018,N_24220,N_24331);
or U26019 (N_26019,N_25584,N_24304);
and U26020 (N_26020,N_24838,N_24406);
and U26021 (N_26021,N_24137,N_25253);
xnor U26022 (N_26022,N_24549,N_24488);
or U26023 (N_26023,N_25744,N_25921);
nor U26024 (N_26024,N_24172,N_25570);
nor U26025 (N_26025,N_24811,N_25305);
and U26026 (N_26026,N_24767,N_25931);
or U26027 (N_26027,N_25052,N_25455);
nand U26028 (N_26028,N_24093,N_24698);
or U26029 (N_26029,N_24746,N_25060);
and U26030 (N_26030,N_24719,N_25502);
and U26031 (N_26031,N_25431,N_25743);
nand U26032 (N_26032,N_25473,N_25451);
or U26033 (N_26033,N_25225,N_25950);
nand U26034 (N_26034,N_24777,N_24997);
or U26035 (N_26035,N_25002,N_25365);
or U26036 (N_26036,N_24861,N_25568);
or U26037 (N_26037,N_24471,N_24669);
nand U26038 (N_26038,N_24850,N_25613);
nor U26039 (N_26039,N_25136,N_25849);
nor U26040 (N_26040,N_24706,N_25026);
nand U26041 (N_26041,N_24453,N_25224);
nand U26042 (N_26042,N_24535,N_24183);
nand U26043 (N_26043,N_24551,N_25071);
or U26044 (N_26044,N_25433,N_24055);
and U26045 (N_26045,N_25160,N_24490);
nor U26046 (N_26046,N_24116,N_24950);
and U26047 (N_26047,N_24755,N_24578);
nor U26048 (N_26048,N_24644,N_24849);
and U26049 (N_26049,N_25088,N_24895);
or U26050 (N_26050,N_24608,N_25563);
and U26051 (N_26051,N_24246,N_24084);
nand U26052 (N_26052,N_24605,N_24562);
nand U26053 (N_26053,N_25289,N_25191);
or U26054 (N_26054,N_25092,N_24648);
or U26055 (N_26055,N_24249,N_25620);
and U26056 (N_26056,N_25429,N_25412);
and U26057 (N_26057,N_24796,N_24325);
nor U26058 (N_26058,N_25842,N_25420);
and U26059 (N_26059,N_24790,N_25409);
and U26060 (N_26060,N_25538,N_25287);
and U26061 (N_26061,N_24915,N_25229);
and U26062 (N_26062,N_24374,N_24002);
nand U26063 (N_26063,N_24440,N_24911);
and U26064 (N_26064,N_25690,N_24517);
or U26065 (N_26065,N_25515,N_25549);
or U26066 (N_26066,N_25285,N_24884);
and U26067 (N_26067,N_24897,N_24598);
nor U26068 (N_26068,N_24939,N_24126);
or U26069 (N_26069,N_25128,N_24324);
nand U26070 (N_26070,N_24934,N_24525);
or U26071 (N_26071,N_25423,N_24556);
nand U26072 (N_26072,N_24932,N_24295);
nand U26073 (N_26073,N_24027,N_25017);
nor U26074 (N_26074,N_25664,N_25216);
or U26075 (N_26075,N_25182,N_25134);
nor U26076 (N_26076,N_25028,N_25111);
nor U26077 (N_26077,N_24981,N_24588);
and U26078 (N_26078,N_25361,N_24095);
nor U26079 (N_26079,N_24260,N_25393);
or U26080 (N_26080,N_24774,N_25934);
and U26081 (N_26081,N_24523,N_24500);
nor U26082 (N_26082,N_24107,N_25453);
nand U26083 (N_26083,N_25917,N_24354);
and U26084 (N_26084,N_24048,N_24925);
and U26085 (N_26085,N_25707,N_24253);
nor U26086 (N_26086,N_25773,N_25630);
nor U26087 (N_26087,N_25383,N_25639);
and U26088 (N_26088,N_24582,N_24539);
and U26089 (N_26089,N_24596,N_25345);
nor U26090 (N_26090,N_25476,N_25304);
nand U26091 (N_26091,N_25719,N_24296);
or U26092 (N_26092,N_24070,N_24377);
or U26093 (N_26093,N_24733,N_25790);
or U26094 (N_26094,N_24692,N_24689);
and U26095 (N_26095,N_24128,N_24294);
nor U26096 (N_26096,N_24204,N_25245);
or U26097 (N_26097,N_24052,N_24339);
and U26098 (N_26098,N_25514,N_24185);
nor U26099 (N_26099,N_24627,N_24846);
and U26100 (N_26100,N_25319,N_25546);
or U26101 (N_26101,N_25676,N_24119);
nor U26102 (N_26102,N_24064,N_25588);
or U26103 (N_26103,N_25085,N_24223);
nor U26104 (N_26104,N_24446,N_24457);
nor U26105 (N_26105,N_24099,N_25686);
or U26106 (N_26106,N_24762,N_25054);
and U26107 (N_26107,N_24806,N_25410);
and U26108 (N_26108,N_24795,N_25900);
and U26109 (N_26109,N_24949,N_25145);
nor U26110 (N_26110,N_25807,N_25997);
and U26111 (N_26111,N_24280,N_24964);
or U26112 (N_26112,N_25758,N_25074);
nand U26113 (N_26113,N_25699,N_24851);
and U26114 (N_26114,N_24984,N_25474);
or U26115 (N_26115,N_24786,N_24174);
nor U26116 (N_26116,N_25037,N_25448);
nand U26117 (N_26117,N_24695,N_25382);
or U26118 (N_26118,N_24541,N_25324);
and U26119 (N_26119,N_25467,N_24916);
or U26120 (N_26120,N_25941,N_25327);
nand U26121 (N_26121,N_24839,N_25915);
or U26122 (N_26122,N_25955,N_24388);
and U26123 (N_26123,N_25137,N_24216);
and U26124 (N_26124,N_25192,N_24342);
nand U26125 (N_26125,N_24952,N_24211);
or U26126 (N_26126,N_25219,N_25101);
and U26127 (N_26127,N_25535,N_24349);
nor U26128 (N_26128,N_25693,N_24222);
nor U26129 (N_26129,N_24251,N_25226);
and U26130 (N_26130,N_24885,N_25206);
or U26131 (N_26131,N_24177,N_24860);
and U26132 (N_26132,N_25601,N_24661);
nand U26133 (N_26133,N_24622,N_25618);
nor U26134 (N_26134,N_24594,N_25466);
and U26135 (N_26135,N_25079,N_24370);
or U26136 (N_26136,N_25746,N_25625);
or U26137 (N_26137,N_25090,N_24269);
or U26138 (N_26138,N_25600,N_24505);
and U26139 (N_26139,N_24455,N_25354);
nor U26140 (N_26140,N_24442,N_25576);
or U26141 (N_26141,N_25927,N_24135);
nand U26142 (N_26142,N_25281,N_25078);
nor U26143 (N_26143,N_24807,N_24266);
or U26144 (N_26144,N_25666,N_25048);
nor U26145 (N_26145,N_25008,N_24219);
or U26146 (N_26146,N_25785,N_25012);
or U26147 (N_26147,N_25933,N_25482);
or U26148 (N_26148,N_25946,N_25631);
nand U26149 (N_26149,N_24003,N_24108);
nand U26150 (N_26150,N_25942,N_25011);
nor U26151 (N_26151,N_24782,N_24164);
or U26152 (N_26152,N_24034,N_25161);
and U26153 (N_26153,N_24142,N_25164);
nand U26154 (N_26154,N_24748,N_24421);
nor U26155 (N_26155,N_24361,N_24470);
nand U26156 (N_26156,N_25893,N_25233);
xnor U26157 (N_26157,N_24158,N_25652);
nand U26158 (N_26158,N_24428,N_24479);
and U26159 (N_26159,N_25125,N_25523);
or U26160 (N_26160,N_24352,N_25745);
or U26161 (N_26161,N_24244,N_25099);
nand U26162 (N_26162,N_24300,N_24937);
nor U26163 (N_26163,N_25042,N_24672);
and U26164 (N_26164,N_25173,N_25958);
nor U26165 (N_26165,N_24392,N_24889);
or U26166 (N_26166,N_25057,N_25391);
and U26167 (N_26167,N_25341,N_25399);
and U26168 (N_26168,N_25885,N_25590);
nor U26169 (N_26169,N_25389,N_25551);
nor U26170 (N_26170,N_25778,N_25905);
nor U26171 (N_26171,N_25606,N_24924);
nand U26172 (N_26172,N_24071,N_25979);
or U26173 (N_26173,N_24350,N_25662);
or U26174 (N_26174,N_24840,N_25633);
nor U26175 (N_26175,N_24679,N_25976);
or U26176 (N_26176,N_25112,N_25829);
and U26177 (N_26177,N_25813,N_25781);
or U26178 (N_26178,N_25575,N_24716);
nor U26179 (N_26179,N_25873,N_24886);
nand U26180 (N_26180,N_25202,N_24521);
nand U26181 (N_26181,N_25834,N_24387);
or U26182 (N_26182,N_25831,N_24379);
nand U26183 (N_26183,N_25679,N_24610);
nand U26184 (N_26184,N_24954,N_25668);
nor U26185 (N_26185,N_24640,N_24496);
nand U26186 (N_26186,N_25572,N_25489);
nand U26187 (N_26187,N_25475,N_24138);
and U26188 (N_26188,N_24678,N_25266);
or U26189 (N_26189,N_24870,N_24499);
nor U26190 (N_26190,N_24394,N_25603);
nand U26191 (N_26191,N_25397,N_25531);
nand U26192 (N_26192,N_25725,N_25189);
or U26193 (N_26193,N_24075,N_24039);
nor U26194 (N_26194,N_25846,N_25106);
and U26195 (N_26195,N_25356,N_24080);
or U26196 (N_26196,N_24732,N_25918);
nand U26197 (N_26197,N_24918,N_25468);
nor U26198 (N_26198,N_24936,N_25646);
nor U26199 (N_26199,N_25322,N_25368);
and U26200 (N_26200,N_24302,N_25208);
or U26201 (N_26201,N_24209,N_24709);
and U26202 (N_26202,N_25770,N_24464);
nand U26203 (N_26203,N_25018,N_25053);
xor U26204 (N_26204,N_25246,N_24473);
and U26205 (N_26205,N_25083,N_25406);
and U26206 (N_26206,N_24017,N_24301);
or U26207 (N_26207,N_24106,N_25146);
nand U26208 (N_26208,N_25714,N_25442);
and U26209 (N_26209,N_25803,N_25424);
or U26210 (N_26210,N_25681,N_24764);
or U26211 (N_26211,N_24234,N_24530);
or U26212 (N_26212,N_24760,N_25395);
or U26213 (N_26213,N_25626,N_24667);
nand U26214 (N_26214,N_24708,N_24182);
nand U26215 (N_26215,N_24254,N_25187);
nor U26216 (N_26216,N_24942,N_24883);
or U26217 (N_26217,N_25267,N_24801);
nand U26218 (N_26218,N_24291,N_24315);
nor U26219 (N_26219,N_25881,N_24194);
and U26220 (N_26220,N_25513,N_25170);
or U26221 (N_26221,N_24843,N_25874);
xnor U26222 (N_26222,N_25236,N_25297);
nand U26223 (N_26223,N_25908,N_24237);
nor U26224 (N_26224,N_25116,N_25821);
nand U26225 (N_26225,N_24891,N_25670);
nand U26226 (N_26226,N_25038,N_24654);
nor U26227 (N_26227,N_24687,N_25392);
nand U26228 (N_26228,N_24639,N_24122);
and U26229 (N_26229,N_24112,N_24023);
or U26230 (N_26230,N_25867,N_24109);
nor U26231 (N_26231,N_25437,N_24805);
nand U26232 (N_26232,N_24789,N_24299);
or U26233 (N_26233,N_25086,N_24011);
or U26234 (N_26234,N_25162,N_24540);
and U26235 (N_26235,N_24662,N_24066);
nand U26236 (N_26236,N_25854,N_25027);
nor U26237 (N_26237,N_24550,N_25463);
nor U26238 (N_26238,N_25459,N_24180);
nor U26239 (N_26239,N_24726,N_25998);
or U26240 (N_26240,N_25511,N_24329);
and U26241 (N_26241,N_24413,N_25082);
nor U26242 (N_26242,N_24262,N_24877);
and U26243 (N_26243,N_24157,N_24928);
and U26244 (N_26244,N_24265,N_24365);
and U26245 (N_26245,N_24263,N_25194);
nand U26246 (N_26246,N_24247,N_24279);
or U26247 (N_26247,N_25274,N_24033);
and U26248 (N_26248,N_25869,N_25520);
nor U26249 (N_26249,N_25396,N_24512);
and U26250 (N_26250,N_24974,N_24469);
nor U26251 (N_26251,N_25861,N_25709);
nand U26252 (N_26252,N_25186,N_24548);
nand U26253 (N_26253,N_25866,N_25408);
nor U26254 (N_26254,N_25375,N_25848);
nor U26255 (N_26255,N_24345,N_25460);
nor U26256 (N_26256,N_24935,N_25619);
nand U26257 (N_26257,N_24176,N_25720);
or U26258 (N_26258,N_24120,N_25573);
nand U26259 (N_26259,N_24799,N_24491);
or U26260 (N_26260,N_24520,N_24553);
or U26261 (N_26261,N_24922,N_25107);
nand U26262 (N_26262,N_24771,N_24403);
and U26263 (N_26263,N_25031,N_25615);
nand U26264 (N_26264,N_25087,N_24962);
or U26265 (N_26265,N_25857,N_24831);
or U26266 (N_26266,N_25529,N_25553);
or U26267 (N_26267,N_25723,N_24865);
nand U26268 (N_26268,N_25418,N_24863);
or U26269 (N_26269,N_24409,N_24959);
and U26270 (N_26270,N_24401,N_25932);
and U26271 (N_26271,N_24624,N_24783);
and U26272 (N_26272,N_25215,N_25493);
and U26273 (N_26273,N_25847,N_25608);
nand U26274 (N_26274,N_25728,N_24163);
nand U26275 (N_26275,N_24923,N_25764);
or U26276 (N_26276,N_25385,N_24983);
or U26277 (N_26277,N_25342,N_25098);
or U26278 (N_26278,N_24871,N_24825);
nand U26279 (N_26279,N_25667,N_25248);
and U26280 (N_26280,N_24019,N_25642);
and U26281 (N_26281,N_24542,N_25738);
nor U26282 (N_26282,N_24178,N_25349);
nand U26283 (N_26283,N_25817,N_25005);
nand U26284 (N_26284,N_25228,N_24310);
and U26285 (N_26285,N_24444,N_25935);
xnor U26286 (N_26286,N_24134,N_24902);
or U26287 (N_26287,N_25954,N_24398);
or U26288 (N_26288,N_24054,N_25748);
nand U26289 (N_26289,N_25692,N_24483);
and U26290 (N_26290,N_24433,N_25120);
and U26291 (N_26291,N_25825,N_24381);
nand U26292 (N_26292,N_24083,N_25566);
and U26293 (N_26293,N_24368,N_24498);
and U26294 (N_26294,N_25255,N_25655);
and U26295 (N_26295,N_24230,N_25040);
nand U26296 (N_26296,N_24493,N_25860);
nand U26297 (N_26297,N_24511,N_25755);
nand U26298 (N_26298,N_25826,N_24256);
and U26299 (N_26299,N_24396,N_25961);
nor U26300 (N_26300,N_25496,N_25163);
nand U26301 (N_26301,N_24098,N_25717);
and U26302 (N_26302,N_25405,N_24705);
or U26303 (N_26303,N_24334,N_24371);
nor U26304 (N_26304,N_25323,N_25757);
nor U26305 (N_26305,N_24252,N_24887);
and U26306 (N_26306,N_25970,N_25114);
nand U26307 (N_26307,N_25540,N_25278);
nand U26308 (N_26308,N_25230,N_25996);
nor U26309 (N_26309,N_25461,N_25550);
and U26310 (N_26310,N_24665,N_25045);
nor U26311 (N_26311,N_25490,N_25318);
nand U26312 (N_26312,N_24975,N_25659);
nor U26313 (N_26313,N_25141,N_24492);
nand U26314 (N_26314,N_24196,N_25547);
or U26315 (N_26315,N_25730,N_25295);
xor U26316 (N_26316,N_24318,N_25528);
nand U26317 (N_26317,N_24615,N_25200);
or U26318 (N_26318,N_25441,N_24173);
or U26319 (N_26319,N_24264,N_24042);
or U26320 (N_26320,N_24830,N_24650);
or U26321 (N_26321,N_24287,N_24292);
and U26322 (N_26322,N_24327,N_25149);
nor U26323 (N_26323,N_25945,N_25198);
nor U26324 (N_26324,N_25280,N_24992);
nor U26325 (N_26325,N_25279,N_25221);
nor U26326 (N_26326,N_24441,N_25403);
or U26327 (N_26327,N_25579,N_25828);
nor U26328 (N_26328,N_25810,N_25795);
and U26329 (N_26329,N_25413,N_24058);
or U26330 (N_26330,N_25239,N_24638);
and U26331 (N_26331,N_25272,N_24125);
and U26332 (N_26332,N_25113,N_25640);
nor U26333 (N_26333,N_25390,N_24637);
and U26334 (N_26334,N_24044,N_25641);
or U26335 (N_26335,N_24103,N_24664);
nand U26336 (N_26336,N_24569,N_25812);
nand U26337 (N_26337,N_25928,N_24810);
nor U26338 (N_26338,N_24366,N_25916);
xor U26339 (N_26339,N_25559,N_25320);
and U26340 (N_26340,N_25268,N_25205);
and U26341 (N_26341,N_24544,N_24979);
nor U26342 (N_26342,N_25338,N_24241);
and U26343 (N_26343,N_24367,N_24725);
and U26344 (N_26344,N_25814,N_25981);
nor U26345 (N_26345,N_24791,N_25839);
nand U26346 (N_26346,N_25858,N_24652);
or U26347 (N_26347,N_25595,N_24372);
and U26348 (N_26348,N_25484,N_25702);
nand U26349 (N_26349,N_25241,N_24880);
and U26350 (N_26350,N_25789,N_25288);
and U26351 (N_26351,N_25154,N_24853);
or U26352 (N_26352,N_24127,N_25220);
nor U26353 (N_26353,N_25591,N_25358);
or U26354 (N_26354,N_24040,N_25721);
and U26355 (N_26355,N_25912,N_25033);
nor U26356 (N_26356,N_24606,N_24857);
and U26357 (N_26357,N_24697,N_24018);
nand U26358 (N_26358,N_24429,N_25792);
nand U26359 (N_26359,N_24035,N_25334);
nor U26360 (N_26360,N_24397,N_25706);
xnor U26361 (N_26361,N_25081,N_25276);
or U26362 (N_26362,N_25308,N_24319);
and U26363 (N_26363,N_24438,N_25974);
or U26364 (N_26364,N_24259,N_25147);
nand U26365 (N_26365,N_25436,N_25610);
and U26366 (N_26366,N_24224,N_24758);
and U26367 (N_26367,N_24326,N_24110);
or U26368 (N_26368,N_24205,N_25172);
nor U26369 (N_26369,N_24730,N_24020);
nand U26370 (N_26370,N_24270,N_25555);
or U26371 (N_26371,N_24522,N_25171);
or U26372 (N_26372,N_25047,N_25377);
nand U26373 (N_26373,N_25627,N_25021);
nor U26374 (N_26374,N_25232,N_24854);
and U26375 (N_26375,N_25350,N_25663);
or U26376 (N_26376,N_25936,N_24423);
or U26377 (N_26377,N_25283,N_25836);
nand U26378 (N_26378,N_24422,N_25920);
nor U26379 (N_26379,N_24570,N_24856);
and U26380 (N_26380,N_25895,N_24978);
nand U26381 (N_26381,N_25727,N_25526);
or U26382 (N_26382,N_24798,N_24675);
or U26383 (N_26383,N_25593,N_24621);
and U26384 (N_26384,N_25117,N_24242);
or U26385 (N_26385,N_24425,N_24408);
and U26386 (N_26386,N_24898,N_24920);
nand U26387 (N_26387,N_24633,N_25894);
nor U26388 (N_26388,N_24448,N_25574);
or U26389 (N_26389,N_25010,N_25614);
nor U26390 (N_26390,N_25635,N_24834);
or U26391 (N_26391,N_25450,N_25426);
and U26392 (N_26392,N_25337,N_25628);
nand U26393 (N_26393,N_25649,N_25330);
nand U26394 (N_26394,N_25910,N_25492);
or U26395 (N_26395,N_24199,N_24817);
xnor U26396 (N_26396,N_25750,N_25612);
or U26397 (N_26397,N_24674,N_24090);
nor U26398 (N_26398,N_24486,N_24769);
nand U26399 (N_26399,N_25359,N_24673);
and U26400 (N_26400,N_25995,N_24228);
or U26401 (N_26401,N_25167,N_25222);
or U26402 (N_26402,N_24351,N_25798);
nand U26403 (N_26403,N_24671,N_24841);
nor U26404 (N_26404,N_25937,N_25104);
or U26405 (N_26405,N_24495,N_24961);
or U26406 (N_26406,N_24595,N_25592);
and U26407 (N_26407,N_25035,N_25091);
and U26408 (N_26408,N_25806,N_25919);
and U26409 (N_26409,N_24461,N_25583);
or U26410 (N_26410,N_24411,N_24572);
nand U26411 (N_26411,N_24827,N_25193);
or U26412 (N_26412,N_24072,N_25065);
or U26413 (N_26413,N_25661,N_25794);
or U26414 (N_26414,N_24552,N_25335);
xor U26415 (N_26415,N_24714,N_25703);
nor U26416 (N_26416,N_24970,N_25367);
nand U26417 (N_26417,N_24658,N_25131);
nor U26418 (N_26418,N_25472,N_24794);
and U26419 (N_26419,N_25325,N_24958);
and U26420 (N_26420,N_25957,N_24063);
or U26421 (N_26421,N_25043,N_24344);
nand U26422 (N_26422,N_24316,N_25533);
or U26423 (N_26423,N_24298,N_25796);
nor U26424 (N_26424,N_25066,N_24038);
nand U26425 (N_26425,N_24907,N_25971);
and U26426 (N_26426,N_25800,N_25889);
nor U26427 (N_26427,N_24235,N_25548);
nor U26428 (N_26428,N_24768,N_25736);
or U26429 (N_26429,N_25159,N_25316);
and U26430 (N_26430,N_25291,N_25369);
and U26431 (N_26431,N_25203,N_25366);
nor U26432 (N_26432,N_24617,N_24663);
or U26433 (N_26433,N_24696,N_25199);
nor U26434 (N_26434,N_24908,N_25762);
nor U26435 (N_26435,N_24286,N_25594);
or U26436 (N_26436,N_25830,N_25975);
xor U26437 (N_26437,N_25710,N_24994);
and U26438 (N_26438,N_24956,N_24581);
nand U26439 (N_26439,N_25004,N_24557);
nor U26440 (N_26440,N_25604,N_25914);
nor U26441 (N_26441,N_24508,N_25622);
and U26442 (N_26442,N_24025,N_25597);
nor U26443 (N_26443,N_25373,N_24745);
nand U26444 (N_26444,N_25793,N_25599);
nand U26445 (N_26445,N_25959,N_24015);
nor U26446 (N_26446,N_24045,N_25657);
or U26447 (N_26447,N_25471,N_25771);
nor U26448 (N_26448,N_24162,N_25150);
and U26449 (N_26449,N_24221,N_24547);
and U26450 (N_26450,N_24929,N_25363);
nor U26451 (N_26451,N_24001,N_24583);
nor U26452 (N_26452,N_25168,N_25741);
or U26453 (N_26453,N_24792,N_25315);
nand U26454 (N_26454,N_24901,N_24655);
or U26455 (N_26455,N_24969,N_24601);
nor U26456 (N_26456,N_25680,N_24101);
nand U26457 (N_26457,N_25336,N_25249);
nand U26458 (N_26458,N_25015,N_25811);
or U26459 (N_26459,N_25580,N_24376);
and U26460 (N_26460,N_24195,N_24536);
and U26461 (N_26461,N_25063,N_24945);
and U26462 (N_26462,N_25486,N_25747);
or U26463 (N_26463,N_24463,N_25903);
and U26464 (N_26464,N_24380,N_24378);
nor U26465 (N_26465,N_24681,N_25275);
or U26466 (N_26466,N_25415,N_25080);
and U26467 (N_26467,N_24451,N_25013);
nor U26468 (N_26468,N_25469,N_25695);
nand U26469 (N_26469,N_24593,N_24619);
and U26470 (N_26470,N_24207,N_25704);
nand U26471 (N_26471,N_24272,N_24597);
nor U26472 (N_26472,N_25252,N_25705);
nand U26473 (N_26473,N_25510,N_25326);
nand U26474 (N_26474,N_24145,N_24362);
or U26475 (N_26475,N_25530,N_24718);
or U26476 (N_26476,N_25444,N_25636);
nor U26477 (N_26477,N_25123,N_24129);
and U26478 (N_26478,N_24684,N_24078);
xnor U26479 (N_26479,N_25296,N_25494);
and U26480 (N_26480,N_24587,N_25264);
nand U26481 (N_26481,N_25557,N_25132);
or U26482 (N_26482,N_25855,N_24743);
and U26483 (N_26483,N_24699,N_25605);
xor U26484 (N_26484,N_24159,N_24460);
and U26485 (N_26485,N_24032,N_24268);
nand U26486 (N_26486,N_24029,N_24141);
nor U26487 (N_26487,N_25019,N_24577);
nand U26488 (N_26488,N_24369,N_24821);
nand U26489 (N_26489,N_25506,N_24636);
nor U26490 (N_26490,N_24772,N_25020);
or U26491 (N_26491,N_24478,N_24609);
or U26492 (N_26492,N_25298,N_24067);
or U26493 (N_26493,N_24056,N_25545);
and U26494 (N_26494,N_25300,N_24462);
or U26495 (N_26495,N_24628,N_25644);
nand U26496 (N_26496,N_25891,N_25977);
nand U26497 (N_26497,N_25749,N_24503);
nand U26498 (N_26498,N_24004,N_24828);
or U26499 (N_26499,N_24757,N_25478);
nor U26500 (N_26500,N_25301,N_25598);
nor U26501 (N_26501,N_25840,N_24113);
nor U26502 (N_26502,N_25783,N_24416);
nand U26503 (N_26503,N_25788,N_25930);
nor U26504 (N_26504,N_24049,N_24154);
and U26505 (N_26505,N_24212,N_25508);
and U26506 (N_26506,N_25838,N_25949);
or U26507 (N_26507,N_24424,N_25537);
or U26508 (N_26508,N_25299,N_25944);
nor U26509 (N_26509,N_25371,N_25339);
nor U26510 (N_26510,N_25969,N_24393);
or U26511 (N_26511,N_24797,N_25009);
nor U26512 (N_26512,N_24166,N_24559);
or U26513 (N_26513,N_25833,N_24707);
and U26514 (N_26514,N_24649,N_25994);
and U26515 (N_26515,N_24563,N_24136);
nand U26516 (N_26516,N_24712,N_25217);
or U26517 (N_26517,N_25364,N_24206);
and U26518 (N_26518,N_25953,N_25753);
nor U26519 (N_26519,N_24686,N_25210);
nand U26520 (N_26520,N_24061,N_24407);
or U26521 (N_26521,N_24389,N_24643);
and U26522 (N_26522,N_25967,N_25003);
nor U26523 (N_26523,N_25561,N_24432);
nor U26524 (N_26524,N_25419,N_24819);
and U26525 (N_26525,N_25331,N_24021);
nor U26526 (N_26526,N_24215,N_24501);
or U26527 (N_26527,N_25660,N_25733);
nor U26528 (N_26528,N_25925,N_25972);
or U26529 (N_26529,N_25211,N_24656);
nor U26530 (N_26530,N_25902,N_24190);
nand U26531 (N_26531,N_25487,N_24285);
nor U26532 (N_26532,N_24904,N_24073);
nor U26533 (N_26533,N_25731,N_24631);
and U26534 (N_26534,N_25684,N_25344);
nand U26535 (N_26535,N_24927,N_24519);
and U26536 (N_26536,N_24087,N_24872);
nor U26537 (N_26537,N_24170,N_24965);
xnor U26538 (N_26538,N_25780,N_25070);
nor U26539 (N_26539,N_24188,N_24642);
and U26540 (N_26540,N_25564,N_24014);
nand U26541 (N_26541,N_24917,N_25871);
and U26542 (N_26542,N_24288,N_24437);
or U26543 (N_26543,N_25766,N_24878);
and U26544 (N_26544,N_24753,N_24169);
and U26545 (N_26545,N_25638,N_24740);
or U26546 (N_26546,N_25178,N_25956);
or U26547 (N_26547,N_24427,N_24802);
or U26548 (N_26548,N_25643,N_24243);
and U26549 (N_26549,N_25355,N_24585);
nor U26550 (N_26550,N_25870,N_25212);
or U26551 (N_26551,N_25039,N_24653);
or U26552 (N_26552,N_25329,N_24208);
and U26553 (N_26553,N_25270,N_24412);
nor U26554 (N_26554,N_24102,N_24990);
nor U26555 (N_26555,N_25380,N_24773);
nand U26556 (N_26556,N_24504,N_25376);
nor U26557 (N_26557,N_24852,N_24321);
nor U26558 (N_26558,N_24657,N_25244);
or U26559 (N_26559,N_24703,N_24348);
xnor U26560 (N_26560,N_24683,N_25439);
or U26561 (N_26561,N_25634,N_24590);
or U26562 (N_26562,N_24955,N_25983);
or U26563 (N_26563,N_25077,N_25623);
nor U26564 (N_26564,N_24395,N_25980);
and U26565 (N_26565,N_25585,N_25386);
nand U26566 (N_26566,N_25025,N_25582);
or U26567 (N_26567,N_24893,N_24193);
and U26568 (N_26568,N_24328,N_24813);
and U26569 (N_26569,N_24290,N_24599);
and U26570 (N_26570,N_24431,N_24513);
or U26571 (N_26571,N_24982,N_25853);
and U26572 (N_26572,N_24963,N_24820);
and U26573 (N_26573,N_25716,N_24502);
and U26574 (N_26574,N_25140,N_24565);
nor U26575 (N_26575,N_25127,N_24144);
or U26576 (N_26576,N_25844,N_24837);
nor U26577 (N_26577,N_24737,N_25948);
xor U26578 (N_26578,N_25779,N_24452);
and U26579 (N_26579,N_25293,N_25400);
nand U26580 (N_26580,N_25898,N_24940);
nand U26581 (N_26581,N_25751,N_24013);
xor U26582 (N_26582,N_24905,N_24761);
and U26583 (N_26583,N_25665,N_25387);
or U26584 (N_26584,N_24487,N_25481);
and U26585 (N_26585,N_25094,N_25156);
and U26586 (N_26586,N_24289,N_25051);
and U26587 (N_26587,N_24335,N_25209);
or U26588 (N_26588,N_24766,N_24531);
or U26589 (N_26589,N_25978,N_24823);
nor U26590 (N_26590,N_25122,N_25824);
nand U26591 (N_26591,N_25787,N_25675);
and U26592 (N_26592,N_24414,N_24614);
nor U26593 (N_26593,N_24780,N_24735);
nand U26594 (N_26594,N_25103,N_25006);
or U26595 (N_26595,N_25888,N_25678);
nor U26596 (N_26596,N_24226,N_24386);
nor U26597 (N_26597,N_24729,N_25029);
nand U26598 (N_26598,N_25863,N_25872);
nor U26599 (N_26599,N_24514,N_24694);
nor U26600 (N_26600,N_25064,N_25632);
and U26601 (N_26601,N_24434,N_24168);
nand U26602 (N_26602,N_24008,N_25843);
and U26603 (N_26603,N_25454,N_24353);
and U26604 (N_26604,N_24332,N_25257);
nor U26605 (N_26605,N_24738,N_25718);
nor U26606 (N_26606,N_24873,N_25181);
and U26607 (N_26607,N_25000,N_25560);
nand U26608 (N_26608,N_25204,N_24467);
or U26609 (N_26609,N_24938,N_25761);
and U26610 (N_26610,N_24973,N_25589);
nand U26611 (N_26611,N_24972,N_25569);
nand U26612 (N_26612,N_25062,N_24472);
nor U26613 (N_26613,N_24527,N_24130);
nor U26614 (N_26614,N_24384,N_24515);
nor U26615 (N_26615,N_25554,N_24360);
xor U26616 (N_26616,N_24921,N_25808);
nor U26617 (N_26617,N_24892,N_24776);
nor U26618 (N_26618,N_25503,N_24888);
nor U26619 (N_26619,N_25577,N_25799);
or U26620 (N_26620,N_25034,N_24560);
nand U26621 (N_26621,N_25041,N_24507);
and U26622 (N_26622,N_24816,N_24274);
and U26623 (N_26623,N_25075,N_24271);
nor U26624 (N_26624,N_24814,N_25713);
nand U26625 (N_26625,N_25427,N_24155);
or U26626 (N_26626,N_24187,N_25587);
and U26627 (N_26627,N_25907,N_24443);
nand U26628 (N_26628,N_25314,N_25990);
and U26629 (N_26629,N_24225,N_25879);
and U26630 (N_26630,N_24069,N_25651);
nor U26631 (N_26631,N_24031,N_25518);
or U26632 (N_26632,N_24815,N_24089);
and U26633 (N_26633,N_25841,N_24736);
nor U26634 (N_26634,N_24485,N_24143);
or U26635 (N_26635,N_25694,N_25247);
nor U26636 (N_26636,N_25477,N_24148);
or U26637 (N_26637,N_25672,N_24214);
nand U26638 (N_26638,N_24347,N_24132);
and U26639 (N_26639,N_25562,N_25742);
nor U26640 (N_26640,N_25890,N_25801);
nand U26641 (N_26641,N_25404,N_25394);
nor U26642 (N_26642,N_24081,N_24724);
and U26643 (N_26643,N_25152,N_25231);
or U26644 (N_26644,N_24731,N_25068);
or U26645 (N_26645,N_25966,N_25852);
nand U26646 (N_26646,N_25196,N_24778);
nand U26647 (N_26647,N_25133,N_25819);
or U26648 (N_26648,N_25521,N_25987);
and U26649 (N_26649,N_24297,N_24385);
nand U26650 (N_26650,N_25754,N_25507);
and U26651 (N_26651,N_25722,N_24613);
nor U26652 (N_26652,N_24047,N_25786);
or U26653 (N_26653,N_24589,N_24765);
nor U26654 (N_26654,N_24357,N_25001);
nand U26655 (N_26655,N_24338,N_24210);
or U26656 (N_26656,N_24314,N_24236);
nand U26657 (N_26657,N_25856,N_25165);
xnor U26658 (N_26658,N_25698,N_25940);
and U26659 (N_26659,N_25685,N_25056);
xor U26660 (N_26660,N_24046,N_25772);
nor U26661 (N_26661,N_24275,N_25536);
xnor U26662 (N_26662,N_25271,N_25126);
nand U26663 (N_26663,N_25804,N_25023);
and U26664 (N_26664,N_24477,N_24848);
or U26665 (N_26665,N_24481,N_25964);
nand U26666 (N_26666,N_25177,N_24879);
and U26667 (N_26667,N_25256,N_24899);
nor U26668 (N_26668,N_24092,N_25687);
nand U26669 (N_26669,N_25179,N_25097);
and U26670 (N_26670,N_24131,N_24826);
nor U26671 (N_26671,N_24435,N_24784);
nor U26672 (N_26672,N_24323,N_25157);
or U26673 (N_26673,N_25791,N_24281);
nand U26674 (N_26674,N_25965,N_25362);
nand U26675 (N_26675,N_25541,N_25732);
nand U26676 (N_26676,N_24240,N_24405);
nor U26677 (N_26677,N_25456,N_25174);
or U26678 (N_26678,N_25261,N_25677);
or U26679 (N_26679,N_25862,N_25581);
and U26680 (N_26680,N_25818,N_24739);
nor U26681 (N_26681,N_24231,N_25290);
or U26682 (N_26682,N_24160,N_25782);
nand U26683 (N_26683,N_25311,N_25739);
or U26684 (N_26684,N_24233,N_24273);
nand U26685 (N_26685,N_24742,N_25175);
xnor U26686 (N_26686,N_24124,N_24690);
nand U26687 (N_26687,N_24363,N_25552);
nand U26688 (N_26688,N_25195,N_25169);
or U26689 (N_26689,N_24869,N_25734);
and U26690 (N_26690,N_25139,N_25809);
or U26691 (N_26691,N_25602,N_25135);
nor U26692 (N_26692,N_24320,N_25184);
nor U26693 (N_26693,N_24824,N_24149);
nor U26694 (N_26694,N_25876,N_24293);
nand U26695 (N_26695,N_24584,N_25735);
and U26696 (N_26696,N_24800,N_24691);
or U26697 (N_26697,N_24635,N_25445);
or U26698 (N_26698,N_24303,N_25378);
nand U26699 (N_26699,N_24082,N_24604);
nor U26700 (N_26700,N_25273,N_25310);
and U26701 (N_26701,N_25968,N_25282);
nor U26702 (N_26702,N_24079,N_25343);
or U26703 (N_26703,N_24867,N_25485);
or U26704 (N_26704,N_25414,N_24641);
or U26705 (N_26705,N_24568,N_24571);
nand U26706 (N_26706,N_25024,N_24007);
and U26707 (N_26707,N_25105,N_24909);
or U26708 (N_26708,N_24931,N_25823);
and U26709 (N_26709,N_24400,N_24171);
nand U26710 (N_26710,N_25254,N_24977);
and U26711 (N_26711,N_25654,N_24333);
or U26712 (N_26712,N_25973,N_25102);
nand U26713 (N_26713,N_24763,N_25213);
and U26714 (N_26714,N_24629,N_24991);
or U26715 (N_26715,N_25235,N_24459);
nand U26716 (N_26716,N_24028,N_25708);
nand U26717 (N_26717,N_24516,N_24759);
or U26718 (N_26718,N_25578,N_24744);
or U26719 (N_26719,N_25321,N_24181);
nor U26720 (N_26720,N_24494,N_25682);
and U26721 (N_26721,N_24489,N_24133);
or U26722 (N_26722,N_25653,N_24191);
nor U26723 (N_26723,N_25227,N_25218);
nand U26724 (N_26724,N_25611,N_25960);
or U26725 (N_26725,N_24449,N_24161);
xor U26726 (N_26726,N_24261,N_24012);
and U26727 (N_26727,N_24770,N_25190);
or U26728 (N_26728,N_24532,N_25234);
nor U26729 (N_26729,N_25845,N_24375);
nand U26730 (N_26730,N_24312,N_24043);
nor U26731 (N_26731,N_24537,N_24202);
or U26732 (N_26732,N_25076,N_25887);
and U26733 (N_26733,N_24151,N_25938);
nor U26734 (N_26734,N_24041,N_25904);
or U26735 (N_26735,N_25756,N_24906);
or U26736 (N_26736,N_25558,N_25658);
nor U26737 (N_26737,N_24713,N_24580);
nand U26738 (N_26738,N_24715,N_25498);
or U26739 (N_26739,N_24651,N_25089);
xnor U26740 (N_26740,N_25360,N_25250);
nor U26741 (N_26741,N_24833,N_24309);
and U26742 (N_26742,N_25989,N_25014);
and U26743 (N_26743,N_24117,N_25144);
nor U26744 (N_26744,N_25328,N_24074);
and U26745 (N_26745,N_24524,N_24701);
nand U26746 (N_26746,N_24200,N_24747);
nor U26747 (N_26747,N_24835,N_25166);
or U26748 (N_26748,N_24844,N_25882);
or U26749 (N_26749,N_24022,N_24111);
nand U26750 (N_26750,N_24430,N_25084);
or U26751 (N_26751,N_25805,N_25422);
nand U26752 (N_26752,N_24567,N_25073);
and U26753 (N_26753,N_25689,N_25542);
and U26754 (N_26754,N_25899,N_25951);
nand U26755 (N_26755,N_25121,N_24307);
nand U26756 (N_26756,N_24659,N_24526);
or U26757 (N_26757,N_24623,N_24051);
and U26758 (N_26758,N_24953,N_24646);
xor U26759 (N_26759,N_25242,N_25539);
or U26760 (N_26760,N_25534,N_24036);
and U26761 (N_26761,N_24988,N_24257);
nor U26762 (N_26762,N_25130,N_25351);
and U26763 (N_26763,N_25332,N_25629);
nor U26764 (N_26764,N_25340,N_24573);
nor U26765 (N_26765,N_25401,N_24611);
nand U26766 (N_26766,N_24711,N_24620);
or U26767 (N_26767,N_25243,N_24804);
nand U26768 (N_26768,N_24484,N_25384);
and U26769 (N_26769,N_24088,N_25851);
nor U26770 (N_26770,N_24999,N_24575);
or U26771 (N_26771,N_24630,N_24809);
or U26772 (N_26772,N_25865,N_24175);
or U26773 (N_26773,N_24890,N_24751);
or U26774 (N_26774,N_25100,N_25504);
nand U26775 (N_26775,N_25470,N_25095);
and U26776 (N_26776,N_24618,N_25886);
and U26777 (N_26777,N_25884,N_25372);
nand U26778 (N_26778,N_24091,N_24121);
and U26779 (N_26779,N_24450,N_25647);
or U26780 (N_26780,N_25381,N_25883);
nand U26781 (N_26781,N_25875,N_24152);
nor U26782 (N_26782,N_25617,N_24793);
and U26783 (N_26783,N_24186,N_25407);
nor U26784 (N_26784,N_24313,N_24734);
or U26785 (N_26785,N_25609,N_25425);
nor U26786 (N_26786,N_24203,N_25302);
nand U26787 (N_26787,N_24787,N_24009);
nor U26788 (N_26788,N_24016,N_24968);
and U26789 (N_26789,N_25430,N_24704);
and U26790 (N_26790,N_25452,N_24139);
nor U26791 (N_26791,N_25223,N_24987);
nor U26792 (N_26792,N_24602,N_25607);
nor U26793 (N_26793,N_25512,N_24317);
and U26794 (N_26794,N_24359,N_25645);
nor U26795 (N_26795,N_25108,N_25180);
nand U26796 (N_26796,N_24104,N_24995);
nor U26797 (N_26797,N_24914,N_24382);
or U26798 (N_26798,N_25265,N_25993);
or U26799 (N_26799,N_24976,N_25309);
and U26800 (N_26800,N_24114,N_24085);
nor U26801 (N_26801,N_24229,N_25656);
nor U26802 (N_26802,N_25878,N_25479);
nand U26803 (N_26803,N_24779,N_25258);
nand U26804 (N_26804,N_25827,N_24439);
nor U26805 (N_26805,N_24832,N_25050);
and U26806 (N_26806,N_25388,N_25061);
nand U26807 (N_26807,N_25251,N_25988);
nor U26808 (N_26808,N_25911,N_25347);
or U26809 (N_26809,N_24688,N_25434);
nand U26810 (N_26810,N_24418,N_24876);
or U26811 (N_26811,N_25525,N_25715);
nor U26812 (N_26812,N_24967,N_24741);
or U26813 (N_26813,N_24258,N_24913);
xor U26814 (N_26814,N_25864,N_25571);
and U26815 (N_26815,N_25499,N_24410);
or U26816 (N_26816,N_25096,N_24933);
or U26817 (N_26817,N_25464,N_25352);
xor U26818 (N_26818,N_25457,N_25674);
nand U26819 (N_26819,N_25992,N_25701);
and U26820 (N_26820,N_25348,N_25501);
nor U26821 (N_26821,N_24722,N_25505);
nor U26822 (N_26822,N_25913,N_24818);
nor U26823 (N_26823,N_24179,N_25650);
or U26824 (N_26824,N_25982,N_25765);
and U26825 (N_26825,N_25802,N_24576);
and U26826 (N_26826,N_24717,N_24277);
and U26827 (N_26827,N_24346,N_24616);
and U26828 (N_26828,N_25777,N_25465);
xor U26829 (N_26829,N_24591,N_24447);
and U26830 (N_26830,N_24574,N_24670);
nand U26831 (N_26831,N_25984,N_24097);
nand U26832 (N_26832,N_24426,N_24866);
nand U26833 (N_26833,N_24480,N_24053);
nand U26834 (N_26834,N_24586,N_24068);
nand U26835 (N_26835,N_24284,N_25671);
or U26836 (N_26836,N_24903,N_25763);
nor U26837 (N_26837,N_25432,N_25353);
and U26838 (N_26838,N_25402,N_25260);
and U26839 (N_26839,N_24197,N_24217);
nor U26840 (N_26840,N_24785,N_25292);
and U26841 (N_26841,N_24189,N_24720);
nor U26842 (N_26842,N_25556,N_24096);
nand U26843 (N_26843,N_25909,N_24875);
nand U26844 (N_26844,N_24812,N_24926);
nor U26845 (N_26845,N_25421,N_24118);
nand U26846 (N_26846,N_24238,N_25016);
nand U26847 (N_26847,N_24026,N_25142);
and U26848 (N_26848,N_24476,N_25207);
nand U26849 (N_26849,N_24458,N_25307);
nand U26850 (N_26850,N_25901,N_24881);
and U26851 (N_26851,N_25370,N_25696);
and U26852 (N_26852,N_25449,N_25616);
and U26853 (N_26853,N_24558,N_25740);
nand U26854 (N_26854,N_25188,N_24561);
nand U26855 (N_26855,N_24842,N_24006);
or U26856 (N_26856,N_25411,N_25527);
nor U26857 (N_26857,N_25416,N_24951);
and U26858 (N_26858,N_24192,N_25868);
or U26859 (N_26859,N_24966,N_25567);
and U26860 (N_26860,N_25509,N_24944);
nand U26861 (N_26861,N_25952,N_24728);
nand U26862 (N_26862,N_24030,N_24894);
or U26863 (N_26863,N_25176,N_25532);
nor U26864 (N_26864,N_25458,N_25357);
or U26865 (N_26865,N_24634,N_25822);
and U26866 (N_26866,N_24466,N_24727);
nand U26867 (N_26867,N_24948,N_24960);
nor U26868 (N_26868,N_25022,N_24752);
and U26869 (N_26869,N_25688,N_24625);
or U26870 (N_26870,N_24123,N_24248);
nand U26871 (N_26871,N_24989,N_25417);
and U26872 (N_26872,N_25691,N_24543);
or U26873 (N_26873,N_24980,N_24533);
nand U26874 (N_26874,N_24445,N_24140);
nor U26875 (N_26875,N_24213,N_25832);
or U26876 (N_26876,N_24399,N_25447);
and U26877 (N_26877,N_25032,N_24693);
and U26878 (N_26878,N_24276,N_25109);
nand U26879 (N_26879,N_25269,N_24912);
nor U26880 (N_26880,N_24358,N_24554);
nor U26881 (N_26881,N_25197,N_24781);
and U26882 (N_26882,N_24474,N_25007);
or U26883 (N_26883,N_24874,N_24626);
nor U26884 (N_26884,N_24510,N_24721);
and U26885 (N_26885,N_25947,N_25201);
nor U26886 (N_26886,N_24862,N_24417);
nand U26887 (N_26887,N_25435,N_25596);
nor U26888 (N_26888,N_24910,N_25906);
or U26889 (N_26889,N_25238,N_25153);
or U26890 (N_26890,N_24373,N_24998);
or U26891 (N_26891,N_24153,N_25859);
or U26892 (N_26892,N_24676,N_24509);
or U26893 (N_26893,N_25240,N_24941);
or U26894 (N_26894,N_24383,N_24919);
nand U26895 (N_26895,N_24355,N_24282);
or U26896 (N_26896,N_25759,N_25143);
nand U26897 (N_26897,N_24239,N_25030);
and U26898 (N_26898,N_25524,N_24858);
nand U26899 (N_26899,N_25673,N_24037);
and U26900 (N_26900,N_25440,N_25317);
nand U26901 (N_26901,N_24059,N_25046);
and U26902 (N_26902,N_25488,N_24677);
and U26903 (N_26903,N_24702,N_25072);
nor U26904 (N_26904,N_24454,N_24545);
or U26905 (N_26905,N_25669,N_24278);
and U26906 (N_26906,N_25737,N_24647);
nor U26907 (N_26907,N_25443,N_24415);
or U26908 (N_26908,N_25624,N_25543);
and U26909 (N_26909,N_25922,N_24337);
nor U26910 (N_26910,N_24436,N_24456);
xor U26911 (N_26911,N_24986,N_24077);
or U26912 (N_26912,N_25943,N_25820);
or U26913 (N_26913,N_24847,N_25259);
or U26914 (N_26914,N_25036,N_24754);
or U26915 (N_26915,N_25119,N_24788);
or U26916 (N_26916,N_24710,N_25495);
nand U26917 (N_26917,N_24882,N_25516);
nor U26918 (N_26918,N_24756,N_24836);
or U26919 (N_26919,N_25313,N_25058);
and U26920 (N_26920,N_24050,N_24468);
and U26921 (N_26921,N_24005,N_24245);
and U26922 (N_26922,N_25850,N_24147);
nand U26923 (N_26923,N_24668,N_24146);
nor U26924 (N_26924,N_24564,N_24775);
or U26925 (N_26925,N_25929,N_24518);
nor U26926 (N_26926,N_24000,N_24947);
nor U26927 (N_26927,N_24167,N_24896);
and U26928 (N_26928,N_25586,N_24930);
nand U26929 (N_26929,N_25333,N_24060);
and U26930 (N_26930,N_24723,N_25939);
nor U26931 (N_26931,N_25500,N_24218);
nand U26932 (N_26932,N_24308,N_25262);
nor U26933 (N_26933,N_25483,N_24201);
and U26934 (N_26934,N_25237,N_25214);
and U26935 (N_26935,N_25519,N_25185);
or U26936 (N_26936,N_24115,N_24845);
nand U26937 (N_26937,N_24024,N_25158);
and U26938 (N_26938,N_25991,N_25724);
nand U26939 (N_26939,N_24680,N_25962);
or U26940 (N_26940,N_25286,N_24343);
nor U26941 (N_26941,N_24855,N_25379);
nor U26942 (N_26942,N_24340,N_24010);
and U26943 (N_26943,N_25462,N_25999);
nor U26944 (N_26944,N_25880,N_24749);
or U26945 (N_26945,N_24566,N_24255);
nand U26946 (N_26946,N_24497,N_25985);
and U26947 (N_26947,N_25697,N_25896);
nor U26948 (N_26948,N_24311,N_25769);
nand U26949 (N_26949,N_25155,N_25446);
or U26950 (N_26950,N_25776,N_25049);
nor U26951 (N_26951,N_25837,N_25284);
nand U26952 (N_26952,N_25760,N_25124);
and U26953 (N_26953,N_25151,N_24985);
nand U26954 (N_26954,N_24305,N_25767);
nor U26955 (N_26955,N_24971,N_25774);
nor U26956 (N_26956,N_24062,N_24996);
nand U26957 (N_26957,N_25055,N_25712);
or U26958 (N_26958,N_25700,N_25897);
nand U26959 (N_26959,N_24750,N_24612);
nor U26960 (N_26960,N_25784,N_25374);
xor U26961 (N_26961,N_25129,N_24660);
nand U26962 (N_26962,N_25621,N_24404);
nand U26963 (N_26963,N_24391,N_25346);
nor U26964 (N_26964,N_25775,N_24868);
or U26965 (N_26965,N_24156,N_25892);
and U26966 (N_26966,N_24100,N_24603);
and U26967 (N_26967,N_24682,N_24592);
nand U26968 (N_26968,N_24390,N_24057);
and U26969 (N_26969,N_24993,N_24232);
and U26970 (N_26970,N_25069,N_24685);
or U26971 (N_26971,N_24829,N_25044);
and U26972 (N_26972,N_25544,N_25926);
and U26973 (N_26973,N_24105,N_24283);
or U26974 (N_26974,N_24420,N_25138);
nor U26975 (N_26975,N_25565,N_24227);
nor U26976 (N_26976,N_25768,N_24094);
nand U26977 (N_26977,N_25986,N_24076);
nand U26978 (N_26978,N_24943,N_25924);
nor U26979 (N_26979,N_24579,N_25294);
nor U26980 (N_26980,N_25110,N_24546);
and U26981 (N_26981,N_25183,N_25517);
nand U26982 (N_26982,N_24198,N_24859);
and U26983 (N_26983,N_24538,N_24645);
or U26984 (N_26984,N_25816,N_25648);
nor U26985 (N_26985,N_24534,N_24528);
nor U26986 (N_26986,N_25497,N_24419);
nand U26987 (N_26987,N_25637,N_24666);
and U26988 (N_26988,N_24322,N_24506);
and U26989 (N_26989,N_25059,N_25963);
and U26990 (N_26990,N_24306,N_24165);
and U26991 (N_26991,N_24555,N_24336);
xor U26992 (N_26992,N_25726,N_25729);
or U26993 (N_26993,N_24529,N_25815);
nand U26994 (N_26994,N_24250,N_25306);
nand U26995 (N_26995,N_25923,N_25398);
nand U26996 (N_26996,N_25277,N_25683);
or U26997 (N_26997,N_24330,N_24808);
nor U26998 (N_26998,N_25303,N_25877);
nand U26999 (N_26999,N_25093,N_24465);
and U27000 (N_27000,N_25887,N_24281);
nand U27001 (N_27001,N_24403,N_24232);
or U27002 (N_27002,N_25291,N_24836);
nand U27003 (N_27003,N_25838,N_24029);
nand U27004 (N_27004,N_24688,N_24497);
or U27005 (N_27005,N_25953,N_24143);
or U27006 (N_27006,N_25374,N_24994);
nor U27007 (N_27007,N_25703,N_25401);
nand U27008 (N_27008,N_24718,N_24997);
or U27009 (N_27009,N_25793,N_24684);
xnor U27010 (N_27010,N_25630,N_24158);
nor U27011 (N_27011,N_25028,N_25139);
or U27012 (N_27012,N_25579,N_25344);
nand U27013 (N_27013,N_24669,N_25267);
nand U27014 (N_27014,N_24208,N_25247);
and U27015 (N_27015,N_25288,N_25498);
or U27016 (N_27016,N_24019,N_25778);
nor U27017 (N_27017,N_24727,N_24215);
nor U27018 (N_27018,N_25198,N_24636);
or U27019 (N_27019,N_25330,N_25553);
nor U27020 (N_27020,N_25209,N_24719);
nand U27021 (N_27021,N_25706,N_24477);
or U27022 (N_27022,N_25972,N_25109);
nor U27023 (N_27023,N_24451,N_25344);
or U27024 (N_27024,N_25879,N_25593);
and U27025 (N_27025,N_24645,N_25635);
nor U27026 (N_27026,N_24950,N_24616);
or U27027 (N_27027,N_24562,N_24877);
and U27028 (N_27028,N_25320,N_25105);
nand U27029 (N_27029,N_25079,N_24252);
and U27030 (N_27030,N_24326,N_25842);
or U27031 (N_27031,N_24130,N_25764);
nand U27032 (N_27032,N_25477,N_24300);
or U27033 (N_27033,N_25445,N_24942);
nor U27034 (N_27034,N_25938,N_25164);
or U27035 (N_27035,N_25447,N_25806);
nor U27036 (N_27036,N_25411,N_24126);
nor U27037 (N_27037,N_25781,N_25761);
and U27038 (N_27038,N_24941,N_24358);
nand U27039 (N_27039,N_25606,N_25464);
and U27040 (N_27040,N_25958,N_24505);
nand U27041 (N_27041,N_25724,N_25967);
or U27042 (N_27042,N_25369,N_24190);
nor U27043 (N_27043,N_24523,N_25217);
and U27044 (N_27044,N_24193,N_24536);
or U27045 (N_27045,N_25025,N_25785);
and U27046 (N_27046,N_25166,N_25060);
and U27047 (N_27047,N_24420,N_24656);
nor U27048 (N_27048,N_25631,N_24371);
and U27049 (N_27049,N_24937,N_24516);
nor U27050 (N_27050,N_25190,N_25598);
nand U27051 (N_27051,N_25976,N_24887);
nor U27052 (N_27052,N_25644,N_24140);
or U27053 (N_27053,N_24120,N_24745);
nor U27054 (N_27054,N_24407,N_24516);
nand U27055 (N_27055,N_25750,N_24480);
nand U27056 (N_27056,N_24335,N_24526);
or U27057 (N_27057,N_25627,N_25989);
nand U27058 (N_27058,N_24280,N_24397);
and U27059 (N_27059,N_24114,N_24000);
nand U27060 (N_27060,N_24966,N_25027);
and U27061 (N_27061,N_24407,N_25185);
nand U27062 (N_27062,N_24061,N_24330);
and U27063 (N_27063,N_25592,N_25376);
or U27064 (N_27064,N_25960,N_24028);
nor U27065 (N_27065,N_25124,N_25741);
nor U27066 (N_27066,N_25355,N_24521);
nand U27067 (N_27067,N_25007,N_25744);
and U27068 (N_27068,N_24493,N_25924);
and U27069 (N_27069,N_24525,N_25695);
nand U27070 (N_27070,N_25672,N_25894);
xnor U27071 (N_27071,N_25291,N_24700);
or U27072 (N_27072,N_24411,N_25040);
or U27073 (N_27073,N_25280,N_25046);
or U27074 (N_27074,N_25362,N_25644);
and U27075 (N_27075,N_24359,N_25545);
or U27076 (N_27076,N_25838,N_24950);
or U27077 (N_27077,N_24686,N_25203);
or U27078 (N_27078,N_25524,N_24918);
and U27079 (N_27079,N_24265,N_25825);
or U27080 (N_27080,N_24823,N_25414);
nor U27081 (N_27081,N_24099,N_25622);
nor U27082 (N_27082,N_24810,N_24729);
and U27083 (N_27083,N_25430,N_24995);
nor U27084 (N_27084,N_25308,N_25792);
nand U27085 (N_27085,N_25692,N_24220);
xnor U27086 (N_27086,N_25810,N_24892);
nor U27087 (N_27087,N_24179,N_24941);
nor U27088 (N_27088,N_25948,N_24043);
nand U27089 (N_27089,N_25690,N_24372);
or U27090 (N_27090,N_25701,N_24133);
nor U27091 (N_27091,N_24499,N_25540);
nand U27092 (N_27092,N_25797,N_25811);
nand U27093 (N_27093,N_25591,N_25893);
nor U27094 (N_27094,N_24239,N_24192);
or U27095 (N_27095,N_24337,N_25447);
and U27096 (N_27096,N_25121,N_24951);
nor U27097 (N_27097,N_25512,N_25375);
nand U27098 (N_27098,N_24772,N_24059);
nand U27099 (N_27099,N_25586,N_24862);
or U27100 (N_27100,N_25737,N_24633);
nor U27101 (N_27101,N_25125,N_24004);
or U27102 (N_27102,N_24750,N_25927);
nor U27103 (N_27103,N_24696,N_25740);
or U27104 (N_27104,N_24101,N_25631);
or U27105 (N_27105,N_24821,N_24123);
nor U27106 (N_27106,N_24979,N_24214);
nor U27107 (N_27107,N_25762,N_24816);
or U27108 (N_27108,N_24649,N_24183);
and U27109 (N_27109,N_24409,N_24930);
and U27110 (N_27110,N_25616,N_24938);
and U27111 (N_27111,N_24268,N_25182);
nand U27112 (N_27112,N_24451,N_24828);
nand U27113 (N_27113,N_25512,N_24367);
and U27114 (N_27114,N_25252,N_24862);
nand U27115 (N_27115,N_24826,N_25871);
or U27116 (N_27116,N_25262,N_25147);
nor U27117 (N_27117,N_24298,N_25211);
or U27118 (N_27118,N_25681,N_25209);
or U27119 (N_27119,N_25851,N_24905);
or U27120 (N_27120,N_24372,N_24452);
or U27121 (N_27121,N_25338,N_25679);
and U27122 (N_27122,N_24264,N_25519);
nor U27123 (N_27123,N_24060,N_25513);
and U27124 (N_27124,N_25752,N_24004);
nand U27125 (N_27125,N_25797,N_24809);
nand U27126 (N_27126,N_25673,N_24839);
and U27127 (N_27127,N_25678,N_24044);
nand U27128 (N_27128,N_24631,N_24716);
xor U27129 (N_27129,N_24174,N_25123);
and U27130 (N_27130,N_25666,N_25678);
and U27131 (N_27131,N_25133,N_25764);
or U27132 (N_27132,N_24444,N_24835);
nor U27133 (N_27133,N_24064,N_24179);
nand U27134 (N_27134,N_25751,N_24293);
nor U27135 (N_27135,N_24075,N_24913);
nand U27136 (N_27136,N_25072,N_25467);
nand U27137 (N_27137,N_24603,N_25694);
nor U27138 (N_27138,N_24981,N_24073);
nand U27139 (N_27139,N_24752,N_24424);
or U27140 (N_27140,N_24921,N_25934);
nand U27141 (N_27141,N_24384,N_25078);
nand U27142 (N_27142,N_24570,N_24482);
nor U27143 (N_27143,N_24195,N_25986);
nand U27144 (N_27144,N_25087,N_24870);
and U27145 (N_27145,N_25034,N_25947);
and U27146 (N_27146,N_24357,N_25569);
nor U27147 (N_27147,N_25377,N_24178);
nor U27148 (N_27148,N_24754,N_24554);
nor U27149 (N_27149,N_24330,N_25084);
nand U27150 (N_27150,N_24881,N_25564);
nor U27151 (N_27151,N_24767,N_24864);
nand U27152 (N_27152,N_24951,N_24671);
or U27153 (N_27153,N_25458,N_24296);
and U27154 (N_27154,N_24883,N_25598);
or U27155 (N_27155,N_25887,N_25358);
or U27156 (N_27156,N_24088,N_24106);
and U27157 (N_27157,N_25534,N_24967);
or U27158 (N_27158,N_24078,N_24500);
and U27159 (N_27159,N_25085,N_24084);
or U27160 (N_27160,N_24528,N_24904);
nor U27161 (N_27161,N_25298,N_25629);
nor U27162 (N_27162,N_24623,N_24437);
nand U27163 (N_27163,N_25103,N_25766);
and U27164 (N_27164,N_25351,N_24333);
nor U27165 (N_27165,N_25692,N_24284);
and U27166 (N_27166,N_25755,N_25108);
nand U27167 (N_27167,N_24432,N_25097);
nor U27168 (N_27168,N_25915,N_24287);
and U27169 (N_27169,N_24641,N_25147);
nor U27170 (N_27170,N_24096,N_25018);
and U27171 (N_27171,N_24950,N_25756);
nor U27172 (N_27172,N_24576,N_25219);
or U27173 (N_27173,N_25739,N_24654);
or U27174 (N_27174,N_25220,N_24140);
and U27175 (N_27175,N_25922,N_24850);
or U27176 (N_27176,N_24721,N_24145);
nand U27177 (N_27177,N_25014,N_24345);
nand U27178 (N_27178,N_25995,N_24315);
nand U27179 (N_27179,N_25148,N_25269);
nand U27180 (N_27180,N_24796,N_24952);
nand U27181 (N_27181,N_24637,N_24485);
and U27182 (N_27182,N_24103,N_25435);
nor U27183 (N_27183,N_25636,N_25536);
nor U27184 (N_27184,N_24771,N_24475);
or U27185 (N_27185,N_25552,N_25679);
and U27186 (N_27186,N_25018,N_25196);
or U27187 (N_27187,N_25202,N_25757);
xor U27188 (N_27188,N_25979,N_24131);
and U27189 (N_27189,N_24574,N_25648);
and U27190 (N_27190,N_25044,N_25376);
nand U27191 (N_27191,N_24516,N_24213);
and U27192 (N_27192,N_24328,N_24866);
nor U27193 (N_27193,N_24026,N_25183);
nor U27194 (N_27194,N_24781,N_25885);
nand U27195 (N_27195,N_25523,N_25285);
nand U27196 (N_27196,N_24507,N_24900);
nand U27197 (N_27197,N_24038,N_24658);
or U27198 (N_27198,N_25094,N_24105);
xor U27199 (N_27199,N_25012,N_25936);
nor U27200 (N_27200,N_25118,N_24307);
and U27201 (N_27201,N_25904,N_24362);
nor U27202 (N_27202,N_25401,N_24149);
nor U27203 (N_27203,N_24628,N_25447);
xnor U27204 (N_27204,N_25449,N_25869);
nor U27205 (N_27205,N_25715,N_25391);
or U27206 (N_27206,N_24919,N_25176);
nor U27207 (N_27207,N_25146,N_24551);
and U27208 (N_27208,N_25889,N_24859);
nand U27209 (N_27209,N_25433,N_24036);
nand U27210 (N_27210,N_25760,N_24989);
or U27211 (N_27211,N_25765,N_24568);
nor U27212 (N_27212,N_24032,N_25278);
nor U27213 (N_27213,N_24487,N_25955);
or U27214 (N_27214,N_25720,N_24747);
or U27215 (N_27215,N_25329,N_24878);
nor U27216 (N_27216,N_24117,N_25485);
and U27217 (N_27217,N_25002,N_25307);
and U27218 (N_27218,N_25709,N_25763);
and U27219 (N_27219,N_25861,N_25634);
nor U27220 (N_27220,N_24331,N_24255);
and U27221 (N_27221,N_24917,N_24214);
nor U27222 (N_27222,N_24109,N_24731);
and U27223 (N_27223,N_25861,N_24370);
nand U27224 (N_27224,N_25772,N_24767);
nor U27225 (N_27225,N_25832,N_25587);
and U27226 (N_27226,N_25288,N_24746);
and U27227 (N_27227,N_25394,N_24878);
or U27228 (N_27228,N_24807,N_25946);
nor U27229 (N_27229,N_25018,N_24697);
or U27230 (N_27230,N_24620,N_25052);
nor U27231 (N_27231,N_24345,N_25586);
and U27232 (N_27232,N_25695,N_24953);
xor U27233 (N_27233,N_24648,N_24485);
and U27234 (N_27234,N_24675,N_25831);
or U27235 (N_27235,N_25308,N_25914);
nand U27236 (N_27236,N_24161,N_24577);
nor U27237 (N_27237,N_25079,N_24162);
and U27238 (N_27238,N_24281,N_25231);
and U27239 (N_27239,N_25998,N_24394);
nor U27240 (N_27240,N_24745,N_25420);
nor U27241 (N_27241,N_24493,N_25748);
or U27242 (N_27242,N_25102,N_25595);
and U27243 (N_27243,N_25569,N_24392);
or U27244 (N_27244,N_25657,N_24382);
nor U27245 (N_27245,N_24530,N_24280);
or U27246 (N_27246,N_25846,N_24775);
nand U27247 (N_27247,N_24748,N_25814);
and U27248 (N_27248,N_24343,N_24166);
or U27249 (N_27249,N_24022,N_25304);
and U27250 (N_27250,N_24973,N_25576);
nand U27251 (N_27251,N_24089,N_25725);
and U27252 (N_27252,N_25285,N_24844);
nand U27253 (N_27253,N_24691,N_25212);
xor U27254 (N_27254,N_24746,N_25189);
or U27255 (N_27255,N_24495,N_25475);
nand U27256 (N_27256,N_24513,N_25482);
nand U27257 (N_27257,N_25716,N_24673);
or U27258 (N_27258,N_24162,N_25987);
nand U27259 (N_27259,N_25077,N_25662);
or U27260 (N_27260,N_24699,N_24745);
and U27261 (N_27261,N_24063,N_25066);
nor U27262 (N_27262,N_24444,N_25395);
or U27263 (N_27263,N_25980,N_25264);
nor U27264 (N_27264,N_24453,N_25001);
nand U27265 (N_27265,N_25429,N_24433);
nand U27266 (N_27266,N_24898,N_25860);
nor U27267 (N_27267,N_25123,N_24220);
or U27268 (N_27268,N_24586,N_24938);
nand U27269 (N_27269,N_24833,N_24580);
nand U27270 (N_27270,N_25629,N_24943);
xor U27271 (N_27271,N_25285,N_24686);
nand U27272 (N_27272,N_25993,N_25540);
nand U27273 (N_27273,N_24175,N_24035);
and U27274 (N_27274,N_24300,N_25005);
xnor U27275 (N_27275,N_25980,N_25114);
or U27276 (N_27276,N_24567,N_25230);
and U27277 (N_27277,N_25854,N_24058);
nor U27278 (N_27278,N_24111,N_24410);
and U27279 (N_27279,N_24062,N_24900);
or U27280 (N_27280,N_25616,N_24437);
nor U27281 (N_27281,N_24837,N_25928);
nand U27282 (N_27282,N_25765,N_25439);
or U27283 (N_27283,N_25948,N_24554);
nand U27284 (N_27284,N_25568,N_24082);
or U27285 (N_27285,N_25209,N_24269);
nor U27286 (N_27286,N_24216,N_25505);
nor U27287 (N_27287,N_25014,N_24085);
nand U27288 (N_27288,N_24666,N_24705);
nand U27289 (N_27289,N_24262,N_25592);
nand U27290 (N_27290,N_24373,N_25752);
nor U27291 (N_27291,N_24891,N_24860);
nor U27292 (N_27292,N_25249,N_25154);
nor U27293 (N_27293,N_24581,N_25617);
nor U27294 (N_27294,N_25324,N_25451);
and U27295 (N_27295,N_24257,N_24276);
or U27296 (N_27296,N_24212,N_25040);
nand U27297 (N_27297,N_24476,N_25592);
nand U27298 (N_27298,N_24340,N_25152);
or U27299 (N_27299,N_25999,N_24613);
and U27300 (N_27300,N_25236,N_24751);
or U27301 (N_27301,N_24467,N_25745);
or U27302 (N_27302,N_24351,N_24954);
or U27303 (N_27303,N_25434,N_25234);
nor U27304 (N_27304,N_25898,N_25971);
xnor U27305 (N_27305,N_24711,N_24673);
and U27306 (N_27306,N_25321,N_24895);
nand U27307 (N_27307,N_24718,N_24883);
nand U27308 (N_27308,N_24714,N_24283);
nand U27309 (N_27309,N_24400,N_25755);
or U27310 (N_27310,N_25708,N_24422);
nor U27311 (N_27311,N_24235,N_25502);
nor U27312 (N_27312,N_24557,N_24983);
and U27313 (N_27313,N_25957,N_24008);
or U27314 (N_27314,N_24481,N_25943);
or U27315 (N_27315,N_24633,N_25046);
or U27316 (N_27316,N_25848,N_24485);
nand U27317 (N_27317,N_24006,N_25616);
nor U27318 (N_27318,N_24468,N_25890);
or U27319 (N_27319,N_24298,N_24069);
nor U27320 (N_27320,N_24593,N_25537);
and U27321 (N_27321,N_25624,N_25222);
nor U27322 (N_27322,N_25260,N_24723);
xnor U27323 (N_27323,N_24355,N_25340);
or U27324 (N_27324,N_25029,N_24437);
or U27325 (N_27325,N_25533,N_24701);
and U27326 (N_27326,N_24930,N_25330);
nand U27327 (N_27327,N_24393,N_25448);
nand U27328 (N_27328,N_25955,N_25085);
nand U27329 (N_27329,N_24398,N_25450);
or U27330 (N_27330,N_25121,N_25194);
or U27331 (N_27331,N_24396,N_24552);
nand U27332 (N_27332,N_25252,N_24370);
xor U27333 (N_27333,N_24075,N_24772);
and U27334 (N_27334,N_24561,N_25430);
nor U27335 (N_27335,N_25442,N_24637);
xor U27336 (N_27336,N_24346,N_24017);
nand U27337 (N_27337,N_25513,N_25292);
or U27338 (N_27338,N_25903,N_25254);
nor U27339 (N_27339,N_25070,N_24729);
or U27340 (N_27340,N_25025,N_25506);
nor U27341 (N_27341,N_25443,N_24880);
nand U27342 (N_27342,N_25864,N_25806);
nor U27343 (N_27343,N_25132,N_25386);
nor U27344 (N_27344,N_24305,N_25603);
nand U27345 (N_27345,N_24079,N_24163);
and U27346 (N_27346,N_25305,N_25794);
xnor U27347 (N_27347,N_25379,N_24410);
and U27348 (N_27348,N_24733,N_25190);
and U27349 (N_27349,N_24356,N_25808);
nand U27350 (N_27350,N_24257,N_24238);
nand U27351 (N_27351,N_25726,N_25668);
or U27352 (N_27352,N_25258,N_25130);
and U27353 (N_27353,N_25324,N_24254);
nand U27354 (N_27354,N_25985,N_25418);
nor U27355 (N_27355,N_24253,N_25573);
and U27356 (N_27356,N_25350,N_24140);
or U27357 (N_27357,N_24627,N_24936);
nand U27358 (N_27358,N_24615,N_25232);
and U27359 (N_27359,N_25802,N_24111);
or U27360 (N_27360,N_24583,N_24613);
and U27361 (N_27361,N_25407,N_25157);
nand U27362 (N_27362,N_24331,N_25495);
and U27363 (N_27363,N_24136,N_25331);
and U27364 (N_27364,N_24041,N_24640);
nor U27365 (N_27365,N_25425,N_24657);
xor U27366 (N_27366,N_24546,N_24081);
or U27367 (N_27367,N_25119,N_24556);
and U27368 (N_27368,N_24797,N_24066);
and U27369 (N_27369,N_25374,N_25788);
or U27370 (N_27370,N_24420,N_25210);
or U27371 (N_27371,N_24406,N_25362);
or U27372 (N_27372,N_25406,N_25305);
xor U27373 (N_27373,N_25301,N_25462);
nor U27374 (N_27374,N_25774,N_24905);
and U27375 (N_27375,N_25075,N_25685);
and U27376 (N_27376,N_25560,N_25199);
or U27377 (N_27377,N_24675,N_24587);
and U27378 (N_27378,N_25877,N_25126);
nand U27379 (N_27379,N_24491,N_25148);
nor U27380 (N_27380,N_24421,N_25869);
nand U27381 (N_27381,N_24566,N_25428);
nand U27382 (N_27382,N_24549,N_25842);
or U27383 (N_27383,N_25358,N_24169);
or U27384 (N_27384,N_24942,N_24736);
nor U27385 (N_27385,N_24395,N_24322);
and U27386 (N_27386,N_25533,N_25835);
nor U27387 (N_27387,N_24218,N_25680);
or U27388 (N_27388,N_25301,N_25957);
nand U27389 (N_27389,N_24128,N_25771);
nand U27390 (N_27390,N_25338,N_25436);
and U27391 (N_27391,N_25428,N_24399);
and U27392 (N_27392,N_24511,N_25839);
xor U27393 (N_27393,N_25784,N_24089);
nand U27394 (N_27394,N_24015,N_24992);
and U27395 (N_27395,N_25790,N_24388);
nor U27396 (N_27396,N_24443,N_25597);
or U27397 (N_27397,N_24375,N_24107);
and U27398 (N_27398,N_25516,N_25680);
nand U27399 (N_27399,N_24195,N_24712);
nand U27400 (N_27400,N_24524,N_25411);
nand U27401 (N_27401,N_24846,N_25535);
and U27402 (N_27402,N_24481,N_25844);
nor U27403 (N_27403,N_25882,N_24641);
nand U27404 (N_27404,N_25497,N_25466);
or U27405 (N_27405,N_25940,N_24031);
nand U27406 (N_27406,N_24085,N_24404);
nor U27407 (N_27407,N_25384,N_25550);
and U27408 (N_27408,N_24866,N_25665);
or U27409 (N_27409,N_24748,N_25710);
or U27410 (N_27410,N_25719,N_24390);
nand U27411 (N_27411,N_24032,N_24552);
or U27412 (N_27412,N_24191,N_25140);
nand U27413 (N_27413,N_25822,N_25096);
or U27414 (N_27414,N_24290,N_25607);
and U27415 (N_27415,N_25911,N_25821);
nor U27416 (N_27416,N_24710,N_25695);
nand U27417 (N_27417,N_24885,N_24557);
or U27418 (N_27418,N_25964,N_24947);
nor U27419 (N_27419,N_24901,N_24627);
nor U27420 (N_27420,N_25686,N_24358);
nor U27421 (N_27421,N_24335,N_25311);
and U27422 (N_27422,N_25767,N_25832);
nand U27423 (N_27423,N_25272,N_24023);
nor U27424 (N_27424,N_25408,N_24318);
nor U27425 (N_27425,N_24176,N_24023);
and U27426 (N_27426,N_24341,N_25795);
nor U27427 (N_27427,N_25079,N_25467);
nand U27428 (N_27428,N_25210,N_24213);
and U27429 (N_27429,N_25366,N_25088);
or U27430 (N_27430,N_25537,N_24888);
nor U27431 (N_27431,N_25755,N_24500);
nor U27432 (N_27432,N_25111,N_24152);
nor U27433 (N_27433,N_25009,N_24566);
xor U27434 (N_27434,N_25378,N_25901);
nand U27435 (N_27435,N_25701,N_25954);
or U27436 (N_27436,N_25011,N_24097);
or U27437 (N_27437,N_25328,N_24759);
or U27438 (N_27438,N_25108,N_25455);
and U27439 (N_27439,N_24647,N_25293);
nand U27440 (N_27440,N_25630,N_25528);
and U27441 (N_27441,N_25448,N_25623);
or U27442 (N_27442,N_25625,N_24975);
nor U27443 (N_27443,N_25041,N_25314);
nand U27444 (N_27444,N_25026,N_24970);
or U27445 (N_27445,N_25559,N_25867);
and U27446 (N_27446,N_24351,N_24305);
nand U27447 (N_27447,N_24802,N_25609);
and U27448 (N_27448,N_24899,N_24518);
or U27449 (N_27449,N_25615,N_24620);
and U27450 (N_27450,N_25445,N_24850);
or U27451 (N_27451,N_25266,N_25014);
nor U27452 (N_27452,N_25085,N_25626);
nor U27453 (N_27453,N_24107,N_24385);
xnor U27454 (N_27454,N_24148,N_24299);
or U27455 (N_27455,N_25807,N_24776);
and U27456 (N_27456,N_24964,N_25942);
and U27457 (N_27457,N_25099,N_24995);
nor U27458 (N_27458,N_25421,N_24514);
nand U27459 (N_27459,N_25789,N_25497);
nand U27460 (N_27460,N_25286,N_24076);
nor U27461 (N_27461,N_25483,N_25344);
or U27462 (N_27462,N_25480,N_25962);
nand U27463 (N_27463,N_25265,N_24832);
and U27464 (N_27464,N_25658,N_24380);
and U27465 (N_27465,N_25454,N_25919);
or U27466 (N_27466,N_24777,N_25906);
nor U27467 (N_27467,N_24268,N_25597);
nor U27468 (N_27468,N_25667,N_25204);
and U27469 (N_27469,N_25022,N_24074);
or U27470 (N_27470,N_24446,N_24681);
nor U27471 (N_27471,N_24223,N_24483);
and U27472 (N_27472,N_25172,N_24501);
nand U27473 (N_27473,N_25780,N_25741);
and U27474 (N_27474,N_24708,N_25077);
and U27475 (N_27475,N_25030,N_25720);
nor U27476 (N_27476,N_24663,N_24388);
or U27477 (N_27477,N_25936,N_24364);
nand U27478 (N_27478,N_25776,N_25404);
nand U27479 (N_27479,N_24497,N_25692);
or U27480 (N_27480,N_25187,N_24909);
and U27481 (N_27481,N_24665,N_24529);
nand U27482 (N_27482,N_24309,N_24194);
and U27483 (N_27483,N_24607,N_25995);
or U27484 (N_27484,N_25581,N_25096);
and U27485 (N_27485,N_24029,N_25973);
nor U27486 (N_27486,N_25084,N_24217);
nor U27487 (N_27487,N_25885,N_25552);
and U27488 (N_27488,N_24978,N_25707);
and U27489 (N_27489,N_25083,N_24160);
nand U27490 (N_27490,N_24170,N_25423);
nor U27491 (N_27491,N_25458,N_25062);
nand U27492 (N_27492,N_25997,N_24200);
nor U27493 (N_27493,N_25443,N_25762);
nor U27494 (N_27494,N_25527,N_25553);
nand U27495 (N_27495,N_25410,N_25859);
or U27496 (N_27496,N_25522,N_24235);
nand U27497 (N_27497,N_25270,N_24704);
nor U27498 (N_27498,N_24553,N_24755);
and U27499 (N_27499,N_25834,N_24891);
and U27500 (N_27500,N_25390,N_24732);
nand U27501 (N_27501,N_24240,N_25272);
xnor U27502 (N_27502,N_24721,N_24428);
nand U27503 (N_27503,N_25138,N_24961);
and U27504 (N_27504,N_24634,N_24966);
and U27505 (N_27505,N_25898,N_24490);
and U27506 (N_27506,N_25016,N_25048);
nand U27507 (N_27507,N_25963,N_25356);
nand U27508 (N_27508,N_25205,N_25207);
or U27509 (N_27509,N_25807,N_25014);
xnor U27510 (N_27510,N_24546,N_24031);
nor U27511 (N_27511,N_25178,N_25655);
nand U27512 (N_27512,N_24748,N_25732);
or U27513 (N_27513,N_25297,N_24381);
and U27514 (N_27514,N_25736,N_24196);
nor U27515 (N_27515,N_24123,N_25671);
nor U27516 (N_27516,N_25331,N_25883);
and U27517 (N_27517,N_25790,N_25440);
nor U27518 (N_27518,N_24740,N_25640);
or U27519 (N_27519,N_25064,N_25814);
xor U27520 (N_27520,N_25558,N_25463);
nand U27521 (N_27521,N_25904,N_24233);
nand U27522 (N_27522,N_24075,N_24334);
or U27523 (N_27523,N_25036,N_24632);
or U27524 (N_27524,N_24123,N_24046);
nand U27525 (N_27525,N_25218,N_24211);
or U27526 (N_27526,N_25898,N_25924);
and U27527 (N_27527,N_25831,N_24705);
or U27528 (N_27528,N_25233,N_24872);
and U27529 (N_27529,N_24194,N_24142);
or U27530 (N_27530,N_25904,N_24495);
and U27531 (N_27531,N_25937,N_24956);
or U27532 (N_27532,N_24688,N_24313);
or U27533 (N_27533,N_24145,N_25753);
nor U27534 (N_27534,N_24773,N_25269);
nand U27535 (N_27535,N_25460,N_24737);
xnor U27536 (N_27536,N_25707,N_25204);
and U27537 (N_27537,N_25641,N_24348);
and U27538 (N_27538,N_25200,N_24582);
or U27539 (N_27539,N_25770,N_25671);
nor U27540 (N_27540,N_25969,N_25983);
or U27541 (N_27541,N_25997,N_25740);
and U27542 (N_27542,N_24558,N_25828);
nand U27543 (N_27543,N_25368,N_24599);
or U27544 (N_27544,N_25201,N_24208);
or U27545 (N_27545,N_24106,N_25635);
nand U27546 (N_27546,N_25155,N_24955);
and U27547 (N_27547,N_24918,N_25177);
or U27548 (N_27548,N_25838,N_25241);
nor U27549 (N_27549,N_25883,N_24601);
nand U27550 (N_27550,N_24120,N_25535);
nor U27551 (N_27551,N_24106,N_24779);
and U27552 (N_27552,N_25775,N_25885);
and U27553 (N_27553,N_25817,N_25693);
nor U27554 (N_27554,N_24170,N_25929);
and U27555 (N_27555,N_25639,N_24347);
nand U27556 (N_27556,N_25295,N_24549);
or U27557 (N_27557,N_25570,N_25016);
and U27558 (N_27558,N_25754,N_25453);
and U27559 (N_27559,N_25611,N_24111);
or U27560 (N_27560,N_25355,N_25989);
xnor U27561 (N_27561,N_24807,N_25562);
xor U27562 (N_27562,N_25164,N_25415);
nor U27563 (N_27563,N_25691,N_24873);
nor U27564 (N_27564,N_25243,N_25767);
and U27565 (N_27565,N_24541,N_24642);
or U27566 (N_27566,N_24330,N_24375);
nand U27567 (N_27567,N_24938,N_24854);
nor U27568 (N_27568,N_24156,N_25878);
nand U27569 (N_27569,N_24213,N_24971);
nand U27570 (N_27570,N_25458,N_24806);
and U27571 (N_27571,N_24648,N_25537);
nor U27572 (N_27572,N_24726,N_24509);
and U27573 (N_27573,N_25776,N_25657);
nor U27574 (N_27574,N_24419,N_24071);
or U27575 (N_27575,N_24162,N_25570);
or U27576 (N_27576,N_24380,N_24271);
nand U27577 (N_27577,N_25446,N_25061);
and U27578 (N_27578,N_24362,N_24696);
or U27579 (N_27579,N_25975,N_25756);
or U27580 (N_27580,N_25678,N_25402);
or U27581 (N_27581,N_25862,N_25880);
nand U27582 (N_27582,N_25769,N_24291);
or U27583 (N_27583,N_25772,N_25610);
nand U27584 (N_27584,N_24737,N_25347);
nand U27585 (N_27585,N_24715,N_25870);
xor U27586 (N_27586,N_25737,N_24833);
and U27587 (N_27587,N_25677,N_24449);
and U27588 (N_27588,N_25541,N_24831);
or U27589 (N_27589,N_25136,N_25549);
nand U27590 (N_27590,N_25328,N_25207);
nor U27591 (N_27591,N_24109,N_24606);
nor U27592 (N_27592,N_25121,N_25751);
nor U27593 (N_27593,N_25472,N_25709);
or U27594 (N_27594,N_25684,N_24672);
nor U27595 (N_27595,N_24770,N_25517);
and U27596 (N_27596,N_25698,N_24972);
nor U27597 (N_27597,N_24327,N_24699);
and U27598 (N_27598,N_25877,N_25078);
and U27599 (N_27599,N_25871,N_25348);
and U27600 (N_27600,N_24815,N_24612);
or U27601 (N_27601,N_25490,N_25834);
and U27602 (N_27602,N_25306,N_25572);
and U27603 (N_27603,N_25732,N_25294);
and U27604 (N_27604,N_25303,N_24147);
and U27605 (N_27605,N_25062,N_25490);
nand U27606 (N_27606,N_25578,N_24994);
nand U27607 (N_27607,N_25004,N_25339);
or U27608 (N_27608,N_25592,N_24982);
and U27609 (N_27609,N_25715,N_25696);
nor U27610 (N_27610,N_24015,N_25142);
or U27611 (N_27611,N_25229,N_25317);
and U27612 (N_27612,N_24301,N_25011);
nand U27613 (N_27613,N_25115,N_24623);
nand U27614 (N_27614,N_24673,N_24790);
nor U27615 (N_27615,N_24132,N_24229);
or U27616 (N_27616,N_25658,N_25817);
nand U27617 (N_27617,N_25610,N_25833);
or U27618 (N_27618,N_25662,N_24346);
nor U27619 (N_27619,N_24489,N_25117);
or U27620 (N_27620,N_25373,N_25433);
nand U27621 (N_27621,N_24969,N_25021);
and U27622 (N_27622,N_24599,N_24516);
or U27623 (N_27623,N_25032,N_25933);
nor U27624 (N_27624,N_25984,N_25522);
or U27625 (N_27625,N_25469,N_25906);
and U27626 (N_27626,N_24043,N_24047);
nand U27627 (N_27627,N_25210,N_24316);
and U27628 (N_27628,N_25622,N_25326);
or U27629 (N_27629,N_24350,N_24168);
and U27630 (N_27630,N_24363,N_25306);
nor U27631 (N_27631,N_25416,N_24581);
or U27632 (N_27632,N_25383,N_25067);
and U27633 (N_27633,N_25738,N_25955);
and U27634 (N_27634,N_25372,N_24347);
and U27635 (N_27635,N_25177,N_24947);
nand U27636 (N_27636,N_24682,N_25007);
nand U27637 (N_27637,N_24046,N_25622);
or U27638 (N_27638,N_24538,N_25948);
and U27639 (N_27639,N_25223,N_25766);
or U27640 (N_27640,N_24010,N_24111);
nand U27641 (N_27641,N_25160,N_24334);
or U27642 (N_27642,N_25826,N_24195);
or U27643 (N_27643,N_25410,N_25397);
or U27644 (N_27644,N_24270,N_24018);
nand U27645 (N_27645,N_25066,N_25586);
nand U27646 (N_27646,N_24430,N_24108);
or U27647 (N_27647,N_25682,N_25620);
nand U27648 (N_27648,N_25804,N_24326);
xnor U27649 (N_27649,N_24961,N_24070);
xnor U27650 (N_27650,N_25495,N_24773);
nor U27651 (N_27651,N_24570,N_24604);
nor U27652 (N_27652,N_25989,N_25176);
or U27653 (N_27653,N_25318,N_25371);
nand U27654 (N_27654,N_24615,N_24130);
nand U27655 (N_27655,N_24560,N_24975);
nand U27656 (N_27656,N_24485,N_24815);
and U27657 (N_27657,N_25751,N_25447);
or U27658 (N_27658,N_24930,N_24506);
nor U27659 (N_27659,N_24982,N_25521);
xor U27660 (N_27660,N_25685,N_24077);
or U27661 (N_27661,N_24916,N_24258);
nand U27662 (N_27662,N_24362,N_24631);
nor U27663 (N_27663,N_24743,N_25548);
nand U27664 (N_27664,N_25942,N_24124);
nor U27665 (N_27665,N_25456,N_24401);
nand U27666 (N_27666,N_25878,N_25354);
nand U27667 (N_27667,N_24704,N_25369);
xnor U27668 (N_27668,N_24509,N_24394);
or U27669 (N_27669,N_24880,N_25710);
nor U27670 (N_27670,N_25852,N_24841);
nor U27671 (N_27671,N_24130,N_24719);
nor U27672 (N_27672,N_25341,N_24008);
and U27673 (N_27673,N_25096,N_25708);
or U27674 (N_27674,N_24582,N_25264);
nor U27675 (N_27675,N_24807,N_25183);
nor U27676 (N_27676,N_25596,N_25372);
and U27677 (N_27677,N_25523,N_25984);
nor U27678 (N_27678,N_24259,N_25804);
nor U27679 (N_27679,N_24469,N_25086);
and U27680 (N_27680,N_25893,N_25155);
and U27681 (N_27681,N_25339,N_24960);
and U27682 (N_27682,N_24817,N_25701);
nor U27683 (N_27683,N_25641,N_24029);
nand U27684 (N_27684,N_24753,N_25257);
and U27685 (N_27685,N_24824,N_24340);
or U27686 (N_27686,N_25920,N_24355);
and U27687 (N_27687,N_25602,N_24775);
nor U27688 (N_27688,N_24850,N_25563);
or U27689 (N_27689,N_24611,N_24590);
nand U27690 (N_27690,N_24926,N_24399);
or U27691 (N_27691,N_25257,N_25242);
nor U27692 (N_27692,N_24762,N_24163);
and U27693 (N_27693,N_24732,N_25877);
nor U27694 (N_27694,N_24245,N_24517);
nand U27695 (N_27695,N_24396,N_24635);
nand U27696 (N_27696,N_25652,N_24086);
or U27697 (N_27697,N_24773,N_24247);
nor U27698 (N_27698,N_25169,N_25527);
or U27699 (N_27699,N_24018,N_25112);
or U27700 (N_27700,N_24868,N_25889);
or U27701 (N_27701,N_24692,N_25548);
nor U27702 (N_27702,N_25122,N_25668);
nand U27703 (N_27703,N_24741,N_24018);
and U27704 (N_27704,N_25832,N_24308);
nand U27705 (N_27705,N_24747,N_24886);
or U27706 (N_27706,N_24810,N_25394);
or U27707 (N_27707,N_24874,N_25459);
nor U27708 (N_27708,N_24354,N_25288);
and U27709 (N_27709,N_24197,N_24100);
xnor U27710 (N_27710,N_25936,N_25565);
nor U27711 (N_27711,N_25961,N_24101);
nand U27712 (N_27712,N_24638,N_25160);
and U27713 (N_27713,N_25106,N_24916);
or U27714 (N_27714,N_24800,N_24225);
nand U27715 (N_27715,N_25088,N_24510);
nand U27716 (N_27716,N_24609,N_24874);
or U27717 (N_27717,N_24519,N_25920);
nand U27718 (N_27718,N_25695,N_24615);
nor U27719 (N_27719,N_25799,N_25010);
or U27720 (N_27720,N_25652,N_24149);
nor U27721 (N_27721,N_25882,N_24479);
and U27722 (N_27722,N_25497,N_25175);
xor U27723 (N_27723,N_25208,N_25096);
nand U27724 (N_27724,N_24100,N_25350);
or U27725 (N_27725,N_25000,N_24719);
or U27726 (N_27726,N_25179,N_25731);
and U27727 (N_27727,N_25666,N_25341);
nor U27728 (N_27728,N_24447,N_25007);
nand U27729 (N_27729,N_25152,N_25824);
and U27730 (N_27730,N_24582,N_24437);
nand U27731 (N_27731,N_24068,N_24393);
nor U27732 (N_27732,N_24103,N_24994);
nor U27733 (N_27733,N_24021,N_24104);
nor U27734 (N_27734,N_25734,N_24278);
or U27735 (N_27735,N_24889,N_24478);
or U27736 (N_27736,N_25614,N_24142);
xnor U27737 (N_27737,N_25448,N_24644);
or U27738 (N_27738,N_25469,N_24631);
nand U27739 (N_27739,N_24490,N_25830);
nor U27740 (N_27740,N_25300,N_24696);
nor U27741 (N_27741,N_25234,N_25331);
nor U27742 (N_27742,N_24101,N_24169);
nor U27743 (N_27743,N_24457,N_24231);
nand U27744 (N_27744,N_24028,N_25527);
and U27745 (N_27745,N_24587,N_25773);
or U27746 (N_27746,N_24529,N_25379);
nor U27747 (N_27747,N_24507,N_24330);
nor U27748 (N_27748,N_24895,N_25891);
nor U27749 (N_27749,N_24731,N_25071);
nand U27750 (N_27750,N_24636,N_24104);
nand U27751 (N_27751,N_24572,N_24813);
or U27752 (N_27752,N_25807,N_24402);
and U27753 (N_27753,N_24967,N_24942);
and U27754 (N_27754,N_24987,N_25385);
or U27755 (N_27755,N_25057,N_25739);
nand U27756 (N_27756,N_24186,N_24372);
xnor U27757 (N_27757,N_24610,N_24524);
or U27758 (N_27758,N_24421,N_25876);
or U27759 (N_27759,N_24047,N_24418);
nor U27760 (N_27760,N_24896,N_25821);
or U27761 (N_27761,N_24542,N_24083);
nor U27762 (N_27762,N_25719,N_24792);
nand U27763 (N_27763,N_25907,N_25612);
and U27764 (N_27764,N_25815,N_25306);
or U27765 (N_27765,N_24062,N_24552);
and U27766 (N_27766,N_25422,N_25895);
and U27767 (N_27767,N_25438,N_25563);
or U27768 (N_27768,N_24219,N_24972);
and U27769 (N_27769,N_24612,N_24738);
nor U27770 (N_27770,N_25902,N_24984);
nor U27771 (N_27771,N_24439,N_24253);
or U27772 (N_27772,N_24819,N_24683);
nor U27773 (N_27773,N_24544,N_24115);
nor U27774 (N_27774,N_24328,N_25969);
nand U27775 (N_27775,N_25595,N_25761);
and U27776 (N_27776,N_25070,N_25151);
nor U27777 (N_27777,N_24098,N_24120);
nand U27778 (N_27778,N_25158,N_25469);
or U27779 (N_27779,N_25573,N_24433);
nand U27780 (N_27780,N_25100,N_24458);
and U27781 (N_27781,N_24712,N_24150);
nor U27782 (N_27782,N_25391,N_25035);
or U27783 (N_27783,N_24903,N_24748);
nand U27784 (N_27784,N_25741,N_24221);
xnor U27785 (N_27785,N_24192,N_25752);
nand U27786 (N_27786,N_24090,N_25327);
nor U27787 (N_27787,N_24430,N_25269);
or U27788 (N_27788,N_25184,N_24217);
nand U27789 (N_27789,N_24202,N_24005);
nand U27790 (N_27790,N_24621,N_24708);
or U27791 (N_27791,N_24516,N_25235);
nor U27792 (N_27792,N_24088,N_24783);
nor U27793 (N_27793,N_24106,N_25428);
or U27794 (N_27794,N_24926,N_25097);
and U27795 (N_27795,N_25079,N_24578);
and U27796 (N_27796,N_25764,N_25774);
nand U27797 (N_27797,N_24391,N_24173);
nor U27798 (N_27798,N_25895,N_24234);
or U27799 (N_27799,N_24742,N_25906);
nor U27800 (N_27800,N_24775,N_24262);
nand U27801 (N_27801,N_25922,N_25183);
and U27802 (N_27802,N_24099,N_25873);
nor U27803 (N_27803,N_25945,N_24690);
nand U27804 (N_27804,N_25276,N_25877);
or U27805 (N_27805,N_25973,N_25734);
nor U27806 (N_27806,N_25787,N_24916);
or U27807 (N_27807,N_24340,N_24679);
nand U27808 (N_27808,N_25949,N_25595);
nor U27809 (N_27809,N_25673,N_24726);
and U27810 (N_27810,N_24376,N_24545);
nor U27811 (N_27811,N_25152,N_24729);
or U27812 (N_27812,N_24569,N_24828);
or U27813 (N_27813,N_25189,N_25103);
nand U27814 (N_27814,N_24384,N_24576);
or U27815 (N_27815,N_25479,N_24268);
nand U27816 (N_27816,N_25940,N_25713);
or U27817 (N_27817,N_25797,N_24681);
or U27818 (N_27818,N_25391,N_25673);
nor U27819 (N_27819,N_25550,N_24957);
nand U27820 (N_27820,N_24577,N_25247);
or U27821 (N_27821,N_25927,N_25877);
nand U27822 (N_27822,N_24689,N_24087);
or U27823 (N_27823,N_24716,N_24133);
xnor U27824 (N_27824,N_25452,N_25588);
and U27825 (N_27825,N_24015,N_24791);
nor U27826 (N_27826,N_24999,N_25567);
and U27827 (N_27827,N_25132,N_25848);
nor U27828 (N_27828,N_25847,N_24196);
or U27829 (N_27829,N_25189,N_24671);
and U27830 (N_27830,N_24477,N_24069);
and U27831 (N_27831,N_25102,N_24097);
nand U27832 (N_27832,N_25098,N_24228);
or U27833 (N_27833,N_25606,N_24423);
and U27834 (N_27834,N_24495,N_25371);
and U27835 (N_27835,N_24889,N_25562);
nor U27836 (N_27836,N_25085,N_24995);
and U27837 (N_27837,N_24174,N_25821);
nor U27838 (N_27838,N_24406,N_24191);
nand U27839 (N_27839,N_24449,N_24238);
and U27840 (N_27840,N_25968,N_24393);
and U27841 (N_27841,N_25843,N_24038);
nor U27842 (N_27842,N_25751,N_24531);
or U27843 (N_27843,N_25677,N_24592);
nor U27844 (N_27844,N_24059,N_25090);
and U27845 (N_27845,N_25852,N_25675);
nand U27846 (N_27846,N_24717,N_24610);
nand U27847 (N_27847,N_25699,N_25514);
nor U27848 (N_27848,N_24898,N_24306);
nor U27849 (N_27849,N_25704,N_25211);
nor U27850 (N_27850,N_25120,N_24683);
or U27851 (N_27851,N_24862,N_24743);
nand U27852 (N_27852,N_24738,N_25040);
and U27853 (N_27853,N_25855,N_24670);
or U27854 (N_27854,N_25701,N_25046);
nand U27855 (N_27855,N_24217,N_24957);
and U27856 (N_27856,N_25343,N_24350);
or U27857 (N_27857,N_25613,N_25717);
and U27858 (N_27858,N_24643,N_24105);
or U27859 (N_27859,N_25586,N_24573);
nand U27860 (N_27860,N_24266,N_24826);
nand U27861 (N_27861,N_25764,N_25478);
nand U27862 (N_27862,N_24074,N_24610);
nor U27863 (N_27863,N_25841,N_25154);
and U27864 (N_27864,N_24632,N_25260);
nand U27865 (N_27865,N_24527,N_24016);
or U27866 (N_27866,N_25645,N_24049);
and U27867 (N_27867,N_25044,N_24509);
nand U27868 (N_27868,N_25928,N_24786);
nor U27869 (N_27869,N_24561,N_25363);
or U27870 (N_27870,N_24191,N_24680);
and U27871 (N_27871,N_24321,N_24449);
nand U27872 (N_27872,N_25911,N_24269);
nor U27873 (N_27873,N_25302,N_24338);
or U27874 (N_27874,N_25606,N_25322);
nand U27875 (N_27875,N_25447,N_24170);
nor U27876 (N_27876,N_24485,N_25065);
or U27877 (N_27877,N_24725,N_25824);
nand U27878 (N_27878,N_24053,N_24331);
xnor U27879 (N_27879,N_25722,N_24172);
nor U27880 (N_27880,N_25508,N_25509);
nand U27881 (N_27881,N_24401,N_25890);
nor U27882 (N_27882,N_24660,N_25071);
nand U27883 (N_27883,N_25347,N_24604);
nor U27884 (N_27884,N_24501,N_24799);
and U27885 (N_27885,N_25212,N_25104);
and U27886 (N_27886,N_25175,N_25386);
nor U27887 (N_27887,N_25751,N_25527);
or U27888 (N_27888,N_25211,N_25546);
or U27889 (N_27889,N_24007,N_24416);
or U27890 (N_27890,N_25974,N_24651);
nand U27891 (N_27891,N_25950,N_24805);
and U27892 (N_27892,N_24801,N_24840);
nand U27893 (N_27893,N_24828,N_24420);
nand U27894 (N_27894,N_25078,N_24037);
and U27895 (N_27895,N_24008,N_25618);
nand U27896 (N_27896,N_25761,N_25452);
nand U27897 (N_27897,N_25586,N_24619);
nand U27898 (N_27898,N_24095,N_24688);
nor U27899 (N_27899,N_24047,N_25523);
and U27900 (N_27900,N_25445,N_25709);
nor U27901 (N_27901,N_24343,N_24466);
and U27902 (N_27902,N_24717,N_24351);
nor U27903 (N_27903,N_25594,N_25399);
and U27904 (N_27904,N_24606,N_24584);
and U27905 (N_27905,N_24470,N_25061);
and U27906 (N_27906,N_25539,N_25817);
nand U27907 (N_27907,N_25204,N_24006);
and U27908 (N_27908,N_25581,N_25516);
nor U27909 (N_27909,N_24470,N_24836);
or U27910 (N_27910,N_25341,N_25234);
and U27911 (N_27911,N_24697,N_24731);
nor U27912 (N_27912,N_24292,N_24915);
or U27913 (N_27913,N_24148,N_25012);
and U27914 (N_27914,N_25316,N_25269);
nor U27915 (N_27915,N_24040,N_25369);
and U27916 (N_27916,N_25698,N_25787);
and U27917 (N_27917,N_25789,N_24485);
xnor U27918 (N_27918,N_24555,N_24800);
or U27919 (N_27919,N_24505,N_24881);
and U27920 (N_27920,N_24204,N_25187);
nand U27921 (N_27921,N_24949,N_24763);
or U27922 (N_27922,N_25099,N_25038);
or U27923 (N_27923,N_24468,N_24332);
xor U27924 (N_27924,N_24089,N_25007);
nor U27925 (N_27925,N_25672,N_25239);
and U27926 (N_27926,N_25010,N_24720);
or U27927 (N_27927,N_25416,N_24622);
nor U27928 (N_27928,N_24171,N_25933);
nand U27929 (N_27929,N_24296,N_24645);
nand U27930 (N_27930,N_25676,N_24906);
nand U27931 (N_27931,N_24835,N_24664);
nand U27932 (N_27932,N_25068,N_25858);
nand U27933 (N_27933,N_25269,N_24408);
or U27934 (N_27934,N_24891,N_24008);
or U27935 (N_27935,N_24546,N_25538);
or U27936 (N_27936,N_24587,N_24087);
nor U27937 (N_27937,N_24969,N_24335);
nand U27938 (N_27938,N_24129,N_25025);
or U27939 (N_27939,N_25720,N_24528);
or U27940 (N_27940,N_24790,N_25573);
or U27941 (N_27941,N_25500,N_24455);
or U27942 (N_27942,N_25545,N_24461);
nand U27943 (N_27943,N_25965,N_24520);
nand U27944 (N_27944,N_24518,N_24152);
xor U27945 (N_27945,N_25880,N_25720);
and U27946 (N_27946,N_24549,N_25119);
or U27947 (N_27947,N_24542,N_25820);
nor U27948 (N_27948,N_24191,N_24550);
and U27949 (N_27949,N_25374,N_25750);
nor U27950 (N_27950,N_25005,N_24537);
nor U27951 (N_27951,N_25411,N_24914);
or U27952 (N_27952,N_25543,N_24457);
nand U27953 (N_27953,N_25360,N_25444);
and U27954 (N_27954,N_25949,N_24909);
nand U27955 (N_27955,N_25008,N_24779);
or U27956 (N_27956,N_24812,N_24600);
nand U27957 (N_27957,N_25107,N_24616);
nand U27958 (N_27958,N_25127,N_24254);
nand U27959 (N_27959,N_25293,N_25289);
nor U27960 (N_27960,N_24359,N_25360);
or U27961 (N_27961,N_25962,N_25461);
nand U27962 (N_27962,N_24727,N_24435);
nand U27963 (N_27963,N_25363,N_25124);
and U27964 (N_27964,N_24516,N_25672);
and U27965 (N_27965,N_24724,N_25230);
and U27966 (N_27966,N_24143,N_24059);
or U27967 (N_27967,N_24481,N_24346);
or U27968 (N_27968,N_24547,N_25168);
or U27969 (N_27969,N_25993,N_24038);
nand U27970 (N_27970,N_25018,N_25540);
or U27971 (N_27971,N_24707,N_25953);
nor U27972 (N_27972,N_25193,N_25434);
nor U27973 (N_27973,N_24810,N_24241);
nand U27974 (N_27974,N_24739,N_25576);
or U27975 (N_27975,N_24412,N_25159);
nand U27976 (N_27976,N_24053,N_24679);
nor U27977 (N_27977,N_25086,N_24800);
or U27978 (N_27978,N_25120,N_25530);
nand U27979 (N_27979,N_24942,N_24207);
and U27980 (N_27980,N_25967,N_25643);
nor U27981 (N_27981,N_24428,N_24946);
nand U27982 (N_27982,N_25411,N_24936);
xnor U27983 (N_27983,N_25323,N_24359);
nor U27984 (N_27984,N_25753,N_24013);
nor U27985 (N_27985,N_25939,N_24874);
or U27986 (N_27986,N_25993,N_24293);
nand U27987 (N_27987,N_24775,N_24522);
nand U27988 (N_27988,N_24506,N_24381);
nor U27989 (N_27989,N_24738,N_24219);
nand U27990 (N_27990,N_25638,N_24191);
or U27991 (N_27991,N_24884,N_25959);
nand U27992 (N_27992,N_24992,N_24808);
nor U27993 (N_27993,N_25371,N_24773);
xor U27994 (N_27994,N_24818,N_25069);
nand U27995 (N_27995,N_25047,N_25830);
nand U27996 (N_27996,N_24167,N_24979);
nor U27997 (N_27997,N_24384,N_25205);
and U27998 (N_27998,N_24046,N_25292);
nand U27999 (N_27999,N_25871,N_24324);
or U28000 (N_28000,N_27295,N_26953);
nand U28001 (N_28001,N_27349,N_26231);
or U28002 (N_28002,N_26508,N_27701);
xor U28003 (N_28003,N_26187,N_27046);
nand U28004 (N_28004,N_26076,N_26634);
or U28005 (N_28005,N_27641,N_26489);
and U28006 (N_28006,N_27655,N_27103);
and U28007 (N_28007,N_26123,N_27040);
and U28008 (N_28008,N_26128,N_26176);
and U28009 (N_28009,N_27534,N_26906);
nand U28010 (N_28010,N_27512,N_26770);
nand U28011 (N_28011,N_26055,N_26334);
nor U28012 (N_28012,N_27278,N_27780);
nand U28013 (N_28013,N_27174,N_27665);
or U28014 (N_28014,N_26855,N_27000);
and U28015 (N_28015,N_27399,N_27260);
nand U28016 (N_28016,N_26926,N_27925);
and U28017 (N_28017,N_27685,N_27269);
and U28018 (N_28018,N_27517,N_27853);
and U28019 (N_28019,N_27307,N_26667);
nand U28020 (N_28020,N_26956,N_26848);
or U28021 (N_28021,N_27463,N_26645);
and U28022 (N_28022,N_27352,N_27537);
nand U28023 (N_28023,N_27870,N_26539);
nor U28024 (N_28024,N_26309,N_27603);
xor U28025 (N_28025,N_26476,N_27956);
or U28026 (N_28026,N_26918,N_26138);
nor U28027 (N_28027,N_27614,N_26766);
nand U28028 (N_28028,N_26612,N_26842);
nor U28029 (N_28029,N_26199,N_26390);
nor U28030 (N_28030,N_27508,N_27973);
or U28031 (N_28031,N_27860,N_26499);
or U28032 (N_28032,N_27112,N_27808);
or U28033 (N_28033,N_26198,N_26074);
nand U28034 (N_28034,N_27520,N_26229);
and U28035 (N_28035,N_27358,N_26980);
nor U28036 (N_28036,N_27444,N_26912);
or U28037 (N_28037,N_26638,N_27494);
or U28038 (N_28038,N_26541,N_26393);
or U28039 (N_28039,N_26023,N_26837);
and U28040 (N_28040,N_27228,N_27716);
nand U28041 (N_28041,N_26321,N_26678);
nor U28042 (N_28042,N_27108,N_27284);
or U28043 (N_28043,N_27903,N_26360);
xnor U28044 (N_28044,N_26226,N_26751);
nand U28045 (N_28045,N_27626,N_26028);
or U28046 (N_28046,N_27505,N_26600);
and U28047 (N_28047,N_26915,N_27457);
and U28048 (N_28048,N_26069,N_26119);
and U28049 (N_28049,N_27281,N_27674);
xor U28050 (N_28050,N_26440,N_26588);
nand U28051 (N_28051,N_27114,N_27948);
nand U28052 (N_28052,N_26181,N_26898);
and U28053 (N_28053,N_26991,N_26790);
and U28054 (N_28054,N_27985,N_26474);
nand U28055 (N_28055,N_26978,N_26479);
or U28056 (N_28056,N_27210,N_26594);
or U28057 (N_28057,N_26486,N_27793);
and U28058 (N_28058,N_27316,N_27382);
or U28059 (N_28059,N_27299,N_27207);
nand U28060 (N_28060,N_26903,N_27042);
nand U28061 (N_28061,N_27197,N_27468);
or U28062 (N_28062,N_26428,N_26294);
nor U28063 (N_28063,N_27335,N_27462);
or U28064 (N_28064,N_26758,N_26787);
and U28065 (N_28065,N_26523,N_26773);
and U28066 (N_28066,N_26937,N_26133);
or U28067 (N_28067,N_27863,N_26989);
and U28068 (N_28068,N_27240,N_26732);
or U28069 (N_28069,N_26129,N_27740);
or U28070 (N_28070,N_26884,N_27699);
and U28071 (N_28071,N_26386,N_26747);
and U28072 (N_28072,N_26931,N_27830);
or U28073 (N_28073,N_26739,N_27972);
nor U28074 (N_28074,N_27157,N_27497);
and U28075 (N_28075,N_26689,N_27642);
nand U28076 (N_28076,N_26228,N_26603);
nand U28077 (N_28077,N_26968,N_26994);
or U28078 (N_28078,N_26312,N_27688);
and U28079 (N_28079,N_26344,N_27540);
or U28080 (N_28080,N_26418,N_26168);
nor U28081 (N_28081,N_26308,N_27082);
and U28082 (N_28082,N_27552,N_26992);
nor U28083 (N_28083,N_26972,N_27049);
and U28084 (N_28084,N_27730,N_27158);
nor U28085 (N_28085,N_26338,N_27110);
or U28086 (N_28086,N_26748,N_26870);
and U28087 (N_28087,N_27017,N_26147);
and U28088 (N_28088,N_27785,N_27181);
nand U28089 (N_28089,N_27484,N_26429);
nand U28090 (N_28090,N_26781,N_26840);
xor U28091 (N_28091,N_26565,N_27448);
nor U28092 (N_28092,N_27589,N_27951);
nor U28093 (N_28093,N_27450,N_27563);
nand U28094 (N_28094,N_27579,N_26871);
and U28095 (N_28095,N_27900,N_26144);
or U28096 (N_28096,N_27731,N_27081);
xor U28097 (N_28097,N_27729,N_26013);
nand U28098 (N_28098,N_26711,N_26712);
or U28099 (N_28099,N_27962,N_27694);
nor U28100 (N_28100,N_26544,N_27053);
nor U28101 (N_28101,N_26679,N_27050);
nand U28102 (N_28102,N_27713,N_27193);
nand U28103 (N_28103,N_27543,N_26714);
nor U28104 (N_28104,N_27763,N_26530);
and U28105 (N_28105,N_27464,N_27979);
nand U28106 (N_28106,N_26412,N_26111);
nand U28107 (N_28107,N_27089,N_27211);
nand U28108 (N_28108,N_27811,N_27127);
and U28109 (N_28109,N_26369,N_27850);
or U28110 (N_28110,N_27954,N_27375);
nor U28111 (N_28111,N_26396,N_27213);
and U28112 (N_28112,N_27815,N_27798);
and U28113 (N_28113,N_27647,N_26527);
and U28114 (N_28114,N_26613,N_26987);
nand U28115 (N_28115,N_26012,N_27254);
nor U28116 (N_28116,N_26681,N_26222);
nand U28117 (N_28117,N_26365,N_26126);
nand U28118 (N_28118,N_26949,N_27721);
and U28119 (N_28119,N_26162,N_26720);
nand U28120 (N_28120,N_27249,N_26045);
nand U28121 (N_28121,N_26608,N_26815);
nand U28122 (N_28122,N_26173,N_27212);
or U28123 (N_28123,N_26165,N_26546);
nor U28124 (N_28124,N_26290,N_26626);
nand U28125 (N_28125,N_27714,N_27059);
or U28126 (N_28126,N_26889,N_27670);
or U28127 (N_28127,N_26340,N_27624);
or U28128 (N_28128,N_27341,N_26876);
or U28129 (N_28129,N_27995,N_26079);
xor U28130 (N_28130,N_26110,N_26826);
nand U28131 (N_28131,N_27509,N_26155);
or U28132 (N_28132,N_26450,N_27649);
nand U28133 (N_28133,N_27290,N_27007);
nand U28134 (N_28134,N_26291,N_27594);
or U28135 (N_28135,N_26952,N_26736);
and U28136 (N_28136,N_27504,N_26057);
nor U28137 (N_28137,N_26413,N_27009);
nand U28138 (N_28138,N_26256,N_26172);
nor U28139 (N_28139,N_27220,N_27291);
xor U28140 (N_28140,N_27364,N_26621);
and U28141 (N_28141,N_26142,N_26472);
nand U28142 (N_28142,N_27136,N_27828);
and U28143 (N_28143,N_27266,N_27897);
xnor U28144 (N_28144,N_27935,N_27315);
nand U28145 (N_28145,N_26282,N_27218);
nor U28146 (N_28146,N_27003,N_27086);
nand U28147 (N_28147,N_26467,N_26190);
and U28148 (N_28148,N_26669,N_26922);
nor U28149 (N_28149,N_27918,N_27816);
or U28150 (N_28150,N_26037,N_26267);
nand U28151 (N_28151,N_27060,N_26402);
or U28152 (N_28152,N_26897,N_26847);
nor U28153 (N_28153,N_27423,N_26461);
and U28154 (N_28154,N_26097,N_26117);
nand U28155 (N_28155,N_26742,N_26027);
nor U28156 (N_28156,N_27123,N_27597);
nand U28157 (N_28157,N_27585,N_27156);
or U28158 (N_28158,N_27809,N_27404);
nand U28159 (N_28159,N_27433,N_27263);
nor U28160 (N_28160,N_27654,N_27131);
nand U28161 (N_28161,N_26895,N_27424);
nand U28162 (N_28162,N_26026,N_26211);
or U28163 (N_28163,N_26288,N_27090);
and U28164 (N_28164,N_27340,N_27877);
nand U28165 (N_28165,N_26925,N_26813);
and U28166 (N_28166,N_27247,N_27481);
or U28167 (N_28167,N_26596,N_27888);
nand U28168 (N_28168,N_26259,N_27309);
nor U28169 (N_28169,N_27803,N_27631);
or U28170 (N_28170,N_27664,N_26171);
or U28171 (N_28171,N_26475,N_27311);
nor U28172 (N_28172,N_26439,N_26379);
nor U28173 (N_28173,N_27313,N_26136);
nor U28174 (N_28174,N_27736,N_27273);
and U28175 (N_28175,N_26272,N_26219);
or U28176 (N_28176,N_26096,N_27297);
nor U28177 (N_28177,N_26954,N_27582);
xor U28178 (N_28178,N_27396,N_26820);
and U28179 (N_28179,N_26341,N_27025);
nand U28180 (N_28180,N_27405,N_27357);
or U28181 (N_28181,N_27370,N_27326);
and U28182 (N_28182,N_27936,N_26075);
nor U28183 (N_28183,N_27184,N_27195);
or U28184 (N_28184,N_27486,N_26618);
nand U28185 (N_28185,N_27715,N_27078);
or U28186 (N_28186,N_27401,N_27970);
nor U28187 (N_28187,N_26010,N_27071);
nand U28188 (N_28188,N_27539,N_27513);
nor U28189 (N_28189,N_27101,N_27922);
and U28190 (N_28190,N_27518,N_26002);
or U28191 (N_28191,N_27696,N_26682);
nor U28192 (N_28192,N_27104,N_27248);
nor U28193 (N_28193,N_26447,N_26981);
nor U28194 (N_28194,N_27703,N_26389);
or U28195 (N_28195,N_26754,N_27282);
and U28196 (N_28196,N_27591,N_27035);
nor U28197 (N_28197,N_27532,N_27933);
or U28198 (N_28198,N_26904,N_27366);
and U28199 (N_28199,N_27039,N_27876);
or U28200 (N_28200,N_27971,N_27430);
xnor U28201 (N_28201,N_26623,N_27931);
nor U28202 (N_28202,N_26283,N_26929);
nor U28203 (N_28203,N_27362,N_26407);
or U28204 (N_28204,N_27294,N_26109);
nor U28205 (N_28205,N_26217,N_27140);
or U28206 (N_28206,N_27554,N_27030);
or U28207 (N_28207,N_26798,N_26209);
and U28208 (N_28208,N_26319,N_26342);
nor U28209 (N_28209,N_27690,N_26349);
nand U28210 (N_28210,N_27545,N_27343);
and U28211 (N_28211,N_26462,N_26072);
nor U28212 (N_28212,N_26204,N_26299);
and U28213 (N_28213,N_27635,N_27223);
or U28214 (N_28214,N_26031,N_26350);
nor U28215 (N_28215,N_27515,N_27121);
or U28216 (N_28216,N_27879,N_26210);
or U28217 (N_28217,N_26230,N_27460);
or U28218 (N_28218,N_27923,N_26392);
nand U28219 (N_28219,N_27363,N_27076);
and U28220 (N_28220,N_26131,N_27700);
nor U28221 (N_28221,N_26320,N_27596);
or U28222 (N_28222,N_27243,N_26627);
nor U28223 (N_28223,N_26426,N_26652);
and U28224 (N_28224,N_26080,N_27774);
or U28225 (N_28225,N_26504,N_26744);
nor U28226 (N_28226,N_27332,N_26697);
xor U28227 (N_28227,N_26394,N_27638);
and U28228 (N_28228,N_27998,N_26124);
nand U28229 (N_28229,N_27365,N_26297);
nor U28230 (N_28230,N_27560,N_27800);
nor U28231 (N_28231,N_27781,N_27441);
nand U28232 (N_28232,N_26060,N_26240);
and U28233 (N_28233,N_27408,N_26725);
nor U28234 (N_28234,N_26997,N_27788);
or U28235 (N_28235,N_26969,N_27394);
nand U28236 (N_28236,N_27361,N_27572);
nand U28237 (N_28237,N_26641,N_26692);
nor U28238 (N_28238,N_27675,N_27252);
or U28239 (N_28239,N_26373,N_26347);
nor U28240 (N_28240,N_27821,N_27976);
or U28241 (N_28241,N_26914,N_26572);
nor U28242 (N_28242,N_27264,N_26177);
or U28243 (N_28243,N_26322,N_26841);
or U28244 (N_28244,N_27452,N_26540);
nor U28245 (N_28245,N_26965,N_27420);
nand U28246 (N_28246,N_27344,N_26693);
nor U28247 (N_28247,N_27584,N_26445);
and U28248 (N_28248,N_26470,N_27190);
nor U28249 (N_28249,N_26366,N_27529);
nand U28250 (N_28250,N_26427,N_26468);
nand U28251 (N_28251,N_27899,N_26990);
nor U28252 (N_28252,N_26574,N_27232);
and U28253 (N_28253,N_26056,N_26705);
nor U28254 (N_28254,N_26478,N_26963);
nor U28255 (N_28255,N_27199,N_27029);
nor U28256 (N_28256,N_27824,N_27262);
or U28257 (N_28257,N_26849,N_26242);
or U28258 (N_28258,N_27546,N_26044);
and U28259 (N_28259,N_27728,N_27338);
nor U28260 (N_28260,N_27753,N_26633);
or U28261 (N_28261,N_27246,N_26276);
nor U28262 (N_28262,N_27975,N_26254);
and U28263 (N_28263,N_26303,N_26713);
and U28264 (N_28264,N_27272,N_27153);
or U28265 (N_28265,N_27322,N_26146);
nand U28266 (N_28266,N_26823,N_27478);
and U28267 (N_28267,N_26831,N_27531);
nand U28268 (N_28268,N_27627,N_27439);
nor U28269 (N_28269,N_27967,N_26514);
nor U28270 (N_28270,N_27706,N_27864);
or U28271 (N_28271,N_27194,N_27469);
or U28272 (N_28272,N_26616,N_27818);
or U28273 (N_28273,N_27856,N_26318);
nor U28274 (N_28274,N_27477,N_27611);
nor U28275 (N_28275,N_26502,N_27301);
or U28276 (N_28276,N_26213,N_27575);
nor U28277 (N_28277,N_26068,N_26493);
nand U28278 (N_28278,N_26277,N_26717);
nand U28279 (N_28279,N_26708,N_26300);
nand U28280 (N_28280,N_26431,N_27306);
nor U28281 (N_28281,N_26971,N_26970);
nor U28282 (N_28282,N_26535,N_27491);
xnor U28283 (N_28283,N_27680,N_27710);
and U28284 (N_28284,N_26246,N_26496);
nor U28285 (N_28285,N_26672,N_27937);
nand U28286 (N_28286,N_26515,N_26212);
nand U28287 (N_28287,N_26545,N_26160);
or U28288 (N_28288,N_27606,N_26030);
nor U28289 (N_28289,N_27372,N_27737);
and U28290 (N_28290,N_26356,N_26585);
and U28291 (N_28291,N_27427,N_26786);
and U28292 (N_28292,N_27259,N_27063);
nor U28293 (N_28293,N_27835,N_27229);
nor U28294 (N_28294,N_27032,N_26785);
nor U28295 (N_28295,N_27744,N_27727);
nor U28296 (N_28296,N_26551,N_26036);
and U28297 (N_28297,N_27473,N_26803);
nor U28298 (N_28298,N_26215,N_27077);
and U28299 (N_28299,N_26016,N_27607);
nor U28300 (N_28300,N_27887,N_26580);
or U28301 (N_28301,N_26568,N_26206);
nor U28302 (N_28302,N_27432,N_26384);
or U28303 (N_28303,N_26631,N_26879);
nand U28304 (N_28304,N_27650,N_27910);
or U28305 (N_28305,N_26741,N_27447);
nor U28306 (N_28306,N_27549,N_26067);
or U28307 (N_28307,N_26833,N_26579);
nand U28308 (N_28308,N_26361,N_27455);
and U28309 (N_28309,N_26999,N_26017);
nand U28310 (N_28310,N_26995,N_26930);
and U28311 (N_28311,N_26329,N_26856);
nor U28312 (N_28312,N_27048,N_27506);
nor U28313 (N_28313,N_27791,N_26159);
nand U28314 (N_28314,N_27734,N_26643);
nor U28315 (N_28315,N_26690,N_27709);
and U28316 (N_28316,N_26114,N_26404);
or U28317 (N_28317,N_26196,N_27746);
nand U28318 (N_28318,N_27356,N_27339);
nor U28319 (N_28319,N_27932,N_26182);
nor U28320 (N_28320,N_26385,N_26250);
and U28321 (N_28321,N_26140,N_27390);
or U28322 (N_28322,N_27732,N_27304);
nand U28323 (N_28323,N_27135,N_27601);
and U28324 (N_28324,N_27276,N_27386);
and U28325 (N_28325,N_26087,N_26622);
and U28326 (N_28326,N_26314,N_27541);
or U28327 (N_28327,N_27946,N_27350);
nor U28328 (N_28328,N_27720,N_27057);
and U28329 (N_28329,N_27538,N_26490);
or U28330 (N_28330,N_26592,N_26305);
xor U28331 (N_28331,N_27329,N_27012);
or U28332 (N_28332,N_27833,N_27268);
or U28333 (N_28333,N_26867,N_26039);
nand U28334 (N_28334,N_26919,N_26169);
and U28335 (N_28335,N_26924,N_26738);
and U28336 (N_28336,N_26619,N_26607);
nand U28337 (N_28337,N_27799,N_26553);
nor U28338 (N_28338,N_26083,N_26481);
and U28339 (N_28339,N_26722,N_27718);
and U28340 (N_28340,N_26591,N_26666);
nand U28341 (N_28341,N_26839,N_26157);
nor U28342 (N_28342,N_27558,N_27418);
nand U28343 (N_28343,N_26101,N_26827);
nand U28344 (N_28344,N_27843,N_26853);
nand U28345 (N_28345,N_26896,N_26830);
nand U28346 (N_28346,N_26756,N_27258);
nand U28347 (N_28347,N_26153,N_27625);
nor U28348 (N_28348,N_26704,N_27656);
or U28349 (N_28349,N_26043,N_27742);
and U28350 (N_28350,N_26698,N_26917);
or U28351 (N_28351,N_26106,N_27070);
and U28352 (N_28352,N_27697,N_27143);
or U28353 (N_28353,N_26865,N_26960);
and U28354 (N_28354,N_26485,N_27996);
or U28355 (N_28355,N_26108,N_26085);
nand U28356 (N_28356,N_27412,N_26292);
or U28357 (N_28357,N_27615,N_27187);
and U28358 (N_28358,N_26885,N_26636);
or U28359 (N_28359,N_27109,N_27292);
xnor U28360 (N_28360,N_27959,N_26033);
nor U28361 (N_28361,N_26503,N_26042);
nor U28362 (N_28362,N_26014,N_27988);
nor U28363 (N_28363,N_27653,N_27839);
nor U28364 (N_28364,N_26730,N_27978);
nor U28365 (N_28365,N_26348,N_26691);
and U28366 (N_28366,N_26007,N_27526);
and U28367 (N_28367,N_26234,N_26542);
nand U28368 (N_28368,N_26710,N_26000);
nand U28369 (N_28369,N_26941,N_27846);
nand U28370 (N_28370,N_27704,N_27501);
or U28371 (N_28371,N_27137,N_27723);
and U28372 (N_28372,N_26330,N_27741);
nand U28373 (N_28373,N_26979,N_26644);
nand U28374 (N_28374,N_27283,N_27286);
nand U28375 (N_28375,N_26307,N_27421);
and U28376 (N_28376,N_27355,N_26845);
nand U28377 (N_28377,N_26838,N_27165);
xor U28378 (N_28378,N_26665,N_26208);
or U28379 (N_28379,N_26265,N_27810);
or U28380 (N_28380,N_27021,N_26642);
or U28381 (N_28381,N_27852,N_27392);
and U28382 (N_28382,N_27321,N_27639);
nand U28383 (N_28383,N_27771,N_26422);
nand U28384 (N_28384,N_26964,N_27941);
nand U28385 (N_28385,N_26733,N_27886);
and U28386 (N_28386,N_27488,N_27023);
xor U28387 (N_28387,N_27074,N_26421);
and U28388 (N_28388,N_27861,N_27991);
nand U28389 (N_28389,N_26150,N_27202);
or U28390 (N_28390,N_26374,N_27175);
nor U28391 (N_28391,N_27573,N_27043);
or U28392 (N_28392,N_27872,N_26189);
nand U28393 (N_28393,N_26658,N_27735);
nand U28394 (N_28394,N_27566,N_26498);
and U28395 (N_28395,N_26279,N_26345);
or U28396 (N_28396,N_27588,N_27679);
or U28397 (N_28397,N_27844,N_27397);
nor U28398 (N_28398,N_27323,N_27208);
nand U28399 (N_28399,N_26492,N_27777);
xnor U28400 (N_28400,N_26762,N_27275);
nor U28401 (N_28401,N_26576,N_27673);
and U28402 (N_28402,N_27419,N_27454);
or U28403 (N_28403,N_26151,N_27055);
or U28404 (N_28404,N_26081,N_26872);
nand U28405 (N_28405,N_26050,N_26724);
nor U28406 (N_28406,N_27682,N_27466);
and U28407 (N_28407,N_26175,N_27073);
nor U28408 (N_28408,N_27461,N_27916);
and U28409 (N_28409,N_27548,N_26416);
nand U28410 (N_28410,N_26337,N_27822);
nor U28411 (N_28411,N_27801,N_27265);
and U28412 (N_28412,N_27241,N_27535);
and U28413 (N_28413,N_26289,N_26235);
nor U28414 (N_28414,N_26777,N_27556);
or U28415 (N_28415,N_26238,N_27166);
and U28416 (N_28416,N_26737,N_27425);
xnor U28417 (N_28417,N_27891,N_27001);
nor U28418 (N_28418,N_26935,N_27676);
and U28419 (N_28419,N_26604,N_27128);
nand U28420 (N_28420,N_27237,N_27928);
nor U28421 (N_28421,N_26236,N_26400);
nor U28422 (N_28422,N_26112,N_27745);
or U28423 (N_28423,N_27929,N_26590);
and U28424 (N_28424,N_27256,N_27085);
or U28425 (N_28425,N_26866,N_26537);
nor U28426 (N_28426,N_26048,N_26145);
nand U28427 (N_28427,N_27942,N_26232);
and U28428 (N_28428,N_27231,N_26166);
nor U28429 (N_28429,N_27832,N_26561);
nand U28430 (N_28430,N_27407,N_26339);
xnor U28431 (N_28431,N_27317,N_26332);
nand U28432 (N_28432,N_26624,N_27686);
or U28433 (N_28433,N_26721,N_26452);
nor U28434 (N_28434,N_26411,N_26587);
and U28435 (N_28435,N_27692,N_27431);
or U28436 (N_28436,N_26846,N_26005);
or U28437 (N_28437,N_26148,N_26245);
nor U28438 (N_28438,N_27672,N_27551);
nor U28439 (N_28439,N_27475,N_27052);
or U28440 (N_28440,N_26528,N_26873);
nor U28441 (N_28441,N_27097,N_26788);
nor U28442 (N_28442,N_27126,N_26632);
nand U28443 (N_28443,N_27161,N_26441);
or U28444 (N_28444,N_26098,N_27150);
and U28445 (N_28445,N_26094,N_27755);
nor U28446 (N_28446,N_26547,N_26273);
and U28447 (N_28447,N_27075,N_27955);
nand U28448 (N_28448,N_27889,N_27609);
nor U28449 (N_28449,N_26651,N_27377);
nand U28450 (N_28450,N_26327,N_26252);
and U28451 (N_28451,N_27005,N_26734);
nor U28452 (N_28452,N_27510,N_27422);
or U28453 (N_28453,N_27761,N_27482);
nand U28454 (N_28454,N_27279,N_27987);
or U28455 (N_28455,N_27391,N_27428);
or U28456 (N_28456,N_26403,N_26188);
and U28457 (N_28457,N_27099,N_27794);
or U28458 (N_28458,N_27024,N_26609);
xor U28459 (N_28459,N_26296,N_26483);
or U28460 (N_28460,N_27930,N_27100);
nand U28461 (N_28461,N_27400,N_27470);
nor U28462 (N_28462,N_27395,N_26118);
and U28463 (N_28463,N_26832,N_26650);
or U28464 (N_28464,N_27695,N_27031);
or U28465 (N_28465,N_27434,N_27406);
nand U28466 (N_28466,N_27637,N_27847);
nand U28467 (N_28467,N_26313,N_27388);
or U28468 (N_28468,N_27837,N_26051);
nand U28469 (N_28469,N_26791,N_26671);
nand U28470 (N_28470,N_26868,N_26457);
xor U28471 (N_28471,N_26996,N_26548);
or U28472 (N_28472,N_26220,N_27608);
nor U28473 (N_28473,N_26167,N_26191);
nor U28474 (N_28474,N_27236,N_26436);
nand U28475 (N_28475,N_26046,N_26891);
nor U28476 (N_28476,N_26662,N_27331);
and U28477 (N_28477,N_26280,N_26363);
and U28478 (N_28478,N_27947,N_26967);
nand U28479 (N_28479,N_26778,N_26554);
or U28480 (N_28480,N_26518,N_27330);
and U28481 (N_28481,N_26598,N_27107);
nand U28482 (N_28482,N_27026,N_26983);
or U28483 (N_28483,N_26253,N_26668);
nor U28484 (N_28484,N_27173,N_27221);
nor U28485 (N_28485,N_26648,N_26193);
nand U28486 (N_28486,N_26243,N_26531);
and U28487 (N_28487,N_27587,N_26765);
nand U28488 (N_28488,N_26597,N_26371);
nand U28489 (N_28489,N_27130,N_26420);
nor U28490 (N_28490,N_27965,N_26707);
nor U28491 (N_28491,N_26041,N_26516);
or U28492 (N_28492,N_27881,N_26464);
or U28493 (N_28493,N_26982,N_27623);
or U28494 (N_28494,N_27974,N_27308);
nor U28495 (N_28495,N_26814,N_26566);
nand U28496 (N_28496,N_27209,N_26444);
and U28497 (N_28497,N_26586,N_27969);
nand U28498 (N_28498,N_26664,N_26378);
nor U28499 (N_28499,N_26993,N_27142);
xnor U28500 (N_28500,N_27940,N_26794);
nand U28501 (N_28501,N_26006,N_26617);
and U28502 (N_28502,N_26909,N_27047);
and U28503 (N_28503,N_27743,N_26854);
nor U28504 (N_28504,N_26507,N_26434);
or U28505 (N_28505,N_27519,N_26536);
or U28506 (N_28506,N_26410,N_26122);
or U28507 (N_28507,N_27612,N_27367);
nor U28508 (N_28508,N_27095,N_27346);
or U28509 (N_28509,N_26024,N_27449);
nor U28510 (N_28510,N_26388,N_27376);
nor U28511 (N_28511,N_26053,N_27192);
or U28512 (N_28512,N_27878,N_26357);
nor U28513 (N_28513,N_27056,N_26463);
and U28514 (N_28514,N_27848,N_26397);
and U28515 (N_28515,N_26225,N_26916);
nor U28516 (N_28516,N_27119,N_27374);
nand U28517 (N_28517,N_27592,N_26449);
nand U28518 (N_28518,N_27953,N_26850);
or U28519 (N_28519,N_27598,N_26495);
nand U28520 (N_28520,N_27250,N_26984);
nor U28521 (N_28521,N_27144,N_27476);
nand U28522 (N_28522,N_27414,N_26207);
nand U28523 (N_28523,N_26911,N_27002);
and U28524 (N_28524,N_26581,N_27018);
and U28525 (N_28525,N_27880,N_27066);
nor U28526 (N_28526,N_26201,N_26829);
and U28527 (N_28527,N_27458,N_26602);
or U28528 (N_28528,N_26726,N_27989);
nand U28529 (N_28529,N_27858,N_27022);
nor U28530 (N_28530,N_26899,N_26974);
nor U28531 (N_28531,N_26456,N_26377);
nor U28532 (N_28532,N_27567,N_27200);
nand U28533 (N_28533,N_27807,N_26780);
and U28534 (N_28534,N_27347,N_27580);
nand U28535 (N_28535,N_26886,N_26433);
and U28536 (N_28536,N_27787,N_27651);
nor U28537 (N_28537,N_26680,N_26316);
nor U28538 (N_28538,N_26801,N_27230);
or U28539 (N_28539,N_26735,N_26583);
and U28540 (N_28540,N_26615,N_27038);
and U28541 (N_28541,N_27171,N_26772);
nand U28542 (N_28542,N_26874,N_27113);
and U28543 (N_28543,N_27708,N_26380);
nand U28544 (N_28544,N_27660,N_27921);
nor U28545 (N_28545,N_27442,N_27176);
or U28546 (N_28546,N_27576,N_27581);
nor U28547 (N_28547,N_27904,N_26301);
or U28548 (N_28548,N_26324,N_26674);
and U28549 (N_28549,N_26399,N_27617);
nor U28550 (N_28550,N_26501,N_26779);
nand U28551 (N_28551,N_26716,N_27182);
nand U28552 (N_28552,N_27901,N_26806);
or U28553 (N_28553,N_26834,N_26715);
xnor U28554 (N_28554,N_27909,N_26782);
nor U28555 (N_28555,N_27522,N_26152);
nand U28556 (N_28556,N_27764,N_26432);
nand U28557 (N_28557,N_26343,N_26920);
and U28558 (N_28558,N_27986,N_26809);
and U28559 (N_28559,N_27536,N_27725);
nor U28560 (N_28560,N_27253,N_27141);
and U28561 (N_28561,N_26353,N_26049);
or U28562 (N_28562,N_26263,N_27216);
nor U28563 (N_28563,N_27646,N_27353);
and U28564 (N_28564,N_27817,N_26661);
nand U28565 (N_28565,N_26861,N_27892);
nand U28566 (N_28566,N_26800,N_26706);
or U28567 (N_28567,N_26797,N_26270);
nand U28568 (N_28568,N_27739,N_27977);
or U28569 (N_28569,N_27643,N_27905);
and U28570 (N_28570,N_27154,N_26946);
nor U28571 (N_28571,N_27765,N_26251);
and U28572 (N_28572,N_26593,N_26654);
and U28573 (N_28573,N_26975,N_26487);
nor U28574 (N_28574,N_26768,N_27854);
and U28575 (N_28575,N_26093,N_26694);
or U28576 (N_28576,N_26893,N_27779);
or U28577 (N_28577,N_26559,N_26740);
nand U28578 (N_28578,N_26021,N_26843);
or U28579 (N_28579,N_27640,N_27514);
nand U28580 (N_28580,N_27722,N_26372);
nor U28581 (N_28581,N_26810,N_26858);
nand U28582 (N_28582,N_26775,N_26453);
and U28583 (N_28583,N_27287,N_26473);
nor U28584 (N_28584,N_26558,N_26022);
and U28585 (N_28585,N_26943,N_27170);
nand U28586 (N_28586,N_27179,N_26538);
or U28587 (N_28587,N_26158,N_27750);
and U28588 (N_28588,N_27271,N_26677);
nand U28589 (N_28589,N_27620,N_27618);
and U28590 (N_28590,N_27726,N_26628);
nor U28591 (N_28591,N_27274,N_26529);
and U28592 (N_28592,N_26882,N_27719);
nand U28593 (N_28593,N_27079,N_27198);
or U28594 (N_28594,N_26584,N_26352);
nand U28595 (N_28595,N_27490,N_26367);
and U28596 (N_28596,N_27255,N_27507);
and U28597 (N_28597,N_26249,N_27034);
nor U28598 (N_28598,N_26718,N_27096);
and U28599 (N_28599,N_27919,N_27094);
and U28600 (N_28600,N_26783,N_26223);
nand U28601 (N_28601,N_26351,N_27496);
nand U28602 (N_28602,N_27403,N_26640);
and U28603 (N_28603,N_27751,N_27530);
or U28604 (N_28604,N_26913,N_26900);
nor U28605 (N_28605,N_27471,N_27139);
nand U28606 (N_28606,N_27147,N_27527);
and U28607 (N_28607,N_26471,N_27409);
nand U28608 (N_28608,N_26819,N_26443);
and U28609 (N_28609,N_27770,N_26746);
or U28610 (N_28610,N_27037,N_27756);
and U28611 (N_28611,N_26610,N_26805);
nor U28612 (N_28612,N_26355,N_26986);
and U28613 (N_28613,N_26599,N_26237);
nor U28614 (N_28614,N_26120,N_26425);
nand U28615 (N_28615,N_27845,N_26078);
nand U28616 (N_28616,N_27172,N_26034);
or U28617 (N_28617,N_27502,N_26278);
nor U28618 (N_28618,N_27542,N_26928);
or U28619 (N_28619,N_27305,N_26202);
or U28620 (N_28620,N_26239,N_27678);
nand U28621 (N_28621,N_26614,N_26258);
or U28622 (N_28622,N_26719,N_27118);
nand U28623 (N_28623,N_26359,N_27325);
xnor U28624 (N_28624,N_26563,N_27648);
and U28625 (N_28625,N_27312,N_26179);
nand U28626 (N_28626,N_26637,N_27604);
or U28627 (N_28627,N_27759,N_27629);
nand U28628 (N_28628,N_27829,N_27926);
xor U28629 (N_28629,N_26625,N_26073);
nand U28630 (N_28630,N_26125,N_27222);
and U28631 (N_28631,N_27632,N_27480);
and U28632 (N_28632,N_26310,N_26875);
or U28633 (N_28633,N_27819,N_27245);
nand U28634 (N_28634,N_27570,N_27945);
and U28635 (N_28635,N_27474,N_26567);
and U28636 (N_28636,N_27242,N_26381);
and U28637 (N_28637,N_26105,N_27058);
and U28638 (N_28638,N_26266,N_27958);
nand U28639 (N_28639,N_26759,N_26029);
nor U28640 (N_28640,N_26534,N_26446);
nand U28641 (N_28641,N_26676,N_27016);
nand U28642 (N_28642,N_26387,N_27724);
nor U28643 (N_28643,N_26860,N_26709);
nand U28644 (N_28644,N_26685,N_27280);
nor U28645 (N_28645,N_26376,N_26760);
nand U28646 (N_28646,N_27105,N_27162);
nand U28647 (N_28647,N_26688,N_26835);
nand U28648 (N_28648,N_27004,N_27645);
nand U28649 (N_28649,N_26549,N_26019);
xor U28650 (N_28650,N_26647,N_26293);
or U28651 (N_28651,N_26058,N_26491);
nor U28652 (N_28652,N_26500,N_27533);
and U28653 (N_28653,N_27658,N_27516);
nand U28654 (N_28654,N_27795,N_26795);
nand U28655 (N_28655,N_26825,N_27521);
nand U28656 (N_28656,N_27234,N_27896);
nand U28657 (N_28657,N_26940,N_26214);
and U28658 (N_28658,N_27911,N_27851);
or U28659 (N_28659,N_26375,N_26564);
nor U28660 (N_28660,N_27657,N_27320);
and U28661 (N_28661,N_27555,N_26095);
or U28662 (N_28662,N_26521,N_27334);
nand U28663 (N_28663,N_27993,N_26437);
xnor U28664 (N_28664,N_26336,N_27705);
nor U28665 (N_28665,N_27873,N_27116);
nor U28666 (N_28666,N_27069,N_27336);
nand U28667 (N_28667,N_27483,N_27871);
nand U28668 (N_28668,N_26156,N_26406);
xnor U28669 (N_28669,N_26287,N_26961);
and U28670 (N_28670,N_27416,N_27472);
nand U28671 (N_28671,N_27681,N_26090);
nor U28672 (N_28672,N_27451,N_27825);
nand U28673 (N_28673,N_27797,N_27963);
nor U28674 (N_28674,N_27296,N_27383);
nand U28675 (N_28675,N_26100,N_27912);
nor U28676 (N_28676,N_27796,N_26763);
or U28677 (N_28677,N_26828,N_26185);
nand U28678 (N_28678,N_27189,N_26414);
nor U28679 (N_28679,N_26701,N_26025);
nor U28680 (N_28680,N_26139,N_27398);
and U28681 (N_28681,N_27733,N_26469);
nor U28682 (N_28682,N_26519,N_27758);
xor U28683 (N_28683,N_26001,N_27767);
nand U28684 (N_28684,N_26511,N_27802);
nand U28685 (N_28685,N_26391,N_26137);
or U28686 (N_28686,N_26793,N_27593);
xnor U28687 (N_28687,N_26362,N_27616);
and U28688 (N_28688,N_27138,N_27359);
and U28689 (N_28689,N_27578,N_27302);
nand U28690 (N_28690,N_27524,N_27950);
xor U28691 (N_28691,N_26550,N_27186);
nor U28692 (N_28692,N_26789,N_26942);
nand U28693 (N_28693,N_27805,N_27738);
nor U28694 (N_28694,N_27413,N_26660);
and U28695 (N_28695,N_26059,N_27949);
and U28696 (N_28696,N_27550,N_27495);
nand U28697 (N_28697,N_26731,N_27062);
or U28698 (N_28698,N_26877,N_26933);
nand U28699 (N_28699,N_27983,N_26064);
nand U28700 (N_28700,N_27188,N_26163);
and U28701 (N_28701,N_26807,N_27776);
or U28702 (N_28702,N_26774,N_26656);
nor U28703 (N_28703,N_26052,N_26180);
nor U28704 (N_28704,N_26032,N_27677);
xnor U28705 (N_28705,N_27219,N_26921);
nand U28706 (N_28706,N_27961,N_26639);
and U28707 (N_28707,N_26723,N_26932);
nand U28708 (N_28708,N_26959,N_27812);
and U28709 (N_28709,N_27087,N_26451);
nand U28710 (N_28710,N_26264,N_27155);
nand U28711 (N_28711,N_27622,N_26601);
nand U28712 (N_28712,N_26696,N_26944);
and U28713 (N_28713,N_26066,N_27014);
nand U28714 (N_28714,N_26836,N_27051);
nor U28715 (N_28715,N_26824,N_27328);
nor U28716 (N_28716,N_26040,N_26764);
nand U28717 (N_28717,N_27915,N_26121);
nand U28718 (N_28718,N_26200,N_27426);
or U28719 (N_28719,N_27859,N_27747);
or U28720 (N_28720,N_27564,N_27164);
and U28721 (N_28721,N_27789,N_27084);
or U28722 (N_28722,N_26227,N_27351);
or U28723 (N_28723,N_26513,N_26070);
and U28724 (N_28724,N_27882,N_26776);
or U28725 (N_28725,N_27083,N_27559);
and U28726 (N_28726,N_26822,N_27380);
nor U28727 (N_28727,N_26104,N_27485);
xnor U28728 (N_28728,N_27125,N_26520);
nor U28729 (N_28729,N_26082,N_27054);
nand U28730 (N_28730,N_27238,N_27124);
nand U28731 (N_28731,N_26728,N_26894);
and U28732 (N_28732,N_26315,N_27446);
and U28733 (N_28733,N_27634,N_27010);
nand U28734 (N_28734,N_26195,N_27525);
nand U28735 (N_28735,N_27064,N_26130);
or U28736 (N_28736,N_26792,N_26143);
nand U28737 (N_28737,N_27997,N_27205);
nand U28738 (N_28738,N_26883,N_26973);
nand U28739 (N_28739,N_27065,N_27214);
nand U28740 (N_28740,N_26761,N_26164);
or U28741 (N_28741,N_26311,N_27613);
or U28742 (N_28742,N_27990,N_27178);
or U28743 (N_28743,N_26753,N_27191);
and U28744 (N_28744,N_26881,N_27757);
nor U28745 (N_28745,N_27288,N_27102);
and U28746 (N_28746,N_26512,N_26401);
nand U28747 (N_28747,N_26966,N_27668);
nor U28748 (N_28748,N_26408,N_27410);
or U28749 (N_28749,N_26011,N_26784);
nand U28750 (N_28750,N_26368,N_26174);
nor U28751 (N_28751,N_26532,N_26255);
nand U28752 (N_28752,N_27389,N_27453);
nor U28753 (N_28753,N_26241,N_27760);
nand U28754 (N_28754,N_27898,N_27443);
nand U28755 (N_28755,N_26103,N_26435);
or U28756 (N_28756,N_26415,N_26221);
nand U28757 (N_28757,N_27215,N_26482);
and U28758 (N_28758,N_27605,N_26947);
and U28759 (N_28759,N_27999,N_26657);
nor U28760 (N_28760,N_26557,N_26092);
or U28761 (N_28761,N_26089,N_26945);
nand U28762 (N_28762,N_27994,N_26649);
and U28763 (N_28763,N_27120,N_27285);
or U28764 (N_28764,N_27599,N_26488);
and U28765 (N_28765,N_26998,N_27938);
or U28766 (N_28766,N_27748,N_27298);
nor U28767 (N_28767,N_27565,N_27111);
or U28768 (N_28768,N_26326,N_27841);
nand U28769 (N_28769,N_27561,N_26497);
and U28770 (N_28770,N_27630,N_27091);
and U28771 (N_28771,N_26562,N_27159);
or U28772 (N_28772,N_26655,N_27849);
nand U28773 (N_28773,N_27149,N_26099);
nand U28774 (N_28774,N_27769,N_27571);
nand U28775 (N_28775,N_26285,N_26465);
nor U28776 (N_28776,N_26905,N_27467);
or U28777 (N_28777,N_27169,N_26755);
and U28778 (N_28778,N_27033,N_26364);
or U28779 (N_28779,N_27920,N_26620);
or U28780 (N_28780,N_26522,N_26880);
and U28781 (N_28781,N_26088,N_26268);
or U28782 (N_28782,N_26178,N_26767);
or U28783 (N_28783,N_27385,N_26328);
nor U28784 (N_28784,N_26257,N_27239);
nand U28785 (N_28785,N_27917,N_27456);
nand U28786 (N_28786,N_26218,N_27465);
nor U28787 (N_28787,N_27180,N_26405);
nand U28788 (N_28788,N_26552,N_27289);
nor U28789 (N_28789,N_26844,N_27957);
nor U28790 (N_28790,N_27122,N_27310);
nand U28791 (N_28791,N_26569,N_26086);
xnor U28792 (N_28792,N_26962,N_27224);
xor U28793 (N_28793,N_27894,N_27712);
nand U28794 (N_28794,N_27934,N_27944);
or U28795 (N_28795,N_26224,N_27577);
or U28796 (N_28796,N_26743,N_27867);
nor U28797 (N_28797,N_26205,N_27368);
and U28798 (N_28798,N_27960,N_26675);
nand U28799 (N_28799,N_27129,N_26134);
nor U28800 (N_28800,N_26354,N_27227);
nand U28801 (N_28801,N_26459,N_26749);
or U28802 (N_28802,N_27277,N_26442);
or U28803 (N_28803,N_27028,N_27146);
or U28804 (N_28804,N_27500,N_27303);
nor U28805 (N_28805,N_26197,N_26702);
and U28806 (N_28806,N_26004,N_27666);
nand U28807 (N_28807,N_27132,N_26460);
nor U28808 (N_28808,N_26939,N_26084);
and U28809 (N_28809,N_27226,N_26141);
and U28810 (N_28810,N_27117,N_26670);
and U28811 (N_28811,N_26808,N_26852);
or U28812 (N_28812,N_26653,N_27784);
and U28813 (N_28813,N_26526,N_27768);
nand U28814 (N_28814,N_27183,N_27943);
nor U28815 (N_28815,N_27498,N_27827);
and U28816 (N_28816,N_26578,N_27883);
or U28817 (N_28817,N_27908,N_26102);
and U28818 (N_28818,N_26149,N_26335);
nor U28819 (N_28819,N_26262,N_27523);
or U28820 (N_28820,N_27586,N_27402);
and U28821 (N_28821,N_26727,N_26008);
nand U28822 (N_28822,N_26009,N_27707);
or U28823 (N_28823,N_27671,N_26077);
or U28824 (N_28824,N_27257,N_26985);
nor U28825 (N_28825,N_27984,N_27820);
or U28826 (N_28826,N_27528,N_27992);
xnor U28827 (N_28827,N_26864,N_26065);
nand U28828 (N_28828,N_26556,N_27092);
or U28829 (N_28829,N_27814,N_26769);
and U28830 (N_28830,N_27217,N_27020);
or U28831 (N_28831,N_27044,N_26859);
or U28832 (N_28832,N_27233,N_26560);
nor U28833 (N_28833,N_27619,N_27327);
or U28834 (N_28834,N_27373,N_27884);
and U28835 (N_28835,N_27371,N_26466);
nor U28836 (N_28836,N_26907,N_27225);
or U28837 (N_28837,N_27437,N_27663);
or U28838 (N_28838,N_26071,N_26194);
or U28839 (N_28839,N_26659,N_26015);
or U28840 (N_28840,N_26611,N_27914);
nor U28841 (N_28841,N_27806,N_27324);
nor U28842 (N_28842,N_27684,N_27106);
nor U28843 (N_28843,N_27621,N_26018);
nor U28844 (N_28844,N_27927,N_27762);
and U28845 (N_28845,N_27196,N_26281);
or U28846 (N_28846,N_26306,N_27628);
nor U28847 (N_28847,N_26295,N_27752);
and U28848 (N_28848,N_26771,N_27669);
or U28849 (N_28849,N_26091,N_27602);
and U28850 (N_28850,N_26729,N_27823);
nand U28851 (N_28851,N_26851,N_27345);
nand U28852 (N_28852,N_26248,N_27067);
nor U28853 (N_28853,N_27691,N_26417);
nand U28854 (N_28854,N_26977,N_26358);
or U28855 (N_28855,N_26976,N_26509);
or U28856 (N_28856,N_26062,N_27203);
or U28857 (N_28857,N_27342,N_27479);
or U28858 (N_28858,N_27360,N_27088);
and U28859 (N_28859,N_26458,N_27610);
nand U28860 (N_28860,N_26510,N_27417);
and U28861 (N_28861,N_27766,N_27966);
nor U28862 (N_28862,N_27893,N_26673);
nor U28863 (N_28863,N_27826,N_26687);
or U28864 (N_28864,N_27711,N_27145);
nor U28865 (N_28865,N_27061,N_27134);
nand U28866 (N_28866,N_26629,N_26395);
nand U28867 (N_28867,N_27842,N_27251);
or U28868 (N_28868,N_26700,N_26818);
or U28869 (N_28869,N_27862,N_26382);
and U28870 (N_28870,N_27393,N_26455);
nor U28871 (N_28871,N_26370,N_26934);
nand U28872 (N_28872,N_26115,N_26863);
nor U28873 (N_28873,N_27011,N_26484);
nand U28874 (N_28874,N_27890,N_26686);
nor U28875 (N_28875,N_27590,N_27415);
nand U28876 (N_28876,N_26955,N_26304);
nor U28877 (N_28877,N_27435,N_26695);
nand U28878 (N_28878,N_26260,N_27152);
or U28879 (N_28879,N_26107,N_26448);
nand U28880 (N_28880,N_26275,N_27148);
nand U28881 (N_28881,N_27503,N_27429);
nor U28882 (N_28882,N_27045,N_27968);
nor U28883 (N_28883,N_26757,N_27980);
or U28884 (N_28884,N_26419,N_26869);
nor U28885 (N_28885,N_27924,N_26524);
and U28886 (N_28886,N_27749,N_26573);
or U28887 (N_28887,N_26423,N_27318);
or U28888 (N_28888,N_26325,N_27702);
or U28889 (N_28889,N_26950,N_27261);
and U28890 (N_28890,N_27792,N_26936);
nand U28891 (N_28891,N_26555,N_27773);
or U28892 (N_28892,N_27836,N_26958);
or U28893 (N_28893,N_27201,N_26116);
nor U28894 (N_28894,N_26938,N_27865);
and U28895 (N_28895,N_27952,N_26890);
and U28896 (N_28896,N_26284,N_27574);
xnor U28897 (N_28897,N_27006,N_26663);
nand U28898 (N_28898,N_26796,N_27293);
or U28899 (N_28899,N_27790,N_26517);
nand U28900 (N_28900,N_26170,N_27838);
or U28901 (N_28901,N_27235,N_26951);
or U28902 (N_28902,N_27270,N_27659);
and U28903 (N_28903,N_27687,N_26752);
nand U28904 (N_28904,N_27167,N_27600);
nand U28905 (N_28905,N_26154,N_26020);
nand U28906 (N_28906,N_27981,N_27866);
nor U28907 (N_28907,N_26575,N_26132);
and U28908 (N_28908,N_27244,N_26745);
or U28909 (N_28909,N_26816,N_27041);
nand U28910 (N_28910,N_26135,N_26595);
or U28911 (N_28911,N_26186,N_26409);
or U28912 (N_28912,N_26630,N_27557);
nand U28913 (N_28913,N_26454,N_26821);
or U28914 (N_28914,N_27775,N_27445);
nor U28915 (N_28915,N_27778,N_27786);
or U28916 (N_28916,N_26113,N_26383);
and U28917 (N_28917,N_27644,N_26438);
or U28918 (N_28918,N_27027,N_26047);
or U28919 (N_28919,N_26203,N_26857);
or U28920 (N_28920,N_27015,N_26244);
nor U28921 (N_28921,N_26799,N_26888);
or U28922 (N_28922,N_27772,N_26570);
nand U28923 (N_28923,N_27874,N_26887);
or U28924 (N_28924,N_27869,N_27693);
and U28925 (N_28925,N_27019,N_27168);
nor U28926 (N_28926,N_26346,N_26703);
nand U28927 (N_28927,N_27319,N_27068);
nor U28928 (N_28928,N_27804,N_27964);
and U28929 (N_28929,N_27583,N_27163);
nand U28930 (N_28930,N_26477,N_26192);
or U28931 (N_28931,N_27652,N_27982);
or U28932 (N_28932,N_27151,N_27493);
or U28933 (N_28933,N_27782,N_26957);
or U28934 (N_28934,N_27314,N_26286);
nor U28935 (N_28935,N_26646,N_26317);
or U28936 (N_28936,N_27547,N_26910);
or U28937 (N_28937,N_26505,N_26061);
nand U28938 (N_28938,N_26901,N_26216);
nor U28939 (N_28939,N_26506,N_27906);
and U28940 (N_28940,N_26750,N_26533);
and U28941 (N_28941,N_27008,N_26398);
nand U28942 (N_28942,N_26582,N_27013);
or U28943 (N_28943,N_27754,N_27411);
nor U28944 (N_28944,N_27133,N_27783);
or U28945 (N_28945,N_27595,N_27511);
or U28946 (N_28946,N_26802,N_27907);
and U28947 (N_28947,N_27499,N_27185);
nor U28948 (N_28948,N_27553,N_27868);
nor U28949 (N_28949,N_26184,N_27381);
and U28950 (N_28950,N_26684,N_27544);
nand U28951 (N_28951,N_27206,N_27813);
and U28952 (N_28952,N_27098,N_26543);
nor U28953 (N_28953,N_27080,N_27855);
or U28954 (N_28954,N_26038,N_27204);
or U28955 (N_28955,N_27487,N_26577);
or U28956 (N_28956,N_27562,N_27354);
and U28957 (N_28957,N_26127,N_27379);
and U28958 (N_28958,N_27662,N_26571);
or U28959 (N_28959,N_27902,N_26331);
nor U28960 (N_28960,N_26063,N_26183);
nor U28961 (N_28961,N_26035,N_26878);
and U28962 (N_28962,N_27459,N_27072);
nor U28963 (N_28963,N_26161,N_27438);
or U28964 (N_28964,N_27661,N_26812);
nor U28965 (N_28965,N_26480,N_26902);
nand U28966 (N_28966,N_27857,N_27436);
nand U28967 (N_28967,N_26430,N_27683);
nor U28968 (N_28968,N_27633,N_27384);
or U28969 (N_28969,N_26269,N_26271);
or U28970 (N_28970,N_26589,N_27489);
nand U28971 (N_28971,N_27378,N_26494);
nor U28972 (N_28972,N_27300,N_26302);
and U28973 (N_28973,N_27267,N_26606);
nor U28974 (N_28974,N_26862,N_26892);
or U28975 (N_28975,N_27093,N_26683);
or U28976 (N_28976,N_26699,N_27834);
nor U28977 (N_28977,N_27895,N_26233);
xor U28978 (N_28978,N_26988,N_26424);
or U28979 (N_28979,N_27177,N_27036);
or U28980 (N_28980,N_26525,N_27569);
and U28981 (N_28981,N_26605,N_26817);
and U28982 (N_28982,N_26948,N_26003);
and U28983 (N_28983,N_27840,N_27939);
nor U28984 (N_28984,N_26908,N_27698);
or U28985 (N_28985,N_27875,N_27636);
nor U28986 (N_28986,N_26635,N_26923);
and U28987 (N_28987,N_27717,N_27913);
or U28988 (N_28988,N_26247,N_27667);
or U28989 (N_28989,N_27440,N_26054);
nor U28990 (N_28990,N_26298,N_27387);
nor U28991 (N_28991,N_26927,N_26274);
nand U28992 (N_28992,N_27333,N_26811);
xnor U28993 (N_28993,N_27337,N_27369);
nor U28994 (N_28994,N_27831,N_26804);
nand U28995 (N_28995,N_27160,N_26261);
nand U28996 (N_28996,N_27568,N_26323);
nor U28997 (N_28997,N_27492,N_26333);
nand U28998 (N_28998,N_27115,N_27348);
or U28999 (N_28999,N_27885,N_27689);
nor U29000 (N_29000,N_27267,N_27234);
nor U29001 (N_29001,N_26994,N_27320);
and U29002 (N_29002,N_27932,N_26342);
nor U29003 (N_29003,N_26475,N_26760);
nand U29004 (N_29004,N_27233,N_26437);
or U29005 (N_29005,N_27004,N_26213);
xnor U29006 (N_29006,N_27624,N_27251);
nor U29007 (N_29007,N_27581,N_27975);
nor U29008 (N_29008,N_26726,N_26713);
or U29009 (N_29009,N_27641,N_27163);
nand U29010 (N_29010,N_27476,N_27004);
nand U29011 (N_29011,N_27350,N_26197);
and U29012 (N_29012,N_26475,N_27147);
or U29013 (N_29013,N_26072,N_26209);
xor U29014 (N_29014,N_26951,N_26503);
nor U29015 (N_29015,N_26092,N_26515);
nand U29016 (N_29016,N_26001,N_27204);
and U29017 (N_29017,N_26562,N_26792);
and U29018 (N_29018,N_27127,N_27542);
or U29019 (N_29019,N_27934,N_27196);
or U29020 (N_29020,N_27045,N_27516);
or U29021 (N_29021,N_26213,N_26569);
and U29022 (N_29022,N_26274,N_26177);
and U29023 (N_29023,N_26734,N_26263);
nand U29024 (N_29024,N_27720,N_27964);
and U29025 (N_29025,N_26057,N_27900);
nand U29026 (N_29026,N_27901,N_27298);
and U29027 (N_29027,N_27459,N_26996);
and U29028 (N_29028,N_26968,N_27282);
and U29029 (N_29029,N_26648,N_26849);
and U29030 (N_29030,N_26255,N_27690);
or U29031 (N_29031,N_26432,N_27717);
nand U29032 (N_29032,N_26335,N_26022);
and U29033 (N_29033,N_27086,N_26011);
nand U29034 (N_29034,N_26001,N_26033);
or U29035 (N_29035,N_26853,N_26119);
or U29036 (N_29036,N_27632,N_27453);
nor U29037 (N_29037,N_27512,N_26875);
or U29038 (N_29038,N_27805,N_26553);
and U29039 (N_29039,N_26205,N_27656);
or U29040 (N_29040,N_26295,N_26857);
or U29041 (N_29041,N_26944,N_27276);
nand U29042 (N_29042,N_27941,N_27421);
or U29043 (N_29043,N_26520,N_26228);
and U29044 (N_29044,N_27782,N_27145);
nor U29045 (N_29045,N_26302,N_27244);
nand U29046 (N_29046,N_27350,N_27676);
and U29047 (N_29047,N_27288,N_27976);
and U29048 (N_29048,N_27804,N_27033);
and U29049 (N_29049,N_26997,N_27945);
and U29050 (N_29050,N_26673,N_27422);
or U29051 (N_29051,N_26144,N_26320);
or U29052 (N_29052,N_27707,N_26793);
or U29053 (N_29053,N_27026,N_27567);
and U29054 (N_29054,N_27450,N_26169);
and U29055 (N_29055,N_26481,N_26493);
or U29056 (N_29056,N_27728,N_26484);
nor U29057 (N_29057,N_26435,N_26351);
and U29058 (N_29058,N_27335,N_26683);
and U29059 (N_29059,N_27825,N_26964);
nor U29060 (N_29060,N_27267,N_26276);
nand U29061 (N_29061,N_26929,N_27238);
and U29062 (N_29062,N_27385,N_26476);
xor U29063 (N_29063,N_27338,N_27083);
nor U29064 (N_29064,N_27750,N_27973);
nand U29065 (N_29065,N_26827,N_26372);
or U29066 (N_29066,N_27339,N_27291);
nand U29067 (N_29067,N_27888,N_27691);
or U29068 (N_29068,N_26215,N_27446);
and U29069 (N_29069,N_26691,N_27110);
and U29070 (N_29070,N_27407,N_27005);
and U29071 (N_29071,N_27060,N_27555);
nor U29072 (N_29072,N_27615,N_27607);
nor U29073 (N_29073,N_27385,N_26647);
nand U29074 (N_29074,N_27131,N_26562);
nor U29075 (N_29075,N_27990,N_26497);
and U29076 (N_29076,N_27650,N_26825);
nor U29077 (N_29077,N_27207,N_26301);
or U29078 (N_29078,N_27922,N_27257);
nor U29079 (N_29079,N_26197,N_27232);
and U29080 (N_29080,N_27472,N_27687);
and U29081 (N_29081,N_26642,N_27889);
and U29082 (N_29082,N_26564,N_26710);
nand U29083 (N_29083,N_26228,N_26213);
and U29084 (N_29084,N_26281,N_27280);
nor U29085 (N_29085,N_27001,N_26680);
and U29086 (N_29086,N_27624,N_26137);
nand U29087 (N_29087,N_26781,N_27631);
nor U29088 (N_29088,N_26282,N_26065);
and U29089 (N_29089,N_27258,N_26090);
nand U29090 (N_29090,N_26153,N_26425);
and U29091 (N_29091,N_27021,N_27507);
nor U29092 (N_29092,N_26611,N_26731);
and U29093 (N_29093,N_26202,N_26560);
nor U29094 (N_29094,N_27651,N_27756);
nor U29095 (N_29095,N_27800,N_26263);
and U29096 (N_29096,N_27642,N_27708);
and U29097 (N_29097,N_26475,N_26400);
nand U29098 (N_29098,N_26429,N_26018);
and U29099 (N_29099,N_27455,N_26904);
nand U29100 (N_29100,N_26925,N_27803);
nand U29101 (N_29101,N_27772,N_27521);
or U29102 (N_29102,N_27489,N_26102);
and U29103 (N_29103,N_26201,N_26968);
or U29104 (N_29104,N_26324,N_26771);
nor U29105 (N_29105,N_27712,N_26718);
or U29106 (N_29106,N_26382,N_26190);
or U29107 (N_29107,N_27971,N_27201);
and U29108 (N_29108,N_27780,N_26997);
or U29109 (N_29109,N_27572,N_27720);
nor U29110 (N_29110,N_27117,N_26904);
nand U29111 (N_29111,N_27915,N_26291);
or U29112 (N_29112,N_26897,N_27522);
nand U29113 (N_29113,N_27909,N_26934);
nand U29114 (N_29114,N_27595,N_27604);
or U29115 (N_29115,N_26418,N_27774);
and U29116 (N_29116,N_27830,N_27610);
and U29117 (N_29117,N_26846,N_27306);
nand U29118 (N_29118,N_26042,N_27683);
or U29119 (N_29119,N_26129,N_27378);
nor U29120 (N_29120,N_27454,N_26393);
and U29121 (N_29121,N_27098,N_27339);
nor U29122 (N_29122,N_26195,N_27463);
nor U29123 (N_29123,N_26171,N_26153);
nor U29124 (N_29124,N_26566,N_26955);
or U29125 (N_29125,N_26535,N_26729);
nor U29126 (N_29126,N_27693,N_26959);
and U29127 (N_29127,N_27058,N_27606);
nand U29128 (N_29128,N_26331,N_26252);
and U29129 (N_29129,N_27432,N_27653);
nand U29130 (N_29130,N_26379,N_26767);
xor U29131 (N_29131,N_26692,N_27948);
or U29132 (N_29132,N_26986,N_27834);
and U29133 (N_29133,N_27276,N_26130);
or U29134 (N_29134,N_27455,N_26333);
or U29135 (N_29135,N_26562,N_26016);
and U29136 (N_29136,N_26406,N_27309);
or U29137 (N_29137,N_26226,N_27250);
nand U29138 (N_29138,N_27896,N_27641);
and U29139 (N_29139,N_27767,N_26882);
nand U29140 (N_29140,N_26673,N_26066);
nand U29141 (N_29141,N_27126,N_27105);
nor U29142 (N_29142,N_26648,N_26679);
nor U29143 (N_29143,N_26025,N_27492);
nand U29144 (N_29144,N_27115,N_26356);
nand U29145 (N_29145,N_27806,N_27914);
or U29146 (N_29146,N_26705,N_26640);
nand U29147 (N_29147,N_27322,N_26522);
nand U29148 (N_29148,N_27720,N_26423);
or U29149 (N_29149,N_26365,N_26771);
nor U29150 (N_29150,N_27933,N_27821);
nor U29151 (N_29151,N_27914,N_27823);
nand U29152 (N_29152,N_27171,N_27711);
and U29153 (N_29153,N_27058,N_26461);
and U29154 (N_29154,N_26129,N_27863);
nor U29155 (N_29155,N_27504,N_27860);
nor U29156 (N_29156,N_27583,N_26448);
nor U29157 (N_29157,N_27868,N_26131);
or U29158 (N_29158,N_27926,N_26972);
or U29159 (N_29159,N_26005,N_27711);
nor U29160 (N_29160,N_27444,N_27966);
nor U29161 (N_29161,N_26255,N_26433);
nand U29162 (N_29162,N_26859,N_27791);
nor U29163 (N_29163,N_27298,N_26310);
nor U29164 (N_29164,N_27043,N_27858);
nand U29165 (N_29165,N_26077,N_26963);
or U29166 (N_29166,N_27792,N_26100);
and U29167 (N_29167,N_27720,N_26639);
or U29168 (N_29168,N_27290,N_26431);
or U29169 (N_29169,N_27595,N_27519);
and U29170 (N_29170,N_26842,N_26933);
nor U29171 (N_29171,N_26718,N_26833);
and U29172 (N_29172,N_26883,N_26304);
nor U29173 (N_29173,N_26654,N_27729);
nor U29174 (N_29174,N_26914,N_27005);
and U29175 (N_29175,N_27789,N_26484);
or U29176 (N_29176,N_27064,N_26185);
nor U29177 (N_29177,N_26640,N_27273);
nand U29178 (N_29178,N_27034,N_26861);
or U29179 (N_29179,N_27716,N_27730);
nor U29180 (N_29180,N_27410,N_26608);
nand U29181 (N_29181,N_27764,N_26228);
or U29182 (N_29182,N_27817,N_26586);
nand U29183 (N_29183,N_27900,N_27608);
nand U29184 (N_29184,N_27895,N_27487);
nand U29185 (N_29185,N_26585,N_26293);
nand U29186 (N_29186,N_26326,N_27005);
and U29187 (N_29187,N_27849,N_26453);
nor U29188 (N_29188,N_27489,N_26057);
and U29189 (N_29189,N_27042,N_27657);
and U29190 (N_29190,N_27966,N_26020);
nand U29191 (N_29191,N_26672,N_26481);
nand U29192 (N_29192,N_26177,N_26808);
and U29193 (N_29193,N_26550,N_27986);
or U29194 (N_29194,N_26889,N_26625);
nand U29195 (N_29195,N_26550,N_27934);
or U29196 (N_29196,N_27252,N_27008);
and U29197 (N_29197,N_26163,N_26766);
nand U29198 (N_29198,N_27066,N_26326);
or U29199 (N_29199,N_26142,N_26940);
nor U29200 (N_29200,N_27371,N_27770);
nand U29201 (N_29201,N_27911,N_27105);
or U29202 (N_29202,N_26374,N_26711);
xnor U29203 (N_29203,N_26004,N_27013);
or U29204 (N_29204,N_27372,N_26431);
nor U29205 (N_29205,N_26529,N_26114);
and U29206 (N_29206,N_27932,N_26942);
nand U29207 (N_29207,N_26339,N_26415);
or U29208 (N_29208,N_27691,N_27138);
nand U29209 (N_29209,N_27758,N_27943);
nand U29210 (N_29210,N_26631,N_26598);
nand U29211 (N_29211,N_26764,N_27189);
or U29212 (N_29212,N_27809,N_26666);
and U29213 (N_29213,N_26548,N_27799);
and U29214 (N_29214,N_27116,N_26280);
and U29215 (N_29215,N_27450,N_27024);
nand U29216 (N_29216,N_27818,N_26668);
nor U29217 (N_29217,N_26683,N_26793);
or U29218 (N_29218,N_27406,N_27693);
and U29219 (N_29219,N_27900,N_27341);
and U29220 (N_29220,N_27486,N_27735);
nand U29221 (N_29221,N_27410,N_27791);
or U29222 (N_29222,N_27656,N_27966);
or U29223 (N_29223,N_27798,N_27524);
and U29224 (N_29224,N_26305,N_27913);
xor U29225 (N_29225,N_26783,N_27544);
or U29226 (N_29226,N_27227,N_27642);
or U29227 (N_29227,N_26805,N_26695);
and U29228 (N_29228,N_26543,N_27192);
and U29229 (N_29229,N_27526,N_27244);
and U29230 (N_29230,N_27721,N_26167);
xor U29231 (N_29231,N_27489,N_27073);
and U29232 (N_29232,N_27615,N_26389);
or U29233 (N_29233,N_26909,N_27115);
and U29234 (N_29234,N_27094,N_27051);
xor U29235 (N_29235,N_26061,N_27904);
or U29236 (N_29236,N_27831,N_27519);
nand U29237 (N_29237,N_26835,N_27859);
nand U29238 (N_29238,N_26365,N_27059);
nor U29239 (N_29239,N_26546,N_27280);
nor U29240 (N_29240,N_26752,N_27849);
nor U29241 (N_29241,N_27333,N_27894);
and U29242 (N_29242,N_26226,N_26865);
nand U29243 (N_29243,N_26697,N_26954);
nor U29244 (N_29244,N_27131,N_27566);
or U29245 (N_29245,N_26878,N_26078);
nor U29246 (N_29246,N_27762,N_27358);
nor U29247 (N_29247,N_27234,N_27313);
nand U29248 (N_29248,N_26606,N_27989);
nor U29249 (N_29249,N_27095,N_26315);
nor U29250 (N_29250,N_26008,N_27218);
and U29251 (N_29251,N_26629,N_27919);
and U29252 (N_29252,N_27249,N_26645);
or U29253 (N_29253,N_27785,N_27909);
and U29254 (N_29254,N_27097,N_26755);
or U29255 (N_29255,N_27014,N_27796);
and U29256 (N_29256,N_27547,N_27366);
nand U29257 (N_29257,N_27236,N_27899);
nor U29258 (N_29258,N_26667,N_27450);
or U29259 (N_29259,N_27566,N_26628);
nor U29260 (N_29260,N_26061,N_26182);
nand U29261 (N_29261,N_26120,N_26945);
nand U29262 (N_29262,N_26527,N_27896);
or U29263 (N_29263,N_27276,N_26382);
nor U29264 (N_29264,N_27984,N_26646);
or U29265 (N_29265,N_26623,N_27061);
nor U29266 (N_29266,N_27044,N_27562);
nor U29267 (N_29267,N_27298,N_26831);
nand U29268 (N_29268,N_26238,N_26808);
nor U29269 (N_29269,N_27664,N_26606);
and U29270 (N_29270,N_26160,N_26202);
xnor U29271 (N_29271,N_26009,N_27686);
and U29272 (N_29272,N_27996,N_26612);
or U29273 (N_29273,N_27048,N_26916);
and U29274 (N_29274,N_26491,N_27794);
nand U29275 (N_29275,N_26178,N_26288);
nor U29276 (N_29276,N_26823,N_27379);
xor U29277 (N_29277,N_26145,N_26178);
and U29278 (N_29278,N_27537,N_27507);
and U29279 (N_29279,N_27965,N_27171);
nor U29280 (N_29280,N_27241,N_26144);
and U29281 (N_29281,N_26665,N_26436);
or U29282 (N_29282,N_27418,N_27542);
nor U29283 (N_29283,N_26092,N_26861);
or U29284 (N_29284,N_26239,N_26177);
or U29285 (N_29285,N_27239,N_26869);
nand U29286 (N_29286,N_27363,N_27091);
nand U29287 (N_29287,N_27098,N_26077);
nor U29288 (N_29288,N_26377,N_26256);
nand U29289 (N_29289,N_27658,N_27359);
nor U29290 (N_29290,N_27466,N_27833);
or U29291 (N_29291,N_26441,N_26713);
nand U29292 (N_29292,N_26983,N_27740);
or U29293 (N_29293,N_27198,N_26913);
or U29294 (N_29294,N_26240,N_27897);
or U29295 (N_29295,N_26394,N_27693);
and U29296 (N_29296,N_27622,N_27493);
and U29297 (N_29297,N_27581,N_26164);
and U29298 (N_29298,N_26559,N_27295);
or U29299 (N_29299,N_27787,N_26617);
and U29300 (N_29300,N_26807,N_26117);
or U29301 (N_29301,N_27799,N_27520);
nor U29302 (N_29302,N_27933,N_26892);
or U29303 (N_29303,N_27252,N_27745);
nand U29304 (N_29304,N_26554,N_26243);
nand U29305 (N_29305,N_26372,N_27478);
nand U29306 (N_29306,N_27463,N_27214);
nand U29307 (N_29307,N_27915,N_26980);
nor U29308 (N_29308,N_26830,N_26096);
and U29309 (N_29309,N_26836,N_26792);
or U29310 (N_29310,N_27581,N_26147);
nor U29311 (N_29311,N_26590,N_27961);
or U29312 (N_29312,N_27229,N_27783);
nor U29313 (N_29313,N_27720,N_26026);
and U29314 (N_29314,N_27294,N_26957);
nor U29315 (N_29315,N_27595,N_27128);
and U29316 (N_29316,N_27844,N_26546);
and U29317 (N_29317,N_26306,N_26747);
nor U29318 (N_29318,N_27851,N_27859);
or U29319 (N_29319,N_26472,N_27304);
and U29320 (N_29320,N_26091,N_26708);
or U29321 (N_29321,N_27507,N_27541);
and U29322 (N_29322,N_27441,N_26468);
nor U29323 (N_29323,N_27040,N_26893);
and U29324 (N_29324,N_27591,N_26247);
and U29325 (N_29325,N_27078,N_26750);
nand U29326 (N_29326,N_26384,N_26834);
nor U29327 (N_29327,N_27109,N_26987);
or U29328 (N_29328,N_27641,N_26043);
nand U29329 (N_29329,N_26815,N_26671);
and U29330 (N_29330,N_27638,N_26170);
nor U29331 (N_29331,N_27426,N_27567);
nand U29332 (N_29332,N_27294,N_26101);
nor U29333 (N_29333,N_26380,N_26377);
nand U29334 (N_29334,N_26078,N_26145);
nor U29335 (N_29335,N_26752,N_27866);
or U29336 (N_29336,N_27632,N_27493);
or U29337 (N_29337,N_26002,N_27952);
nor U29338 (N_29338,N_26298,N_27362);
nor U29339 (N_29339,N_27380,N_27350);
and U29340 (N_29340,N_27803,N_26378);
and U29341 (N_29341,N_27623,N_27532);
nor U29342 (N_29342,N_27245,N_26427);
and U29343 (N_29343,N_26172,N_26385);
nand U29344 (N_29344,N_26855,N_27596);
or U29345 (N_29345,N_26929,N_26602);
nor U29346 (N_29346,N_26908,N_27750);
nand U29347 (N_29347,N_27956,N_27301);
or U29348 (N_29348,N_27559,N_26145);
and U29349 (N_29349,N_26275,N_26900);
nor U29350 (N_29350,N_26956,N_26155);
or U29351 (N_29351,N_26833,N_26226);
and U29352 (N_29352,N_26165,N_27940);
or U29353 (N_29353,N_26279,N_26393);
and U29354 (N_29354,N_26095,N_27489);
nor U29355 (N_29355,N_26240,N_26935);
and U29356 (N_29356,N_26364,N_26109);
nor U29357 (N_29357,N_26835,N_26626);
or U29358 (N_29358,N_27349,N_26687);
nand U29359 (N_29359,N_27963,N_27419);
nor U29360 (N_29360,N_26296,N_26680);
and U29361 (N_29361,N_27050,N_27730);
and U29362 (N_29362,N_27882,N_26409);
and U29363 (N_29363,N_27130,N_27031);
nor U29364 (N_29364,N_27974,N_26688);
nand U29365 (N_29365,N_26856,N_26474);
or U29366 (N_29366,N_26554,N_26759);
nand U29367 (N_29367,N_27592,N_27017);
nand U29368 (N_29368,N_26731,N_26593);
nand U29369 (N_29369,N_26070,N_27746);
nor U29370 (N_29370,N_27296,N_26259);
and U29371 (N_29371,N_26036,N_27305);
or U29372 (N_29372,N_26125,N_26349);
nor U29373 (N_29373,N_27907,N_27734);
or U29374 (N_29374,N_26069,N_27620);
nor U29375 (N_29375,N_27338,N_27534);
nand U29376 (N_29376,N_26558,N_26675);
nor U29377 (N_29377,N_27423,N_27603);
nand U29378 (N_29378,N_26129,N_26903);
and U29379 (N_29379,N_26991,N_27437);
nor U29380 (N_29380,N_26910,N_26814);
nor U29381 (N_29381,N_27349,N_27867);
nor U29382 (N_29382,N_27126,N_27057);
and U29383 (N_29383,N_26384,N_26103);
nand U29384 (N_29384,N_26754,N_27089);
nand U29385 (N_29385,N_26234,N_27918);
or U29386 (N_29386,N_26332,N_26392);
nand U29387 (N_29387,N_26735,N_27971);
nand U29388 (N_29388,N_26366,N_26716);
nand U29389 (N_29389,N_26687,N_27388);
nand U29390 (N_29390,N_27957,N_27482);
nor U29391 (N_29391,N_27401,N_26888);
or U29392 (N_29392,N_26373,N_26496);
nand U29393 (N_29393,N_27965,N_27162);
nand U29394 (N_29394,N_27232,N_27875);
nand U29395 (N_29395,N_26059,N_27105);
or U29396 (N_29396,N_27521,N_26491);
and U29397 (N_29397,N_26322,N_27732);
and U29398 (N_29398,N_27506,N_26477);
nand U29399 (N_29399,N_27901,N_27491);
or U29400 (N_29400,N_26571,N_27123);
and U29401 (N_29401,N_26984,N_26510);
nand U29402 (N_29402,N_26359,N_27567);
or U29403 (N_29403,N_26861,N_26590);
nand U29404 (N_29404,N_27748,N_27027);
or U29405 (N_29405,N_26076,N_26996);
nand U29406 (N_29406,N_26388,N_26169);
nor U29407 (N_29407,N_27223,N_27064);
or U29408 (N_29408,N_26857,N_26454);
nand U29409 (N_29409,N_26205,N_27402);
nand U29410 (N_29410,N_27589,N_26048);
or U29411 (N_29411,N_27220,N_27251);
nand U29412 (N_29412,N_26035,N_27756);
nand U29413 (N_29413,N_26977,N_26005);
or U29414 (N_29414,N_27094,N_27047);
or U29415 (N_29415,N_27695,N_27523);
or U29416 (N_29416,N_26395,N_26043);
xor U29417 (N_29417,N_26033,N_27741);
nand U29418 (N_29418,N_27264,N_26201);
nor U29419 (N_29419,N_27186,N_27874);
nor U29420 (N_29420,N_26875,N_26362);
and U29421 (N_29421,N_27939,N_27203);
and U29422 (N_29422,N_27740,N_26808);
or U29423 (N_29423,N_27213,N_27356);
nand U29424 (N_29424,N_26657,N_26561);
and U29425 (N_29425,N_27616,N_26042);
nor U29426 (N_29426,N_26469,N_26899);
nand U29427 (N_29427,N_27016,N_27317);
nand U29428 (N_29428,N_27561,N_26038);
and U29429 (N_29429,N_27055,N_26906);
and U29430 (N_29430,N_26727,N_27069);
or U29431 (N_29431,N_26671,N_26737);
and U29432 (N_29432,N_26418,N_26936);
nor U29433 (N_29433,N_26813,N_27559);
nand U29434 (N_29434,N_26351,N_26823);
or U29435 (N_29435,N_27225,N_26445);
nor U29436 (N_29436,N_27580,N_26967);
nor U29437 (N_29437,N_26636,N_26307);
or U29438 (N_29438,N_26878,N_26263);
or U29439 (N_29439,N_26779,N_26493);
and U29440 (N_29440,N_26515,N_27283);
nand U29441 (N_29441,N_27104,N_27637);
and U29442 (N_29442,N_26895,N_27768);
and U29443 (N_29443,N_27270,N_27024);
and U29444 (N_29444,N_26255,N_27563);
or U29445 (N_29445,N_26214,N_27893);
nand U29446 (N_29446,N_26853,N_26700);
or U29447 (N_29447,N_26135,N_26272);
and U29448 (N_29448,N_27046,N_26544);
nand U29449 (N_29449,N_27854,N_26001);
nand U29450 (N_29450,N_27680,N_26346);
nor U29451 (N_29451,N_27776,N_27872);
or U29452 (N_29452,N_27518,N_26569);
nor U29453 (N_29453,N_27203,N_27185);
and U29454 (N_29454,N_26557,N_27791);
or U29455 (N_29455,N_26423,N_27800);
and U29456 (N_29456,N_27750,N_26645);
nand U29457 (N_29457,N_27493,N_27876);
and U29458 (N_29458,N_26625,N_27839);
and U29459 (N_29459,N_27791,N_26751);
nand U29460 (N_29460,N_26365,N_26900);
nand U29461 (N_29461,N_27238,N_26630);
nor U29462 (N_29462,N_26820,N_27854);
nor U29463 (N_29463,N_26033,N_27005);
or U29464 (N_29464,N_27622,N_26151);
and U29465 (N_29465,N_26403,N_26752);
nor U29466 (N_29466,N_26508,N_26252);
nand U29467 (N_29467,N_27447,N_27684);
or U29468 (N_29468,N_26671,N_27920);
and U29469 (N_29469,N_27126,N_27709);
nor U29470 (N_29470,N_27691,N_26330);
nor U29471 (N_29471,N_27238,N_26875);
nor U29472 (N_29472,N_27197,N_27651);
nand U29473 (N_29473,N_26867,N_27588);
or U29474 (N_29474,N_26055,N_27255);
and U29475 (N_29475,N_26996,N_27136);
or U29476 (N_29476,N_27263,N_26356);
and U29477 (N_29477,N_26896,N_26563);
nand U29478 (N_29478,N_27039,N_26081);
or U29479 (N_29479,N_27702,N_27549);
or U29480 (N_29480,N_27333,N_27382);
or U29481 (N_29481,N_26991,N_26870);
nand U29482 (N_29482,N_27152,N_26872);
or U29483 (N_29483,N_27535,N_26518);
and U29484 (N_29484,N_26814,N_27111);
nand U29485 (N_29485,N_27448,N_27495);
and U29486 (N_29486,N_27859,N_26094);
nor U29487 (N_29487,N_26104,N_27938);
or U29488 (N_29488,N_26174,N_26451);
or U29489 (N_29489,N_27125,N_27345);
nor U29490 (N_29490,N_26064,N_26301);
nor U29491 (N_29491,N_26297,N_27007);
nand U29492 (N_29492,N_26540,N_27535);
nand U29493 (N_29493,N_26877,N_27653);
nor U29494 (N_29494,N_27213,N_27431);
nor U29495 (N_29495,N_27948,N_26228);
and U29496 (N_29496,N_26882,N_27507);
xor U29497 (N_29497,N_26032,N_27014);
and U29498 (N_29498,N_27117,N_26979);
nand U29499 (N_29499,N_27523,N_27067);
or U29500 (N_29500,N_26600,N_27091);
and U29501 (N_29501,N_26123,N_26227);
nand U29502 (N_29502,N_27498,N_26615);
and U29503 (N_29503,N_26246,N_27697);
or U29504 (N_29504,N_26169,N_26612);
nand U29505 (N_29505,N_26741,N_27709);
xnor U29506 (N_29506,N_27909,N_27168);
and U29507 (N_29507,N_27492,N_27129);
nor U29508 (N_29508,N_26305,N_27977);
and U29509 (N_29509,N_26707,N_26471);
and U29510 (N_29510,N_27881,N_27552);
or U29511 (N_29511,N_26581,N_26629);
or U29512 (N_29512,N_26734,N_27940);
or U29513 (N_29513,N_26817,N_26774);
nand U29514 (N_29514,N_26873,N_27707);
nor U29515 (N_29515,N_26228,N_27748);
and U29516 (N_29516,N_27331,N_27102);
or U29517 (N_29517,N_27829,N_27930);
and U29518 (N_29518,N_26592,N_27140);
and U29519 (N_29519,N_27158,N_26676);
nand U29520 (N_29520,N_27370,N_26514);
nand U29521 (N_29521,N_27949,N_26922);
nand U29522 (N_29522,N_26834,N_26010);
nand U29523 (N_29523,N_26296,N_26115);
nor U29524 (N_29524,N_27980,N_26266);
nand U29525 (N_29525,N_27063,N_26647);
and U29526 (N_29526,N_27851,N_27210);
or U29527 (N_29527,N_26458,N_27590);
and U29528 (N_29528,N_27941,N_26934);
nor U29529 (N_29529,N_27665,N_27473);
and U29530 (N_29530,N_27299,N_27467);
and U29531 (N_29531,N_26183,N_26833);
and U29532 (N_29532,N_26809,N_26782);
or U29533 (N_29533,N_27358,N_26432);
and U29534 (N_29534,N_27244,N_26094);
and U29535 (N_29535,N_26032,N_26894);
or U29536 (N_29536,N_27496,N_27852);
or U29537 (N_29537,N_27133,N_26193);
and U29538 (N_29538,N_26396,N_26841);
or U29539 (N_29539,N_26917,N_27812);
nor U29540 (N_29540,N_26771,N_26467);
or U29541 (N_29541,N_27073,N_27912);
nor U29542 (N_29542,N_26844,N_27584);
or U29543 (N_29543,N_27569,N_27657);
or U29544 (N_29544,N_26118,N_26102);
xor U29545 (N_29545,N_27318,N_26916);
nor U29546 (N_29546,N_26255,N_27642);
or U29547 (N_29547,N_26761,N_27128);
nand U29548 (N_29548,N_27046,N_26618);
and U29549 (N_29549,N_26928,N_27722);
nand U29550 (N_29550,N_26068,N_26749);
nor U29551 (N_29551,N_26022,N_26899);
nor U29552 (N_29552,N_26423,N_27809);
or U29553 (N_29553,N_26767,N_26342);
or U29554 (N_29554,N_26779,N_27774);
and U29555 (N_29555,N_26955,N_26477);
and U29556 (N_29556,N_27097,N_27472);
nand U29557 (N_29557,N_26223,N_26118);
nor U29558 (N_29558,N_26621,N_26993);
or U29559 (N_29559,N_26197,N_27736);
and U29560 (N_29560,N_26153,N_26968);
or U29561 (N_29561,N_26898,N_27303);
or U29562 (N_29562,N_27757,N_26570);
nor U29563 (N_29563,N_27521,N_26590);
or U29564 (N_29564,N_26879,N_26899);
or U29565 (N_29565,N_26333,N_27312);
and U29566 (N_29566,N_27365,N_27265);
nor U29567 (N_29567,N_26616,N_27317);
and U29568 (N_29568,N_27216,N_27888);
nor U29569 (N_29569,N_26809,N_26889);
nand U29570 (N_29570,N_26245,N_27633);
nand U29571 (N_29571,N_26204,N_27426);
and U29572 (N_29572,N_26292,N_27855);
nand U29573 (N_29573,N_26747,N_26121);
or U29574 (N_29574,N_26545,N_27920);
nor U29575 (N_29575,N_26608,N_27071);
or U29576 (N_29576,N_27300,N_26041);
or U29577 (N_29577,N_27120,N_27150);
nor U29578 (N_29578,N_27575,N_27639);
and U29579 (N_29579,N_27878,N_27285);
and U29580 (N_29580,N_27368,N_27340);
or U29581 (N_29581,N_26068,N_27051);
nand U29582 (N_29582,N_27016,N_26200);
or U29583 (N_29583,N_27824,N_26780);
and U29584 (N_29584,N_26929,N_26187);
nand U29585 (N_29585,N_26391,N_27205);
nor U29586 (N_29586,N_27652,N_26264);
and U29587 (N_29587,N_26869,N_27463);
nor U29588 (N_29588,N_27188,N_26145);
and U29589 (N_29589,N_26760,N_27391);
and U29590 (N_29590,N_26593,N_27511);
or U29591 (N_29591,N_26605,N_26625);
nor U29592 (N_29592,N_26808,N_27235);
or U29593 (N_29593,N_27738,N_26709);
and U29594 (N_29594,N_26695,N_27466);
or U29595 (N_29595,N_27005,N_26876);
or U29596 (N_29596,N_26428,N_26610);
or U29597 (N_29597,N_26194,N_26586);
and U29598 (N_29598,N_26282,N_26479);
and U29599 (N_29599,N_27334,N_26576);
nor U29600 (N_29600,N_27951,N_27451);
xor U29601 (N_29601,N_26216,N_26469);
nor U29602 (N_29602,N_26255,N_27260);
or U29603 (N_29603,N_27306,N_26708);
or U29604 (N_29604,N_27357,N_26317);
and U29605 (N_29605,N_26614,N_27955);
xor U29606 (N_29606,N_27764,N_26287);
and U29607 (N_29607,N_26390,N_27404);
nor U29608 (N_29608,N_27187,N_27802);
and U29609 (N_29609,N_26928,N_27583);
nor U29610 (N_29610,N_27435,N_26460);
and U29611 (N_29611,N_26970,N_26547);
xor U29612 (N_29612,N_26236,N_26285);
or U29613 (N_29613,N_27171,N_27446);
nor U29614 (N_29614,N_26686,N_26131);
and U29615 (N_29615,N_26231,N_26514);
or U29616 (N_29616,N_27961,N_26919);
nand U29617 (N_29617,N_27260,N_26307);
nor U29618 (N_29618,N_26342,N_26251);
nand U29619 (N_29619,N_26274,N_27195);
nand U29620 (N_29620,N_26442,N_26074);
nand U29621 (N_29621,N_27560,N_26803);
nor U29622 (N_29622,N_27280,N_26908);
nand U29623 (N_29623,N_26322,N_26981);
and U29624 (N_29624,N_26588,N_27107);
nand U29625 (N_29625,N_26061,N_27445);
nand U29626 (N_29626,N_26961,N_26092);
or U29627 (N_29627,N_27604,N_26419);
nand U29628 (N_29628,N_26721,N_27584);
nor U29629 (N_29629,N_27168,N_26001);
nor U29630 (N_29630,N_26304,N_26092);
and U29631 (N_29631,N_27631,N_27041);
and U29632 (N_29632,N_27686,N_27477);
nor U29633 (N_29633,N_26300,N_27287);
and U29634 (N_29634,N_27824,N_27079);
and U29635 (N_29635,N_27070,N_27684);
nand U29636 (N_29636,N_27105,N_26348);
nor U29637 (N_29637,N_27262,N_27599);
and U29638 (N_29638,N_27833,N_27521);
nand U29639 (N_29639,N_27194,N_26124);
nand U29640 (N_29640,N_26307,N_27619);
and U29641 (N_29641,N_26779,N_27778);
nor U29642 (N_29642,N_26035,N_27819);
nand U29643 (N_29643,N_26350,N_26152);
nand U29644 (N_29644,N_26996,N_26387);
and U29645 (N_29645,N_27966,N_27229);
or U29646 (N_29646,N_26206,N_26048);
nand U29647 (N_29647,N_26779,N_26129);
or U29648 (N_29648,N_27770,N_26272);
nor U29649 (N_29649,N_27416,N_26529);
xor U29650 (N_29650,N_26118,N_27931);
xnor U29651 (N_29651,N_27541,N_26866);
nand U29652 (N_29652,N_27448,N_27033);
and U29653 (N_29653,N_26851,N_26891);
nand U29654 (N_29654,N_27298,N_27775);
nor U29655 (N_29655,N_26747,N_27062);
nor U29656 (N_29656,N_27599,N_27152);
nor U29657 (N_29657,N_27178,N_27583);
nand U29658 (N_29658,N_27386,N_26417);
or U29659 (N_29659,N_27776,N_26314);
or U29660 (N_29660,N_26358,N_27261);
and U29661 (N_29661,N_27074,N_26789);
or U29662 (N_29662,N_27558,N_26327);
and U29663 (N_29663,N_26367,N_27445);
nand U29664 (N_29664,N_27126,N_27794);
or U29665 (N_29665,N_27608,N_26311);
nor U29666 (N_29666,N_27652,N_27752);
nand U29667 (N_29667,N_27991,N_27771);
xnor U29668 (N_29668,N_27685,N_26773);
or U29669 (N_29669,N_27837,N_27450);
xor U29670 (N_29670,N_27272,N_27352);
nor U29671 (N_29671,N_27800,N_26914);
or U29672 (N_29672,N_26355,N_27355);
and U29673 (N_29673,N_26082,N_26440);
nor U29674 (N_29674,N_27636,N_26828);
nor U29675 (N_29675,N_27903,N_27775);
and U29676 (N_29676,N_27571,N_26511);
nand U29677 (N_29677,N_27119,N_27182);
nand U29678 (N_29678,N_26033,N_26782);
and U29679 (N_29679,N_26044,N_27367);
nor U29680 (N_29680,N_27284,N_27627);
nor U29681 (N_29681,N_26026,N_27198);
nor U29682 (N_29682,N_27506,N_27358);
or U29683 (N_29683,N_26895,N_27904);
and U29684 (N_29684,N_27032,N_27070);
nand U29685 (N_29685,N_27027,N_27170);
nand U29686 (N_29686,N_27207,N_26071);
or U29687 (N_29687,N_27883,N_26734);
and U29688 (N_29688,N_27823,N_27628);
nor U29689 (N_29689,N_27671,N_26053);
or U29690 (N_29690,N_27167,N_26767);
nand U29691 (N_29691,N_26575,N_27711);
nand U29692 (N_29692,N_26986,N_27932);
nor U29693 (N_29693,N_27667,N_27896);
nand U29694 (N_29694,N_26610,N_27908);
nand U29695 (N_29695,N_26153,N_26111);
nand U29696 (N_29696,N_26401,N_27087);
nand U29697 (N_29697,N_26686,N_26782);
or U29698 (N_29698,N_27859,N_27423);
and U29699 (N_29699,N_26904,N_26674);
nor U29700 (N_29700,N_26213,N_26758);
nor U29701 (N_29701,N_27052,N_27508);
or U29702 (N_29702,N_27201,N_26541);
nand U29703 (N_29703,N_26858,N_27940);
or U29704 (N_29704,N_27513,N_27230);
nand U29705 (N_29705,N_27711,N_26847);
xnor U29706 (N_29706,N_26693,N_27095);
and U29707 (N_29707,N_26939,N_26136);
and U29708 (N_29708,N_26134,N_27641);
or U29709 (N_29709,N_26840,N_26904);
or U29710 (N_29710,N_27133,N_27990);
nor U29711 (N_29711,N_26195,N_26379);
nand U29712 (N_29712,N_27015,N_26312);
nand U29713 (N_29713,N_27933,N_27550);
nand U29714 (N_29714,N_26746,N_26137);
nor U29715 (N_29715,N_27350,N_26610);
or U29716 (N_29716,N_26182,N_26320);
nand U29717 (N_29717,N_27817,N_26291);
nor U29718 (N_29718,N_26046,N_27853);
and U29719 (N_29719,N_26798,N_26068);
or U29720 (N_29720,N_27118,N_27924);
and U29721 (N_29721,N_26157,N_27511);
or U29722 (N_29722,N_26611,N_26434);
nor U29723 (N_29723,N_27598,N_26801);
nand U29724 (N_29724,N_27777,N_26870);
nand U29725 (N_29725,N_26808,N_27523);
and U29726 (N_29726,N_27576,N_27574);
or U29727 (N_29727,N_26633,N_27233);
nor U29728 (N_29728,N_27531,N_26983);
nand U29729 (N_29729,N_26495,N_27154);
nor U29730 (N_29730,N_26921,N_27120);
nor U29731 (N_29731,N_27113,N_27739);
nor U29732 (N_29732,N_26778,N_27849);
or U29733 (N_29733,N_27326,N_26034);
and U29734 (N_29734,N_27678,N_27763);
and U29735 (N_29735,N_27678,N_26582);
nand U29736 (N_29736,N_27784,N_27926);
nand U29737 (N_29737,N_27391,N_27783);
xor U29738 (N_29738,N_27072,N_26041);
nand U29739 (N_29739,N_26662,N_27388);
nor U29740 (N_29740,N_27910,N_27909);
and U29741 (N_29741,N_27266,N_27967);
nand U29742 (N_29742,N_26983,N_27598);
nand U29743 (N_29743,N_27820,N_26694);
nand U29744 (N_29744,N_27885,N_27573);
and U29745 (N_29745,N_26051,N_27504);
nand U29746 (N_29746,N_26142,N_26786);
or U29747 (N_29747,N_27737,N_26468);
and U29748 (N_29748,N_27043,N_26903);
and U29749 (N_29749,N_27915,N_26979);
and U29750 (N_29750,N_26439,N_26569);
or U29751 (N_29751,N_26604,N_26870);
nand U29752 (N_29752,N_27649,N_26401);
xnor U29753 (N_29753,N_27140,N_26355);
nand U29754 (N_29754,N_27662,N_26958);
or U29755 (N_29755,N_26670,N_27340);
nand U29756 (N_29756,N_26782,N_27700);
or U29757 (N_29757,N_27043,N_27490);
nand U29758 (N_29758,N_27109,N_27911);
nor U29759 (N_29759,N_27290,N_27939);
or U29760 (N_29760,N_27812,N_27995);
or U29761 (N_29761,N_27397,N_26187);
or U29762 (N_29762,N_27902,N_26549);
and U29763 (N_29763,N_27770,N_26858);
nand U29764 (N_29764,N_26770,N_27059);
nor U29765 (N_29765,N_26372,N_27515);
nand U29766 (N_29766,N_26853,N_26382);
nand U29767 (N_29767,N_27987,N_27452);
and U29768 (N_29768,N_26890,N_27178);
and U29769 (N_29769,N_26858,N_26812);
xnor U29770 (N_29770,N_27218,N_26272);
xor U29771 (N_29771,N_27544,N_26521);
and U29772 (N_29772,N_27733,N_26258);
nand U29773 (N_29773,N_26477,N_27668);
nor U29774 (N_29774,N_26399,N_27824);
nand U29775 (N_29775,N_26002,N_26341);
or U29776 (N_29776,N_26031,N_26788);
or U29777 (N_29777,N_26647,N_27064);
or U29778 (N_29778,N_26897,N_27989);
nand U29779 (N_29779,N_26742,N_26594);
nand U29780 (N_29780,N_26564,N_26745);
and U29781 (N_29781,N_27054,N_27118);
or U29782 (N_29782,N_27994,N_27313);
xor U29783 (N_29783,N_27691,N_27268);
nor U29784 (N_29784,N_27487,N_27525);
nor U29785 (N_29785,N_26246,N_26010);
or U29786 (N_29786,N_26735,N_26827);
nand U29787 (N_29787,N_27641,N_26872);
nand U29788 (N_29788,N_26824,N_26308);
and U29789 (N_29789,N_26749,N_26473);
or U29790 (N_29790,N_27090,N_27535);
nor U29791 (N_29791,N_26859,N_27571);
nor U29792 (N_29792,N_27869,N_27676);
and U29793 (N_29793,N_27435,N_26078);
nand U29794 (N_29794,N_27887,N_27347);
nand U29795 (N_29795,N_26158,N_27547);
and U29796 (N_29796,N_26264,N_27122);
nor U29797 (N_29797,N_27199,N_27221);
or U29798 (N_29798,N_27982,N_26692);
nor U29799 (N_29799,N_26611,N_27359);
and U29800 (N_29800,N_27384,N_26038);
nor U29801 (N_29801,N_27908,N_27742);
and U29802 (N_29802,N_26516,N_26776);
xnor U29803 (N_29803,N_27621,N_27983);
nor U29804 (N_29804,N_27093,N_26054);
nand U29805 (N_29805,N_27857,N_26858);
and U29806 (N_29806,N_27933,N_26779);
nand U29807 (N_29807,N_26623,N_26273);
nand U29808 (N_29808,N_27656,N_26562);
and U29809 (N_29809,N_26721,N_27083);
nand U29810 (N_29810,N_26983,N_27205);
nand U29811 (N_29811,N_26216,N_26502);
nor U29812 (N_29812,N_26505,N_26125);
and U29813 (N_29813,N_27513,N_26595);
or U29814 (N_29814,N_27288,N_27948);
nor U29815 (N_29815,N_26043,N_27913);
and U29816 (N_29816,N_27345,N_26654);
and U29817 (N_29817,N_27835,N_26294);
nor U29818 (N_29818,N_26032,N_26957);
and U29819 (N_29819,N_27774,N_26184);
and U29820 (N_29820,N_26332,N_27445);
or U29821 (N_29821,N_26510,N_26350);
nor U29822 (N_29822,N_26432,N_26009);
xor U29823 (N_29823,N_26166,N_26432);
nor U29824 (N_29824,N_26315,N_27672);
nand U29825 (N_29825,N_27553,N_26991);
and U29826 (N_29826,N_27823,N_27447);
nand U29827 (N_29827,N_27069,N_27267);
nand U29828 (N_29828,N_27049,N_26650);
or U29829 (N_29829,N_26835,N_27161);
or U29830 (N_29830,N_27649,N_26843);
nor U29831 (N_29831,N_27120,N_26202);
and U29832 (N_29832,N_27334,N_26468);
nor U29833 (N_29833,N_27451,N_26956);
or U29834 (N_29834,N_26552,N_27974);
or U29835 (N_29835,N_26492,N_27182);
or U29836 (N_29836,N_26171,N_26989);
nand U29837 (N_29837,N_26481,N_26085);
or U29838 (N_29838,N_26462,N_27206);
nand U29839 (N_29839,N_27696,N_27083);
and U29840 (N_29840,N_26198,N_27081);
nor U29841 (N_29841,N_27737,N_27075);
nand U29842 (N_29842,N_27402,N_27135);
or U29843 (N_29843,N_26420,N_26533);
or U29844 (N_29844,N_26265,N_27410);
or U29845 (N_29845,N_26360,N_27411);
nor U29846 (N_29846,N_26951,N_27959);
or U29847 (N_29847,N_26639,N_26191);
and U29848 (N_29848,N_27040,N_27277);
xnor U29849 (N_29849,N_27556,N_27053);
xnor U29850 (N_29850,N_26843,N_27379);
nor U29851 (N_29851,N_26009,N_27190);
nand U29852 (N_29852,N_26158,N_26254);
or U29853 (N_29853,N_27285,N_26867);
xor U29854 (N_29854,N_26045,N_27615);
and U29855 (N_29855,N_27805,N_26378);
nand U29856 (N_29856,N_26113,N_27653);
or U29857 (N_29857,N_26277,N_26088);
and U29858 (N_29858,N_27505,N_27733);
and U29859 (N_29859,N_27483,N_27920);
xnor U29860 (N_29860,N_26795,N_27874);
or U29861 (N_29861,N_26340,N_26352);
nand U29862 (N_29862,N_27680,N_26518);
and U29863 (N_29863,N_26569,N_27411);
and U29864 (N_29864,N_27788,N_27271);
nand U29865 (N_29865,N_26404,N_27903);
and U29866 (N_29866,N_27632,N_27430);
nor U29867 (N_29867,N_26287,N_27786);
and U29868 (N_29868,N_26109,N_27497);
and U29869 (N_29869,N_27014,N_26715);
or U29870 (N_29870,N_27649,N_26906);
nor U29871 (N_29871,N_27360,N_27981);
or U29872 (N_29872,N_26577,N_26122);
nor U29873 (N_29873,N_27817,N_27062);
nand U29874 (N_29874,N_26922,N_27872);
nor U29875 (N_29875,N_26146,N_27325);
or U29876 (N_29876,N_26890,N_27146);
and U29877 (N_29877,N_27545,N_26874);
or U29878 (N_29878,N_26313,N_27987);
nor U29879 (N_29879,N_26233,N_26319);
nor U29880 (N_29880,N_26988,N_27389);
and U29881 (N_29881,N_27380,N_27405);
nand U29882 (N_29882,N_26935,N_27829);
nor U29883 (N_29883,N_27470,N_26148);
and U29884 (N_29884,N_27281,N_27393);
nand U29885 (N_29885,N_27760,N_27690);
or U29886 (N_29886,N_27435,N_26741);
nand U29887 (N_29887,N_26199,N_26513);
nor U29888 (N_29888,N_26747,N_27267);
and U29889 (N_29889,N_26744,N_26126);
nor U29890 (N_29890,N_27965,N_26415);
or U29891 (N_29891,N_27856,N_26682);
xor U29892 (N_29892,N_27668,N_27071);
or U29893 (N_29893,N_26126,N_26293);
nor U29894 (N_29894,N_27201,N_27262);
nor U29895 (N_29895,N_27106,N_26318);
nor U29896 (N_29896,N_27368,N_27649);
and U29897 (N_29897,N_26315,N_26213);
nor U29898 (N_29898,N_27050,N_26911);
nor U29899 (N_29899,N_26829,N_26847);
nand U29900 (N_29900,N_27980,N_26583);
and U29901 (N_29901,N_27280,N_27469);
or U29902 (N_29902,N_26460,N_27930);
nor U29903 (N_29903,N_26099,N_26276);
and U29904 (N_29904,N_26542,N_26740);
nand U29905 (N_29905,N_27097,N_26079);
nor U29906 (N_29906,N_26284,N_26616);
and U29907 (N_29907,N_26082,N_26227);
nand U29908 (N_29908,N_27926,N_26815);
nand U29909 (N_29909,N_27558,N_26487);
or U29910 (N_29910,N_27161,N_27540);
nand U29911 (N_29911,N_26294,N_26698);
and U29912 (N_29912,N_27820,N_26436);
and U29913 (N_29913,N_26663,N_27926);
and U29914 (N_29914,N_27019,N_27565);
nand U29915 (N_29915,N_27732,N_26206);
nor U29916 (N_29916,N_27728,N_27229);
nand U29917 (N_29917,N_27510,N_26754);
and U29918 (N_29918,N_27836,N_27317);
and U29919 (N_29919,N_27666,N_27050);
nand U29920 (N_29920,N_26515,N_26957);
and U29921 (N_29921,N_27502,N_27421);
or U29922 (N_29922,N_26956,N_26839);
nor U29923 (N_29923,N_26215,N_26681);
and U29924 (N_29924,N_27131,N_27636);
nand U29925 (N_29925,N_26764,N_26133);
nor U29926 (N_29926,N_26861,N_26134);
or U29927 (N_29927,N_26308,N_26996);
and U29928 (N_29928,N_26789,N_26378);
or U29929 (N_29929,N_27210,N_27700);
or U29930 (N_29930,N_27541,N_27367);
nor U29931 (N_29931,N_26663,N_26569);
and U29932 (N_29932,N_27023,N_26208);
nor U29933 (N_29933,N_27405,N_26813);
nand U29934 (N_29934,N_26459,N_27016);
or U29935 (N_29935,N_27533,N_27178);
or U29936 (N_29936,N_26357,N_26328);
and U29937 (N_29937,N_26014,N_26602);
or U29938 (N_29938,N_26429,N_26370);
nor U29939 (N_29939,N_27108,N_26368);
xnor U29940 (N_29940,N_27364,N_27748);
or U29941 (N_29941,N_26168,N_27437);
nor U29942 (N_29942,N_27535,N_27126);
and U29943 (N_29943,N_26095,N_26519);
and U29944 (N_29944,N_27407,N_27015);
and U29945 (N_29945,N_27119,N_27125);
nand U29946 (N_29946,N_26563,N_27177);
nor U29947 (N_29947,N_26983,N_26511);
nand U29948 (N_29948,N_27451,N_26097);
and U29949 (N_29949,N_27641,N_26736);
nor U29950 (N_29950,N_26811,N_27602);
or U29951 (N_29951,N_26592,N_26759);
or U29952 (N_29952,N_27034,N_26831);
or U29953 (N_29953,N_27075,N_26246);
nand U29954 (N_29954,N_27894,N_27414);
and U29955 (N_29955,N_27004,N_26170);
nor U29956 (N_29956,N_27726,N_27954);
xnor U29957 (N_29957,N_27031,N_27648);
or U29958 (N_29958,N_26975,N_26264);
nand U29959 (N_29959,N_27889,N_26306);
nor U29960 (N_29960,N_27430,N_26890);
and U29961 (N_29961,N_26740,N_26307);
or U29962 (N_29962,N_27040,N_26062);
nand U29963 (N_29963,N_26326,N_26156);
or U29964 (N_29964,N_27333,N_27591);
and U29965 (N_29965,N_27265,N_26685);
and U29966 (N_29966,N_27818,N_26988);
nor U29967 (N_29967,N_27676,N_27667);
nand U29968 (N_29968,N_27682,N_26094);
or U29969 (N_29969,N_26671,N_26904);
nand U29970 (N_29970,N_27663,N_27545);
nand U29971 (N_29971,N_27774,N_26334);
nor U29972 (N_29972,N_26076,N_27020);
xor U29973 (N_29973,N_27238,N_26852);
nand U29974 (N_29974,N_26589,N_27374);
or U29975 (N_29975,N_27860,N_26860);
and U29976 (N_29976,N_27112,N_26768);
nor U29977 (N_29977,N_26163,N_26524);
nor U29978 (N_29978,N_26043,N_27128);
and U29979 (N_29979,N_26038,N_27441);
nand U29980 (N_29980,N_26574,N_27745);
nand U29981 (N_29981,N_26259,N_26324);
nand U29982 (N_29982,N_26243,N_27871);
and U29983 (N_29983,N_26302,N_27450);
nor U29984 (N_29984,N_26617,N_27132);
nor U29985 (N_29985,N_26801,N_26810);
or U29986 (N_29986,N_27605,N_27828);
nand U29987 (N_29987,N_27099,N_27607);
or U29988 (N_29988,N_26748,N_27225);
nor U29989 (N_29989,N_27533,N_26004);
nor U29990 (N_29990,N_27538,N_26957);
nor U29991 (N_29991,N_26997,N_27994);
or U29992 (N_29992,N_27117,N_27579);
and U29993 (N_29993,N_27780,N_26428);
or U29994 (N_29994,N_27100,N_27461);
and U29995 (N_29995,N_26040,N_27741);
and U29996 (N_29996,N_27837,N_27355);
nor U29997 (N_29997,N_26445,N_26868);
nand U29998 (N_29998,N_27740,N_27119);
or U29999 (N_29999,N_27361,N_26220);
and U30000 (N_30000,N_28345,N_29089);
nor U30001 (N_30001,N_28754,N_28927);
nor U30002 (N_30002,N_28426,N_28178);
nand U30003 (N_30003,N_29015,N_28903);
nand U30004 (N_30004,N_29468,N_29627);
or U30005 (N_30005,N_29977,N_28886);
or U30006 (N_30006,N_29360,N_29511);
nor U30007 (N_30007,N_29751,N_28817);
or U30008 (N_30008,N_29621,N_29731);
or U30009 (N_30009,N_28733,N_28298);
nand U30010 (N_30010,N_28648,N_28931);
xor U30011 (N_30011,N_29316,N_28845);
and U30012 (N_30012,N_29113,N_29782);
or U30013 (N_30013,N_28271,N_29382);
or U30014 (N_30014,N_28210,N_28892);
nand U30015 (N_30015,N_29629,N_29713);
nand U30016 (N_30016,N_28166,N_29309);
or U30017 (N_30017,N_29573,N_29454);
nor U30018 (N_30018,N_29153,N_28299);
or U30019 (N_30019,N_29609,N_29144);
or U30020 (N_30020,N_28380,N_28326);
and U30021 (N_30021,N_29825,N_28861);
nor U30022 (N_30022,N_28971,N_29487);
nand U30023 (N_30023,N_29680,N_29997);
nand U30024 (N_30024,N_29881,N_28910);
nor U30025 (N_30025,N_29444,N_29306);
nor U30026 (N_30026,N_29325,N_29778);
nor U30027 (N_30027,N_28394,N_29310);
or U30028 (N_30028,N_29994,N_29385);
nor U30029 (N_30029,N_28300,N_29167);
or U30030 (N_30030,N_29707,N_28690);
nand U30031 (N_30031,N_28372,N_29636);
nand U30032 (N_30032,N_29995,N_28292);
nor U30033 (N_30033,N_29357,N_28431);
nor U30034 (N_30034,N_29319,N_29358);
nand U30035 (N_30035,N_29570,N_28093);
nor U30036 (N_30036,N_29507,N_29117);
nand U30037 (N_30037,N_29038,N_29384);
nor U30038 (N_30038,N_28740,N_28900);
nand U30039 (N_30039,N_29893,N_29365);
and U30040 (N_30040,N_28608,N_28712);
nor U30041 (N_30041,N_29361,N_29499);
or U30042 (N_30042,N_28446,N_28416);
and U30043 (N_30043,N_29483,N_29830);
or U30044 (N_30044,N_29470,N_29069);
nand U30045 (N_30045,N_28260,N_29971);
xnor U30046 (N_30046,N_28441,N_29286);
nand U30047 (N_30047,N_29908,N_28484);
nor U30048 (N_30048,N_28790,N_28400);
and U30049 (N_30049,N_28947,N_28647);
nand U30050 (N_30050,N_28053,N_28666);
and U30051 (N_30051,N_28638,N_29135);
and U30052 (N_30052,N_28285,N_28987);
nand U30053 (N_30053,N_28350,N_28730);
and U30054 (N_30054,N_29019,N_29773);
and U30055 (N_30055,N_28286,N_28640);
and U30056 (N_30056,N_28098,N_29281);
nor U30057 (N_30057,N_29345,N_29052);
or U30058 (N_30058,N_28370,N_29809);
nand U30059 (N_30059,N_29689,N_29540);
and U30060 (N_30060,N_29603,N_28766);
nand U30061 (N_30061,N_29222,N_28948);
nand U30062 (N_30062,N_28836,N_28376);
or U30063 (N_30063,N_28874,N_29072);
nor U30064 (N_30064,N_29127,N_29161);
nand U30065 (N_30065,N_28953,N_28095);
or U30066 (N_30066,N_29170,N_28813);
and U30067 (N_30067,N_28170,N_29269);
or U30068 (N_30068,N_29710,N_28348);
and U30069 (N_30069,N_28004,N_29930);
or U30070 (N_30070,N_29101,N_28173);
nor U30071 (N_30071,N_28430,N_28842);
or U30072 (N_30072,N_29983,N_29386);
nor U30073 (N_30073,N_28551,N_29756);
nand U30074 (N_30074,N_29327,N_28448);
and U30075 (N_30075,N_28857,N_28725);
nor U30076 (N_30076,N_28807,N_29683);
and U30077 (N_30077,N_28154,N_29461);
nor U30078 (N_30078,N_28691,N_28851);
and U30079 (N_30079,N_28552,N_28782);
nand U30080 (N_30080,N_29863,N_28600);
and U30081 (N_30081,N_28133,N_29473);
or U30082 (N_30082,N_28720,N_29133);
nor U30083 (N_30083,N_28082,N_28025);
nor U30084 (N_30084,N_29060,N_28989);
nand U30085 (N_30085,N_29786,N_28103);
nand U30086 (N_30086,N_28655,N_29377);
or U30087 (N_30087,N_29688,N_29498);
or U30088 (N_30088,N_28447,N_29864);
nor U30089 (N_30089,N_28320,N_28988);
nor U30090 (N_30090,N_28627,N_29404);
and U30091 (N_30091,N_28214,N_28227);
nand U30092 (N_30092,N_28205,N_29673);
nor U30093 (N_30093,N_29560,N_28250);
or U30094 (N_30094,N_28556,N_29427);
nor U30095 (N_30095,N_28657,N_29951);
or U30096 (N_30096,N_28662,N_29624);
or U30097 (N_30097,N_29542,N_28429);
and U30098 (N_30098,N_28709,N_29899);
nand U30099 (N_30099,N_28768,N_29594);
and U30100 (N_30100,N_28715,N_28054);
xnor U30101 (N_30101,N_29040,N_28080);
nand U30102 (N_30102,N_29036,N_29438);
nor U30103 (N_30103,N_29595,N_29942);
nor U30104 (N_30104,N_29264,N_28179);
or U30105 (N_30105,N_29248,N_29581);
nor U30106 (N_30106,N_28839,N_28065);
nor U30107 (N_30107,N_28658,N_29156);
and U30108 (N_30108,N_29564,N_28891);
nor U30109 (N_30109,N_28788,N_28741);
and U30110 (N_30110,N_29582,N_28496);
and U30111 (N_30111,N_29589,N_28010);
or U30112 (N_30112,N_28324,N_28256);
and U30113 (N_30113,N_28219,N_29142);
nor U30114 (N_30114,N_29650,N_28506);
nand U30115 (N_30115,N_28387,N_29270);
xnor U30116 (N_30116,N_28689,N_28963);
nor U30117 (N_30117,N_29279,N_29042);
nor U30118 (N_30118,N_28304,N_28682);
nor U30119 (N_30119,N_29146,N_28873);
nand U30120 (N_30120,N_29734,N_28120);
or U30121 (N_30121,N_28038,N_29642);
or U30122 (N_30122,N_28195,N_28625);
and U30123 (N_30123,N_28273,N_29293);
nand U30124 (N_30124,N_28193,N_28465);
and U30125 (N_30125,N_29652,N_28194);
or U30126 (N_30126,N_29716,N_28478);
nor U30127 (N_30127,N_28486,N_28843);
nor U30128 (N_30128,N_28140,N_29867);
or U30129 (N_30129,N_29157,N_28505);
or U30130 (N_30130,N_28611,N_29768);
nand U30131 (N_30131,N_28895,N_29972);
nand U30132 (N_30132,N_29800,N_28485);
nand U30133 (N_30133,N_28435,N_29634);
and U30134 (N_30134,N_29579,N_29393);
or U30135 (N_30135,N_29148,N_28353);
and U30136 (N_30136,N_29744,N_28616);
xnor U30137 (N_30137,N_28453,N_28583);
nor U30138 (N_30138,N_28223,N_29583);
and U30139 (N_30139,N_28096,N_28808);
or U30140 (N_30140,N_28379,N_28112);
nand U30141 (N_30141,N_28185,N_29267);
nand U30142 (N_30142,N_29124,N_29115);
or U30143 (N_30143,N_29261,N_29512);
or U30144 (N_30144,N_29077,N_28381);
nand U30145 (N_30145,N_29096,N_28489);
nor U30146 (N_30146,N_29685,N_29805);
nand U30147 (N_30147,N_28359,N_29178);
nor U30148 (N_30148,N_28050,N_29505);
nor U30149 (N_30149,N_28247,N_29120);
or U30150 (N_30150,N_29243,N_28143);
nor U30151 (N_30151,N_28301,N_28646);
nand U30152 (N_30152,N_28239,N_28509);
xor U30153 (N_30153,N_28528,N_28795);
nand U30154 (N_30154,N_28156,N_28076);
and U30155 (N_30155,N_29987,N_29730);
or U30156 (N_30156,N_28644,N_29383);
nand U30157 (N_30157,N_28091,N_29063);
nand U30158 (N_30158,N_28203,N_28705);
nand U30159 (N_30159,N_29350,N_28252);
and U30160 (N_30160,N_28762,N_29034);
nor U30161 (N_30161,N_29719,N_29336);
or U30162 (N_30162,N_29048,N_28405);
or U30163 (N_30163,N_28183,N_29846);
nor U30164 (N_30164,N_29200,N_28029);
nand U30165 (N_30165,N_29870,N_28118);
nor U30166 (N_30166,N_29390,N_28582);
and U30167 (N_30167,N_29901,N_28546);
nand U30168 (N_30168,N_28984,N_29418);
nand U30169 (N_30169,N_28840,N_29495);
and U30170 (N_30170,N_28169,N_28311);
nand U30171 (N_30171,N_29412,N_29099);
or U30172 (N_30172,N_29442,N_28277);
nand U30173 (N_30173,N_29802,N_28966);
nand U30174 (N_30174,N_29571,N_29790);
or U30175 (N_30175,N_29532,N_28366);
nand U30176 (N_30176,N_28511,N_29533);
nor U30177 (N_30177,N_29408,N_28264);
and U30178 (N_30178,N_28187,N_29307);
nand U30179 (N_30179,N_29858,N_28667);
and U30180 (N_30180,N_28375,N_28630);
or U30181 (N_30181,N_28064,N_29931);
nand U30182 (N_30182,N_29607,N_29294);
and U30183 (N_30183,N_29417,N_29586);
and U30184 (N_30184,N_28898,N_29939);
and U30185 (N_30185,N_28999,N_29013);
nand U30186 (N_30186,N_29047,N_28675);
and U30187 (N_30187,N_29321,N_28867);
nand U30188 (N_30188,N_28731,N_29812);
and U30189 (N_30189,N_29185,N_29789);
and U30190 (N_30190,N_29422,N_29154);
or U30191 (N_30191,N_28579,N_29329);
nand U30192 (N_30192,N_28174,N_29763);
nor U30193 (N_30193,N_29897,N_29572);
xor U30194 (N_30194,N_28821,N_28336);
and U30195 (N_30195,N_29152,N_28973);
and U30196 (N_30196,N_28540,N_28581);
or U30197 (N_30197,N_29679,N_28779);
nor U30198 (N_30198,N_29678,N_29810);
and U30199 (N_30199,N_29921,N_29181);
nor U30200 (N_30200,N_28883,N_28207);
nand U30201 (N_30201,N_28665,N_29781);
nor U30202 (N_30202,N_28933,N_29198);
nand U30203 (N_30203,N_28949,N_28890);
or U30204 (N_30204,N_29330,N_29242);
nand U30205 (N_30205,N_28742,N_29999);
nand U30206 (N_30206,N_28357,N_28364);
nand U30207 (N_30207,N_29797,N_28427);
or U30208 (N_30208,N_29339,N_29903);
nor U30209 (N_30209,N_29323,N_28211);
or U30210 (N_30210,N_28234,N_28932);
nor U30211 (N_30211,N_29104,N_28610);
nand U30212 (N_30212,N_29474,N_29909);
and U30213 (N_30213,N_28176,N_29302);
or U30214 (N_30214,N_29290,N_28959);
nand U30215 (N_30215,N_28363,N_28946);
nor U30216 (N_30216,N_29381,N_29966);
and U30217 (N_30217,N_29484,N_29503);
and U30218 (N_30218,N_28823,N_29861);
nor U30219 (N_30219,N_29132,N_28015);
nor U30220 (N_30220,N_29202,N_29876);
nand U30221 (N_30221,N_28902,N_28908);
or U30222 (N_30222,N_28549,N_29717);
and U30223 (N_30223,N_28673,N_29742);
or U30224 (N_30224,N_29945,N_28312);
nor U30225 (N_30225,N_28000,N_28554);
and U30226 (N_30226,N_28339,N_29428);
nand U30227 (N_30227,N_29150,N_29410);
nor U30228 (N_30228,N_29039,N_29326);
nand U30229 (N_30229,N_29064,N_29136);
xnor U30230 (N_30230,N_29733,N_28637);
nand U30231 (N_30231,N_29380,N_28434);
or U30232 (N_30232,N_29643,N_28668);
or U30233 (N_30233,N_28349,N_28774);
and U30234 (N_30234,N_28199,N_29788);
nor U30235 (N_30235,N_29979,N_29806);
or U30236 (N_30236,N_28124,N_28274);
nor U30237 (N_30237,N_28555,N_28736);
nor U30238 (N_30238,N_29456,N_28164);
or U30239 (N_30239,N_29915,N_29758);
nor U30240 (N_30240,N_28165,N_28472);
nand U30241 (N_30241,N_29873,N_29414);
or U30242 (N_30242,N_28729,N_28745);
and U30243 (N_30243,N_29280,N_29088);
xnor U30244 (N_30244,N_28115,N_28329);
nand U30245 (N_30245,N_29522,N_28197);
nand U30246 (N_30246,N_29845,N_28149);
or U30247 (N_30247,N_29221,N_28443);
or U30248 (N_30248,N_28026,N_28759);
or U30249 (N_30249,N_29389,N_29406);
and U30250 (N_30250,N_29165,N_29684);
nor U30251 (N_30251,N_29320,N_28418);
nand U30252 (N_30252,N_28512,N_29282);
nor U30253 (N_30253,N_29552,N_29098);
nor U30254 (N_30254,N_28020,N_28683);
nand U30255 (N_30255,N_29993,N_29044);
and U30256 (N_30256,N_28802,N_28809);
or U30257 (N_30257,N_28590,N_29284);
nand U30258 (N_30258,N_29842,N_28226);
nor U30259 (N_30259,N_29125,N_29801);
or U30260 (N_30260,N_28805,N_28944);
and U30261 (N_30261,N_29990,N_28635);
or U30262 (N_30262,N_28500,N_28834);
and U30263 (N_30263,N_29547,N_28222);
or U30264 (N_30264,N_28323,N_29655);
or U30265 (N_30265,N_29940,N_29086);
or U30266 (N_30266,N_29538,N_28229);
or U30267 (N_30267,N_28367,N_29254);
nor U30268 (N_30268,N_29054,N_29189);
and U30269 (N_30269,N_29046,N_29919);
nand U30270 (N_30270,N_28424,N_28151);
nand U30271 (N_30271,N_29392,N_28454);
and U30272 (N_30272,N_29215,N_28884);
nand U30273 (N_30273,N_29567,N_29767);
or U30274 (N_30274,N_29947,N_29450);
and U30275 (N_30275,N_28351,N_28235);
nor U30276 (N_30276,N_29526,N_29158);
or U30277 (N_30277,N_28083,N_29738);
nor U30278 (N_30278,N_29451,N_28992);
nand U30279 (N_30279,N_29188,N_29396);
or U30280 (N_30280,N_28284,N_28965);
and U30281 (N_30281,N_28826,N_28738);
or U30282 (N_30282,N_28473,N_29265);
nand U30283 (N_30283,N_29424,N_29531);
xor U30284 (N_30284,N_28954,N_28775);
nor U30285 (N_30285,N_28464,N_29301);
and U30286 (N_30286,N_29482,N_29693);
or U30287 (N_30287,N_28138,N_29886);
or U30288 (N_30288,N_28444,N_28039);
and U30289 (N_30289,N_29159,N_28440);
xnor U30290 (N_30290,N_28152,N_28664);
or U30291 (N_30291,N_28893,N_28592);
and U30292 (N_30292,N_28455,N_29619);
nand U30293 (N_30293,N_29967,N_29796);
nand U30294 (N_30294,N_28837,N_28526);
nand U30295 (N_30295,N_29637,N_29653);
nor U30296 (N_30296,N_29944,N_29394);
and U30297 (N_30297,N_29035,N_28981);
nand U30298 (N_30298,N_29694,N_29725);
nor U30299 (N_30299,N_28934,N_29885);
nand U30300 (N_30300,N_29565,N_29421);
and U30301 (N_30301,N_29364,N_29895);
nor U30302 (N_30302,N_28393,N_28119);
nor U30303 (N_30303,N_28679,N_29866);
nand U30304 (N_30304,N_29398,N_28463);
nand U30305 (N_30305,N_29804,N_29601);
nor U30306 (N_30306,N_28043,N_28692);
nor U30307 (N_30307,N_29235,N_28184);
nor U30308 (N_30308,N_28468,N_29065);
nor U30309 (N_30309,N_28924,N_28501);
nand U30310 (N_30310,N_28938,N_29366);
nor U30311 (N_30311,N_28642,N_28342);
nand U30312 (N_30312,N_28798,N_28939);
or U30313 (N_30313,N_29014,N_29193);
nor U30314 (N_30314,N_29798,N_29577);
nor U30315 (N_30315,N_28626,N_28586);
nand U30316 (N_30316,N_29859,N_29819);
and U30317 (N_30317,N_29935,N_28678);
nor U30318 (N_30318,N_28404,N_28215);
nand U30319 (N_30319,N_28302,N_28780);
or U30320 (N_30320,N_28397,N_28797);
and U30321 (N_30321,N_28389,N_28694);
and U30322 (N_30322,N_29195,N_28778);
xnor U30323 (N_30323,N_28003,N_28585);
xnor U30324 (N_30324,N_29030,N_28421);
and U30325 (N_30325,N_28040,N_28700);
nor U30326 (N_30326,N_28728,N_29545);
and U30327 (N_30327,N_29105,N_28707);
and U30328 (N_30328,N_28068,N_28519);
nor U30329 (N_30329,N_29537,N_28520);
nor U30330 (N_30330,N_28570,N_29701);
and U30331 (N_30331,N_29510,N_28727);
or U30332 (N_30332,N_29433,N_28245);
nor U30333 (N_30333,N_29605,N_28882);
nor U30334 (N_30334,N_28597,N_29555);
nand U30335 (N_30335,N_28906,N_29068);
nor U30336 (N_30336,N_28483,N_28534);
and U30337 (N_30337,N_29183,N_29743);
or U30338 (N_30338,N_29016,N_29658);
nand U30339 (N_30339,N_28522,N_29628);
nand U30340 (N_30340,N_28052,N_29911);
nor U30341 (N_30341,N_28401,N_28539);
or U30342 (N_30342,N_29896,N_29184);
nand U30343 (N_30343,N_28792,N_28887);
nand U30344 (N_30344,N_29388,N_29449);
xnor U30345 (N_30345,N_28408,N_29862);
or U30346 (N_30346,N_28975,N_29766);
and U30347 (N_30347,N_28018,N_29349);
nor U30348 (N_30348,N_28009,N_29711);
nor U30349 (N_30349,N_28072,N_29578);
or U30350 (N_30350,N_28200,N_29667);
and U30351 (N_30351,N_28283,N_29022);
nor U30352 (N_30352,N_29949,N_28769);
nor U30353 (N_30353,N_29287,N_28261);
nor U30354 (N_30354,N_29980,N_29663);
or U30355 (N_30355,N_29107,N_28061);
or U30356 (N_30356,N_28021,N_29080);
nand U30357 (N_30357,N_28192,N_28110);
nor U30358 (N_30358,N_29925,N_29258);
nor U30359 (N_30359,N_28764,N_29479);
or U30360 (N_30360,N_29544,N_29775);
nand U30361 (N_30361,N_29648,N_29268);
or U30362 (N_30362,N_29783,N_29878);
or U30363 (N_30363,N_29837,N_28327);
nor U30364 (N_30364,N_29891,N_28417);
or U30365 (N_30365,N_28825,N_28848);
and U30366 (N_30366,N_29430,N_28221);
nor U30367 (N_30367,N_29962,N_29900);
or U30368 (N_30368,N_29140,N_29602);
or U30369 (N_30369,N_28022,N_29003);
or U30370 (N_30370,N_28280,N_28204);
or U30371 (N_30371,N_29839,N_29121);
nand U30372 (N_30372,N_28943,N_28624);
nand U30373 (N_30373,N_28132,N_29288);
nor U30374 (N_30374,N_29405,N_29210);
nand U30375 (N_30375,N_29640,N_29073);
or U30376 (N_30376,N_29793,N_29702);
and U30377 (N_30377,N_28952,N_28494);
nand U30378 (N_30378,N_28101,N_28550);
nor U30379 (N_30379,N_28598,N_29613);
or U30380 (N_30380,N_29434,N_28153);
nand U30381 (N_30381,N_29724,N_28623);
nand U30382 (N_30382,N_28693,N_28508);
nand U30383 (N_30383,N_29562,N_28785);
or U30384 (N_30384,N_29727,N_29238);
and U30385 (N_30385,N_29204,N_29056);
xor U30386 (N_30386,N_28876,N_29753);
nor U30387 (N_30387,N_29934,N_28543);
or U30388 (N_30388,N_28862,N_29587);
and U30389 (N_30389,N_29436,N_29612);
nor U30390 (N_30390,N_29807,N_29965);
or U30391 (N_30391,N_28530,N_28282);
nand U30392 (N_30392,N_29982,N_28889);
and U30393 (N_30393,N_28716,N_28097);
nor U30394 (N_30394,N_28308,N_29854);
and U30395 (N_30395,N_28746,N_28594);
nor U30396 (N_30396,N_28386,N_28645);
or U30397 (N_30397,N_29081,N_29413);
or U30398 (N_30398,N_28711,N_29536);
and U30399 (N_30399,N_29423,N_29465);
nand U30400 (N_30400,N_28136,N_29978);
and U30401 (N_30401,N_29907,N_29160);
and U30402 (N_30402,N_29872,N_29403);
nor U30403 (N_30403,N_28107,N_28621);
nor U30404 (N_30404,N_28071,N_28783);
nand U30405 (N_30405,N_29008,N_29025);
or U30406 (N_30406,N_28913,N_29084);
nand U30407 (N_30407,N_29362,N_29657);
nand U30408 (N_30408,N_29848,N_28079);
and U30409 (N_30409,N_29466,N_29341);
and U30410 (N_30410,N_29737,N_29236);
nand U30411 (N_30411,N_28333,N_28537);
nor U30412 (N_30412,N_28027,N_28743);
nand U30413 (N_30413,N_29169,N_28744);
and U30414 (N_30414,N_29554,N_28925);
or U30415 (N_30415,N_29898,N_29219);
nor U30416 (N_30416,N_28047,N_29974);
or U30417 (N_30417,N_28752,N_29528);
and U30418 (N_30418,N_29654,N_29969);
or U30419 (N_30419,N_29757,N_29246);
nand U30420 (N_30420,N_29656,N_29440);
and U30421 (N_30421,N_28158,N_29151);
and U30422 (N_30422,N_28684,N_29173);
or U30423 (N_30423,N_29524,N_28710);
nor U30424 (N_30424,N_29431,N_29066);
and U30425 (N_30425,N_28328,N_29660);
nor U30426 (N_30426,N_28314,N_29278);
nor U30427 (N_30427,N_29633,N_29076);
and U30428 (N_30428,N_29563,N_28017);
nand U30429 (N_30429,N_29062,N_29457);
nor U30430 (N_30430,N_29735,N_28904);
nor U30431 (N_30431,N_29373,N_28654);
and U30432 (N_30432,N_28104,N_28249);
nand U30433 (N_30433,N_29163,N_29289);
nand U30434 (N_30434,N_29058,N_28618);
nand U30435 (N_30435,N_29816,N_28753);
nand U30436 (N_30436,N_28270,N_28595);
nand U30437 (N_30437,N_29708,N_28269);
or U30438 (N_30438,N_29253,N_28206);
nand U30439 (N_30439,N_29715,N_29695);
nand U30440 (N_30440,N_29166,N_29292);
or U30441 (N_30441,N_28388,N_29776);
nand U30442 (N_30442,N_28816,N_28411);
or U30443 (N_30443,N_28332,N_28620);
nor U30444 (N_30444,N_29853,N_28117);
or U30445 (N_30445,N_29051,N_28121);
nand U30446 (N_30446,N_29649,N_28246);
and U30447 (N_30447,N_28915,N_29055);
or U30448 (N_30448,N_29588,N_28688);
nor U30449 (N_30449,N_28310,N_29028);
or U30450 (N_30450,N_28631,N_29824);
nor U30451 (N_30451,N_29959,N_28827);
nand U30452 (N_30452,N_29283,N_28863);
and U30453 (N_30453,N_28799,N_29622);
nand U30454 (N_30454,N_29827,N_29213);
nand U30455 (N_30455,N_28676,N_28069);
or U30456 (N_30456,N_29225,N_28190);
nor U30457 (N_30457,N_29475,N_29129);
or U30458 (N_30458,N_29196,N_28036);
nand U30459 (N_30459,N_28392,N_29543);
or U30460 (N_30460,N_29860,N_28482);
nand U30461 (N_30461,N_29666,N_29550);
nand U30462 (N_30462,N_29256,N_29517);
nand U30463 (N_30463,N_28749,N_29374);
nand U30464 (N_30464,N_29342,N_29199);
nor U30465 (N_30465,N_28492,N_29266);
nand U30466 (N_30466,N_29006,N_29255);
nor U30467 (N_30467,N_28172,N_28056);
and U30468 (N_30468,N_28703,N_28704);
nor U30469 (N_30469,N_29083,N_29143);
or U30470 (N_30470,N_28317,N_28495);
nand U30471 (N_30471,N_28875,N_29122);
or U30472 (N_30472,N_29749,N_29750);
and U30473 (N_30473,N_28319,N_28578);
nor U30474 (N_30474,N_28111,N_29892);
and U30475 (N_30475,N_28002,N_29324);
nand U30476 (N_30476,N_29500,N_28831);
or U30477 (N_30477,N_29670,N_28601);
or U30478 (N_30478,N_28343,N_29918);
and U30479 (N_30479,N_29443,N_29850);
nand U30480 (N_30480,N_28423,N_29765);
or U30481 (N_30481,N_28812,N_29399);
nand U30482 (N_30482,N_28671,N_28962);
and U30483 (N_30483,N_29933,N_28955);
and U30484 (N_30484,N_28599,N_28242);
or U30485 (N_30485,N_28060,N_29913);
nor U30486 (N_30486,N_28961,N_28860);
nor U30487 (N_30487,N_28128,N_28402);
or U30488 (N_30488,N_28516,N_28672);
nand U30489 (N_30489,N_29228,N_29604);
nand U30490 (N_30490,N_28089,N_29446);
nor U30491 (N_30491,N_29795,N_29920);
nor U30492 (N_30492,N_29368,N_28565);
and U30493 (N_30493,N_28175,N_29676);
and U30494 (N_30494,N_28373,N_29464);
nor U30495 (N_30495,N_28498,N_29187);
nand U30496 (N_30496,N_29297,N_29492);
and U30497 (N_30497,N_29638,N_29662);
and U30498 (N_30498,N_29722,N_28086);
nor U30499 (N_30499,N_29985,N_28756);
xnor U30500 (N_30500,N_29723,N_28196);
nor U30501 (N_30501,N_29114,N_28577);
or U30502 (N_30502,N_29369,N_28263);
or U30503 (N_30503,N_28538,N_29340);
xor U30504 (N_30504,N_28681,N_29271);
nand U30505 (N_30505,N_29843,N_28929);
nor U30506 (N_30506,N_28067,N_28046);
nand U30507 (N_30507,N_29067,N_28362);
or U30508 (N_30508,N_29771,N_29904);
or U30509 (N_30509,N_29180,N_28428);
or U30510 (N_30510,N_29518,N_28739);
or U30511 (N_30511,N_28399,N_29343);
nand U30512 (N_30512,N_29370,N_29905);
or U30513 (N_30513,N_28695,N_29346);
and U30514 (N_30514,N_29071,N_29448);
nand U30515 (N_30515,N_29462,N_29785);
nor U30516 (N_30516,N_29375,N_28847);
and U30517 (N_30517,N_28872,N_28462);
nor U30518 (N_30518,N_29247,N_29946);
or U30519 (N_30519,N_28789,N_28659);
nand U30520 (N_30520,N_29871,N_28801);
nand U30521 (N_30521,N_28708,N_29435);
nor U30522 (N_30522,N_28562,N_28177);
nor U30523 (N_30523,N_28171,N_28041);
or U30524 (N_30524,N_29739,N_28643);
nor U30525 (N_30525,N_29616,N_29879);
and U30526 (N_30526,N_29354,N_28497);
and U30527 (N_30527,N_28613,N_28105);
xor U30528 (N_30528,N_28532,N_28057);
nor U30529 (N_30529,N_29890,N_29664);
nand U30530 (N_30530,N_28853,N_28293);
and U30531 (N_30531,N_29049,N_28008);
and U30532 (N_30532,N_28917,N_28918);
xor U30533 (N_30533,N_29110,N_29041);
and U30534 (N_30534,N_28490,N_29480);
nand U30535 (N_30535,N_28571,N_28515);
or U30536 (N_30536,N_28238,N_28123);
or U30537 (N_30537,N_28480,N_28034);
nor U30538 (N_30538,N_29787,N_28236);
nor U30539 (N_30539,N_28033,N_29762);
and U30540 (N_30540,N_28614,N_28383);
or U30541 (N_30541,N_29141,N_29932);
or U30542 (N_30542,N_28901,N_29857);
and U30543 (N_30543,N_28751,N_29831);
and U30544 (N_30544,N_29111,N_29761);
and U30545 (N_30545,N_29748,N_28084);
nand U30546 (N_30546,N_28305,N_28819);
nand U30547 (N_30547,N_29497,N_28275);
and U30548 (N_30548,N_29696,N_28287);
nand U30549 (N_30549,N_28281,N_28810);
nand U30550 (N_30550,N_29815,N_29155);
nor U30551 (N_30551,N_29777,N_28794);
nor U30552 (N_30552,N_28722,N_29610);
nand U30553 (N_30553,N_29257,N_28513);
nand U30554 (N_30554,N_29004,N_28972);
nor U30555 (N_30555,N_29220,N_29472);
or U30556 (N_30556,N_29162,N_29961);
and U30557 (N_30557,N_28055,N_28460);
or U30558 (N_30558,N_29274,N_28669);
nor U30559 (N_30559,N_28070,N_28603);
or U30560 (N_30560,N_28407,N_29740);
or U30561 (N_30561,N_28575,N_28670);
nor U30562 (N_30562,N_29305,N_28914);
nor U30563 (N_30563,N_28467,N_29566);
nand U30564 (N_30564,N_29337,N_28639);
nor U30565 (N_30565,N_29400,N_28653);
nor U30566 (N_30566,N_29331,N_28950);
nor U30567 (N_30567,N_28502,N_28770);
or U30568 (N_30568,N_29608,N_28721);
or U30569 (N_30569,N_28713,N_29635);
nand U30570 (N_30570,N_28456,N_29425);
or U30571 (N_30571,N_29712,N_28391);
or U30572 (N_30572,N_28450,N_28718);
and U30573 (N_30573,N_29888,N_29665);
and U30574 (N_30574,N_29347,N_29452);
nor U30575 (N_30575,N_29355,N_29296);
or U30576 (N_30576,N_29304,N_29794);
nand U30577 (N_30577,N_29397,N_29322);
and U30578 (N_30578,N_28622,N_28786);
nand U30579 (N_30579,N_29856,N_29244);
nand U30580 (N_30580,N_29924,N_28701);
nand U30581 (N_30581,N_28589,N_28894);
and U30582 (N_30582,N_28566,N_29519);
nor U30583 (N_30583,N_29700,N_29623);
and U30584 (N_30584,N_29792,N_29118);
nor U30585 (N_30585,N_29832,N_28865);
nand U30586 (N_30586,N_28523,N_29770);
or U30587 (N_30587,N_29902,N_28940);
and U30588 (N_30588,N_28584,N_29865);
or U30589 (N_30589,N_29432,N_28871);
nor U30590 (N_30590,N_29799,N_28148);
and U30591 (N_30591,N_28188,N_29937);
and U30592 (N_30592,N_29916,N_28800);
and U30593 (N_30593,N_29690,N_28088);
or U30594 (N_30594,N_28536,N_28262);
nand U30595 (N_30595,N_28748,N_29353);
and U30596 (N_30596,N_28023,N_29299);
nor U30597 (N_30597,N_29191,N_29395);
nand U30598 (N_30598,N_28186,N_29363);
xnor U30599 (N_30599,N_28031,N_29259);
nor U30600 (N_30600,N_29529,N_28442);
and U30601 (N_30601,N_29174,N_28650);
and U30602 (N_30602,N_28116,N_29303);
nor U30603 (N_30603,N_29631,N_29617);
and U30604 (N_30604,N_28838,N_28771);
and U30605 (N_30605,N_29277,N_29504);
nor U30606 (N_30606,N_29379,N_28996);
nor U30607 (N_30607,N_29883,N_28168);
and U30608 (N_30608,N_28878,N_29409);
and U30609 (N_30609,N_29208,N_28338);
and U30610 (N_30610,N_29559,N_28967);
nor U30611 (N_30611,N_29928,N_29333);
nand U30612 (N_30612,N_29420,N_28157);
nand U30613 (N_30613,N_29240,N_29126);
nor U30614 (N_30614,N_28477,N_29836);
nor U30615 (N_30615,N_28852,N_28699);
nor U30616 (N_30616,N_28337,N_29043);
nand U30617 (N_30617,N_29721,N_28833);
nand U30618 (N_30618,N_28451,N_29953);
and U30619 (N_30619,N_28145,N_28757);
or U30620 (N_30620,N_29108,N_29535);
nor U30621 (N_30621,N_29645,N_29045);
or U30622 (N_30622,N_29882,N_28619);
nand U30623 (N_30623,N_29755,N_29596);
and U30624 (N_30624,N_28390,N_28059);
nor U30625 (N_30625,N_29912,N_28290);
nand U30626 (N_30626,N_29000,N_28518);
nand U30627 (N_30627,N_28942,N_29838);
and U30628 (N_30628,N_29549,N_29216);
nor U30629 (N_30629,N_29082,N_28503);
or U30630 (N_30630,N_28677,N_28232);
nand U30631 (N_30631,N_28935,N_28228);
and U30632 (N_30632,N_28958,N_29441);
and U30633 (N_30633,N_28517,N_28763);
xor U30634 (N_30634,N_28606,N_29772);
nand U30635 (N_30635,N_28617,N_29416);
nor U30636 (N_30636,N_28628,N_29736);
or U30637 (N_30637,N_28991,N_29387);
nor U30638 (N_30638,N_29960,N_29851);
nand U30639 (N_30639,N_29823,N_28964);
nand U30640 (N_30640,N_29754,N_28102);
and U30641 (N_30641,N_28045,N_29027);
and U30642 (N_30642,N_29548,N_28007);
nor U30643 (N_30643,N_28881,N_29661);
nor U30644 (N_30644,N_29514,N_29102);
and U30645 (N_30645,N_28396,N_28979);
nor U30646 (N_30646,N_28352,N_29206);
or U30647 (N_30647,N_29541,N_28094);
nand U30648 (N_30648,N_28896,N_28560);
nand U30649 (N_30649,N_29948,N_29952);
or U30650 (N_30650,N_29097,N_29176);
or U30651 (N_30651,N_29359,N_28265);
or U30652 (N_30652,N_28968,N_29906);
or U30653 (N_30653,N_29976,N_28413);
or U30654 (N_30654,N_29371,N_28403);
and U30655 (N_30655,N_29553,N_28573);
nor U30656 (N_30656,N_29508,N_29975);
or U30657 (N_30657,N_28385,N_28212);
and U30658 (N_30658,N_29991,N_29033);
nand U30659 (N_30659,N_29298,N_28732);
nand U30660 (N_30660,N_28824,N_29164);
and U30661 (N_30661,N_28828,N_28796);
nor U30662 (N_30662,N_29205,N_29936);
nand U30663 (N_30663,N_29426,N_28445);
or U30664 (N_30664,N_28719,N_28557);
xor U30665 (N_30665,N_28723,N_29295);
and U30666 (N_30666,N_28330,N_28433);
nand U30667 (N_30667,N_29059,N_28734);
nor U30668 (N_30668,N_28346,N_28340);
or U30669 (N_30669,N_29597,N_29012);
nand U30670 (N_30670,N_29632,N_28024);
or U30671 (N_30671,N_29938,N_29032);
or U30672 (N_30672,N_29546,N_28019);
xor U30673 (N_30673,N_29681,N_28044);
and U30674 (N_30674,N_28368,N_28106);
and U30675 (N_30675,N_29813,N_28970);
nand U30676 (N_30676,N_28276,N_29308);
nor U30677 (N_30677,N_29615,N_28325);
or U30678 (N_30678,N_28977,N_28218);
nand U30679 (N_30679,N_28986,N_28461);
nand U30680 (N_30680,N_29001,N_28354);
nor U30681 (N_30681,N_29250,N_29644);
and U30682 (N_30682,N_29989,N_28814);
and U30683 (N_30683,N_28189,N_29300);
and U30684 (N_30684,N_29671,N_28344);
nand U30685 (N_30685,N_28702,N_28013);
or U30686 (N_30686,N_29509,N_28303);
nand U30687 (N_30687,N_29179,N_28470);
and U30688 (N_30688,N_28371,N_29021);
nand U30689 (N_30689,N_28905,N_28499);
nand U30690 (N_30690,N_29453,N_28854);
or U30691 (N_30691,N_29172,N_28297);
nand U30692 (N_30692,N_29691,N_29651);
or U30693 (N_30693,N_28612,N_28167);
and U30694 (N_30694,N_28360,N_29720);
or U30695 (N_30695,N_29988,N_29556);
and U30696 (N_30696,N_29502,N_28633);
nand U30697 (N_30697,N_28661,N_28698);
or U30698 (N_30698,N_29732,N_28945);
and U30699 (N_30699,N_28976,N_29849);
nand U30700 (N_30700,N_29585,N_28998);
and U30701 (N_30701,N_28201,N_28466);
nor U30702 (N_30702,N_29968,N_29123);
nand U30703 (N_30703,N_28980,N_28974);
nand U30704 (N_30704,N_29010,N_29970);
or U30705 (N_30705,N_29593,N_28155);
xor U30706 (N_30706,N_29501,N_29714);
nand U30707 (N_30707,N_29252,N_29943);
nand U30708 (N_30708,N_29697,N_28006);
nor U30709 (N_30709,N_29090,N_28806);
nor U30710 (N_30710,N_28533,N_28781);
nor U30711 (N_30711,N_29625,N_29175);
nor U30712 (N_30712,N_28398,N_28258);
and U30713 (N_30713,N_28607,N_28811);
and U30714 (N_30714,N_29614,N_28474);
and U30715 (N_30715,N_29481,N_28267);
nor U30716 (N_30716,N_29139,N_28251);
nor U30717 (N_30717,N_29729,N_28982);
and U30718 (N_30718,N_28237,N_28288);
and U30719 (N_30719,N_29477,N_29087);
nor U30720 (N_30720,N_28092,N_28358);
or U30721 (N_30721,N_28134,N_28928);
nor U30722 (N_30722,N_29402,N_29874);
nand U30723 (N_30723,N_28099,N_28425);
nand U30724 (N_30724,N_29209,N_29057);
or U30725 (N_30725,N_29312,N_28035);
or U30726 (N_30726,N_29458,N_28773);
xor U30727 (N_30727,N_28160,N_29241);
and U30728 (N_30728,N_28378,N_28983);
and U30729 (N_30729,N_28075,N_29826);
or U30730 (N_30730,N_28374,N_28248);
nor U30731 (N_30731,N_28437,N_29779);
and U30732 (N_30732,N_29197,N_29820);
nor U30733 (N_30733,N_29182,N_29647);
nor U30734 (N_30734,N_29950,N_29031);
nor U30735 (N_30735,N_28995,N_29569);
nand U30736 (N_30736,N_28077,N_28244);
or U30737 (N_30737,N_28395,N_29835);
xnor U30738 (N_30738,N_28198,N_28476);
xnor U30739 (N_30739,N_29941,N_28531);
nor U30740 (N_30740,N_28514,N_28051);
or U30741 (N_30741,N_28829,N_28146);
nor U30742 (N_30742,N_28580,N_29131);
nor U30743 (N_30743,N_29317,N_28163);
or U30744 (N_30744,N_28548,N_28651);
nor U30745 (N_30745,N_29557,N_29351);
xor U30746 (N_30746,N_28815,N_28331);
or U30747 (N_30747,N_29828,N_28161);
and U30748 (N_30748,N_28568,N_28306);
nor U30749 (N_30749,N_29668,N_29007);
nand U30750 (N_30750,N_29611,N_29592);
nand U30751 (N_30751,N_29618,N_28230);
or U30752 (N_30752,N_29318,N_29207);
or U30753 (N_30753,N_28253,N_28930);
and U30754 (N_30754,N_28356,N_29551);
nor U30755 (N_30755,N_29018,N_29437);
and U30756 (N_30756,N_28142,N_28048);
nand U30757 (N_30757,N_28558,N_28969);
nand U30758 (N_30758,N_28960,N_29493);
or U30759 (N_30759,N_28085,N_29214);
or U30760 (N_30760,N_29231,N_29534);
and U30761 (N_30761,N_29620,N_29927);
nand U30762 (N_30762,N_29245,N_28772);
and U30763 (N_30763,N_28202,N_28545);
and U30764 (N_30764,N_28803,N_29476);
or U30765 (N_30765,N_28561,N_29061);
nand U30766 (N_30766,N_29230,N_29926);
or U30767 (N_30767,N_28266,N_28291);
nand U30768 (N_30768,N_28855,N_29276);
nor U30769 (N_30769,N_29709,N_28254);
nand U30770 (N_30770,N_29203,N_29759);
or U30771 (N_30771,N_29411,N_29116);
and U30772 (N_30772,N_29429,N_29460);
and U30773 (N_30773,N_29525,N_29401);
and U30774 (N_30774,N_28535,N_29378);
or U30775 (N_30775,N_28714,N_28994);
nand U30776 (N_30776,N_29646,N_28510);
and U30777 (N_30777,N_29079,N_29194);
nand U30778 (N_30778,N_29527,N_28144);
nor U30779 (N_30779,N_29367,N_28129);
and U30780 (N_30780,N_28919,N_28180);
xor U30781 (N_30781,N_29704,N_29026);
or U30782 (N_30782,N_29539,N_28587);
or U30783 (N_30783,N_28941,N_28870);
nor U30784 (N_30784,N_28049,N_29352);
and U30785 (N_30785,N_28361,N_29211);
nor U30786 (N_30786,N_28559,N_28341);
and U30787 (N_30787,N_29168,N_28042);
and U30788 (N_30788,N_29568,N_29078);
nand U30789 (N_30789,N_28576,N_29922);
nand U30790 (N_30790,N_28012,N_29130);
nand U30791 (N_30791,N_28491,N_29910);
nand U30792 (N_30792,N_29868,N_28131);
and U30793 (N_30793,N_28844,N_28951);
nor U30794 (N_30794,N_29272,N_29530);
and U30795 (N_30795,N_28309,N_29699);
nand U30796 (N_30796,N_29344,N_29273);
and U30797 (N_30797,N_29598,N_28347);
and U30798 (N_30798,N_29705,N_29515);
nand U30799 (N_30799,N_29855,N_29249);
and U30800 (N_30800,N_29138,N_29314);
nand U30801 (N_30801,N_28697,N_28090);
and U30802 (N_30802,N_29372,N_29639);
or U30803 (N_30803,N_29177,N_28032);
nor U30804 (N_30804,N_28866,N_29877);
nor U30805 (N_30805,N_28382,N_28641);
and U30806 (N_30806,N_28469,N_29760);
nor U30807 (N_30807,N_28793,N_29574);
nor U30808 (N_30808,N_28058,N_29050);
nand U30809 (N_30809,N_29005,N_28880);
or U30810 (N_30810,N_28217,N_28377);
and U30811 (N_30811,N_29728,N_28912);
nand U30812 (N_30812,N_29774,N_28296);
nand U30813 (N_30813,N_29106,N_29328);
and U30814 (N_30814,N_28087,N_28078);
and U30815 (N_30815,N_28135,N_28066);
nand U30816 (N_30816,N_28907,N_29260);
and U30817 (N_30817,N_28758,N_29513);
nor U30818 (N_30818,N_29190,N_28567);
nor U30819 (N_30819,N_28680,N_28422);
and U30820 (N_30820,N_29998,N_29407);
or U30821 (N_30821,N_28504,N_28412);
nand U30822 (N_30822,N_29829,N_28820);
and U30823 (N_30823,N_28294,N_29626);
nand U30824 (N_30824,N_29232,N_29251);
nand U30825 (N_30825,N_28122,N_28384);
or U30826 (N_30826,N_28438,N_28127);
or U30827 (N_30827,N_28850,N_29332);
nor U30828 (N_30828,N_29313,N_29840);
nor U30829 (N_30829,N_28791,N_29112);
and U30830 (N_30830,N_29285,N_29692);
nor U30831 (N_30831,N_28126,N_28755);
and U30832 (N_30832,N_28369,N_28649);
nand U30833 (N_30833,N_29338,N_28660);
nor U30834 (N_30834,N_28014,N_29822);
and U30835 (N_30835,N_28859,N_29811);
nor U30836 (N_30836,N_29455,N_29808);
nor U30837 (N_30837,N_28268,N_28956);
and U30838 (N_30838,N_29964,N_29923);
or U30839 (N_30839,N_28685,N_29391);
or U30840 (N_30840,N_28481,N_28225);
and U30841 (N_30841,N_29764,N_29070);
nand U30842 (N_30842,N_28937,N_28615);
and U30843 (N_30843,N_29791,N_29706);
nand U30844 (N_30844,N_28858,N_28696);
nand U30845 (N_30845,N_28735,N_28150);
nor U30846 (N_30846,N_28541,N_28335);
and U30847 (N_30847,N_29192,N_29672);
nand U30848 (N_30848,N_28717,N_29017);
nand U30849 (N_30849,N_28355,N_28869);
and U30850 (N_30850,N_29963,N_28074);
or U30851 (N_30851,N_29224,N_28208);
or U30852 (N_30852,N_28596,N_29880);
or U30853 (N_30853,N_28182,N_29954);
nor U30854 (N_30854,N_28936,N_28985);
and U30855 (N_30855,N_28804,N_29262);
nor U30856 (N_30856,N_29682,N_29955);
nor U30857 (N_30857,N_29356,N_29521);
or U30858 (N_30858,N_28272,N_28897);
or U30859 (N_30859,N_28307,N_28830);
nor U30860 (N_30860,N_28569,N_28591);
nand U30861 (N_30861,N_29490,N_28130);
and U30862 (N_30862,N_29335,N_28588);
nor U30863 (N_30863,N_28922,N_29091);
and U30864 (N_30864,N_29478,N_28547);
and U30865 (N_30865,N_29523,N_29981);
and U30866 (N_30866,N_29703,N_28737);
nor U30867 (N_30867,N_29002,N_29875);
or U30868 (N_30868,N_28479,N_29584);
nor U30869 (N_30869,N_28213,N_29957);
nor U30870 (N_30870,N_28313,N_28776);
or U30871 (N_30871,N_29984,N_29516);
xnor U30872 (N_30872,N_29687,N_28864);
and U30873 (N_30873,N_28028,N_28278);
nor U30874 (N_30874,N_28856,N_29669);
nand U30875 (N_30875,N_29686,N_29485);
nand U30876 (N_30876,N_28005,N_29134);
and U30877 (N_30877,N_29074,N_28220);
xor U30878 (N_30878,N_28037,N_28652);
or U30879 (N_30879,N_29869,N_28406);
nand U30880 (N_30880,N_29291,N_29752);
nor U30881 (N_30881,N_28159,N_29147);
and U30882 (N_30882,N_28001,N_28295);
nand U30883 (N_30883,N_28885,N_29471);
nor U30884 (N_30884,N_29488,N_28414);
and U30885 (N_30885,N_28879,N_28521);
nor U30886 (N_30886,N_28572,N_29100);
nand U30887 (N_30887,N_29227,N_28108);
nand U30888 (N_30888,N_28073,N_28322);
or U30889 (N_30889,N_29606,N_29009);
nand U30890 (N_30890,N_29011,N_29841);
nand U30891 (N_30891,N_28634,N_29092);
or U30892 (N_30892,N_28767,N_29520);
or U30893 (N_30893,N_28993,N_28527);
nor U30894 (N_30894,N_28240,N_28832);
nand U30895 (N_30895,N_28724,N_28835);
or U30896 (N_30896,N_29741,N_29263);
nor U30897 (N_30897,N_29894,N_28452);
nor U30898 (N_30898,N_29847,N_29149);
nor U30899 (N_30899,N_28334,N_29784);
nand U30900 (N_30900,N_28784,N_28706);
or U30901 (N_30901,N_28321,N_28899);
and U30902 (N_30902,N_28978,N_29024);
nor U30903 (N_30903,N_29746,N_28544);
nand U30904 (N_30904,N_28822,N_28609);
nor U30905 (N_30905,N_29917,N_29852);
or U30906 (N_30906,N_28663,N_28686);
or U30907 (N_30907,N_28459,N_29956);
or U30908 (N_30908,N_29491,N_29575);
or U30909 (N_30909,N_29677,N_28109);
nand U30910 (N_30910,N_29212,N_29817);
nor U30911 (N_30911,N_28243,N_29630);
and U30912 (N_30912,N_28011,N_29834);
nand U30913 (N_30913,N_28315,N_29489);
nor U30914 (N_30914,N_28787,N_29674);
and U30915 (N_30915,N_28524,N_28081);
xor U30916 (N_30916,N_28920,N_29201);
nor U30917 (N_30917,N_28125,N_28957);
xnor U30918 (N_30918,N_28409,N_28224);
nand U30919 (N_30919,N_28846,N_29844);
nand U30920 (N_30920,N_29419,N_29494);
nor U30921 (N_30921,N_29137,N_28888);
xnor U30922 (N_30922,N_29821,N_29217);
and U30923 (N_30923,N_29641,N_28257);
and U30924 (N_30924,N_29833,N_28141);
nor U30925 (N_30925,N_29818,N_29229);
xnor U30926 (N_30926,N_28016,N_28542);
and U30927 (N_30927,N_29803,N_29311);
nand U30928 (N_30928,N_29145,N_28415);
nand U30929 (N_30929,N_28923,N_28100);
nor U30930 (N_30930,N_29315,N_28432);
and U30931 (N_30931,N_29992,N_28636);
and U30932 (N_30932,N_29496,N_28114);
or U30933 (N_30933,N_29415,N_28439);
or U30934 (N_30934,N_28916,N_28629);
and U30935 (N_30935,N_28162,N_28216);
nor U30936 (N_30936,N_28255,N_28279);
nand U30937 (N_30937,N_28604,N_29023);
nand U30938 (N_30938,N_29085,N_28990);
and U30939 (N_30939,N_28458,N_28436);
nor U30940 (N_30940,N_29506,N_29103);
or U30941 (N_30941,N_28475,N_28231);
and U30942 (N_30942,N_29591,N_28687);
nor U30943 (N_30943,N_28605,N_29348);
xnor U30944 (N_30944,N_28818,N_29447);
or U30945 (N_30945,N_29726,N_29469);
and U30946 (N_30946,N_28760,N_29929);
nand U30947 (N_30947,N_29128,N_28877);
and U30948 (N_30948,N_29889,N_29053);
nand U30949 (N_30949,N_28113,N_29486);
nor U30950 (N_30950,N_29986,N_29459);
or U30951 (N_30951,N_28747,N_28529);
nor U30952 (N_30952,N_28420,N_28926);
nand U30953 (N_30953,N_28563,N_29029);
and U30954 (N_30954,N_29275,N_28841);
and U30955 (N_30955,N_29463,N_28493);
or U30956 (N_30956,N_29914,N_28750);
nor U30957 (N_30957,N_28761,N_29745);
nand U30958 (N_30958,N_28553,N_28318);
and U30959 (N_30959,N_28921,N_28289);
nor U30960 (N_30960,N_29226,N_28365);
or U30961 (N_30961,N_28777,N_28410);
or U30962 (N_30962,N_29698,N_29439);
nand U30963 (N_30963,N_29780,N_29109);
or U30964 (N_30964,N_28030,N_29233);
or U30965 (N_30965,N_28487,N_29037);
or U30966 (N_30966,N_29958,N_29234);
and U30967 (N_30967,N_29769,N_28564);
and U30968 (N_30968,N_28909,N_29675);
and U30969 (N_30969,N_28457,N_29093);
and U30970 (N_30970,N_29996,N_29814);
xnor U30971 (N_30971,N_28911,N_28593);
nand U30972 (N_30972,N_28137,N_29576);
nand U30973 (N_30973,N_29237,N_29094);
or U30974 (N_30974,N_29884,N_28656);
and U30975 (N_30975,N_28419,N_28233);
and U30976 (N_30976,N_28147,N_29376);
nor U30977 (N_30977,N_28602,N_29334);
and U30978 (N_30978,N_29747,N_29590);
nand U30979 (N_30979,N_28507,N_28449);
or U30980 (N_30980,N_28063,N_29718);
nor U30981 (N_30981,N_28062,N_29600);
and U30982 (N_30982,N_28181,N_29020);
nand U30983 (N_30983,N_29467,N_29445);
and U30984 (N_30984,N_29599,N_29973);
nand U30985 (N_30985,N_29171,N_28209);
nor U30986 (N_30986,N_28488,N_29659);
nand U30987 (N_30987,N_29186,N_28868);
nor U30988 (N_30988,N_28726,N_28997);
and U30989 (N_30989,N_28765,N_28241);
nor U30990 (N_30990,N_28849,N_28574);
nand U30991 (N_30991,N_28471,N_29218);
nor U30992 (N_30992,N_29580,N_29239);
and U30993 (N_30993,N_29223,N_28674);
nor U30994 (N_30994,N_28139,N_28191);
or U30995 (N_30995,N_29561,N_28259);
or U30996 (N_30996,N_28525,N_28632);
nand U30997 (N_30997,N_29075,N_29095);
or U30998 (N_30998,N_28316,N_29119);
and U30999 (N_30999,N_29558,N_29887);
nand U31000 (N_31000,N_28175,N_29382);
or U31001 (N_31001,N_29357,N_29722);
or U31002 (N_31002,N_29299,N_28274);
xnor U31003 (N_31003,N_28008,N_28816);
or U31004 (N_31004,N_29897,N_29574);
and U31005 (N_31005,N_29859,N_28455);
or U31006 (N_31006,N_28042,N_29184);
nor U31007 (N_31007,N_28946,N_28681);
nand U31008 (N_31008,N_29616,N_29009);
and U31009 (N_31009,N_28255,N_28725);
and U31010 (N_31010,N_28445,N_29154);
and U31011 (N_31011,N_28113,N_29552);
or U31012 (N_31012,N_29266,N_28561);
nand U31013 (N_31013,N_28237,N_28849);
and U31014 (N_31014,N_29325,N_28853);
or U31015 (N_31015,N_28905,N_29655);
nand U31016 (N_31016,N_28438,N_28641);
nand U31017 (N_31017,N_28309,N_28935);
nand U31018 (N_31018,N_28248,N_29742);
nor U31019 (N_31019,N_28322,N_28395);
nor U31020 (N_31020,N_28531,N_29650);
nor U31021 (N_31021,N_28382,N_28164);
nand U31022 (N_31022,N_28720,N_28004);
and U31023 (N_31023,N_28554,N_29707);
and U31024 (N_31024,N_29313,N_29201);
or U31025 (N_31025,N_29073,N_28762);
and U31026 (N_31026,N_29368,N_29146);
or U31027 (N_31027,N_29803,N_28920);
and U31028 (N_31028,N_28480,N_28462);
or U31029 (N_31029,N_28370,N_28946);
or U31030 (N_31030,N_29284,N_28462);
nor U31031 (N_31031,N_28730,N_29595);
or U31032 (N_31032,N_28792,N_29259);
xor U31033 (N_31033,N_28833,N_29603);
nor U31034 (N_31034,N_28979,N_29151);
nor U31035 (N_31035,N_29375,N_28620);
nor U31036 (N_31036,N_28634,N_28094);
and U31037 (N_31037,N_28696,N_29570);
and U31038 (N_31038,N_28667,N_29665);
or U31039 (N_31039,N_29525,N_28245);
or U31040 (N_31040,N_29836,N_28460);
nor U31041 (N_31041,N_28288,N_28494);
nand U31042 (N_31042,N_28411,N_28690);
and U31043 (N_31043,N_29546,N_28677);
and U31044 (N_31044,N_29777,N_28085);
nand U31045 (N_31045,N_29218,N_28611);
nand U31046 (N_31046,N_28556,N_29274);
and U31047 (N_31047,N_29153,N_28286);
or U31048 (N_31048,N_29940,N_28832);
nand U31049 (N_31049,N_29363,N_29240);
nand U31050 (N_31050,N_29080,N_28317);
nand U31051 (N_31051,N_28853,N_28705);
or U31052 (N_31052,N_29766,N_28130);
nand U31053 (N_31053,N_28574,N_29286);
nor U31054 (N_31054,N_28344,N_28926);
nor U31055 (N_31055,N_29518,N_28244);
nand U31056 (N_31056,N_29054,N_29661);
or U31057 (N_31057,N_28619,N_28966);
nand U31058 (N_31058,N_29810,N_28372);
nor U31059 (N_31059,N_28803,N_29187);
nand U31060 (N_31060,N_28885,N_29306);
or U31061 (N_31061,N_29042,N_28929);
and U31062 (N_31062,N_28281,N_28969);
or U31063 (N_31063,N_29100,N_29608);
nand U31064 (N_31064,N_29699,N_28177);
nor U31065 (N_31065,N_29041,N_28271);
and U31066 (N_31066,N_29860,N_28119);
nor U31067 (N_31067,N_28699,N_28375);
and U31068 (N_31068,N_29014,N_29153);
or U31069 (N_31069,N_29709,N_28136);
and U31070 (N_31070,N_29954,N_29112);
or U31071 (N_31071,N_29440,N_28667);
and U31072 (N_31072,N_28883,N_28537);
and U31073 (N_31073,N_29981,N_28765);
nand U31074 (N_31074,N_29815,N_28060);
nand U31075 (N_31075,N_29784,N_29636);
and U31076 (N_31076,N_28340,N_28767);
and U31077 (N_31077,N_29105,N_29113);
or U31078 (N_31078,N_28384,N_28931);
and U31079 (N_31079,N_29093,N_29763);
nand U31080 (N_31080,N_29240,N_29377);
and U31081 (N_31081,N_28369,N_28817);
or U31082 (N_31082,N_28633,N_28902);
or U31083 (N_31083,N_29281,N_29949);
or U31084 (N_31084,N_29550,N_28533);
nand U31085 (N_31085,N_28285,N_28768);
or U31086 (N_31086,N_28515,N_28959);
or U31087 (N_31087,N_28809,N_29401);
nor U31088 (N_31088,N_28062,N_28599);
nor U31089 (N_31089,N_29969,N_28268);
and U31090 (N_31090,N_29093,N_29285);
nand U31091 (N_31091,N_29157,N_29260);
nor U31092 (N_31092,N_28536,N_28159);
nand U31093 (N_31093,N_28199,N_29152);
nand U31094 (N_31094,N_29822,N_29333);
and U31095 (N_31095,N_28630,N_29535);
nand U31096 (N_31096,N_28888,N_29865);
or U31097 (N_31097,N_28568,N_28065);
nor U31098 (N_31098,N_28617,N_28526);
or U31099 (N_31099,N_29613,N_28499);
nand U31100 (N_31100,N_28841,N_28792);
nor U31101 (N_31101,N_28129,N_29093);
nand U31102 (N_31102,N_29988,N_29867);
nand U31103 (N_31103,N_28743,N_28652);
and U31104 (N_31104,N_28007,N_29136);
or U31105 (N_31105,N_28538,N_28663);
nand U31106 (N_31106,N_29709,N_28589);
nand U31107 (N_31107,N_28180,N_28779);
or U31108 (N_31108,N_29019,N_29710);
and U31109 (N_31109,N_29826,N_29810);
xor U31110 (N_31110,N_29330,N_28401);
and U31111 (N_31111,N_28700,N_28198);
xor U31112 (N_31112,N_29100,N_29854);
nor U31113 (N_31113,N_28143,N_29318);
nand U31114 (N_31114,N_28917,N_29710);
nand U31115 (N_31115,N_29457,N_29823);
nor U31116 (N_31116,N_28241,N_28793);
nor U31117 (N_31117,N_28219,N_29722);
and U31118 (N_31118,N_28043,N_28068);
nor U31119 (N_31119,N_28955,N_29011);
or U31120 (N_31120,N_29119,N_29903);
nor U31121 (N_31121,N_28466,N_28072);
or U31122 (N_31122,N_29267,N_28564);
nand U31123 (N_31123,N_28756,N_29092);
and U31124 (N_31124,N_29270,N_28934);
nand U31125 (N_31125,N_29624,N_29503);
nand U31126 (N_31126,N_29121,N_28296);
nor U31127 (N_31127,N_29612,N_28543);
nand U31128 (N_31128,N_28215,N_28996);
nor U31129 (N_31129,N_29668,N_28412);
nor U31130 (N_31130,N_28353,N_29570);
nand U31131 (N_31131,N_29120,N_28944);
and U31132 (N_31132,N_28777,N_28322);
nand U31133 (N_31133,N_28139,N_29600);
or U31134 (N_31134,N_29851,N_28553);
nor U31135 (N_31135,N_28938,N_29555);
nand U31136 (N_31136,N_29962,N_29837);
nand U31137 (N_31137,N_29521,N_29415);
nand U31138 (N_31138,N_28834,N_28183);
and U31139 (N_31139,N_29509,N_28606);
and U31140 (N_31140,N_28045,N_28541);
and U31141 (N_31141,N_28829,N_28000);
or U31142 (N_31142,N_28060,N_28575);
or U31143 (N_31143,N_28279,N_28498);
nand U31144 (N_31144,N_28924,N_29420);
nand U31145 (N_31145,N_29348,N_29043);
nor U31146 (N_31146,N_28646,N_29462);
and U31147 (N_31147,N_28018,N_29751);
and U31148 (N_31148,N_28635,N_29517);
nand U31149 (N_31149,N_29554,N_29069);
and U31150 (N_31150,N_29925,N_29725);
nor U31151 (N_31151,N_29791,N_29110);
and U31152 (N_31152,N_28708,N_29515);
nor U31153 (N_31153,N_29012,N_28267);
or U31154 (N_31154,N_28518,N_29518);
nand U31155 (N_31155,N_28702,N_29412);
or U31156 (N_31156,N_28367,N_28623);
nand U31157 (N_31157,N_29852,N_29351);
or U31158 (N_31158,N_28045,N_28072);
and U31159 (N_31159,N_28889,N_29349);
nor U31160 (N_31160,N_28757,N_28085);
xnor U31161 (N_31161,N_29805,N_29668);
and U31162 (N_31162,N_29978,N_29870);
or U31163 (N_31163,N_29419,N_28116);
nor U31164 (N_31164,N_28146,N_28803);
xnor U31165 (N_31165,N_29712,N_29973);
nor U31166 (N_31166,N_29059,N_28811);
nor U31167 (N_31167,N_28178,N_29921);
nor U31168 (N_31168,N_28018,N_29769);
or U31169 (N_31169,N_28952,N_29270);
nor U31170 (N_31170,N_29621,N_28682);
nand U31171 (N_31171,N_28376,N_29708);
or U31172 (N_31172,N_28176,N_28040);
nor U31173 (N_31173,N_28439,N_29497);
nand U31174 (N_31174,N_28275,N_29703);
nor U31175 (N_31175,N_28969,N_29404);
or U31176 (N_31176,N_29085,N_28220);
nor U31177 (N_31177,N_28743,N_28994);
or U31178 (N_31178,N_29395,N_29148);
or U31179 (N_31179,N_28672,N_29750);
nor U31180 (N_31180,N_29271,N_29855);
or U31181 (N_31181,N_28374,N_29662);
or U31182 (N_31182,N_28612,N_29226);
and U31183 (N_31183,N_28351,N_28694);
or U31184 (N_31184,N_28569,N_28203);
nand U31185 (N_31185,N_28358,N_28958);
and U31186 (N_31186,N_28943,N_29673);
and U31187 (N_31187,N_28773,N_29973);
nor U31188 (N_31188,N_28564,N_28896);
nand U31189 (N_31189,N_29181,N_29654);
nand U31190 (N_31190,N_28507,N_28889);
nor U31191 (N_31191,N_29346,N_28991);
or U31192 (N_31192,N_28691,N_29541);
nand U31193 (N_31193,N_28647,N_28821);
nor U31194 (N_31194,N_29930,N_29637);
and U31195 (N_31195,N_28966,N_28628);
and U31196 (N_31196,N_28660,N_29587);
nand U31197 (N_31197,N_28032,N_28648);
nor U31198 (N_31198,N_28276,N_29583);
nor U31199 (N_31199,N_28045,N_29007);
nand U31200 (N_31200,N_28199,N_29211);
nand U31201 (N_31201,N_29670,N_29177);
nand U31202 (N_31202,N_29407,N_28202);
nor U31203 (N_31203,N_28831,N_28759);
nor U31204 (N_31204,N_28770,N_29936);
nand U31205 (N_31205,N_28790,N_29251);
nand U31206 (N_31206,N_29766,N_28892);
and U31207 (N_31207,N_28825,N_28816);
or U31208 (N_31208,N_28279,N_29517);
and U31209 (N_31209,N_28942,N_29135);
and U31210 (N_31210,N_29388,N_28138);
nor U31211 (N_31211,N_28948,N_28331);
or U31212 (N_31212,N_29550,N_28412);
and U31213 (N_31213,N_29757,N_29619);
or U31214 (N_31214,N_29484,N_28079);
or U31215 (N_31215,N_28359,N_29125);
nand U31216 (N_31216,N_28039,N_29234);
nand U31217 (N_31217,N_28475,N_28925);
and U31218 (N_31218,N_29321,N_29198);
xor U31219 (N_31219,N_29010,N_28806);
nand U31220 (N_31220,N_28314,N_28342);
nand U31221 (N_31221,N_29748,N_28839);
nand U31222 (N_31222,N_29342,N_28217);
and U31223 (N_31223,N_28463,N_29430);
nor U31224 (N_31224,N_28889,N_29490);
nand U31225 (N_31225,N_29163,N_28673);
and U31226 (N_31226,N_29037,N_29544);
nor U31227 (N_31227,N_29188,N_29574);
nand U31228 (N_31228,N_28023,N_29219);
and U31229 (N_31229,N_29646,N_29526);
nor U31230 (N_31230,N_28408,N_28426);
nand U31231 (N_31231,N_29052,N_28107);
or U31232 (N_31232,N_29916,N_29441);
nand U31233 (N_31233,N_29416,N_29009);
nand U31234 (N_31234,N_28341,N_28706);
nand U31235 (N_31235,N_29512,N_29028);
xnor U31236 (N_31236,N_28276,N_28983);
and U31237 (N_31237,N_29051,N_28617);
nor U31238 (N_31238,N_28722,N_29432);
or U31239 (N_31239,N_28465,N_29095);
nand U31240 (N_31240,N_28429,N_28394);
nor U31241 (N_31241,N_29960,N_28310);
or U31242 (N_31242,N_29703,N_28331);
nand U31243 (N_31243,N_28073,N_29543);
nand U31244 (N_31244,N_28258,N_28892);
or U31245 (N_31245,N_28823,N_28069);
or U31246 (N_31246,N_28964,N_29510);
nor U31247 (N_31247,N_28699,N_29076);
and U31248 (N_31248,N_29357,N_29151);
or U31249 (N_31249,N_28510,N_28749);
nor U31250 (N_31250,N_29065,N_28031);
nand U31251 (N_31251,N_28633,N_29279);
nor U31252 (N_31252,N_29671,N_29206);
and U31253 (N_31253,N_29873,N_29854);
nand U31254 (N_31254,N_29910,N_29911);
and U31255 (N_31255,N_28091,N_29841);
and U31256 (N_31256,N_28383,N_29802);
nand U31257 (N_31257,N_29053,N_28406);
or U31258 (N_31258,N_28416,N_29849);
and U31259 (N_31259,N_29016,N_29497);
and U31260 (N_31260,N_29325,N_28922);
nor U31261 (N_31261,N_28803,N_29432);
nor U31262 (N_31262,N_28860,N_29307);
and U31263 (N_31263,N_29872,N_28768);
and U31264 (N_31264,N_29639,N_28080);
or U31265 (N_31265,N_28416,N_29371);
nor U31266 (N_31266,N_29051,N_29820);
or U31267 (N_31267,N_29790,N_28612);
or U31268 (N_31268,N_28728,N_28500);
and U31269 (N_31269,N_29740,N_29919);
and U31270 (N_31270,N_29013,N_28590);
and U31271 (N_31271,N_28903,N_28177);
nand U31272 (N_31272,N_29865,N_28273);
nor U31273 (N_31273,N_28013,N_28537);
and U31274 (N_31274,N_28616,N_28984);
nand U31275 (N_31275,N_29936,N_28785);
nor U31276 (N_31276,N_28613,N_28463);
nor U31277 (N_31277,N_29766,N_28675);
nor U31278 (N_31278,N_29808,N_29408);
nor U31279 (N_31279,N_29646,N_28600);
nor U31280 (N_31280,N_29782,N_28834);
nor U31281 (N_31281,N_29954,N_29916);
or U31282 (N_31282,N_28040,N_28491);
nor U31283 (N_31283,N_28793,N_29287);
nor U31284 (N_31284,N_28050,N_29719);
nand U31285 (N_31285,N_29664,N_29292);
nor U31286 (N_31286,N_29165,N_28937);
and U31287 (N_31287,N_28887,N_29188);
nand U31288 (N_31288,N_28774,N_29515);
or U31289 (N_31289,N_29444,N_29633);
nand U31290 (N_31290,N_29745,N_28240);
and U31291 (N_31291,N_28297,N_28289);
nor U31292 (N_31292,N_29110,N_28632);
and U31293 (N_31293,N_29479,N_29760);
nand U31294 (N_31294,N_29748,N_28764);
nand U31295 (N_31295,N_28898,N_29005);
and U31296 (N_31296,N_28024,N_29694);
and U31297 (N_31297,N_28194,N_28316);
or U31298 (N_31298,N_29022,N_28788);
nor U31299 (N_31299,N_29651,N_29327);
and U31300 (N_31300,N_28921,N_29440);
or U31301 (N_31301,N_28299,N_28491);
or U31302 (N_31302,N_29073,N_28942);
and U31303 (N_31303,N_29781,N_29550);
nor U31304 (N_31304,N_29915,N_29976);
or U31305 (N_31305,N_29861,N_29625);
and U31306 (N_31306,N_29637,N_28064);
nand U31307 (N_31307,N_29650,N_29137);
or U31308 (N_31308,N_29291,N_29265);
nand U31309 (N_31309,N_28139,N_29419);
xnor U31310 (N_31310,N_28678,N_28482);
and U31311 (N_31311,N_28269,N_29794);
or U31312 (N_31312,N_28916,N_28113);
and U31313 (N_31313,N_28676,N_28754);
nand U31314 (N_31314,N_29941,N_29426);
or U31315 (N_31315,N_28011,N_29370);
and U31316 (N_31316,N_28244,N_29733);
and U31317 (N_31317,N_29739,N_29090);
nand U31318 (N_31318,N_28136,N_28869);
or U31319 (N_31319,N_28089,N_28043);
nand U31320 (N_31320,N_28636,N_29070);
or U31321 (N_31321,N_29033,N_29063);
nand U31322 (N_31322,N_29280,N_29178);
and U31323 (N_31323,N_29326,N_28519);
or U31324 (N_31324,N_28768,N_28262);
or U31325 (N_31325,N_28980,N_28473);
or U31326 (N_31326,N_29147,N_29484);
nand U31327 (N_31327,N_28938,N_29324);
nand U31328 (N_31328,N_28178,N_28889);
nand U31329 (N_31329,N_28002,N_28225);
or U31330 (N_31330,N_29448,N_28170);
or U31331 (N_31331,N_28661,N_28387);
nand U31332 (N_31332,N_28042,N_28905);
nand U31333 (N_31333,N_28901,N_29640);
nand U31334 (N_31334,N_29775,N_28168);
nand U31335 (N_31335,N_28935,N_29803);
or U31336 (N_31336,N_29693,N_29859);
and U31337 (N_31337,N_29983,N_28599);
nor U31338 (N_31338,N_29792,N_28973);
and U31339 (N_31339,N_28112,N_28377);
nor U31340 (N_31340,N_28542,N_28216);
xor U31341 (N_31341,N_29368,N_29087);
nor U31342 (N_31342,N_29455,N_29677);
nand U31343 (N_31343,N_28040,N_28825);
or U31344 (N_31344,N_29379,N_28805);
nor U31345 (N_31345,N_29329,N_29655);
and U31346 (N_31346,N_28647,N_29763);
and U31347 (N_31347,N_29745,N_28722);
or U31348 (N_31348,N_29096,N_28675);
nand U31349 (N_31349,N_28185,N_29539);
nand U31350 (N_31350,N_28586,N_29889);
and U31351 (N_31351,N_28077,N_29812);
or U31352 (N_31352,N_29068,N_28854);
and U31353 (N_31353,N_29999,N_28054);
nor U31354 (N_31354,N_28174,N_29974);
nor U31355 (N_31355,N_29659,N_29745);
nor U31356 (N_31356,N_28885,N_29960);
or U31357 (N_31357,N_29912,N_29309);
and U31358 (N_31358,N_29572,N_28205);
nor U31359 (N_31359,N_28216,N_29323);
and U31360 (N_31360,N_28230,N_28062);
or U31361 (N_31361,N_29405,N_28712);
or U31362 (N_31362,N_28364,N_28542);
nand U31363 (N_31363,N_29390,N_29743);
nand U31364 (N_31364,N_28728,N_29987);
nor U31365 (N_31365,N_29449,N_28209);
nor U31366 (N_31366,N_29993,N_28260);
and U31367 (N_31367,N_28189,N_29365);
and U31368 (N_31368,N_29563,N_29262);
and U31369 (N_31369,N_29231,N_29764);
and U31370 (N_31370,N_29013,N_29786);
nand U31371 (N_31371,N_29543,N_29556);
nor U31372 (N_31372,N_28919,N_28212);
nor U31373 (N_31373,N_28017,N_28846);
nand U31374 (N_31374,N_28158,N_28882);
and U31375 (N_31375,N_29414,N_28284);
and U31376 (N_31376,N_29079,N_29495);
and U31377 (N_31377,N_29945,N_28645);
nor U31378 (N_31378,N_29176,N_29930);
or U31379 (N_31379,N_28372,N_29011);
or U31380 (N_31380,N_29392,N_29653);
and U31381 (N_31381,N_28929,N_28274);
and U31382 (N_31382,N_28697,N_28242);
and U31383 (N_31383,N_29726,N_28791);
nand U31384 (N_31384,N_29914,N_29309);
nor U31385 (N_31385,N_29383,N_29462);
nor U31386 (N_31386,N_28687,N_29153);
and U31387 (N_31387,N_28569,N_28686);
and U31388 (N_31388,N_29379,N_28619);
or U31389 (N_31389,N_29156,N_29841);
nand U31390 (N_31390,N_29779,N_29105);
or U31391 (N_31391,N_29341,N_29101);
nor U31392 (N_31392,N_29535,N_28364);
and U31393 (N_31393,N_29627,N_28146);
or U31394 (N_31394,N_28398,N_28035);
nor U31395 (N_31395,N_29565,N_28500);
and U31396 (N_31396,N_28930,N_29857);
nor U31397 (N_31397,N_29859,N_29132);
nand U31398 (N_31398,N_29806,N_28495);
and U31399 (N_31399,N_29863,N_29795);
nor U31400 (N_31400,N_28712,N_29098);
and U31401 (N_31401,N_28872,N_28165);
or U31402 (N_31402,N_28397,N_28471);
nand U31403 (N_31403,N_28594,N_28462);
and U31404 (N_31404,N_28735,N_28452);
or U31405 (N_31405,N_28956,N_28065);
and U31406 (N_31406,N_29969,N_28684);
nand U31407 (N_31407,N_29981,N_28738);
and U31408 (N_31408,N_29518,N_29834);
or U31409 (N_31409,N_28181,N_28747);
xor U31410 (N_31410,N_28067,N_29870);
nor U31411 (N_31411,N_28839,N_29718);
nor U31412 (N_31412,N_29804,N_29503);
nor U31413 (N_31413,N_28569,N_28530);
and U31414 (N_31414,N_28179,N_29490);
or U31415 (N_31415,N_29837,N_29772);
nand U31416 (N_31416,N_28893,N_29623);
nor U31417 (N_31417,N_29081,N_29571);
or U31418 (N_31418,N_28542,N_28888);
or U31419 (N_31419,N_28796,N_28110);
nor U31420 (N_31420,N_29885,N_28470);
nor U31421 (N_31421,N_29858,N_29200);
or U31422 (N_31422,N_29450,N_29875);
nand U31423 (N_31423,N_29123,N_29942);
or U31424 (N_31424,N_28327,N_29230);
or U31425 (N_31425,N_29773,N_29051);
xor U31426 (N_31426,N_29108,N_28199);
nand U31427 (N_31427,N_28920,N_28475);
nor U31428 (N_31428,N_28289,N_29557);
xor U31429 (N_31429,N_28311,N_29380);
nand U31430 (N_31430,N_29665,N_29643);
nor U31431 (N_31431,N_28667,N_28941);
and U31432 (N_31432,N_29058,N_28602);
or U31433 (N_31433,N_28762,N_28425);
nand U31434 (N_31434,N_29647,N_29862);
nor U31435 (N_31435,N_28556,N_29097);
or U31436 (N_31436,N_29223,N_28768);
xor U31437 (N_31437,N_28644,N_28939);
and U31438 (N_31438,N_29941,N_29896);
nor U31439 (N_31439,N_28201,N_29639);
nand U31440 (N_31440,N_29623,N_29400);
and U31441 (N_31441,N_28038,N_28542);
nand U31442 (N_31442,N_28813,N_29226);
and U31443 (N_31443,N_28895,N_29115);
or U31444 (N_31444,N_28007,N_28845);
nand U31445 (N_31445,N_28818,N_28262);
and U31446 (N_31446,N_29350,N_28651);
nand U31447 (N_31447,N_29941,N_29909);
nor U31448 (N_31448,N_28744,N_29374);
nor U31449 (N_31449,N_28366,N_28828);
nand U31450 (N_31450,N_29179,N_28023);
and U31451 (N_31451,N_28326,N_28786);
and U31452 (N_31452,N_28785,N_28333);
nand U31453 (N_31453,N_28322,N_28849);
or U31454 (N_31454,N_28685,N_29813);
nor U31455 (N_31455,N_29716,N_28638);
and U31456 (N_31456,N_28481,N_29494);
and U31457 (N_31457,N_28490,N_28757);
nand U31458 (N_31458,N_28080,N_28461);
nor U31459 (N_31459,N_29061,N_28892);
nand U31460 (N_31460,N_28540,N_29430);
and U31461 (N_31461,N_28758,N_28040);
and U31462 (N_31462,N_28490,N_28245);
and U31463 (N_31463,N_29845,N_29126);
and U31464 (N_31464,N_28806,N_29695);
or U31465 (N_31465,N_28128,N_28766);
nor U31466 (N_31466,N_28369,N_29436);
nand U31467 (N_31467,N_28824,N_29495);
and U31468 (N_31468,N_28658,N_29681);
nor U31469 (N_31469,N_28843,N_28440);
nand U31470 (N_31470,N_28066,N_29053);
xor U31471 (N_31471,N_28947,N_28938);
or U31472 (N_31472,N_29969,N_28560);
and U31473 (N_31473,N_28109,N_28484);
nor U31474 (N_31474,N_29440,N_28626);
xor U31475 (N_31475,N_28377,N_28394);
and U31476 (N_31476,N_29009,N_29390);
or U31477 (N_31477,N_29553,N_29943);
nand U31478 (N_31478,N_29837,N_28291);
or U31479 (N_31479,N_28991,N_29260);
or U31480 (N_31480,N_29874,N_29259);
xnor U31481 (N_31481,N_28709,N_28943);
or U31482 (N_31482,N_29992,N_28302);
and U31483 (N_31483,N_28929,N_29669);
and U31484 (N_31484,N_29385,N_29303);
and U31485 (N_31485,N_28202,N_28219);
or U31486 (N_31486,N_28343,N_29796);
and U31487 (N_31487,N_29531,N_29273);
nor U31488 (N_31488,N_28349,N_29887);
nor U31489 (N_31489,N_29126,N_29138);
and U31490 (N_31490,N_28248,N_29475);
and U31491 (N_31491,N_28218,N_28346);
nand U31492 (N_31492,N_29650,N_29571);
or U31493 (N_31493,N_28877,N_29777);
nor U31494 (N_31494,N_28036,N_28583);
nand U31495 (N_31495,N_29498,N_29631);
nand U31496 (N_31496,N_29671,N_29151);
nor U31497 (N_31497,N_28306,N_29469);
nor U31498 (N_31498,N_29087,N_29107);
nor U31499 (N_31499,N_29346,N_29749);
nor U31500 (N_31500,N_29249,N_28257);
and U31501 (N_31501,N_29332,N_29488);
and U31502 (N_31502,N_28851,N_29068);
nand U31503 (N_31503,N_28331,N_29462);
nand U31504 (N_31504,N_29801,N_28923);
nor U31505 (N_31505,N_28913,N_29805);
and U31506 (N_31506,N_28620,N_28650);
nor U31507 (N_31507,N_29490,N_28298);
nand U31508 (N_31508,N_28368,N_29197);
nand U31509 (N_31509,N_29236,N_29951);
or U31510 (N_31510,N_28066,N_29100);
nor U31511 (N_31511,N_28498,N_28021);
nor U31512 (N_31512,N_28138,N_29899);
or U31513 (N_31513,N_28168,N_28367);
and U31514 (N_31514,N_28376,N_28051);
or U31515 (N_31515,N_29207,N_28379);
nor U31516 (N_31516,N_29373,N_29602);
nor U31517 (N_31517,N_28518,N_28013);
and U31518 (N_31518,N_28993,N_28068);
and U31519 (N_31519,N_29720,N_28576);
nand U31520 (N_31520,N_28271,N_28116);
or U31521 (N_31521,N_29182,N_28950);
or U31522 (N_31522,N_29992,N_28821);
and U31523 (N_31523,N_29812,N_29928);
nand U31524 (N_31524,N_28679,N_29737);
and U31525 (N_31525,N_29150,N_28798);
nor U31526 (N_31526,N_29492,N_29910);
nand U31527 (N_31527,N_29058,N_28042);
nor U31528 (N_31528,N_29781,N_28104);
or U31529 (N_31529,N_29301,N_29891);
nor U31530 (N_31530,N_28133,N_28848);
xnor U31531 (N_31531,N_29656,N_28322);
nand U31532 (N_31532,N_28336,N_29799);
or U31533 (N_31533,N_28496,N_28607);
nand U31534 (N_31534,N_29383,N_28854);
nand U31535 (N_31535,N_29531,N_28747);
nand U31536 (N_31536,N_28375,N_28354);
nor U31537 (N_31537,N_28494,N_28906);
xor U31538 (N_31538,N_29679,N_28520);
xor U31539 (N_31539,N_28761,N_29128);
or U31540 (N_31540,N_29767,N_28229);
nor U31541 (N_31541,N_28356,N_28197);
or U31542 (N_31542,N_29594,N_29741);
and U31543 (N_31543,N_29196,N_28530);
nor U31544 (N_31544,N_28812,N_28218);
xor U31545 (N_31545,N_29968,N_28030);
and U31546 (N_31546,N_28526,N_28856);
and U31547 (N_31547,N_28704,N_28650);
and U31548 (N_31548,N_28042,N_29484);
nor U31549 (N_31549,N_29089,N_29210);
and U31550 (N_31550,N_29223,N_29192);
and U31551 (N_31551,N_29126,N_29829);
nor U31552 (N_31552,N_28575,N_29187);
and U31553 (N_31553,N_28006,N_29369);
and U31554 (N_31554,N_28085,N_28478);
nor U31555 (N_31555,N_29981,N_29457);
or U31556 (N_31556,N_29965,N_28480);
nor U31557 (N_31557,N_29338,N_29438);
nor U31558 (N_31558,N_28133,N_28676);
nor U31559 (N_31559,N_28835,N_29639);
nor U31560 (N_31560,N_29970,N_29700);
and U31561 (N_31561,N_28412,N_28767);
nor U31562 (N_31562,N_28698,N_29225);
or U31563 (N_31563,N_29282,N_29790);
and U31564 (N_31564,N_29691,N_28135);
nor U31565 (N_31565,N_28799,N_28619);
or U31566 (N_31566,N_29582,N_29747);
or U31567 (N_31567,N_29332,N_29901);
nand U31568 (N_31568,N_29986,N_28339);
nand U31569 (N_31569,N_29877,N_29411);
nand U31570 (N_31570,N_29769,N_29860);
nand U31571 (N_31571,N_28792,N_28638);
or U31572 (N_31572,N_28535,N_29006);
or U31573 (N_31573,N_28217,N_28940);
and U31574 (N_31574,N_28751,N_28817);
or U31575 (N_31575,N_28594,N_29096);
nand U31576 (N_31576,N_28787,N_28653);
nor U31577 (N_31577,N_28161,N_29356);
nand U31578 (N_31578,N_29142,N_29228);
or U31579 (N_31579,N_29035,N_29283);
nor U31580 (N_31580,N_28232,N_28713);
nand U31581 (N_31581,N_28345,N_29879);
and U31582 (N_31582,N_28756,N_29322);
and U31583 (N_31583,N_29777,N_28302);
or U31584 (N_31584,N_29082,N_28993);
and U31585 (N_31585,N_29885,N_28960);
nor U31586 (N_31586,N_28601,N_29804);
nand U31587 (N_31587,N_29741,N_29492);
or U31588 (N_31588,N_28154,N_28019);
nor U31589 (N_31589,N_28484,N_28540);
nor U31590 (N_31590,N_28593,N_28630);
or U31591 (N_31591,N_29922,N_28225);
and U31592 (N_31592,N_29765,N_28162);
nor U31593 (N_31593,N_28353,N_29291);
nor U31594 (N_31594,N_29898,N_28092);
nor U31595 (N_31595,N_29109,N_29347);
nand U31596 (N_31596,N_28602,N_29094);
nand U31597 (N_31597,N_28894,N_29168);
nand U31598 (N_31598,N_29253,N_28112);
nor U31599 (N_31599,N_29308,N_29630);
and U31600 (N_31600,N_29271,N_29998);
nor U31601 (N_31601,N_28608,N_29272);
and U31602 (N_31602,N_29032,N_29780);
or U31603 (N_31603,N_29285,N_28195);
and U31604 (N_31604,N_28498,N_28383);
or U31605 (N_31605,N_29854,N_29130);
or U31606 (N_31606,N_29964,N_29204);
and U31607 (N_31607,N_28585,N_29031);
and U31608 (N_31608,N_29578,N_28265);
nor U31609 (N_31609,N_29787,N_29763);
nand U31610 (N_31610,N_29281,N_29669);
and U31611 (N_31611,N_28305,N_28673);
and U31612 (N_31612,N_29601,N_29819);
xnor U31613 (N_31613,N_28670,N_29836);
and U31614 (N_31614,N_29686,N_28812);
nor U31615 (N_31615,N_28570,N_28340);
or U31616 (N_31616,N_28397,N_29085);
and U31617 (N_31617,N_28358,N_28710);
or U31618 (N_31618,N_28934,N_29823);
nor U31619 (N_31619,N_28346,N_28943);
and U31620 (N_31620,N_28350,N_28463);
nor U31621 (N_31621,N_28840,N_29001);
or U31622 (N_31622,N_28244,N_29018);
or U31623 (N_31623,N_28357,N_28223);
and U31624 (N_31624,N_28693,N_28154);
and U31625 (N_31625,N_29640,N_29013);
nor U31626 (N_31626,N_29650,N_28592);
nor U31627 (N_31627,N_29809,N_28271);
nand U31628 (N_31628,N_28680,N_28536);
nand U31629 (N_31629,N_29443,N_28770);
nor U31630 (N_31630,N_28960,N_29476);
and U31631 (N_31631,N_28555,N_29960);
and U31632 (N_31632,N_29018,N_29833);
and U31633 (N_31633,N_28115,N_28727);
nand U31634 (N_31634,N_29634,N_29998);
and U31635 (N_31635,N_28966,N_28824);
or U31636 (N_31636,N_29458,N_29572);
nand U31637 (N_31637,N_29239,N_29920);
nor U31638 (N_31638,N_29735,N_29957);
nor U31639 (N_31639,N_28276,N_29980);
and U31640 (N_31640,N_29499,N_28857);
or U31641 (N_31641,N_28390,N_28934);
or U31642 (N_31642,N_29213,N_29171);
nand U31643 (N_31643,N_28833,N_28925);
nand U31644 (N_31644,N_29167,N_28601);
and U31645 (N_31645,N_29063,N_29344);
nor U31646 (N_31646,N_29598,N_29884);
or U31647 (N_31647,N_29680,N_29414);
nand U31648 (N_31648,N_29772,N_29908);
and U31649 (N_31649,N_29584,N_28777);
and U31650 (N_31650,N_29681,N_29379);
or U31651 (N_31651,N_29774,N_28458);
nand U31652 (N_31652,N_28148,N_29955);
nand U31653 (N_31653,N_29185,N_29922);
or U31654 (N_31654,N_28747,N_29465);
or U31655 (N_31655,N_28367,N_29687);
nor U31656 (N_31656,N_28789,N_29138);
nor U31657 (N_31657,N_28002,N_29614);
and U31658 (N_31658,N_29090,N_29421);
nand U31659 (N_31659,N_29674,N_29524);
or U31660 (N_31660,N_28115,N_28098);
nor U31661 (N_31661,N_28563,N_29984);
nor U31662 (N_31662,N_28364,N_29596);
and U31663 (N_31663,N_28911,N_29222);
or U31664 (N_31664,N_28207,N_29158);
and U31665 (N_31665,N_28352,N_29607);
nor U31666 (N_31666,N_29758,N_28567);
and U31667 (N_31667,N_29514,N_29562);
or U31668 (N_31668,N_29916,N_28243);
or U31669 (N_31669,N_29028,N_28932);
and U31670 (N_31670,N_28361,N_28098);
nor U31671 (N_31671,N_28615,N_28625);
or U31672 (N_31672,N_29942,N_28612);
nor U31673 (N_31673,N_29618,N_28587);
nor U31674 (N_31674,N_29291,N_29524);
and U31675 (N_31675,N_29141,N_28225);
or U31676 (N_31676,N_29555,N_28426);
and U31677 (N_31677,N_29737,N_28881);
nor U31678 (N_31678,N_28438,N_29912);
nand U31679 (N_31679,N_29356,N_28827);
or U31680 (N_31680,N_28073,N_28081);
xnor U31681 (N_31681,N_29215,N_29820);
and U31682 (N_31682,N_29386,N_28162);
and U31683 (N_31683,N_28990,N_28487);
and U31684 (N_31684,N_29243,N_28724);
nor U31685 (N_31685,N_28145,N_28097);
nand U31686 (N_31686,N_29143,N_28586);
nor U31687 (N_31687,N_29305,N_29407);
nand U31688 (N_31688,N_28500,N_28165);
nand U31689 (N_31689,N_29418,N_29498);
nor U31690 (N_31690,N_28726,N_29368);
xor U31691 (N_31691,N_28931,N_29489);
or U31692 (N_31692,N_29115,N_29631);
nand U31693 (N_31693,N_29263,N_29900);
or U31694 (N_31694,N_28850,N_28273);
or U31695 (N_31695,N_29373,N_28490);
or U31696 (N_31696,N_28204,N_29715);
nor U31697 (N_31697,N_29458,N_29704);
and U31698 (N_31698,N_28584,N_29426);
nor U31699 (N_31699,N_28375,N_29089);
or U31700 (N_31700,N_29108,N_28532);
or U31701 (N_31701,N_29702,N_29824);
nor U31702 (N_31702,N_29401,N_29205);
nand U31703 (N_31703,N_29544,N_28968);
and U31704 (N_31704,N_29159,N_29538);
nor U31705 (N_31705,N_29188,N_28052);
nor U31706 (N_31706,N_29319,N_28609);
nor U31707 (N_31707,N_29502,N_28284);
nor U31708 (N_31708,N_28354,N_28609);
or U31709 (N_31709,N_28041,N_29587);
xnor U31710 (N_31710,N_28096,N_28541);
nor U31711 (N_31711,N_28703,N_28053);
nand U31712 (N_31712,N_28707,N_29575);
xnor U31713 (N_31713,N_28739,N_29026);
nand U31714 (N_31714,N_29034,N_28769);
nand U31715 (N_31715,N_28299,N_28559);
or U31716 (N_31716,N_28537,N_28808);
nand U31717 (N_31717,N_29786,N_29417);
nand U31718 (N_31718,N_29256,N_28553);
or U31719 (N_31719,N_28269,N_28755);
nand U31720 (N_31720,N_29071,N_28862);
nand U31721 (N_31721,N_28105,N_28696);
nand U31722 (N_31722,N_29516,N_28516);
nor U31723 (N_31723,N_29905,N_29687);
or U31724 (N_31724,N_29874,N_28191);
or U31725 (N_31725,N_28310,N_28340);
nand U31726 (N_31726,N_28426,N_29372);
xor U31727 (N_31727,N_29083,N_28171);
nand U31728 (N_31728,N_29344,N_29026);
or U31729 (N_31729,N_29813,N_28189);
or U31730 (N_31730,N_28692,N_29692);
or U31731 (N_31731,N_28580,N_28174);
nand U31732 (N_31732,N_29932,N_29512);
or U31733 (N_31733,N_29010,N_28636);
nand U31734 (N_31734,N_29107,N_29117);
nor U31735 (N_31735,N_28429,N_28183);
or U31736 (N_31736,N_29067,N_28483);
or U31737 (N_31737,N_29266,N_28707);
and U31738 (N_31738,N_28430,N_29185);
nor U31739 (N_31739,N_28284,N_28890);
xor U31740 (N_31740,N_28932,N_29569);
nor U31741 (N_31741,N_28339,N_29567);
xor U31742 (N_31742,N_29522,N_29670);
nand U31743 (N_31743,N_28427,N_29843);
nand U31744 (N_31744,N_28299,N_29261);
nand U31745 (N_31745,N_28156,N_29768);
or U31746 (N_31746,N_29943,N_29503);
nor U31747 (N_31747,N_28712,N_28180);
nand U31748 (N_31748,N_29460,N_28143);
xnor U31749 (N_31749,N_28132,N_28964);
or U31750 (N_31750,N_29818,N_29111);
nor U31751 (N_31751,N_28627,N_28952);
or U31752 (N_31752,N_28520,N_29735);
nand U31753 (N_31753,N_29133,N_29635);
or U31754 (N_31754,N_28161,N_29552);
nor U31755 (N_31755,N_29300,N_29655);
and U31756 (N_31756,N_29199,N_29250);
nor U31757 (N_31757,N_29072,N_29779);
or U31758 (N_31758,N_28303,N_29230);
or U31759 (N_31759,N_28739,N_29549);
and U31760 (N_31760,N_29981,N_28588);
nor U31761 (N_31761,N_28490,N_29663);
or U31762 (N_31762,N_28209,N_28287);
nand U31763 (N_31763,N_28268,N_29635);
nor U31764 (N_31764,N_29896,N_28889);
nand U31765 (N_31765,N_29655,N_29180);
nor U31766 (N_31766,N_28163,N_29263);
nand U31767 (N_31767,N_29163,N_29897);
nand U31768 (N_31768,N_29128,N_28866);
nand U31769 (N_31769,N_28267,N_28143);
and U31770 (N_31770,N_29812,N_28227);
or U31771 (N_31771,N_29773,N_29904);
and U31772 (N_31772,N_28453,N_28714);
nand U31773 (N_31773,N_28190,N_29147);
nand U31774 (N_31774,N_29206,N_29185);
nand U31775 (N_31775,N_28551,N_28393);
nor U31776 (N_31776,N_28821,N_28435);
xor U31777 (N_31777,N_28894,N_29789);
nor U31778 (N_31778,N_28482,N_28443);
or U31779 (N_31779,N_29525,N_29196);
xor U31780 (N_31780,N_29072,N_29173);
or U31781 (N_31781,N_29679,N_28236);
nand U31782 (N_31782,N_28318,N_29012);
and U31783 (N_31783,N_29691,N_28181);
or U31784 (N_31784,N_28806,N_29831);
nand U31785 (N_31785,N_28001,N_28366);
nand U31786 (N_31786,N_29963,N_28245);
or U31787 (N_31787,N_29732,N_28739);
xor U31788 (N_31788,N_28984,N_28116);
or U31789 (N_31789,N_28443,N_28515);
nor U31790 (N_31790,N_29021,N_29397);
nand U31791 (N_31791,N_29719,N_29449);
and U31792 (N_31792,N_28856,N_29453);
and U31793 (N_31793,N_29460,N_28673);
nor U31794 (N_31794,N_28383,N_29534);
or U31795 (N_31795,N_29883,N_28588);
and U31796 (N_31796,N_28779,N_28469);
and U31797 (N_31797,N_28347,N_28817);
or U31798 (N_31798,N_29260,N_29634);
or U31799 (N_31799,N_29069,N_29414);
nand U31800 (N_31800,N_29432,N_28513);
and U31801 (N_31801,N_29566,N_29841);
nand U31802 (N_31802,N_29706,N_29020);
nand U31803 (N_31803,N_29813,N_29522);
and U31804 (N_31804,N_28943,N_28796);
or U31805 (N_31805,N_28130,N_28750);
nor U31806 (N_31806,N_28042,N_28015);
nand U31807 (N_31807,N_28875,N_29040);
nor U31808 (N_31808,N_29608,N_29157);
nor U31809 (N_31809,N_29009,N_28340);
or U31810 (N_31810,N_28919,N_29894);
nor U31811 (N_31811,N_28821,N_28560);
and U31812 (N_31812,N_29446,N_29590);
and U31813 (N_31813,N_29227,N_29789);
and U31814 (N_31814,N_28538,N_29392);
or U31815 (N_31815,N_28370,N_29820);
and U31816 (N_31816,N_29895,N_28721);
nand U31817 (N_31817,N_29030,N_28892);
nor U31818 (N_31818,N_29663,N_29078);
or U31819 (N_31819,N_28415,N_28625);
and U31820 (N_31820,N_28457,N_28618);
or U31821 (N_31821,N_28666,N_28534);
or U31822 (N_31822,N_28141,N_28919);
or U31823 (N_31823,N_29491,N_29942);
and U31824 (N_31824,N_28910,N_28604);
and U31825 (N_31825,N_28125,N_28703);
nand U31826 (N_31826,N_28652,N_28176);
and U31827 (N_31827,N_28456,N_29493);
and U31828 (N_31828,N_28322,N_28495);
and U31829 (N_31829,N_28439,N_29531);
or U31830 (N_31830,N_28217,N_29642);
nand U31831 (N_31831,N_29768,N_28753);
nand U31832 (N_31832,N_28904,N_29199);
nand U31833 (N_31833,N_29193,N_29717);
nor U31834 (N_31834,N_29011,N_29811);
and U31835 (N_31835,N_28326,N_28854);
or U31836 (N_31836,N_29186,N_28912);
or U31837 (N_31837,N_28171,N_29501);
nand U31838 (N_31838,N_29225,N_29228);
or U31839 (N_31839,N_28541,N_28886);
or U31840 (N_31840,N_28052,N_29161);
and U31841 (N_31841,N_28792,N_28535);
nor U31842 (N_31842,N_28131,N_28073);
or U31843 (N_31843,N_29990,N_28193);
and U31844 (N_31844,N_28725,N_28357);
and U31845 (N_31845,N_29315,N_28566);
and U31846 (N_31846,N_28008,N_29235);
nand U31847 (N_31847,N_28428,N_29817);
and U31848 (N_31848,N_28117,N_29477);
nand U31849 (N_31849,N_29504,N_28878);
nand U31850 (N_31850,N_29853,N_28723);
or U31851 (N_31851,N_28242,N_28963);
nand U31852 (N_31852,N_29986,N_29983);
nor U31853 (N_31853,N_29480,N_29919);
nor U31854 (N_31854,N_29039,N_29180);
and U31855 (N_31855,N_28952,N_28778);
and U31856 (N_31856,N_29911,N_29886);
and U31857 (N_31857,N_28038,N_28388);
and U31858 (N_31858,N_29014,N_29539);
nand U31859 (N_31859,N_28142,N_28735);
nand U31860 (N_31860,N_29837,N_28461);
and U31861 (N_31861,N_29764,N_28616);
and U31862 (N_31862,N_28616,N_29727);
or U31863 (N_31863,N_28805,N_28915);
nand U31864 (N_31864,N_28465,N_28412);
and U31865 (N_31865,N_29973,N_28299);
and U31866 (N_31866,N_29216,N_28899);
or U31867 (N_31867,N_28351,N_29886);
nand U31868 (N_31868,N_28771,N_28871);
nand U31869 (N_31869,N_29355,N_29453);
xor U31870 (N_31870,N_28080,N_29484);
or U31871 (N_31871,N_28382,N_29469);
nor U31872 (N_31872,N_28591,N_29439);
or U31873 (N_31873,N_28838,N_29468);
nand U31874 (N_31874,N_28056,N_29831);
nor U31875 (N_31875,N_29781,N_28731);
nand U31876 (N_31876,N_29543,N_29819);
nand U31877 (N_31877,N_28635,N_28069);
and U31878 (N_31878,N_29811,N_29591);
xnor U31879 (N_31879,N_28914,N_29162);
and U31880 (N_31880,N_28121,N_28469);
or U31881 (N_31881,N_29667,N_29202);
nand U31882 (N_31882,N_28148,N_28789);
or U31883 (N_31883,N_28495,N_29544);
or U31884 (N_31884,N_29097,N_29272);
and U31885 (N_31885,N_29001,N_29527);
nor U31886 (N_31886,N_29401,N_29892);
nor U31887 (N_31887,N_29129,N_29065);
or U31888 (N_31888,N_28828,N_28918);
nor U31889 (N_31889,N_28642,N_29107);
nand U31890 (N_31890,N_29812,N_29021);
or U31891 (N_31891,N_29553,N_28601);
nand U31892 (N_31892,N_29770,N_28076);
nor U31893 (N_31893,N_28545,N_29674);
or U31894 (N_31894,N_28503,N_29137);
or U31895 (N_31895,N_29924,N_29931);
nor U31896 (N_31896,N_28111,N_29484);
nand U31897 (N_31897,N_28204,N_28862);
nand U31898 (N_31898,N_28154,N_29442);
or U31899 (N_31899,N_29056,N_28603);
nor U31900 (N_31900,N_29980,N_28842);
and U31901 (N_31901,N_28782,N_29614);
or U31902 (N_31902,N_29004,N_29814);
or U31903 (N_31903,N_28150,N_28789);
nand U31904 (N_31904,N_28334,N_28583);
or U31905 (N_31905,N_29235,N_29614);
nor U31906 (N_31906,N_28003,N_28913);
and U31907 (N_31907,N_28278,N_28340);
nor U31908 (N_31908,N_28890,N_28776);
nand U31909 (N_31909,N_28957,N_29013);
nand U31910 (N_31910,N_28176,N_29142);
and U31911 (N_31911,N_29484,N_28593);
nand U31912 (N_31912,N_29888,N_28036);
nand U31913 (N_31913,N_28317,N_28003);
nor U31914 (N_31914,N_29374,N_29668);
and U31915 (N_31915,N_29042,N_29087);
nand U31916 (N_31916,N_29320,N_28632);
nand U31917 (N_31917,N_28631,N_28910);
nand U31918 (N_31918,N_28848,N_28249);
and U31919 (N_31919,N_28234,N_28771);
nor U31920 (N_31920,N_28024,N_28891);
nor U31921 (N_31921,N_29990,N_29638);
or U31922 (N_31922,N_28064,N_29818);
and U31923 (N_31923,N_29337,N_29447);
and U31924 (N_31924,N_29897,N_29258);
and U31925 (N_31925,N_29755,N_28468);
nand U31926 (N_31926,N_28697,N_28768);
xnor U31927 (N_31927,N_29234,N_28600);
and U31928 (N_31928,N_29084,N_29775);
and U31929 (N_31929,N_28520,N_29389);
or U31930 (N_31930,N_29156,N_28928);
nor U31931 (N_31931,N_28489,N_28947);
nor U31932 (N_31932,N_28495,N_29593);
nor U31933 (N_31933,N_28110,N_29762);
nand U31934 (N_31934,N_28077,N_29339);
and U31935 (N_31935,N_28259,N_28461);
nand U31936 (N_31936,N_29514,N_28356);
nand U31937 (N_31937,N_29152,N_29563);
or U31938 (N_31938,N_28874,N_29004);
and U31939 (N_31939,N_29546,N_28604);
or U31940 (N_31940,N_29091,N_29710);
and U31941 (N_31941,N_28611,N_28961);
nor U31942 (N_31942,N_29913,N_29055);
nor U31943 (N_31943,N_28210,N_28397);
xnor U31944 (N_31944,N_28496,N_28011);
and U31945 (N_31945,N_29074,N_28553);
nand U31946 (N_31946,N_29364,N_28901);
and U31947 (N_31947,N_28498,N_28533);
nor U31948 (N_31948,N_28214,N_29813);
or U31949 (N_31949,N_29260,N_28095);
and U31950 (N_31950,N_28155,N_29401);
nor U31951 (N_31951,N_29549,N_29596);
or U31952 (N_31952,N_28867,N_29974);
nor U31953 (N_31953,N_29755,N_28842);
or U31954 (N_31954,N_29958,N_29629);
or U31955 (N_31955,N_29400,N_29480);
nand U31956 (N_31956,N_28409,N_29630);
or U31957 (N_31957,N_28776,N_29556);
and U31958 (N_31958,N_28555,N_28589);
and U31959 (N_31959,N_28866,N_29554);
or U31960 (N_31960,N_28901,N_28379);
and U31961 (N_31961,N_28631,N_29245);
or U31962 (N_31962,N_28705,N_29389);
nand U31963 (N_31963,N_28367,N_29638);
and U31964 (N_31964,N_29509,N_28473);
nor U31965 (N_31965,N_29804,N_28653);
or U31966 (N_31966,N_29940,N_28999);
nor U31967 (N_31967,N_28580,N_29609);
or U31968 (N_31968,N_28313,N_29902);
and U31969 (N_31969,N_28746,N_28262);
and U31970 (N_31970,N_29123,N_29752);
or U31971 (N_31971,N_29629,N_28542);
nor U31972 (N_31972,N_28266,N_28312);
nor U31973 (N_31973,N_29728,N_29167);
and U31974 (N_31974,N_29439,N_28960);
or U31975 (N_31975,N_28135,N_29886);
or U31976 (N_31976,N_29701,N_28750);
or U31977 (N_31977,N_28423,N_28549);
nor U31978 (N_31978,N_28954,N_29803);
nand U31979 (N_31979,N_29360,N_28838);
and U31980 (N_31980,N_28574,N_28979);
or U31981 (N_31981,N_28581,N_28829);
and U31982 (N_31982,N_28156,N_28760);
nand U31983 (N_31983,N_28294,N_29833);
nor U31984 (N_31984,N_29452,N_29931);
nand U31985 (N_31985,N_29508,N_29983);
nor U31986 (N_31986,N_29266,N_29361);
or U31987 (N_31987,N_29035,N_29267);
nor U31988 (N_31988,N_28532,N_28437);
nor U31989 (N_31989,N_28748,N_29298);
or U31990 (N_31990,N_28826,N_29238);
and U31991 (N_31991,N_28384,N_28999);
and U31992 (N_31992,N_29390,N_28394);
nand U31993 (N_31993,N_28262,N_29864);
and U31994 (N_31994,N_28678,N_29336);
or U31995 (N_31995,N_28141,N_29609);
nand U31996 (N_31996,N_29671,N_29664);
nor U31997 (N_31997,N_28051,N_28625);
and U31998 (N_31998,N_28470,N_29243);
nor U31999 (N_31999,N_28415,N_29754);
nand U32000 (N_32000,N_30661,N_30895);
or U32001 (N_32001,N_31210,N_30864);
and U32002 (N_32002,N_30990,N_30507);
or U32003 (N_32003,N_31494,N_31350);
and U32004 (N_32004,N_31364,N_30922);
or U32005 (N_32005,N_31644,N_30050);
xnor U32006 (N_32006,N_30450,N_30649);
nand U32007 (N_32007,N_30935,N_31400);
or U32008 (N_32008,N_30036,N_31702);
and U32009 (N_32009,N_31427,N_31159);
nor U32010 (N_32010,N_30166,N_31587);
nor U32011 (N_32011,N_31826,N_30349);
nor U32012 (N_32012,N_30213,N_31188);
nand U32013 (N_32013,N_30887,N_31712);
nand U32014 (N_32014,N_30640,N_30360);
and U32015 (N_32015,N_31288,N_31680);
or U32016 (N_32016,N_31733,N_31178);
or U32017 (N_32017,N_30763,N_31757);
or U32018 (N_32018,N_31889,N_30820);
nor U32019 (N_32019,N_30859,N_31546);
or U32020 (N_32020,N_31166,N_30222);
or U32021 (N_32021,N_31609,N_31742);
or U32022 (N_32022,N_31286,N_30765);
or U32023 (N_32023,N_31642,N_31457);
and U32024 (N_32024,N_31984,N_31924);
and U32025 (N_32025,N_31022,N_31670);
nor U32026 (N_32026,N_31219,N_31374);
nand U32027 (N_32027,N_31256,N_31901);
nor U32028 (N_32028,N_31087,N_30303);
or U32029 (N_32029,N_31861,N_31312);
nand U32030 (N_32030,N_31187,N_30719);
nand U32031 (N_32031,N_30483,N_31274);
and U32032 (N_32032,N_31989,N_31968);
and U32033 (N_32033,N_30839,N_31169);
or U32034 (N_32034,N_31255,N_30064);
and U32035 (N_32035,N_31492,N_31948);
nand U32036 (N_32036,N_30834,N_30361);
nor U32037 (N_32037,N_30356,N_30988);
nand U32038 (N_32038,N_30106,N_30494);
or U32039 (N_32039,N_31544,N_31459);
nand U32040 (N_32040,N_30810,N_30761);
nand U32041 (N_32041,N_31025,N_31433);
and U32042 (N_32042,N_30607,N_31152);
or U32043 (N_32043,N_31357,N_31414);
nand U32044 (N_32044,N_30266,N_30319);
nor U32045 (N_32045,N_31165,N_31519);
nor U32046 (N_32046,N_31719,N_30858);
or U32047 (N_32047,N_30353,N_30196);
nor U32048 (N_32048,N_31354,N_31077);
xor U32049 (N_32049,N_31144,N_30556);
nand U32050 (N_32050,N_30328,N_30265);
nand U32051 (N_32051,N_31882,N_31058);
or U32052 (N_32052,N_31634,N_31073);
nor U32053 (N_32053,N_30647,N_31990);
or U32054 (N_32054,N_31645,N_31020);
and U32055 (N_32055,N_31512,N_31460);
and U32056 (N_32056,N_30754,N_31932);
and U32057 (N_32057,N_31233,N_30125);
nor U32058 (N_32058,N_31123,N_30833);
nand U32059 (N_32059,N_30538,N_30415);
nor U32060 (N_32060,N_30431,N_30684);
nand U32061 (N_32061,N_31441,N_30366);
or U32062 (N_32062,N_31780,N_31366);
and U32063 (N_32063,N_30654,N_30174);
nand U32064 (N_32064,N_30562,N_30592);
and U32065 (N_32065,N_31262,N_30283);
nor U32066 (N_32066,N_31395,N_31816);
or U32067 (N_32067,N_31065,N_30263);
nor U32068 (N_32068,N_31061,N_30630);
nor U32069 (N_32069,N_30151,N_30380);
nand U32070 (N_32070,N_30465,N_30245);
nor U32071 (N_32071,N_31379,N_31865);
or U32072 (N_32072,N_31280,N_30101);
or U32073 (N_32073,N_30532,N_30944);
and U32074 (N_32074,N_31359,N_30149);
nand U32075 (N_32075,N_31054,N_30566);
nor U32076 (N_32076,N_31786,N_30629);
nor U32077 (N_32077,N_31408,N_31538);
nand U32078 (N_32078,N_30777,N_30667);
or U32079 (N_32079,N_31088,N_30132);
or U32080 (N_32080,N_31300,N_30796);
nand U32081 (N_32081,N_31755,N_31410);
and U32082 (N_32082,N_31174,N_31583);
or U32083 (N_32083,N_31714,N_31270);
and U32084 (N_32084,N_30376,N_31091);
or U32085 (N_32085,N_31389,N_30013);
nor U32086 (N_32086,N_31533,N_31662);
nand U32087 (N_32087,N_31119,N_31420);
nor U32088 (N_32088,N_30128,N_30209);
and U32089 (N_32089,N_31998,N_31904);
nor U32090 (N_32090,N_30452,N_31037);
and U32091 (N_32091,N_30750,N_30753);
nand U32092 (N_32092,N_31964,N_31192);
nor U32093 (N_32093,N_31935,N_31078);
or U32094 (N_32094,N_31729,N_31694);
or U32095 (N_32095,N_31050,N_31213);
nand U32096 (N_32096,N_31612,N_30786);
and U32097 (N_32097,N_31551,N_31785);
nor U32098 (N_32098,N_31329,N_30042);
nand U32099 (N_32099,N_30330,N_30012);
nand U32100 (N_32100,N_31317,N_31394);
nand U32101 (N_32101,N_31206,N_31774);
and U32102 (N_32102,N_31529,N_30814);
nand U32103 (N_32103,N_31301,N_30716);
nor U32104 (N_32104,N_30893,N_31950);
and U32105 (N_32105,N_31772,N_30425);
or U32106 (N_32106,N_30103,N_31239);
and U32107 (N_32107,N_31204,N_31847);
and U32108 (N_32108,N_30011,N_30454);
nor U32109 (N_32109,N_30412,N_30197);
nand U32110 (N_32110,N_30843,N_30428);
or U32111 (N_32111,N_31008,N_30482);
or U32112 (N_32112,N_30561,N_31074);
or U32113 (N_32113,N_31342,N_30981);
nor U32114 (N_32114,N_30123,N_31334);
nand U32115 (N_32115,N_30779,N_30589);
nor U32116 (N_32116,N_31944,N_30195);
nor U32117 (N_32117,N_31817,N_30108);
and U32118 (N_32118,N_30611,N_31727);
or U32119 (N_32119,N_31766,N_30416);
or U32120 (N_32120,N_30081,N_30698);
nor U32121 (N_32121,N_30652,N_31537);
nor U32122 (N_32122,N_30393,N_31124);
or U32123 (N_32123,N_31346,N_30216);
and U32124 (N_32124,N_31951,N_31142);
or U32125 (N_32125,N_30644,N_31599);
nor U32126 (N_32126,N_31436,N_30138);
nand U32127 (N_32127,N_30717,N_31155);
and U32128 (N_32128,N_31638,N_31507);
or U32129 (N_32129,N_30097,N_30269);
nor U32130 (N_32130,N_31763,N_30359);
nor U32131 (N_32131,N_30917,N_31046);
and U32132 (N_32132,N_31477,N_30329);
nand U32133 (N_32133,N_31722,N_30590);
or U32134 (N_32134,N_31767,N_30066);
and U32135 (N_32135,N_31205,N_31287);
and U32136 (N_32136,N_31409,N_30588);
or U32137 (N_32137,N_31641,N_30911);
nand U32138 (N_32138,N_31672,N_31230);
nor U32139 (N_32139,N_30941,N_30164);
and U32140 (N_32140,N_30254,N_31413);
and U32141 (N_32141,N_30604,N_31311);
nand U32142 (N_32142,N_30563,N_31391);
nand U32143 (N_32143,N_31550,N_30030);
nand U32144 (N_32144,N_30403,N_31560);
nand U32145 (N_32145,N_30519,N_30664);
or U32146 (N_32146,N_31631,N_31606);
or U32147 (N_32147,N_31596,N_31721);
or U32148 (N_32148,N_30565,N_31335);
and U32149 (N_32149,N_30978,N_30200);
and U32150 (N_32150,N_30964,N_30903);
or U32151 (N_32151,N_31115,N_30218);
and U32152 (N_32152,N_30803,N_31376);
or U32153 (N_32153,N_31960,N_31912);
nand U32154 (N_32154,N_31245,N_30345);
nor U32155 (N_32155,N_31126,N_30493);
or U32156 (N_32156,N_31811,N_30660);
and U32157 (N_32157,N_30971,N_30408);
xor U32158 (N_32158,N_31521,N_31853);
nor U32159 (N_32159,N_30547,N_30920);
and U32160 (N_32160,N_30231,N_31024);
nor U32161 (N_32161,N_30861,N_30377);
or U32162 (N_32162,N_30531,N_31591);
or U32163 (N_32163,N_31859,N_30766);
nor U32164 (N_32164,N_30907,N_31568);
xnor U32165 (N_32165,N_31585,N_30734);
nor U32166 (N_32166,N_30188,N_30745);
or U32167 (N_32167,N_30539,N_30104);
or U32168 (N_32168,N_30872,N_30642);
or U32169 (N_32169,N_31820,N_31458);
nand U32170 (N_32170,N_31695,N_30756);
and U32171 (N_32171,N_31535,N_30608);
nor U32172 (N_32172,N_30067,N_30584);
and U32173 (N_32173,N_30982,N_31474);
and U32174 (N_32174,N_31974,N_30657);
and U32175 (N_32175,N_31002,N_30382);
or U32176 (N_32176,N_31897,N_31862);
and U32177 (N_32177,N_31269,N_30790);
nand U32178 (N_32178,N_31850,N_31042);
nor U32179 (N_32179,N_31543,N_31506);
and U32180 (N_32180,N_30958,N_31996);
and U32181 (N_32181,N_31830,N_31909);
and U32182 (N_32182,N_31275,N_30292);
nand U32183 (N_32183,N_30595,N_31014);
and U32184 (N_32184,N_31186,N_31575);
or U32185 (N_32185,N_31231,N_31232);
nand U32186 (N_32186,N_30117,N_30169);
and U32187 (N_32187,N_30606,N_30508);
nor U32188 (N_32188,N_31858,N_31848);
nor U32189 (N_32189,N_30996,N_30258);
or U32190 (N_32190,N_31613,N_30155);
or U32191 (N_32191,N_30825,N_30040);
and U32192 (N_32192,N_31834,N_30543);
and U32193 (N_32193,N_30692,N_30723);
or U32194 (N_32194,N_31650,N_31663);
nor U32195 (N_32195,N_31039,N_30019);
or U32196 (N_32196,N_30923,N_30863);
nor U32197 (N_32197,N_31717,N_30305);
and U32198 (N_32198,N_30732,N_31095);
nor U32199 (N_32199,N_30325,N_30516);
or U32200 (N_32200,N_31915,N_30517);
and U32201 (N_32201,N_31479,N_30241);
or U32202 (N_32202,N_30896,N_30459);
nand U32203 (N_32203,N_30894,N_30367);
xor U32204 (N_32204,N_31803,N_30998);
or U32205 (N_32205,N_31133,N_30114);
and U32206 (N_32206,N_30405,N_31137);
nor U32207 (N_32207,N_30794,N_31369);
nor U32208 (N_32208,N_31327,N_30039);
or U32209 (N_32209,N_30447,N_31668);
or U32210 (N_32210,N_31138,N_30560);
nand U32211 (N_32211,N_30946,N_31682);
nand U32212 (N_32212,N_31316,N_30844);
xor U32213 (N_32213,N_30043,N_31489);
nor U32214 (N_32214,N_31084,N_30107);
nand U32215 (N_32215,N_30130,N_31553);
or U32216 (N_32216,N_30167,N_31325);
nor U32217 (N_32217,N_30928,N_30514);
nor U32218 (N_32218,N_31121,N_31514);
nand U32219 (N_32219,N_30787,N_31781);
or U32220 (N_32220,N_30221,N_31630);
and U32221 (N_32221,N_30486,N_30165);
nor U32222 (N_32222,N_31467,N_31922);
or U32223 (N_32223,N_30409,N_30942);
nor U32224 (N_32224,N_31660,N_31666);
and U32225 (N_32225,N_30774,N_30666);
nor U32226 (N_32226,N_31750,N_30712);
nand U32227 (N_32227,N_31878,N_30441);
nor U32228 (N_32228,N_30386,N_30161);
nand U32229 (N_32229,N_31677,N_30554);
nor U32230 (N_32230,N_30350,N_31236);
and U32231 (N_32231,N_31639,N_30481);
nand U32232 (N_32232,N_30203,N_30223);
nor U32233 (N_32233,N_30967,N_30651);
nand U32234 (N_32234,N_31833,N_31885);
or U32235 (N_32235,N_30580,N_30784);
nor U32236 (N_32236,N_31444,N_30972);
or U32237 (N_32237,N_30212,N_31676);
or U32238 (N_32238,N_30273,N_30160);
and U32239 (N_32239,N_31526,N_30432);
or U32240 (N_32240,N_30413,N_31290);
and U32241 (N_32241,N_31598,N_31954);
and U32242 (N_32242,N_31378,N_30949);
nor U32243 (N_32243,N_31563,N_30384);
nand U32244 (N_32244,N_31829,N_30764);
nor U32245 (N_32245,N_30577,N_30332);
nor U32246 (N_32246,N_30498,N_31111);
nor U32247 (N_32247,N_31463,N_30518);
nor U32248 (N_32248,N_30821,N_30975);
and U32249 (N_32249,N_31083,N_30973);
and U32250 (N_32250,N_30709,N_31293);
or U32251 (N_32251,N_31653,N_30851);
and U32252 (N_32252,N_31782,N_30751);
nor U32253 (N_32253,N_30007,N_31751);
and U32254 (N_32254,N_31099,N_31004);
nor U32255 (N_32255,N_31888,N_30575);
and U32256 (N_32256,N_31023,N_31825);
and U32257 (N_32257,N_31226,N_31818);
or U32258 (N_32258,N_31168,N_31520);
nand U32259 (N_32259,N_30809,N_30237);
nor U32260 (N_32260,N_30980,N_30867);
nand U32261 (N_32261,N_31502,N_30954);
or U32262 (N_32262,N_30747,N_30852);
and U32263 (N_32263,N_30735,N_31821);
and U32264 (N_32264,N_31798,N_30619);
or U32265 (N_32265,N_30082,N_30737);
nor U32266 (N_32266,N_30358,N_30308);
nor U32267 (N_32267,N_31465,N_30715);
nor U32268 (N_32268,N_30799,N_31880);
and U32269 (N_32269,N_30031,N_30049);
nand U32270 (N_32270,N_31572,N_30146);
nand U32271 (N_32271,N_30773,N_30816);
and U32272 (N_32272,N_31298,N_30417);
or U32273 (N_32273,N_31225,N_30801);
nand U32274 (N_32274,N_31985,N_30625);
or U32275 (N_32275,N_31430,N_31835);
and U32276 (N_32276,N_31735,N_30912);
or U32277 (N_32277,N_31920,N_30392);
nor U32278 (N_32278,N_30476,N_31051);
or U32279 (N_32279,N_30181,N_31516);
nor U32280 (N_32280,N_31643,N_31333);
or U32281 (N_32281,N_31658,N_30677);
or U32282 (N_32282,N_31059,N_31918);
or U32283 (N_32283,N_30210,N_31056);
nor U32284 (N_32284,N_30639,N_30778);
and U32285 (N_32285,N_31569,N_31667);
nor U32286 (N_32286,N_30635,N_30211);
nor U32287 (N_32287,N_31125,N_30111);
or U32288 (N_32288,N_30621,N_31340);
nor U32289 (N_32289,N_30437,N_31080);
or U32290 (N_32290,N_31565,N_30419);
or U32291 (N_32291,N_30479,N_30596);
and U32292 (N_32292,N_31986,N_31066);
nand U32293 (N_32293,N_30995,N_30829);
or U32294 (N_32294,N_31692,N_30785);
or U32295 (N_32295,N_31234,N_30850);
nand U32296 (N_32296,N_31992,N_31970);
nand U32297 (N_32297,N_31075,N_31855);
nor U32298 (N_32298,N_30857,N_30572);
nand U32299 (N_32299,N_30620,N_31701);
xnor U32300 (N_32300,N_30855,N_30257);
nand U32301 (N_32301,N_31883,N_30738);
nand U32302 (N_32302,N_30703,N_30477);
and U32303 (N_32303,N_30742,N_31481);
nand U32304 (N_32304,N_31337,N_31132);
and U32305 (N_32305,N_30892,N_31578);
xor U32306 (N_32306,N_30690,N_30669);
and U32307 (N_32307,N_30006,N_31373);
and U32308 (N_32308,N_30931,N_31582);
and U32309 (N_32309,N_31007,N_31372);
and U32310 (N_32310,N_31267,N_30434);
or U32311 (N_32311,N_31697,N_30264);
nand U32312 (N_32312,N_30286,N_30597);
nand U32313 (N_32313,N_30033,N_30243);
or U32314 (N_32314,N_30120,N_31383);
nor U32315 (N_32315,N_31927,N_31562);
or U32316 (N_32316,N_31884,N_31640);
nor U32317 (N_32317,N_30314,N_30618);
and U32318 (N_32318,N_30665,N_30583);
nand U32319 (N_32319,N_30720,N_30804);
and U32320 (N_32320,N_31434,N_31449);
and U32321 (N_32321,N_31832,N_30913);
nand U32322 (N_32322,N_31251,N_31747);
or U32323 (N_32323,N_31509,N_30848);
and U32324 (N_32324,N_30094,N_31431);
or U32325 (N_32325,N_31581,N_31969);
nor U32326 (N_32326,N_30250,N_30573);
and U32327 (N_32327,N_30485,N_30772);
and U32328 (N_32328,N_31405,N_30144);
or U32329 (N_32329,N_30369,N_30961);
nand U32330 (N_32330,N_30840,N_31401);
and U32331 (N_32331,N_30823,N_30046);
nor U32332 (N_32332,N_31845,N_31925);
nor U32333 (N_32333,N_30225,N_31813);
nor U32334 (N_32334,N_30014,N_31898);
and U32335 (N_32335,N_31698,N_30627);
or U32336 (N_32336,N_31272,N_30676);
nand U32337 (N_32337,N_31193,N_30371);
nand U32338 (N_32338,N_30224,N_31902);
or U32339 (N_32339,N_30798,N_31249);
or U32340 (N_32340,N_31044,N_31365);
and U32341 (N_32341,N_30334,N_30933);
and U32342 (N_32342,N_31744,N_30397);
nand U32343 (N_32343,N_30242,N_31800);
or U32344 (N_32344,N_31264,N_30015);
nand U32345 (N_32345,N_30421,N_31905);
and U32346 (N_32346,N_31426,N_30939);
nand U32347 (N_32347,N_31793,N_31860);
nand U32348 (N_32348,N_31958,N_31425);
nand U32349 (N_32349,N_31973,N_30901);
and U32350 (N_32350,N_30455,N_30145);
nand U32351 (N_32351,N_31686,N_30873);
nand U32352 (N_32352,N_30797,N_30157);
or U32353 (N_32353,N_30278,N_30407);
xnor U32354 (N_32354,N_30159,N_31375);
nor U32355 (N_32355,N_31665,N_30347);
nor U32356 (N_32356,N_31386,N_30411);
and U32357 (N_32357,N_30429,N_31552);
or U32358 (N_32358,N_30119,N_31017);
nor U32359 (N_32359,N_30202,N_30856);
nand U32360 (N_32360,N_31198,N_31504);
and U32361 (N_32361,N_30615,N_30687);
or U32362 (N_32362,N_31913,N_31224);
nand U32363 (N_32363,N_31929,N_31768);
nor U32364 (N_32364,N_30143,N_31062);
and U32365 (N_32365,N_31910,N_31157);
nor U32366 (N_32366,N_31556,N_31739);
and U32367 (N_32367,N_30529,N_30948);
nor U32368 (N_32368,N_31900,N_31822);
xor U32369 (N_32369,N_30324,N_30261);
and U32370 (N_32370,N_31574,N_31214);
nor U32371 (N_32371,N_30003,N_31261);
nand U32372 (N_32372,N_31619,N_30449);
nor U32373 (N_32373,N_30187,N_31466);
or U32374 (N_32374,N_30026,N_31594);
nor U32375 (N_32375,N_30500,N_30173);
or U32376 (N_32376,N_30194,N_30527);
or U32377 (N_32377,N_31684,N_31001);
nand U32378 (N_32378,N_31632,N_30849);
or U32379 (N_32379,N_31470,N_30368);
or U32380 (N_32380,N_30541,N_31141);
or U32381 (N_32381,N_31841,N_30689);
xnor U32382 (N_32382,N_30021,N_30400);
and U32383 (N_32383,N_31306,N_31368);
or U32384 (N_32384,N_30398,N_30259);
or U32385 (N_32385,N_30057,N_30636);
and U32386 (N_32386,N_30297,N_30462);
and U32387 (N_32387,N_31435,N_30668);
or U32388 (N_32388,N_31093,N_30528);
and U32389 (N_32389,N_31573,N_31314);
or U32390 (N_32390,N_31309,N_30593);
nand U32391 (N_32391,N_30700,N_31360);
or U32392 (N_32392,N_30337,N_31705);
nor U32393 (N_32393,N_31627,N_30945);
nor U32394 (N_32394,N_30836,N_30071);
and U32395 (N_32395,N_31867,N_30876);
nor U32396 (N_32396,N_31191,N_30150);
or U32397 (N_32397,N_31257,N_30470);
xnor U32398 (N_32398,N_30880,N_30115);
nand U32399 (N_32399,N_30695,N_30535);
nand U32400 (N_32400,N_31485,N_30755);
nand U32401 (N_32401,N_30137,N_30921);
and U32402 (N_32402,N_30312,N_31807);
and U32403 (N_32403,N_31252,N_31542);
nand U32404 (N_32404,N_31713,N_30028);
or U32405 (N_32405,N_31331,N_30379);
or U32406 (N_32406,N_30044,N_31209);
nand U32407 (N_32407,N_31522,N_30316);
nand U32408 (N_32408,N_31656,N_30063);
and U32409 (N_32409,N_31105,N_30578);
and U32410 (N_32410,N_31358,N_30891);
or U32411 (N_32411,N_31764,N_31281);
or U32412 (N_32412,N_30623,N_30875);
nand U32413 (N_32413,N_30355,N_31242);
nand U32414 (N_32414,N_31265,N_30038);
nor U32415 (N_32415,N_31693,N_31802);
xor U32416 (N_32416,N_31179,N_31999);
or U32417 (N_32417,N_31652,N_31728);
nor U32418 (N_32418,N_31103,N_30557);
and U32419 (N_32419,N_30326,N_30591);
or U32420 (N_32420,N_31873,N_30075);
nand U32421 (N_32421,N_31081,N_30722);
or U32422 (N_32422,N_31784,N_30707);
nor U32423 (N_32423,N_31238,N_30862);
and U32424 (N_32424,N_31063,N_31886);
nand U32425 (N_32425,N_31626,N_31052);
xnor U32426 (N_32426,N_30468,N_31291);
or U32427 (N_32427,N_30808,N_31840);
and U32428 (N_32428,N_31068,N_31307);
nand U32429 (N_32429,N_30501,N_30065);
nor U32430 (N_32430,N_31926,N_31158);
nand U32431 (N_32431,N_30645,N_31057);
nor U32432 (N_32432,N_31207,N_31856);
nand U32433 (N_32433,N_31661,N_31319);
and U32434 (N_32434,N_30233,N_31322);
nand U32435 (N_32435,N_31143,N_31864);
and U32436 (N_32436,N_30321,N_30927);
nor U32437 (N_32437,N_30613,N_30029);
nand U32438 (N_32438,N_31445,N_30248);
and U32439 (N_32439,N_31094,N_30095);
nand U32440 (N_32440,N_31153,N_30176);
nand U32441 (N_32441,N_31758,N_31621);
nor U32442 (N_32442,N_31783,N_30634);
or U32443 (N_32443,N_30076,N_31266);
nand U32444 (N_32444,N_30582,N_30694);
nor U32445 (N_32445,N_30348,N_31899);
or U32446 (N_32446,N_31723,N_30724);
nor U32447 (N_32447,N_31382,N_30072);
nand U32448 (N_32448,N_31778,N_31407);
nor U32449 (N_32449,N_30327,N_30986);
nand U32450 (N_32450,N_30586,N_30909);
nor U32451 (N_32451,N_30287,N_31345);
or U32452 (N_32452,N_30375,N_30489);
nand U32453 (N_32453,N_31101,N_30511);
and U32454 (N_32454,N_31978,N_30889);
and U32455 (N_32455,N_31072,N_30086);
nor U32456 (N_32456,N_30926,N_31026);
and U32457 (N_32457,N_30781,N_31725);
nor U32458 (N_32458,N_31525,N_31092);
or U32459 (N_32459,N_31303,N_30533);
or U32460 (N_32460,N_31741,N_31390);
nor U32461 (N_32461,N_31685,N_30394);
nor U32462 (N_32462,N_30674,N_31997);
nor U32463 (N_32463,N_30813,N_31471);
nor U32464 (N_32464,N_31921,N_31476);
nand U32465 (N_32465,N_31175,N_30282);
nand U32466 (N_32466,N_30277,N_31648);
or U32467 (N_32467,N_30189,N_30824);
and U32468 (N_32468,N_31418,N_30553);
or U32469 (N_32469,N_31442,N_31647);
or U32470 (N_32470,N_31181,N_30680);
nand U32471 (N_32471,N_31240,N_30336);
and U32472 (N_32472,N_31679,N_31730);
or U32473 (N_32473,N_31013,N_30739);
or U32474 (N_32474,N_31963,N_31866);
and U32475 (N_32475,N_30113,N_30842);
nand U32476 (N_32476,N_30424,N_31468);
nand U32477 (N_32477,N_30439,N_31049);
nor U32478 (N_32478,N_31381,N_30463);
or U32479 (N_32479,N_31971,N_31036);
nor U32480 (N_32480,N_30035,N_30339);
or U32481 (N_32481,N_31801,N_30060);
nand U32482 (N_32482,N_31217,N_31305);
or U32483 (N_32483,N_31184,N_30997);
and U32484 (N_32484,N_31363,N_30344);
nand U32485 (N_32485,N_31555,N_31748);
and U32486 (N_32486,N_30571,N_31586);
nor U32487 (N_32487,N_30545,N_31437);
or U32488 (N_32488,N_31454,N_30523);
nor U32489 (N_32489,N_31321,N_30898);
nor U32490 (N_32490,N_30490,N_30093);
or U32491 (N_32491,N_31324,N_30730);
and U32492 (N_32492,N_30395,N_30069);
nor U32493 (N_32493,N_31089,N_31769);
nor U32494 (N_32494,N_31961,N_30953);
nor U32495 (N_32495,N_31617,N_30180);
nand U32496 (N_32496,N_31136,N_31952);
nand U32497 (N_32497,N_31464,N_31746);
nor U32498 (N_32498,N_30109,N_30925);
nor U32499 (N_32499,N_31096,N_30299);
and U32500 (N_32500,N_30757,N_30290);
or U32501 (N_32501,N_30711,N_31540);
or U32502 (N_32502,N_31009,N_31870);
and U32503 (N_32503,N_31189,N_30793);
xnor U32504 (N_32504,N_31549,N_30648);
nand U32505 (N_32505,N_30870,N_31940);
nand U32506 (N_32506,N_30341,N_31361);
and U32507 (N_32507,N_30281,N_30168);
or U32508 (N_32508,N_30070,N_31127);
nand U32509 (N_32509,N_30260,N_30389);
or U32510 (N_32510,N_31034,N_30024);
and U32511 (N_32511,N_31812,N_30291);
and U32512 (N_32512,N_30085,N_31432);
nor U32513 (N_32513,N_31943,N_31021);
or U32514 (N_32514,N_30616,N_30385);
and U32515 (N_32515,N_30234,N_31387);
nor U32516 (N_32516,N_30807,N_30924);
nand U32517 (N_32517,N_30633,N_30087);
nor U32518 (N_32518,N_31196,N_30083);
and U32519 (N_32519,N_31819,N_31791);
nand U32520 (N_32520,N_31352,N_30000);
nand U32521 (N_32521,N_30915,N_31134);
nor U32522 (N_32522,N_31045,N_31180);
xor U32523 (N_32523,N_30746,N_31616);
xnor U32524 (N_32524,N_30055,N_31112);
or U32525 (N_32525,N_31341,N_30088);
or U32526 (N_32526,N_30767,N_30826);
nor U32527 (N_32527,N_30228,N_31423);
xnor U32528 (N_32528,N_31965,N_31895);
or U32529 (N_32529,N_30579,N_31086);
nor U32530 (N_32530,N_30663,N_31871);
or U32531 (N_32531,N_30002,N_31842);
and U32532 (N_32532,N_31945,N_30637);
or U32533 (N_32533,N_30238,N_30232);
and U32534 (N_32534,N_30888,N_30343);
nand U32535 (N_32535,N_31559,N_30182);
nand U32536 (N_32536,N_30594,N_31592);
nor U32537 (N_32537,N_31919,N_31491);
nor U32538 (N_32538,N_31032,N_30828);
nor U32539 (N_32539,N_30340,N_30438);
nand U32540 (N_32540,N_30175,N_31177);
and U32541 (N_32541,N_30244,N_30461);
or U32542 (N_32542,N_30987,N_31299);
nand U32543 (N_32543,N_30199,N_30162);
and U32544 (N_32544,N_30934,N_31979);
nand U32545 (N_32545,N_31637,N_31877);
nand U32546 (N_32546,N_31618,N_31947);
nor U32547 (N_32547,N_31939,N_31348);
nor U32548 (N_32548,N_30937,N_30537);
nand U32549 (N_32549,N_30487,N_31711);
and U32550 (N_32550,N_30929,N_30626);
or U32551 (N_32551,N_31456,N_31060);
nor U32552 (N_32552,N_31706,N_30124);
or U32553 (N_32553,N_30567,N_30789);
or U32554 (N_32554,N_30605,N_31875);
nand U32555 (N_32555,N_30505,N_30708);
nand U32556 (N_32556,N_30318,N_31689);
nand U32557 (N_32557,N_31863,N_30435);
and U32558 (N_32558,N_30091,N_31539);
nand U32559 (N_32559,N_31347,N_31681);
nor U32560 (N_32560,N_31478,N_30274);
nand U32561 (N_32561,N_30638,N_31278);
or U32562 (N_32562,N_31005,N_31988);
xnor U32563 (N_32563,N_31461,N_31508);
nand U32564 (N_32564,N_30184,N_30992);
or U32565 (N_32565,N_31019,N_31576);
nand U32566 (N_32566,N_31113,N_31704);
nand U32567 (N_32567,N_31422,N_30731);
and U32568 (N_32568,N_31738,N_30811);
xor U32569 (N_32569,N_31852,N_31731);
and U32570 (N_32570,N_31030,N_30559);
nand U32571 (N_32571,N_30688,N_30860);
nor U32572 (N_32572,N_30262,N_30027);
nand U32573 (N_32573,N_31200,N_31745);
nor U32574 (N_32574,N_30994,N_30304);
or U32575 (N_32575,N_31792,N_31737);
and U32576 (N_32576,N_30158,N_30456);
nor U32577 (N_32577,N_30017,N_31959);
or U32578 (N_32578,N_31429,N_30658);
nand U32579 (N_32579,N_31343,N_30236);
nor U32580 (N_32580,N_30877,N_31284);
and U32581 (N_32581,N_30041,N_31931);
or U32582 (N_32582,N_31923,N_30020);
nand U32583 (N_32583,N_31500,N_30699);
or U32584 (N_32584,N_30854,N_30979);
and U32585 (N_32585,N_30555,N_30208);
or U32586 (N_32586,N_31452,N_31167);
nand U32587 (N_32587,N_31396,N_31691);
nand U32588 (N_32588,N_30696,N_31006);
and U32589 (N_32589,N_31473,N_31622);
nand U32590 (N_32590,N_31505,N_31823);
and U32591 (N_32591,N_30691,N_30871);
nand U32592 (N_32592,N_30552,N_30422);
or U32593 (N_32593,N_31164,N_31109);
nand U32594 (N_32594,N_30374,N_31771);
nand U32595 (N_32595,N_30974,N_31355);
or U32596 (N_32596,N_30240,N_31987);
and U32597 (N_32597,N_30270,N_31227);
nand U32598 (N_32598,N_31523,N_31397);
or U32599 (N_32599,N_30331,N_30288);
or U32600 (N_32600,N_30078,N_30362);
nor U32601 (N_32601,N_31770,N_30148);
and U32602 (N_32602,N_31669,N_30686);
or U32603 (N_32603,N_30296,N_31380);
or U32604 (N_32604,N_30365,N_30499);
nand U32605 (N_32605,N_31218,N_31734);
nand U32606 (N_32606,N_31982,N_30156);
or U32607 (N_32607,N_30675,N_30908);
and U32608 (N_32608,N_31263,N_31908);
nand U32609 (N_32609,N_31893,N_30568);
or U32610 (N_32610,N_31846,N_31446);
nand U32611 (N_32611,N_31743,N_30079);
nand U32612 (N_32612,N_31069,N_31503);
nand U32613 (N_32613,N_31561,N_31674);
or U32614 (N_32614,N_31160,N_31147);
or U32615 (N_32615,N_31749,N_31472);
or U32616 (N_32616,N_30656,N_31903);
nand U32617 (N_32617,N_30492,N_30363);
and U32618 (N_32618,N_31313,N_31336);
nand U32619 (N_32619,N_31283,N_31199);
or U32620 (N_32620,N_30991,N_31118);
or U32621 (N_32621,N_30815,N_30906);
or U32622 (N_32622,N_30206,N_30373);
nand U32623 (N_32623,N_30662,N_30782);
or U32624 (N_32624,N_30985,N_30900);
or U32625 (N_32625,N_30752,N_31487);
or U32626 (N_32626,N_30172,N_31150);
nand U32627 (N_32627,N_31027,N_31805);
nor U32628 (N_32628,N_31402,N_30298);
nor U32629 (N_32629,N_31541,N_30885);
xnor U32630 (N_32630,N_31403,N_31804);
nor U32631 (N_32631,N_31797,N_31752);
nand U32632 (N_32632,N_30736,N_30940);
nand U32633 (N_32633,N_30034,N_31326);
nand U32634 (N_32634,N_31018,N_31259);
and U32635 (N_32635,N_30285,N_30515);
or U32636 (N_32636,N_30938,N_30062);
or U32637 (N_32637,N_31527,N_30959);
nor U32638 (N_32638,N_30726,N_31795);
nand U32639 (N_32639,N_31248,N_30585);
or U32640 (N_32640,N_31195,N_31890);
and U32641 (N_32641,N_31339,N_31760);
nor U32642 (N_32642,N_30280,N_30475);
nor U32643 (N_32643,N_31308,N_31108);
and U32644 (N_32644,N_30976,N_30471);
nor U32645 (N_32645,N_30092,N_30426);
and U32646 (N_32646,N_30139,N_31602);
and U32647 (N_32647,N_31392,N_31683);
nor U32648 (N_32648,N_30378,N_30783);
nor U32649 (N_32649,N_31448,N_30603);
nor U32650 (N_32650,N_31228,N_30320);
or U32651 (N_32651,N_30440,N_31937);
and U32652 (N_32652,N_30788,N_30874);
nand U32653 (N_32653,N_30205,N_30154);
or U32654 (N_32654,N_30253,N_30744);
nor U32655 (N_32655,N_30762,N_30293);
nor U32656 (N_32656,N_30247,N_31536);
nand U32657 (N_32657,N_30322,N_31498);
nor U32658 (N_32658,N_31486,N_30214);
and U32659 (N_32659,N_31398,N_31597);
nand U32660 (N_32660,N_31545,N_30335);
nand U32661 (N_32661,N_31501,N_31330);
nor U32662 (N_32662,N_31172,N_31244);
and U32663 (N_32663,N_30153,N_30963);
xor U32664 (N_32664,N_30183,N_30497);
nand U32665 (N_32665,N_30122,N_30704);
nor U32666 (N_32666,N_30966,N_31304);
nor U32667 (N_32667,N_30256,N_30701);
nor U32668 (N_32668,N_31814,N_30930);
nand U32669 (N_32669,N_30955,N_31353);
and U32670 (N_32670,N_30835,N_30679);
nand U32671 (N_32671,N_31149,N_30749);
and U32672 (N_32672,N_30163,N_31271);
nor U32673 (N_32673,N_31600,N_31241);
nor U32674 (N_32674,N_30977,N_31102);
and U32675 (N_32675,N_30191,N_30569);
and U32676 (N_32676,N_31098,N_31182);
and U32677 (N_32677,N_30905,N_30473);
or U32678 (N_32678,N_31649,N_31716);
xnor U32679 (N_32679,N_30513,N_30217);
nor U32680 (N_32680,N_30878,N_31462);
and U32681 (N_32681,N_31625,N_31824);
and U32682 (N_32682,N_30952,N_30170);
xor U32683 (N_32683,N_30721,N_30989);
xnor U32684 (N_32684,N_30916,N_30883);
nand U32685 (N_32685,N_31991,N_30598);
nor U32686 (N_32686,N_30406,N_30831);
or U32687 (N_32687,N_30219,N_30306);
xnor U32688 (N_32688,N_31332,N_31608);
and U32689 (N_32689,N_30098,N_31732);
or U32690 (N_32690,N_31759,N_30276);
or U32691 (N_32691,N_30881,N_31938);
or U32692 (N_32692,N_30682,N_30201);
nor U32693 (N_32693,N_30748,N_31443);
or U32694 (N_32694,N_31197,N_30338);
or U32695 (N_32695,N_31496,N_30005);
nand U32696 (N_32696,N_31651,N_30502);
nor U32697 (N_32697,N_30957,N_30681);
nand U32698 (N_32698,N_31282,N_30383);
nand U32699 (N_32699,N_31201,N_31208);
and U32700 (N_32700,N_31100,N_30142);
or U32701 (N_32701,N_31876,N_31250);
or U32702 (N_32702,N_30526,N_30246);
nor U32703 (N_32703,N_30558,N_30352);
nand U32704 (N_32704,N_31534,N_30230);
and U32705 (N_32705,N_31416,N_30249);
nor U32706 (N_32706,N_31907,N_31570);
nor U32707 (N_32707,N_30534,N_31595);
and U32708 (N_32708,N_30706,N_31657);
or U32709 (N_32709,N_31808,N_31176);
nand U32710 (N_32710,N_30301,N_30768);
nand U32711 (N_32711,N_30448,N_30023);
or U32712 (N_32712,N_31547,N_31843);
and U32713 (N_32713,N_30460,N_31493);
nand U32714 (N_32714,N_31949,N_30370);
nor U32715 (N_32715,N_31611,N_31928);
nor U32716 (N_32716,N_30333,N_30546);
nor U32717 (N_32717,N_30099,N_30484);
or U32718 (N_32718,N_31482,N_31975);
or U32719 (N_32719,N_31957,N_31377);
nand U32720 (N_32720,N_31156,N_30536);
nand U32721 (N_32721,N_30822,N_31524);
and U32722 (N_32722,N_30444,N_30743);
nand U32723 (N_32723,N_30051,N_31646);
nor U32724 (N_32724,N_31273,N_30178);
and U32725 (N_32725,N_30614,N_30255);
nand U32726 (N_32726,N_31794,N_30759);
or U32727 (N_32727,N_30670,N_30089);
nand U32728 (N_32728,N_30396,N_30530);
or U32729 (N_32729,N_31517,N_31869);
nand U32730 (N_32730,N_30965,N_31490);
nor U32731 (N_32731,N_31736,N_31040);
or U32732 (N_32732,N_31995,N_31636);
or U32733 (N_32733,N_30671,N_30025);
nor U32734 (N_32734,N_30520,N_31579);
or U32735 (N_32735,N_30705,N_31351);
or U32736 (N_32736,N_31000,N_31243);
nor U32737 (N_32737,N_31117,N_30453);
nand U32738 (N_32738,N_31773,N_30442);
or U32739 (N_32739,N_31488,N_31510);
nand U32740 (N_32740,N_30399,N_31624);
nor U32741 (N_32741,N_30207,N_30008);
nor U32742 (N_32742,N_31455,N_31762);
nor U32743 (N_32743,N_30268,N_31967);
and U32744 (N_32744,N_31076,N_31806);
xor U32745 (N_32745,N_31911,N_31810);
or U32746 (N_32746,N_30503,N_30956);
nor U32747 (N_32747,N_30609,N_30812);
or U32748 (N_32748,N_31699,N_30612);
or U32749 (N_32749,N_30445,N_31499);
and U32750 (N_32750,N_31016,N_31302);
or U32751 (N_32751,N_30220,N_31260);
nand U32752 (N_32752,N_31417,N_31874);
nand U32753 (N_32753,N_31844,N_31411);
nand U32754 (N_32754,N_30890,N_30918);
or U32755 (N_32755,N_31495,N_31048);
nor U32756 (N_32756,N_30048,N_31367);
nand U32757 (N_32757,N_31215,N_30544);
nand U32758 (N_32758,N_30904,N_31554);
nand U32759 (N_32759,N_31515,N_30204);
nand U32760 (N_32760,N_31349,N_30999);
nor U32761 (N_32761,N_30646,N_31831);
nand U32762 (N_32762,N_31709,N_30100);
nor U32763 (N_32763,N_30131,N_31033);
nor U32764 (N_32764,N_30819,N_30792);
and U32765 (N_32765,N_31104,N_30045);
nor U32766 (N_32766,N_31917,N_31765);
and U32767 (N_32767,N_30727,N_31296);
and U32768 (N_32768,N_30846,N_30581);
nor U32769 (N_32769,N_30315,N_31708);
nor U32770 (N_32770,N_30284,N_30271);
nor U32771 (N_32771,N_31148,N_30968);
nor U32772 (N_32772,N_31851,N_30897);
and U32773 (N_32773,N_30628,N_30683);
nor U32774 (N_32774,N_31071,N_30960);
or U32775 (N_32775,N_31145,N_31588);
nand U32776 (N_32776,N_31029,N_31754);
and U32777 (N_32777,N_30430,N_30009);
nand U32778 (N_32778,N_30140,N_31440);
or U32779 (N_32779,N_31438,N_31513);
and U32780 (N_32780,N_31497,N_30404);
nor U32781 (N_32781,N_31041,N_31090);
nor U32782 (N_32782,N_31171,N_31120);
nand U32783 (N_32783,N_30116,N_31031);
nor U32784 (N_32784,N_31253,N_30504);
nor U32785 (N_32785,N_31577,N_31140);
xor U32786 (N_32786,N_31906,N_31010);
and U32787 (N_32787,N_30866,N_30817);
nand U32788 (N_32788,N_31406,N_31789);
nand U32789 (N_32789,N_31815,N_31055);
nor U32790 (N_32790,N_31887,N_30192);
nand U32791 (N_32791,N_31664,N_30001);
nand U32792 (N_32792,N_30886,N_31934);
nor U32793 (N_32793,N_31035,N_31216);
and U32794 (N_32794,N_30010,N_31294);
or U32795 (N_32795,N_30133,N_31277);
nand U32796 (N_32796,N_30983,N_30693);
nor U32797 (N_32797,N_30084,N_30401);
nor U32798 (N_32798,N_30919,N_30491);
nor U32799 (N_32799,N_31777,N_30841);
and U32800 (N_32800,N_31775,N_31936);
and U32801 (N_32801,N_31796,N_31371);
nor U32802 (N_32802,N_31659,N_30118);
and U32803 (N_32803,N_31135,N_31836);
nand U32804 (N_32804,N_30077,N_31892);
or U32805 (N_32805,N_30653,N_31106);
nor U32806 (N_32806,N_31593,N_30622);
or U32807 (N_32807,N_30587,N_30436);
or U32808 (N_32808,N_31469,N_30121);
or U32809 (N_32809,N_30740,N_30235);
and U32810 (N_32810,N_30549,N_31548);
nor U32811 (N_32811,N_30171,N_30791);
nand U32812 (N_32812,N_31655,N_30521);
or U32813 (N_32813,N_31202,N_30770);
xor U32814 (N_32814,N_31518,N_31130);
nand U32815 (N_32815,N_31635,N_31285);
or U32816 (N_32816,N_31222,N_31450);
and U32817 (N_32817,N_31344,N_30510);
or U32818 (N_32818,N_31129,N_30943);
or U32819 (N_32819,N_30685,N_31116);
nand U32820 (N_32820,N_30126,N_30641);
nand U32821 (N_32821,N_30080,N_31687);
nand U32822 (N_32822,N_31268,N_31571);
nor U32823 (N_32823,N_31930,N_31128);
nor U32824 (N_32824,N_31977,N_30295);
or U32825 (N_32825,N_31710,N_30391);
and U32826 (N_32826,N_30420,N_30522);
nor U32827 (N_32827,N_30052,N_31276);
and U32828 (N_32828,N_30390,N_30548);
and U32829 (N_32829,N_31718,N_30357);
nor U32830 (N_32830,N_30714,N_31615);
or U32831 (N_32831,N_30865,N_30832);
nor U32832 (N_32832,N_31531,N_30540);
and U32833 (N_32833,N_30198,N_30837);
nand U32834 (N_32834,N_31696,N_30882);
nor U32835 (N_32835,N_31700,N_30252);
nand U32836 (N_32836,N_30127,N_31690);
and U32837 (N_32837,N_30643,N_31289);
nor U32838 (N_32838,N_31220,N_30993);
nand U32839 (N_32839,N_31955,N_30229);
nor U32840 (N_32840,N_30074,N_30551);
nor U32841 (N_32841,N_30061,N_31567);
xor U32842 (N_32842,N_31097,N_30387);
nand U32843 (N_32843,N_31720,N_31799);
nor U32844 (N_32844,N_30718,N_31962);
and U32845 (N_32845,N_31163,N_30054);
and U32846 (N_32846,N_31053,N_30457);
nor U32847 (N_32847,N_30610,N_30110);
and U32848 (N_32848,N_31328,N_30624);
nand U32849 (N_32849,N_31279,N_30059);
or U32850 (N_32850,N_30402,N_31671);
nand U32851 (N_32851,N_31872,N_31511);
nor U32852 (N_32852,N_30725,N_30388);
and U32853 (N_32853,N_31953,N_31254);
and U32854 (N_32854,N_31605,N_31151);
and U32855 (N_32855,N_30372,N_30311);
nor U32856 (N_32856,N_31933,N_31868);
and U32857 (N_32857,N_30602,N_31122);
nand U32858 (N_32858,N_31292,N_30190);
nor U32859 (N_32859,N_30464,N_31623);
or U32860 (N_32860,N_31891,N_31154);
and U32861 (N_32861,N_31246,N_30818);
or U32862 (N_32862,N_30427,N_31237);
nor U32863 (N_32863,N_31675,N_30570);
and U32864 (N_32864,N_30018,N_30239);
nand U32865 (N_32865,N_30710,N_30423);
or U32866 (N_32866,N_30506,N_31673);
nand U32867 (N_32867,N_30838,N_30414);
or U32868 (N_32868,N_30310,N_30800);
nor U32869 (N_32869,N_31190,N_30847);
and U32870 (N_32870,N_30068,N_30525);
or U32871 (N_32871,N_31827,N_30467);
and U32872 (N_32872,N_31688,N_30469);
or U32873 (N_32873,N_30512,N_31318);
or U32874 (N_32874,N_30215,N_31724);
or U32875 (N_32875,N_30058,N_30769);
nor U32876 (N_32876,N_31229,N_30632);
nor U32877 (N_32877,N_30914,N_31447);
nor U32878 (N_32878,N_31589,N_30177);
or U32879 (N_32879,N_31894,N_31221);
nand U32880 (N_32880,N_31370,N_30112);
and U32881 (N_32881,N_31070,N_30433);
xor U32882 (N_32882,N_31601,N_31323);
nand U32883 (N_32883,N_31584,N_31896);
xnor U32884 (N_32884,N_30309,N_30853);
nand U32885 (N_32885,N_30478,N_31480);
nor U32886 (N_32886,N_31067,N_31879);
or U32887 (N_32887,N_31320,N_31946);
and U32888 (N_32888,N_30354,N_30227);
nor U32889 (N_32889,N_31082,N_31566);
nand U32890 (N_32890,N_30410,N_31849);
or U32891 (N_32891,N_30899,N_30186);
nor U32892 (N_32892,N_31756,N_31678);
xnor U32893 (N_32893,N_31047,N_31610);
and U32894 (N_32894,N_30936,N_31110);
nor U32895 (N_32895,N_30509,N_30147);
or U32896 (N_32896,N_30827,N_30141);
nor U32897 (N_32897,N_30951,N_31941);
xnor U32898 (N_32898,N_30845,N_30346);
and U32899 (N_32899,N_31532,N_30135);
or U32900 (N_32900,N_30728,N_30267);
or U32901 (N_32901,N_30313,N_30053);
nor U32902 (N_32902,N_30179,N_31956);
or U32903 (N_32903,N_31428,N_30564);
or U32904 (N_32904,N_30032,N_31857);
nand U32905 (N_32905,N_31564,N_31530);
nor U32906 (N_32906,N_30136,N_30185);
and U32907 (N_32907,N_31942,N_30351);
or U32908 (N_32908,N_30474,N_31310);
nand U32909 (N_32909,N_30102,N_31295);
nand U32910 (N_32910,N_31439,N_31139);
or U32911 (N_32911,N_30950,N_30984);
or U32912 (N_32912,N_31424,N_31211);
nand U32913 (N_32913,N_30771,N_30650);
nand U32914 (N_32914,N_31185,N_30729);
or U32915 (N_32915,N_31114,N_30947);
nand U32916 (N_32916,N_30902,N_31011);
and U32917 (N_32917,N_30702,N_31043);
or U32918 (N_32918,N_30600,N_30307);
nand U32919 (N_32919,N_31966,N_30096);
nor U32920 (N_32920,N_31107,N_31412);
nor U32921 (N_32921,N_30226,N_30056);
and U32922 (N_32922,N_30272,N_31393);
or U32923 (N_32923,N_30300,N_31421);
nand U32924 (N_32924,N_31839,N_31038);
and U32925 (N_32925,N_31475,N_31715);
nor U32926 (N_32926,N_30673,N_30758);
and U32927 (N_32927,N_31223,N_31620);
nand U32928 (N_32928,N_30090,N_30884);
nand U32929 (N_32929,N_31914,N_30599);
nor U32930 (N_32930,N_30342,N_30004);
nand U32931 (N_32931,N_30466,N_30323);
or U32932 (N_32932,N_30047,N_30910);
nor U32933 (N_32933,N_31012,N_31235);
nand U32934 (N_32934,N_31146,N_30472);
nor U32935 (N_32935,N_30458,N_31980);
and U32936 (N_32936,N_31085,N_31203);
nand U32937 (N_32937,N_30105,N_31916);
nand U32938 (N_32938,N_31972,N_31484);
nand U32939 (N_32939,N_30016,N_30542);
nor U32940 (N_32940,N_30302,N_31787);
nor U32941 (N_32941,N_30970,N_30289);
nor U32942 (N_32942,N_31629,N_30576);
and U32943 (N_32943,N_30672,N_30073);
nor U32944 (N_32944,N_31015,N_31079);
and U32945 (N_32945,N_31528,N_30364);
and U32946 (N_32946,N_31790,N_30275);
nand U32947 (N_32947,N_31419,N_31707);
nor U32948 (N_32948,N_31064,N_30775);
nand U32949 (N_32949,N_31212,N_30969);
nand U32950 (N_32950,N_30381,N_30869);
and U32951 (N_32951,N_31628,N_31194);
nor U32952 (N_32952,N_30152,N_31028);
or U32953 (N_32953,N_31362,N_31173);
xnor U32954 (N_32954,N_30488,N_31003);
nand U32955 (N_32955,N_30480,N_30022);
or U32956 (N_32956,N_31162,N_31451);
nor U32957 (N_32957,N_31983,N_30129);
and U32958 (N_32958,N_31453,N_31170);
nand U32959 (N_32959,N_30418,N_31580);
or U32960 (N_32960,N_31828,N_30574);
and U32961 (N_32961,N_30037,N_30741);
and U32962 (N_32962,N_31614,N_31415);
nand U32963 (N_32963,N_31603,N_30795);
nand U32964 (N_32964,N_30830,N_30776);
nand U32965 (N_32965,N_31779,N_31558);
and U32966 (N_32966,N_31604,N_30451);
nand U32967 (N_32967,N_30446,N_31483);
and U32968 (N_32968,N_30806,N_31590);
and U32969 (N_32969,N_30879,N_31993);
nand U32970 (N_32970,N_30868,N_31161);
or U32971 (N_32971,N_30134,N_30697);
nor U32972 (N_32972,N_31981,N_31994);
and U32973 (N_32973,N_30317,N_30655);
and U32974 (N_32974,N_30733,N_31297);
and U32975 (N_32975,N_30279,N_31740);
nand U32976 (N_32976,N_31557,N_31726);
xor U32977 (N_32977,N_30617,N_31183);
and U32978 (N_32978,N_31633,N_31388);
or U32979 (N_32979,N_31881,N_30659);
nor U32980 (N_32980,N_31258,N_31356);
nor U32981 (N_32981,N_30713,N_31385);
and U32982 (N_32982,N_30760,N_31809);
nand U32983 (N_32983,N_30495,N_31838);
nand U32984 (N_32984,N_31753,N_31761);
or U32985 (N_32985,N_31854,N_31399);
and U32986 (N_32986,N_30631,N_30524);
or U32987 (N_32987,N_30802,N_31703);
and U32988 (N_32988,N_30601,N_31607);
nor U32989 (N_32989,N_31976,N_30443);
and U32990 (N_32990,N_30962,N_31404);
and U32991 (N_32991,N_31384,N_31776);
nand U32992 (N_32992,N_31247,N_30678);
xnor U32993 (N_32993,N_30932,N_30294);
and U32994 (N_32994,N_31837,N_30805);
or U32995 (N_32995,N_31338,N_31788);
nand U32996 (N_32996,N_30496,N_30251);
or U32997 (N_32997,N_31654,N_30550);
xor U32998 (N_32998,N_30780,N_30193);
or U32999 (N_32999,N_31131,N_31315);
and U33000 (N_33000,N_31400,N_30192);
and U33001 (N_33001,N_31299,N_30075);
nand U33002 (N_33002,N_31891,N_31097);
and U33003 (N_33003,N_31484,N_30611);
nor U33004 (N_33004,N_30806,N_30862);
and U33005 (N_33005,N_30498,N_31807);
and U33006 (N_33006,N_31678,N_30777);
or U33007 (N_33007,N_30340,N_31376);
nor U33008 (N_33008,N_30026,N_31400);
nand U33009 (N_33009,N_31522,N_30095);
nand U33010 (N_33010,N_31684,N_31466);
nor U33011 (N_33011,N_30610,N_31356);
or U33012 (N_33012,N_31028,N_31528);
nor U33013 (N_33013,N_31168,N_30819);
nand U33014 (N_33014,N_31556,N_30839);
nand U33015 (N_33015,N_30854,N_31855);
xor U33016 (N_33016,N_30404,N_30181);
nand U33017 (N_33017,N_30878,N_30967);
nor U33018 (N_33018,N_31988,N_31142);
nor U33019 (N_33019,N_30679,N_30904);
nand U33020 (N_33020,N_30043,N_31611);
nand U33021 (N_33021,N_30931,N_30448);
and U33022 (N_33022,N_30028,N_30771);
or U33023 (N_33023,N_30689,N_31632);
and U33024 (N_33024,N_31554,N_31504);
and U33025 (N_33025,N_30067,N_31347);
nor U33026 (N_33026,N_30909,N_30644);
nor U33027 (N_33027,N_30969,N_30672);
and U33028 (N_33028,N_30327,N_31186);
nor U33029 (N_33029,N_30309,N_31136);
nand U33030 (N_33030,N_31516,N_30506);
or U33031 (N_33031,N_31131,N_31369);
nor U33032 (N_33032,N_31919,N_30949);
nand U33033 (N_33033,N_31975,N_31446);
and U33034 (N_33034,N_31817,N_31576);
and U33035 (N_33035,N_30903,N_31603);
nor U33036 (N_33036,N_30783,N_30999);
nand U33037 (N_33037,N_31213,N_30171);
or U33038 (N_33038,N_31913,N_30617);
and U33039 (N_33039,N_31779,N_31547);
nor U33040 (N_33040,N_31098,N_30613);
and U33041 (N_33041,N_30647,N_30956);
nor U33042 (N_33042,N_31959,N_30747);
nand U33043 (N_33043,N_30362,N_30411);
and U33044 (N_33044,N_30050,N_31395);
nor U33045 (N_33045,N_31386,N_30150);
nor U33046 (N_33046,N_31910,N_30886);
nor U33047 (N_33047,N_31487,N_30329);
nor U33048 (N_33048,N_31846,N_31947);
and U33049 (N_33049,N_30229,N_30970);
nor U33050 (N_33050,N_31913,N_31961);
nand U33051 (N_33051,N_30599,N_31429);
nand U33052 (N_33052,N_31033,N_31622);
nor U33053 (N_33053,N_31144,N_31740);
or U33054 (N_33054,N_30117,N_31669);
nand U33055 (N_33055,N_31745,N_30456);
or U33056 (N_33056,N_31939,N_31981);
nand U33057 (N_33057,N_30990,N_30179);
nand U33058 (N_33058,N_30303,N_30317);
and U33059 (N_33059,N_30394,N_31422);
or U33060 (N_33060,N_30733,N_30502);
xnor U33061 (N_33061,N_30468,N_30718);
nor U33062 (N_33062,N_31277,N_30651);
nor U33063 (N_33063,N_30465,N_31806);
nor U33064 (N_33064,N_30470,N_31092);
nand U33065 (N_33065,N_31274,N_30570);
nor U33066 (N_33066,N_30212,N_31943);
or U33067 (N_33067,N_30322,N_31965);
nor U33068 (N_33068,N_31315,N_31974);
and U33069 (N_33069,N_30931,N_31212);
nand U33070 (N_33070,N_30652,N_30221);
nand U33071 (N_33071,N_30663,N_30956);
nor U33072 (N_33072,N_30205,N_30053);
and U33073 (N_33073,N_30594,N_30868);
and U33074 (N_33074,N_31187,N_30767);
nand U33075 (N_33075,N_30275,N_31965);
nand U33076 (N_33076,N_31211,N_31936);
or U33077 (N_33077,N_30985,N_30347);
nor U33078 (N_33078,N_30351,N_30059);
and U33079 (N_33079,N_31328,N_31967);
or U33080 (N_33080,N_31020,N_30017);
or U33081 (N_33081,N_31917,N_30259);
nand U33082 (N_33082,N_30029,N_30760);
nor U33083 (N_33083,N_30884,N_31918);
nand U33084 (N_33084,N_31549,N_31100);
nor U33085 (N_33085,N_30682,N_30281);
nand U33086 (N_33086,N_31851,N_30596);
or U33087 (N_33087,N_31387,N_30503);
nor U33088 (N_33088,N_30658,N_30027);
nand U33089 (N_33089,N_31205,N_31622);
or U33090 (N_33090,N_30301,N_30927);
or U33091 (N_33091,N_31125,N_31018);
nor U33092 (N_33092,N_31739,N_30639);
and U33093 (N_33093,N_30993,N_31920);
nor U33094 (N_33094,N_31202,N_30223);
nand U33095 (N_33095,N_30250,N_31507);
or U33096 (N_33096,N_30671,N_31635);
nor U33097 (N_33097,N_30684,N_30408);
nor U33098 (N_33098,N_30027,N_31787);
nand U33099 (N_33099,N_30521,N_30663);
nor U33100 (N_33100,N_30325,N_30617);
nand U33101 (N_33101,N_31172,N_31857);
nor U33102 (N_33102,N_30644,N_31586);
nor U33103 (N_33103,N_30886,N_31501);
nand U33104 (N_33104,N_30188,N_30467);
or U33105 (N_33105,N_30168,N_30942);
nor U33106 (N_33106,N_30539,N_30275);
and U33107 (N_33107,N_31767,N_31203);
nor U33108 (N_33108,N_30018,N_30958);
nor U33109 (N_33109,N_30320,N_30640);
or U33110 (N_33110,N_30521,N_30027);
and U33111 (N_33111,N_30301,N_31386);
and U33112 (N_33112,N_31470,N_30481);
nor U33113 (N_33113,N_31377,N_31459);
nor U33114 (N_33114,N_31281,N_30821);
nand U33115 (N_33115,N_30102,N_30541);
and U33116 (N_33116,N_30317,N_30670);
or U33117 (N_33117,N_30603,N_31137);
or U33118 (N_33118,N_30678,N_30333);
and U33119 (N_33119,N_31653,N_31346);
nor U33120 (N_33120,N_31237,N_30616);
nand U33121 (N_33121,N_30811,N_30482);
and U33122 (N_33122,N_31520,N_30853);
nand U33123 (N_33123,N_30460,N_30173);
nor U33124 (N_33124,N_31751,N_30248);
and U33125 (N_33125,N_31501,N_30775);
xor U33126 (N_33126,N_30999,N_30660);
xnor U33127 (N_33127,N_30031,N_30392);
nand U33128 (N_33128,N_31333,N_31402);
nand U33129 (N_33129,N_31562,N_31494);
nand U33130 (N_33130,N_31268,N_31483);
or U33131 (N_33131,N_30374,N_30986);
and U33132 (N_33132,N_31167,N_30487);
nor U33133 (N_33133,N_31953,N_31942);
nand U33134 (N_33134,N_30867,N_30637);
nand U33135 (N_33135,N_31605,N_31854);
nor U33136 (N_33136,N_30449,N_30516);
or U33137 (N_33137,N_31166,N_31858);
nand U33138 (N_33138,N_31114,N_30827);
or U33139 (N_33139,N_30257,N_31782);
and U33140 (N_33140,N_30183,N_30119);
or U33141 (N_33141,N_30490,N_31154);
and U33142 (N_33142,N_30132,N_30691);
nand U33143 (N_33143,N_30417,N_30789);
or U33144 (N_33144,N_30383,N_31602);
nand U33145 (N_33145,N_31297,N_30155);
nor U33146 (N_33146,N_31017,N_30878);
nor U33147 (N_33147,N_30258,N_31844);
or U33148 (N_33148,N_30389,N_31364);
or U33149 (N_33149,N_31411,N_30314);
or U33150 (N_33150,N_31594,N_31593);
or U33151 (N_33151,N_31195,N_30280);
nand U33152 (N_33152,N_31079,N_31893);
nand U33153 (N_33153,N_31124,N_30562);
and U33154 (N_33154,N_31623,N_31157);
nor U33155 (N_33155,N_30615,N_30843);
and U33156 (N_33156,N_31974,N_31025);
and U33157 (N_33157,N_31297,N_31834);
or U33158 (N_33158,N_31702,N_30034);
nand U33159 (N_33159,N_30806,N_31153);
and U33160 (N_33160,N_31515,N_31754);
nand U33161 (N_33161,N_31034,N_31626);
or U33162 (N_33162,N_30743,N_31356);
nor U33163 (N_33163,N_31623,N_30336);
or U33164 (N_33164,N_31318,N_31665);
and U33165 (N_33165,N_31008,N_31878);
xnor U33166 (N_33166,N_31908,N_31168);
and U33167 (N_33167,N_30861,N_31229);
nand U33168 (N_33168,N_31932,N_30819);
nand U33169 (N_33169,N_30224,N_31513);
and U33170 (N_33170,N_31086,N_30429);
and U33171 (N_33171,N_30259,N_30759);
and U33172 (N_33172,N_31478,N_31872);
nand U33173 (N_33173,N_31135,N_31855);
or U33174 (N_33174,N_30283,N_30783);
nor U33175 (N_33175,N_30192,N_31477);
nor U33176 (N_33176,N_30065,N_30389);
and U33177 (N_33177,N_31457,N_31393);
nor U33178 (N_33178,N_31004,N_30992);
nor U33179 (N_33179,N_30691,N_31688);
or U33180 (N_33180,N_30984,N_30291);
and U33181 (N_33181,N_30525,N_31605);
or U33182 (N_33182,N_31603,N_30524);
nor U33183 (N_33183,N_31985,N_30726);
nand U33184 (N_33184,N_30440,N_30250);
nor U33185 (N_33185,N_31557,N_31423);
or U33186 (N_33186,N_30712,N_31160);
and U33187 (N_33187,N_31787,N_30724);
or U33188 (N_33188,N_31973,N_30077);
or U33189 (N_33189,N_30228,N_31514);
and U33190 (N_33190,N_31032,N_31556);
nand U33191 (N_33191,N_31468,N_31245);
and U33192 (N_33192,N_30214,N_30202);
or U33193 (N_33193,N_31209,N_31792);
nand U33194 (N_33194,N_30394,N_31224);
or U33195 (N_33195,N_30730,N_30210);
or U33196 (N_33196,N_31369,N_30935);
nor U33197 (N_33197,N_31201,N_31884);
nand U33198 (N_33198,N_31848,N_30535);
xor U33199 (N_33199,N_30484,N_30322);
nand U33200 (N_33200,N_31813,N_30955);
and U33201 (N_33201,N_31231,N_30347);
and U33202 (N_33202,N_31405,N_31939);
nand U33203 (N_33203,N_31444,N_31416);
or U33204 (N_33204,N_30432,N_31823);
or U33205 (N_33205,N_31869,N_31580);
nor U33206 (N_33206,N_30220,N_31553);
nand U33207 (N_33207,N_31175,N_30524);
and U33208 (N_33208,N_30194,N_30157);
nand U33209 (N_33209,N_31196,N_30235);
and U33210 (N_33210,N_30426,N_30494);
or U33211 (N_33211,N_31161,N_30993);
and U33212 (N_33212,N_31133,N_30768);
or U33213 (N_33213,N_30224,N_31690);
nor U33214 (N_33214,N_30433,N_31186);
nor U33215 (N_33215,N_31996,N_30689);
nand U33216 (N_33216,N_31039,N_31603);
nor U33217 (N_33217,N_30761,N_31218);
nand U33218 (N_33218,N_31451,N_30276);
nor U33219 (N_33219,N_30558,N_30396);
and U33220 (N_33220,N_30578,N_31917);
and U33221 (N_33221,N_31848,N_30456);
nand U33222 (N_33222,N_31901,N_30455);
nand U33223 (N_33223,N_31176,N_30060);
and U33224 (N_33224,N_30988,N_30499);
nand U33225 (N_33225,N_30993,N_30707);
nor U33226 (N_33226,N_31501,N_31862);
and U33227 (N_33227,N_31471,N_30814);
nand U33228 (N_33228,N_30893,N_31862);
nand U33229 (N_33229,N_30821,N_31418);
or U33230 (N_33230,N_30289,N_30922);
or U33231 (N_33231,N_30737,N_30107);
nand U33232 (N_33232,N_31185,N_31941);
nand U33233 (N_33233,N_30239,N_30251);
nor U33234 (N_33234,N_31662,N_31202);
nand U33235 (N_33235,N_30574,N_30328);
or U33236 (N_33236,N_30779,N_30089);
and U33237 (N_33237,N_31511,N_30738);
and U33238 (N_33238,N_30702,N_31005);
nor U33239 (N_33239,N_30741,N_30267);
nand U33240 (N_33240,N_30373,N_31347);
xnor U33241 (N_33241,N_30455,N_31434);
nor U33242 (N_33242,N_31752,N_30384);
nor U33243 (N_33243,N_30950,N_31381);
nand U33244 (N_33244,N_30636,N_31962);
and U33245 (N_33245,N_31071,N_31481);
and U33246 (N_33246,N_30377,N_30319);
or U33247 (N_33247,N_30347,N_31720);
nand U33248 (N_33248,N_30733,N_30761);
nand U33249 (N_33249,N_31179,N_30514);
nor U33250 (N_33250,N_30896,N_31599);
nor U33251 (N_33251,N_31441,N_31966);
or U33252 (N_33252,N_30206,N_30218);
nor U33253 (N_33253,N_30820,N_30045);
and U33254 (N_33254,N_30879,N_30256);
or U33255 (N_33255,N_30460,N_30382);
xnor U33256 (N_33256,N_31379,N_30511);
and U33257 (N_33257,N_31584,N_31934);
nand U33258 (N_33258,N_30348,N_30176);
or U33259 (N_33259,N_31101,N_30573);
nand U33260 (N_33260,N_30625,N_30474);
nor U33261 (N_33261,N_30067,N_30069);
nand U33262 (N_33262,N_30201,N_30815);
nand U33263 (N_33263,N_30280,N_31398);
nor U33264 (N_33264,N_30149,N_30581);
nor U33265 (N_33265,N_31461,N_31874);
nand U33266 (N_33266,N_30473,N_30790);
nor U33267 (N_33267,N_31691,N_30344);
and U33268 (N_33268,N_31580,N_30015);
and U33269 (N_33269,N_31110,N_31437);
and U33270 (N_33270,N_30362,N_30536);
and U33271 (N_33271,N_30741,N_30997);
or U33272 (N_33272,N_30666,N_31191);
nor U33273 (N_33273,N_31910,N_30340);
or U33274 (N_33274,N_31539,N_31567);
nand U33275 (N_33275,N_31249,N_31688);
or U33276 (N_33276,N_30348,N_31947);
nand U33277 (N_33277,N_31024,N_31285);
and U33278 (N_33278,N_31169,N_31305);
or U33279 (N_33279,N_31231,N_30562);
nand U33280 (N_33280,N_31986,N_30169);
and U33281 (N_33281,N_31215,N_31554);
nor U33282 (N_33282,N_30750,N_30359);
and U33283 (N_33283,N_31467,N_31900);
or U33284 (N_33284,N_31780,N_31383);
nor U33285 (N_33285,N_31573,N_30820);
nor U33286 (N_33286,N_31271,N_31269);
nand U33287 (N_33287,N_30840,N_31887);
or U33288 (N_33288,N_31008,N_30993);
nand U33289 (N_33289,N_31039,N_31838);
nor U33290 (N_33290,N_30558,N_31887);
nand U33291 (N_33291,N_30284,N_30120);
nor U33292 (N_33292,N_31089,N_30961);
and U33293 (N_33293,N_30161,N_30986);
nor U33294 (N_33294,N_30204,N_31454);
and U33295 (N_33295,N_31670,N_30017);
or U33296 (N_33296,N_31530,N_30335);
and U33297 (N_33297,N_30412,N_31620);
or U33298 (N_33298,N_30006,N_30857);
nor U33299 (N_33299,N_31081,N_31953);
nand U33300 (N_33300,N_31748,N_31356);
and U33301 (N_33301,N_30396,N_31845);
nand U33302 (N_33302,N_30238,N_31104);
or U33303 (N_33303,N_30457,N_31004);
and U33304 (N_33304,N_30934,N_31606);
nor U33305 (N_33305,N_30321,N_31153);
xor U33306 (N_33306,N_30142,N_30161);
nor U33307 (N_33307,N_31345,N_31799);
and U33308 (N_33308,N_31038,N_30303);
nor U33309 (N_33309,N_30647,N_30749);
or U33310 (N_33310,N_30996,N_31588);
nand U33311 (N_33311,N_30782,N_31315);
nand U33312 (N_33312,N_31764,N_31272);
nand U33313 (N_33313,N_31214,N_31446);
or U33314 (N_33314,N_31329,N_30376);
nand U33315 (N_33315,N_31571,N_31936);
or U33316 (N_33316,N_30554,N_31980);
or U33317 (N_33317,N_31266,N_30789);
nor U33318 (N_33318,N_31333,N_30854);
nand U33319 (N_33319,N_31666,N_31996);
and U33320 (N_33320,N_31417,N_30940);
or U33321 (N_33321,N_30706,N_31354);
nand U33322 (N_33322,N_31857,N_31737);
or U33323 (N_33323,N_30439,N_30588);
nor U33324 (N_33324,N_31147,N_30498);
or U33325 (N_33325,N_31960,N_31847);
or U33326 (N_33326,N_30793,N_31509);
nor U33327 (N_33327,N_31680,N_31555);
nand U33328 (N_33328,N_31188,N_31902);
or U33329 (N_33329,N_31170,N_30277);
nand U33330 (N_33330,N_31504,N_30931);
nor U33331 (N_33331,N_30532,N_30937);
nor U33332 (N_33332,N_31362,N_30356);
nand U33333 (N_33333,N_30616,N_30217);
and U33334 (N_33334,N_30141,N_30592);
nand U33335 (N_33335,N_30793,N_30745);
or U33336 (N_33336,N_30186,N_31325);
nor U33337 (N_33337,N_30820,N_30870);
and U33338 (N_33338,N_31180,N_31794);
and U33339 (N_33339,N_31036,N_30649);
xnor U33340 (N_33340,N_31948,N_31204);
nor U33341 (N_33341,N_31594,N_30323);
and U33342 (N_33342,N_31005,N_30014);
nor U33343 (N_33343,N_30505,N_30219);
and U33344 (N_33344,N_30894,N_30837);
nor U33345 (N_33345,N_31322,N_30974);
and U33346 (N_33346,N_30133,N_31915);
or U33347 (N_33347,N_31514,N_30671);
nor U33348 (N_33348,N_31712,N_30242);
nor U33349 (N_33349,N_31615,N_31411);
and U33350 (N_33350,N_30109,N_30911);
or U33351 (N_33351,N_30788,N_30402);
nand U33352 (N_33352,N_31297,N_30938);
and U33353 (N_33353,N_30578,N_30582);
nor U33354 (N_33354,N_30786,N_31747);
or U33355 (N_33355,N_30674,N_30753);
and U33356 (N_33356,N_31458,N_30959);
and U33357 (N_33357,N_30413,N_30597);
and U33358 (N_33358,N_30800,N_30044);
nand U33359 (N_33359,N_30988,N_30936);
or U33360 (N_33360,N_31019,N_30204);
nor U33361 (N_33361,N_30203,N_31327);
and U33362 (N_33362,N_30127,N_30012);
nor U33363 (N_33363,N_31933,N_31249);
nand U33364 (N_33364,N_31536,N_30137);
and U33365 (N_33365,N_30303,N_30809);
or U33366 (N_33366,N_31919,N_31398);
or U33367 (N_33367,N_31154,N_30606);
and U33368 (N_33368,N_30757,N_30818);
nand U33369 (N_33369,N_31898,N_31510);
and U33370 (N_33370,N_31334,N_30823);
nor U33371 (N_33371,N_30971,N_30346);
and U33372 (N_33372,N_30927,N_31472);
nand U33373 (N_33373,N_31040,N_31938);
or U33374 (N_33374,N_30067,N_31533);
or U33375 (N_33375,N_30792,N_31386);
nand U33376 (N_33376,N_30776,N_30182);
and U33377 (N_33377,N_30324,N_31067);
or U33378 (N_33378,N_30161,N_31864);
and U33379 (N_33379,N_30071,N_30262);
or U33380 (N_33380,N_31281,N_31871);
nor U33381 (N_33381,N_30586,N_30059);
and U33382 (N_33382,N_30276,N_31886);
and U33383 (N_33383,N_31922,N_31568);
nand U33384 (N_33384,N_31555,N_30329);
and U33385 (N_33385,N_30146,N_30077);
xor U33386 (N_33386,N_31043,N_30868);
nor U33387 (N_33387,N_30373,N_30010);
nor U33388 (N_33388,N_30942,N_31961);
and U33389 (N_33389,N_30444,N_30485);
nor U33390 (N_33390,N_31970,N_30593);
or U33391 (N_33391,N_30905,N_30164);
nor U33392 (N_33392,N_30682,N_30881);
xor U33393 (N_33393,N_30618,N_31383);
and U33394 (N_33394,N_30370,N_30711);
or U33395 (N_33395,N_30753,N_31373);
nand U33396 (N_33396,N_30236,N_31772);
or U33397 (N_33397,N_31247,N_31754);
nor U33398 (N_33398,N_30391,N_31419);
or U33399 (N_33399,N_30229,N_31666);
nand U33400 (N_33400,N_31048,N_31061);
or U33401 (N_33401,N_30879,N_31119);
nor U33402 (N_33402,N_30493,N_31085);
nand U33403 (N_33403,N_31283,N_31487);
nand U33404 (N_33404,N_31226,N_30793);
or U33405 (N_33405,N_31612,N_30104);
and U33406 (N_33406,N_30920,N_31768);
xnor U33407 (N_33407,N_30356,N_30131);
and U33408 (N_33408,N_31330,N_30591);
and U33409 (N_33409,N_30090,N_31286);
and U33410 (N_33410,N_30794,N_30328);
nand U33411 (N_33411,N_31693,N_31909);
nand U33412 (N_33412,N_31773,N_30020);
or U33413 (N_33413,N_31462,N_30039);
nand U33414 (N_33414,N_31492,N_31536);
and U33415 (N_33415,N_31565,N_31170);
nor U33416 (N_33416,N_31562,N_30694);
or U33417 (N_33417,N_30838,N_30074);
nand U33418 (N_33418,N_30454,N_30691);
nor U33419 (N_33419,N_30844,N_31155);
nand U33420 (N_33420,N_31792,N_31528);
and U33421 (N_33421,N_31830,N_30706);
nand U33422 (N_33422,N_30044,N_31557);
nor U33423 (N_33423,N_31501,N_31442);
or U33424 (N_33424,N_30103,N_31834);
and U33425 (N_33425,N_30599,N_31019);
nand U33426 (N_33426,N_31643,N_30335);
xor U33427 (N_33427,N_31170,N_31793);
nor U33428 (N_33428,N_30101,N_31836);
nand U33429 (N_33429,N_31318,N_31936);
and U33430 (N_33430,N_30442,N_30902);
and U33431 (N_33431,N_30982,N_31148);
xor U33432 (N_33432,N_30128,N_30632);
xnor U33433 (N_33433,N_30388,N_30844);
nor U33434 (N_33434,N_31775,N_30664);
nor U33435 (N_33435,N_31848,N_30575);
or U33436 (N_33436,N_31190,N_30570);
nor U33437 (N_33437,N_31877,N_31394);
nand U33438 (N_33438,N_30488,N_31050);
or U33439 (N_33439,N_31856,N_31030);
and U33440 (N_33440,N_30661,N_30536);
or U33441 (N_33441,N_30725,N_30025);
or U33442 (N_33442,N_30809,N_30633);
or U33443 (N_33443,N_30870,N_30547);
and U33444 (N_33444,N_30486,N_30466);
nor U33445 (N_33445,N_31194,N_31228);
or U33446 (N_33446,N_31202,N_30514);
nand U33447 (N_33447,N_30107,N_30209);
nor U33448 (N_33448,N_30540,N_31204);
or U33449 (N_33449,N_31906,N_31156);
and U33450 (N_33450,N_30391,N_30533);
nand U33451 (N_33451,N_31242,N_31644);
and U33452 (N_33452,N_30862,N_30793);
nand U33453 (N_33453,N_31859,N_31049);
nand U33454 (N_33454,N_30118,N_30374);
nand U33455 (N_33455,N_30151,N_30141);
nand U33456 (N_33456,N_31959,N_31169);
or U33457 (N_33457,N_30749,N_31272);
nand U33458 (N_33458,N_31825,N_30306);
nor U33459 (N_33459,N_30187,N_30123);
or U33460 (N_33460,N_31361,N_30310);
nor U33461 (N_33461,N_31956,N_31896);
and U33462 (N_33462,N_30143,N_31804);
nand U33463 (N_33463,N_30123,N_31068);
nor U33464 (N_33464,N_31139,N_31024);
or U33465 (N_33465,N_31238,N_30366);
and U33466 (N_33466,N_31182,N_31569);
and U33467 (N_33467,N_31970,N_30561);
and U33468 (N_33468,N_30013,N_30724);
nor U33469 (N_33469,N_31826,N_30518);
nand U33470 (N_33470,N_31058,N_30242);
or U33471 (N_33471,N_30258,N_31524);
nand U33472 (N_33472,N_30088,N_31009);
and U33473 (N_33473,N_31188,N_30134);
or U33474 (N_33474,N_30744,N_31586);
nor U33475 (N_33475,N_31443,N_31184);
or U33476 (N_33476,N_31672,N_30305);
nand U33477 (N_33477,N_31342,N_30641);
or U33478 (N_33478,N_31081,N_31630);
nand U33479 (N_33479,N_31754,N_30708);
or U33480 (N_33480,N_30836,N_30463);
nand U33481 (N_33481,N_31596,N_30479);
nor U33482 (N_33482,N_31274,N_30492);
nor U33483 (N_33483,N_31506,N_30241);
or U33484 (N_33484,N_30897,N_31211);
and U33485 (N_33485,N_30890,N_31114);
and U33486 (N_33486,N_30663,N_31136);
nor U33487 (N_33487,N_30746,N_30326);
nor U33488 (N_33488,N_31122,N_31651);
nor U33489 (N_33489,N_31289,N_31929);
and U33490 (N_33490,N_31753,N_31615);
nor U33491 (N_33491,N_31992,N_31408);
nor U33492 (N_33492,N_31885,N_31049);
or U33493 (N_33493,N_30751,N_31932);
nand U33494 (N_33494,N_30618,N_30810);
nor U33495 (N_33495,N_31471,N_31395);
and U33496 (N_33496,N_30861,N_30596);
nor U33497 (N_33497,N_30837,N_30380);
or U33498 (N_33498,N_31490,N_31128);
and U33499 (N_33499,N_31436,N_31925);
nor U33500 (N_33500,N_31088,N_30823);
or U33501 (N_33501,N_31684,N_30887);
and U33502 (N_33502,N_31447,N_31314);
or U33503 (N_33503,N_31595,N_30892);
nor U33504 (N_33504,N_31948,N_31750);
nand U33505 (N_33505,N_31792,N_30130);
nor U33506 (N_33506,N_30638,N_31348);
nor U33507 (N_33507,N_30464,N_30606);
nand U33508 (N_33508,N_30600,N_30560);
or U33509 (N_33509,N_31129,N_30932);
and U33510 (N_33510,N_30022,N_30954);
and U33511 (N_33511,N_30901,N_30424);
or U33512 (N_33512,N_31962,N_30310);
and U33513 (N_33513,N_31484,N_30500);
xor U33514 (N_33514,N_31899,N_31296);
and U33515 (N_33515,N_31541,N_30773);
and U33516 (N_33516,N_30425,N_31881);
nand U33517 (N_33517,N_30153,N_30363);
nand U33518 (N_33518,N_30908,N_31402);
nor U33519 (N_33519,N_30770,N_30577);
nand U33520 (N_33520,N_31023,N_30149);
or U33521 (N_33521,N_31900,N_31019);
or U33522 (N_33522,N_30564,N_30562);
nor U33523 (N_33523,N_31856,N_31315);
or U33524 (N_33524,N_31661,N_30584);
nand U33525 (N_33525,N_31935,N_30053);
nand U33526 (N_33526,N_30128,N_30705);
and U33527 (N_33527,N_31512,N_31908);
nand U33528 (N_33528,N_31209,N_30873);
or U33529 (N_33529,N_30688,N_30403);
nand U33530 (N_33530,N_31295,N_30618);
or U33531 (N_33531,N_31962,N_30749);
nor U33532 (N_33532,N_30096,N_30188);
or U33533 (N_33533,N_31749,N_31833);
or U33534 (N_33534,N_30754,N_30317);
xor U33535 (N_33535,N_31221,N_30166);
or U33536 (N_33536,N_31962,N_30485);
and U33537 (N_33537,N_30003,N_31001);
nor U33538 (N_33538,N_30382,N_31657);
nor U33539 (N_33539,N_30954,N_30561);
and U33540 (N_33540,N_30448,N_30597);
or U33541 (N_33541,N_31723,N_30993);
and U33542 (N_33542,N_31020,N_30632);
nor U33543 (N_33543,N_31361,N_31671);
and U33544 (N_33544,N_30882,N_31985);
nor U33545 (N_33545,N_31545,N_31842);
and U33546 (N_33546,N_31330,N_31698);
nand U33547 (N_33547,N_31517,N_31494);
nand U33548 (N_33548,N_31783,N_31213);
nand U33549 (N_33549,N_30007,N_30125);
xor U33550 (N_33550,N_31540,N_31264);
nand U33551 (N_33551,N_30299,N_31536);
and U33552 (N_33552,N_31761,N_30047);
and U33553 (N_33553,N_31335,N_30153);
nor U33554 (N_33554,N_31979,N_31822);
and U33555 (N_33555,N_30472,N_31799);
nor U33556 (N_33556,N_31085,N_30539);
nand U33557 (N_33557,N_30825,N_30681);
or U33558 (N_33558,N_30859,N_31635);
nand U33559 (N_33559,N_31510,N_30217);
nor U33560 (N_33560,N_31388,N_30646);
nand U33561 (N_33561,N_31698,N_30075);
nor U33562 (N_33562,N_30974,N_30845);
and U33563 (N_33563,N_30005,N_31269);
nor U33564 (N_33564,N_31796,N_31611);
nor U33565 (N_33565,N_31246,N_30026);
and U33566 (N_33566,N_30223,N_31430);
or U33567 (N_33567,N_30682,N_31681);
or U33568 (N_33568,N_30318,N_31363);
or U33569 (N_33569,N_30999,N_31012);
and U33570 (N_33570,N_30884,N_30112);
nor U33571 (N_33571,N_31168,N_31495);
nor U33572 (N_33572,N_30748,N_30087);
nor U33573 (N_33573,N_30167,N_31611);
or U33574 (N_33574,N_31038,N_31007);
and U33575 (N_33575,N_31343,N_30160);
nand U33576 (N_33576,N_31888,N_30671);
nand U33577 (N_33577,N_31895,N_30326);
nor U33578 (N_33578,N_30143,N_30121);
or U33579 (N_33579,N_31388,N_31418);
or U33580 (N_33580,N_31144,N_31373);
or U33581 (N_33581,N_31608,N_31377);
nand U33582 (N_33582,N_31170,N_31784);
nand U33583 (N_33583,N_30468,N_30771);
and U33584 (N_33584,N_30320,N_31868);
nor U33585 (N_33585,N_30221,N_30500);
nand U33586 (N_33586,N_31632,N_31930);
or U33587 (N_33587,N_30873,N_30801);
xor U33588 (N_33588,N_30887,N_30789);
or U33589 (N_33589,N_31685,N_30329);
or U33590 (N_33590,N_31740,N_31317);
nor U33591 (N_33591,N_31362,N_30236);
or U33592 (N_33592,N_30044,N_31244);
and U33593 (N_33593,N_30576,N_30476);
or U33594 (N_33594,N_30610,N_30157);
or U33595 (N_33595,N_30298,N_31532);
nor U33596 (N_33596,N_30086,N_31749);
and U33597 (N_33597,N_30293,N_31405);
nand U33598 (N_33598,N_31222,N_30533);
xnor U33599 (N_33599,N_31693,N_31191);
and U33600 (N_33600,N_30371,N_31593);
nor U33601 (N_33601,N_30525,N_31335);
or U33602 (N_33602,N_31850,N_30481);
and U33603 (N_33603,N_31742,N_31635);
nor U33604 (N_33604,N_31984,N_31658);
nor U33605 (N_33605,N_30115,N_31136);
or U33606 (N_33606,N_31583,N_31055);
and U33607 (N_33607,N_30245,N_31932);
and U33608 (N_33608,N_30223,N_30537);
or U33609 (N_33609,N_31144,N_30222);
nor U33610 (N_33610,N_31095,N_31810);
or U33611 (N_33611,N_30009,N_31021);
and U33612 (N_33612,N_30712,N_30309);
nand U33613 (N_33613,N_31262,N_31935);
and U33614 (N_33614,N_31229,N_31811);
and U33615 (N_33615,N_30803,N_31597);
or U33616 (N_33616,N_30577,N_30965);
nor U33617 (N_33617,N_30465,N_31237);
nand U33618 (N_33618,N_31411,N_31100);
nand U33619 (N_33619,N_31041,N_31988);
nand U33620 (N_33620,N_30397,N_30217);
and U33621 (N_33621,N_30468,N_31476);
xnor U33622 (N_33622,N_30764,N_30937);
and U33623 (N_33623,N_30292,N_30740);
and U33624 (N_33624,N_31821,N_30489);
or U33625 (N_33625,N_31167,N_30604);
nand U33626 (N_33626,N_30766,N_31950);
nor U33627 (N_33627,N_30498,N_31632);
nand U33628 (N_33628,N_30190,N_30887);
nand U33629 (N_33629,N_30101,N_31590);
nor U33630 (N_33630,N_30312,N_30442);
xnor U33631 (N_33631,N_31667,N_30631);
xnor U33632 (N_33632,N_30941,N_31926);
nor U33633 (N_33633,N_30684,N_30932);
and U33634 (N_33634,N_31704,N_30863);
and U33635 (N_33635,N_30062,N_31741);
nor U33636 (N_33636,N_31126,N_31893);
nand U33637 (N_33637,N_30979,N_30312);
nor U33638 (N_33638,N_31759,N_30417);
or U33639 (N_33639,N_30400,N_31541);
nor U33640 (N_33640,N_30013,N_31280);
or U33641 (N_33641,N_31383,N_30810);
and U33642 (N_33642,N_30770,N_30482);
and U33643 (N_33643,N_30047,N_31287);
nor U33644 (N_33644,N_31405,N_30169);
nor U33645 (N_33645,N_31919,N_31364);
nor U33646 (N_33646,N_31927,N_31304);
nand U33647 (N_33647,N_31312,N_31326);
nand U33648 (N_33648,N_31964,N_30503);
nor U33649 (N_33649,N_31422,N_30085);
and U33650 (N_33650,N_30740,N_31941);
or U33651 (N_33651,N_30253,N_30778);
and U33652 (N_33652,N_31071,N_30715);
or U33653 (N_33653,N_30829,N_31375);
xor U33654 (N_33654,N_31453,N_31822);
nor U33655 (N_33655,N_30469,N_31610);
and U33656 (N_33656,N_31797,N_30702);
nor U33657 (N_33657,N_30215,N_30241);
or U33658 (N_33658,N_30272,N_30628);
nand U33659 (N_33659,N_31876,N_30823);
and U33660 (N_33660,N_30873,N_30483);
or U33661 (N_33661,N_31185,N_30596);
or U33662 (N_33662,N_30681,N_30863);
nand U33663 (N_33663,N_30248,N_31919);
nand U33664 (N_33664,N_30038,N_30702);
and U33665 (N_33665,N_31207,N_31104);
nor U33666 (N_33666,N_31655,N_31290);
nor U33667 (N_33667,N_31947,N_31819);
and U33668 (N_33668,N_30794,N_31727);
or U33669 (N_33669,N_30673,N_31781);
and U33670 (N_33670,N_31253,N_30305);
nor U33671 (N_33671,N_30000,N_30670);
nand U33672 (N_33672,N_30877,N_31528);
nor U33673 (N_33673,N_30454,N_30953);
nand U33674 (N_33674,N_30505,N_30545);
and U33675 (N_33675,N_30318,N_30776);
xor U33676 (N_33676,N_31437,N_30352);
nand U33677 (N_33677,N_30163,N_31028);
and U33678 (N_33678,N_31924,N_30323);
nand U33679 (N_33679,N_30553,N_30061);
nor U33680 (N_33680,N_31862,N_30827);
or U33681 (N_33681,N_30896,N_30070);
nand U33682 (N_33682,N_30711,N_31799);
and U33683 (N_33683,N_30279,N_31093);
or U33684 (N_33684,N_30287,N_30174);
and U33685 (N_33685,N_30590,N_31864);
and U33686 (N_33686,N_30299,N_31151);
and U33687 (N_33687,N_30768,N_30332);
nor U33688 (N_33688,N_30588,N_31003);
or U33689 (N_33689,N_30238,N_31311);
or U33690 (N_33690,N_31422,N_30723);
and U33691 (N_33691,N_30298,N_30595);
nor U33692 (N_33692,N_30281,N_31526);
nor U33693 (N_33693,N_31633,N_30114);
or U33694 (N_33694,N_30553,N_31116);
nand U33695 (N_33695,N_30590,N_31007);
and U33696 (N_33696,N_30693,N_31740);
nand U33697 (N_33697,N_31761,N_31647);
or U33698 (N_33698,N_31682,N_30604);
nor U33699 (N_33699,N_31420,N_31819);
nand U33700 (N_33700,N_30083,N_31342);
or U33701 (N_33701,N_31227,N_30996);
and U33702 (N_33702,N_30397,N_31822);
nor U33703 (N_33703,N_30513,N_31363);
nor U33704 (N_33704,N_31203,N_31651);
and U33705 (N_33705,N_30973,N_31236);
and U33706 (N_33706,N_30528,N_31194);
and U33707 (N_33707,N_31171,N_31182);
xor U33708 (N_33708,N_31312,N_31931);
or U33709 (N_33709,N_31068,N_31335);
nand U33710 (N_33710,N_31275,N_31695);
and U33711 (N_33711,N_30364,N_30436);
or U33712 (N_33712,N_31173,N_30300);
nand U33713 (N_33713,N_31385,N_31620);
nand U33714 (N_33714,N_31367,N_30384);
and U33715 (N_33715,N_31636,N_31036);
or U33716 (N_33716,N_30185,N_31448);
or U33717 (N_33717,N_31214,N_31036);
and U33718 (N_33718,N_30498,N_30078);
and U33719 (N_33719,N_31611,N_30191);
or U33720 (N_33720,N_30616,N_30483);
and U33721 (N_33721,N_30004,N_31574);
or U33722 (N_33722,N_31490,N_31664);
and U33723 (N_33723,N_30768,N_31323);
or U33724 (N_33724,N_30772,N_31476);
or U33725 (N_33725,N_30660,N_31929);
nand U33726 (N_33726,N_31673,N_31094);
and U33727 (N_33727,N_30931,N_31834);
nor U33728 (N_33728,N_30397,N_31174);
nand U33729 (N_33729,N_30889,N_30515);
or U33730 (N_33730,N_31441,N_31001);
and U33731 (N_33731,N_30908,N_30977);
xnor U33732 (N_33732,N_31975,N_31481);
and U33733 (N_33733,N_31320,N_30590);
nand U33734 (N_33734,N_30162,N_30612);
nor U33735 (N_33735,N_31961,N_30432);
xor U33736 (N_33736,N_30641,N_30176);
or U33737 (N_33737,N_30474,N_30644);
nand U33738 (N_33738,N_30694,N_30288);
and U33739 (N_33739,N_31106,N_30472);
nor U33740 (N_33740,N_30253,N_31653);
nand U33741 (N_33741,N_31459,N_30843);
nand U33742 (N_33742,N_30079,N_30913);
xor U33743 (N_33743,N_30754,N_30514);
nand U33744 (N_33744,N_31358,N_31993);
nor U33745 (N_33745,N_31428,N_30142);
and U33746 (N_33746,N_30100,N_31813);
or U33747 (N_33747,N_30371,N_30911);
and U33748 (N_33748,N_30317,N_30689);
nand U33749 (N_33749,N_31933,N_30268);
nand U33750 (N_33750,N_31605,N_30197);
nor U33751 (N_33751,N_30857,N_30774);
nor U33752 (N_33752,N_31226,N_31559);
and U33753 (N_33753,N_31294,N_30354);
and U33754 (N_33754,N_30210,N_31428);
or U33755 (N_33755,N_31660,N_30726);
nand U33756 (N_33756,N_31763,N_31312);
nand U33757 (N_33757,N_30815,N_30990);
xor U33758 (N_33758,N_30828,N_30289);
and U33759 (N_33759,N_30990,N_30923);
or U33760 (N_33760,N_30256,N_31823);
or U33761 (N_33761,N_31304,N_30856);
xnor U33762 (N_33762,N_31769,N_31212);
and U33763 (N_33763,N_30568,N_30897);
nor U33764 (N_33764,N_31238,N_31336);
nand U33765 (N_33765,N_31174,N_31499);
xnor U33766 (N_33766,N_31991,N_30239);
nor U33767 (N_33767,N_31133,N_30694);
and U33768 (N_33768,N_31561,N_31349);
and U33769 (N_33769,N_31438,N_30305);
and U33770 (N_33770,N_30325,N_30624);
or U33771 (N_33771,N_31209,N_30334);
and U33772 (N_33772,N_30492,N_31439);
or U33773 (N_33773,N_30630,N_31483);
or U33774 (N_33774,N_30195,N_31894);
nor U33775 (N_33775,N_30523,N_30845);
nand U33776 (N_33776,N_30466,N_30456);
and U33777 (N_33777,N_31196,N_31257);
xnor U33778 (N_33778,N_30139,N_30679);
nand U33779 (N_33779,N_31729,N_31071);
or U33780 (N_33780,N_31672,N_30288);
nand U33781 (N_33781,N_31577,N_30301);
nor U33782 (N_33782,N_30562,N_31476);
nand U33783 (N_33783,N_30981,N_31121);
nand U33784 (N_33784,N_30681,N_31731);
nor U33785 (N_33785,N_30298,N_30264);
and U33786 (N_33786,N_31326,N_30427);
and U33787 (N_33787,N_31320,N_31429);
nor U33788 (N_33788,N_31370,N_31747);
and U33789 (N_33789,N_31016,N_31407);
and U33790 (N_33790,N_31261,N_31289);
or U33791 (N_33791,N_30974,N_31739);
or U33792 (N_33792,N_30001,N_31427);
and U33793 (N_33793,N_30842,N_30988);
nor U33794 (N_33794,N_30506,N_30454);
xnor U33795 (N_33795,N_30140,N_31206);
nor U33796 (N_33796,N_30267,N_30998);
and U33797 (N_33797,N_30876,N_31030);
or U33798 (N_33798,N_31533,N_31472);
nand U33799 (N_33799,N_31241,N_31423);
nor U33800 (N_33800,N_30611,N_30864);
nor U33801 (N_33801,N_31925,N_31452);
and U33802 (N_33802,N_31203,N_30040);
nand U33803 (N_33803,N_30285,N_30886);
and U33804 (N_33804,N_31755,N_31179);
nor U33805 (N_33805,N_31680,N_31979);
and U33806 (N_33806,N_30264,N_30287);
and U33807 (N_33807,N_30559,N_31089);
nand U33808 (N_33808,N_30588,N_30905);
nand U33809 (N_33809,N_30042,N_31102);
or U33810 (N_33810,N_30838,N_31948);
and U33811 (N_33811,N_30737,N_31648);
nor U33812 (N_33812,N_30164,N_31792);
and U33813 (N_33813,N_30386,N_30748);
nor U33814 (N_33814,N_31328,N_31432);
nor U33815 (N_33815,N_31521,N_30842);
or U33816 (N_33816,N_31197,N_30411);
nand U33817 (N_33817,N_31315,N_31309);
nand U33818 (N_33818,N_31056,N_31131);
nand U33819 (N_33819,N_30899,N_30972);
nor U33820 (N_33820,N_30610,N_31702);
or U33821 (N_33821,N_30761,N_30714);
and U33822 (N_33822,N_31852,N_31909);
nor U33823 (N_33823,N_31383,N_31815);
nand U33824 (N_33824,N_31686,N_31401);
and U33825 (N_33825,N_30393,N_30830);
or U33826 (N_33826,N_30529,N_30073);
or U33827 (N_33827,N_30375,N_31373);
and U33828 (N_33828,N_31236,N_30659);
nor U33829 (N_33829,N_30112,N_31744);
or U33830 (N_33830,N_31897,N_31817);
or U33831 (N_33831,N_31600,N_30021);
and U33832 (N_33832,N_30815,N_30443);
or U33833 (N_33833,N_31491,N_30657);
nand U33834 (N_33834,N_30696,N_30416);
nand U33835 (N_33835,N_31560,N_30521);
nor U33836 (N_33836,N_30016,N_30717);
nor U33837 (N_33837,N_31670,N_30948);
or U33838 (N_33838,N_31030,N_31849);
and U33839 (N_33839,N_31076,N_31574);
or U33840 (N_33840,N_31263,N_31134);
nor U33841 (N_33841,N_30492,N_31845);
nor U33842 (N_33842,N_31847,N_31870);
nor U33843 (N_33843,N_31809,N_31093);
or U33844 (N_33844,N_31000,N_30672);
and U33845 (N_33845,N_31412,N_31038);
or U33846 (N_33846,N_31493,N_30196);
nand U33847 (N_33847,N_31064,N_30816);
or U33848 (N_33848,N_30090,N_30541);
xnor U33849 (N_33849,N_31477,N_30421);
or U33850 (N_33850,N_30516,N_30790);
or U33851 (N_33851,N_31108,N_31669);
nand U33852 (N_33852,N_31152,N_30129);
nand U33853 (N_33853,N_30600,N_30033);
xor U33854 (N_33854,N_31885,N_30169);
nand U33855 (N_33855,N_30705,N_31997);
or U33856 (N_33856,N_31669,N_31737);
nand U33857 (N_33857,N_30425,N_31933);
nor U33858 (N_33858,N_31816,N_31583);
nand U33859 (N_33859,N_30926,N_30964);
xor U33860 (N_33860,N_31447,N_30989);
and U33861 (N_33861,N_31744,N_30033);
nand U33862 (N_33862,N_31392,N_31909);
or U33863 (N_33863,N_30790,N_30041);
or U33864 (N_33864,N_31211,N_30354);
or U33865 (N_33865,N_30817,N_31500);
nand U33866 (N_33866,N_31418,N_31366);
nand U33867 (N_33867,N_30008,N_31763);
and U33868 (N_33868,N_31758,N_30747);
or U33869 (N_33869,N_30960,N_31152);
or U33870 (N_33870,N_30385,N_31348);
and U33871 (N_33871,N_31217,N_30219);
or U33872 (N_33872,N_30029,N_31117);
and U33873 (N_33873,N_31363,N_30621);
nor U33874 (N_33874,N_30328,N_31861);
nor U33875 (N_33875,N_30767,N_31707);
or U33876 (N_33876,N_31795,N_31150);
or U33877 (N_33877,N_30730,N_30054);
nor U33878 (N_33878,N_30856,N_30084);
nor U33879 (N_33879,N_31461,N_30585);
and U33880 (N_33880,N_30960,N_31772);
nand U33881 (N_33881,N_30288,N_30917);
nand U33882 (N_33882,N_30793,N_31932);
or U33883 (N_33883,N_30715,N_30426);
and U33884 (N_33884,N_31450,N_30893);
nor U33885 (N_33885,N_31410,N_31392);
nand U33886 (N_33886,N_31616,N_30988);
nor U33887 (N_33887,N_30007,N_30118);
nor U33888 (N_33888,N_31042,N_30940);
nand U33889 (N_33889,N_30877,N_31323);
or U33890 (N_33890,N_30595,N_31385);
or U33891 (N_33891,N_31554,N_31287);
and U33892 (N_33892,N_30915,N_31014);
nor U33893 (N_33893,N_31014,N_30500);
and U33894 (N_33894,N_31202,N_31433);
nor U33895 (N_33895,N_30007,N_31557);
nand U33896 (N_33896,N_31063,N_30350);
nand U33897 (N_33897,N_31910,N_31173);
nor U33898 (N_33898,N_31909,N_31496);
or U33899 (N_33899,N_30570,N_31448);
nand U33900 (N_33900,N_30257,N_30377);
xnor U33901 (N_33901,N_31323,N_30709);
and U33902 (N_33902,N_30753,N_31354);
nor U33903 (N_33903,N_31180,N_30837);
nor U33904 (N_33904,N_30071,N_31400);
or U33905 (N_33905,N_31344,N_31670);
or U33906 (N_33906,N_30233,N_31720);
nor U33907 (N_33907,N_30010,N_31698);
or U33908 (N_33908,N_30665,N_30554);
nand U33909 (N_33909,N_31884,N_31470);
and U33910 (N_33910,N_31990,N_31310);
or U33911 (N_33911,N_31303,N_31464);
and U33912 (N_33912,N_31465,N_30840);
and U33913 (N_33913,N_31617,N_30954);
nor U33914 (N_33914,N_30289,N_30619);
nor U33915 (N_33915,N_31860,N_31538);
or U33916 (N_33916,N_31336,N_30148);
nor U33917 (N_33917,N_30349,N_31818);
or U33918 (N_33918,N_30938,N_31436);
nor U33919 (N_33919,N_30452,N_30783);
or U33920 (N_33920,N_30582,N_30940);
and U33921 (N_33921,N_30942,N_31351);
or U33922 (N_33922,N_30533,N_31539);
nor U33923 (N_33923,N_30003,N_31192);
nor U33924 (N_33924,N_31293,N_30120);
nor U33925 (N_33925,N_30345,N_31497);
nand U33926 (N_33926,N_31859,N_30213);
nor U33927 (N_33927,N_31126,N_31233);
nor U33928 (N_33928,N_30530,N_30716);
or U33929 (N_33929,N_31177,N_30302);
or U33930 (N_33930,N_31429,N_31598);
nor U33931 (N_33931,N_31153,N_30645);
or U33932 (N_33932,N_30391,N_31831);
nand U33933 (N_33933,N_30582,N_31890);
nor U33934 (N_33934,N_30984,N_30187);
nor U33935 (N_33935,N_31718,N_31284);
and U33936 (N_33936,N_30936,N_30722);
nand U33937 (N_33937,N_30695,N_31843);
nor U33938 (N_33938,N_31819,N_30981);
and U33939 (N_33939,N_30535,N_31949);
nor U33940 (N_33940,N_31503,N_30226);
and U33941 (N_33941,N_31995,N_30339);
nand U33942 (N_33942,N_30077,N_30838);
nand U33943 (N_33943,N_30704,N_30641);
and U33944 (N_33944,N_31501,N_31950);
nor U33945 (N_33945,N_31466,N_31555);
nand U33946 (N_33946,N_30934,N_30659);
and U33947 (N_33947,N_31563,N_31538);
nor U33948 (N_33948,N_31072,N_31125);
nand U33949 (N_33949,N_31884,N_31063);
nand U33950 (N_33950,N_31320,N_31508);
nand U33951 (N_33951,N_31197,N_30747);
or U33952 (N_33952,N_30277,N_30077);
and U33953 (N_33953,N_30219,N_30650);
and U33954 (N_33954,N_30266,N_30966);
nand U33955 (N_33955,N_30155,N_31350);
nand U33956 (N_33956,N_30062,N_31513);
and U33957 (N_33957,N_31020,N_31060);
nand U33958 (N_33958,N_31003,N_31597);
and U33959 (N_33959,N_30150,N_31067);
or U33960 (N_33960,N_30190,N_30134);
nand U33961 (N_33961,N_31591,N_30272);
nand U33962 (N_33962,N_30497,N_30590);
and U33963 (N_33963,N_30706,N_31165);
nor U33964 (N_33964,N_30333,N_30340);
and U33965 (N_33965,N_30120,N_30704);
nor U33966 (N_33966,N_31543,N_30902);
or U33967 (N_33967,N_30324,N_30525);
and U33968 (N_33968,N_31693,N_30216);
nor U33969 (N_33969,N_31716,N_31148);
nand U33970 (N_33970,N_30032,N_30998);
and U33971 (N_33971,N_30326,N_31708);
or U33972 (N_33972,N_30208,N_30950);
nand U33973 (N_33973,N_31405,N_30017);
or U33974 (N_33974,N_31004,N_30446);
and U33975 (N_33975,N_30374,N_30394);
or U33976 (N_33976,N_31356,N_30339);
nand U33977 (N_33977,N_31281,N_31658);
nand U33978 (N_33978,N_31077,N_31136);
nor U33979 (N_33979,N_30596,N_31056);
xnor U33980 (N_33980,N_31946,N_30488);
nor U33981 (N_33981,N_30991,N_31866);
nand U33982 (N_33982,N_31364,N_31901);
and U33983 (N_33983,N_31394,N_31701);
and U33984 (N_33984,N_30444,N_30122);
nor U33985 (N_33985,N_30241,N_31608);
and U33986 (N_33986,N_30626,N_31383);
nor U33987 (N_33987,N_30189,N_31788);
and U33988 (N_33988,N_30167,N_31877);
nand U33989 (N_33989,N_31310,N_31987);
nand U33990 (N_33990,N_31178,N_31469);
nand U33991 (N_33991,N_30739,N_31057);
or U33992 (N_33992,N_30620,N_30430);
nand U33993 (N_33993,N_30654,N_30226);
nor U33994 (N_33994,N_30931,N_31869);
and U33995 (N_33995,N_30790,N_30997);
or U33996 (N_33996,N_31960,N_31449);
nor U33997 (N_33997,N_30532,N_31223);
nand U33998 (N_33998,N_31689,N_30027);
xor U33999 (N_33999,N_30329,N_31352);
nor U34000 (N_34000,N_32962,N_33478);
and U34001 (N_34001,N_32943,N_33029);
nand U34002 (N_34002,N_33916,N_33419);
and U34003 (N_34003,N_33206,N_32610);
nand U34004 (N_34004,N_33943,N_32029);
and U34005 (N_34005,N_33630,N_33593);
and U34006 (N_34006,N_32115,N_32879);
and U34007 (N_34007,N_32614,N_33234);
and U34008 (N_34008,N_33071,N_32197);
and U34009 (N_34009,N_32308,N_32790);
nand U34010 (N_34010,N_33114,N_33077);
nor U34011 (N_34011,N_32726,N_33698);
and U34012 (N_34012,N_33113,N_32904);
nand U34013 (N_34013,N_32353,N_32512);
or U34014 (N_34014,N_32472,N_33070);
nand U34015 (N_34015,N_33879,N_32698);
nand U34016 (N_34016,N_33209,N_33675);
or U34017 (N_34017,N_33885,N_33602);
nand U34018 (N_34018,N_33066,N_33826);
or U34019 (N_34019,N_33899,N_32084);
nand U34020 (N_34020,N_32156,N_33064);
nor U34021 (N_34021,N_32997,N_32289);
nand U34022 (N_34022,N_33535,N_33996);
nand U34023 (N_34023,N_33597,N_32442);
nand U34024 (N_34024,N_33846,N_32560);
or U34025 (N_34025,N_33398,N_32880);
or U34026 (N_34026,N_33200,N_32515);
and U34027 (N_34027,N_32963,N_32361);
nor U34028 (N_34028,N_32404,N_32129);
and U34029 (N_34029,N_33735,N_32228);
nor U34030 (N_34030,N_32934,N_33924);
nor U34031 (N_34031,N_33133,N_32586);
or U34032 (N_34032,N_32634,N_33495);
nand U34033 (N_34033,N_32875,N_32522);
nand U34034 (N_34034,N_32122,N_32563);
nand U34035 (N_34035,N_32372,N_33811);
or U34036 (N_34036,N_33087,N_33395);
nor U34037 (N_34037,N_33219,N_32518);
and U34038 (N_34038,N_33103,N_32957);
or U34039 (N_34039,N_32544,N_32028);
and U34040 (N_34040,N_32063,N_32300);
nand U34041 (N_34041,N_33659,N_33500);
and U34042 (N_34042,N_33902,N_33834);
or U34043 (N_34043,N_32629,N_32929);
and U34044 (N_34044,N_32124,N_32207);
nor U34045 (N_34045,N_32584,N_33231);
nand U34046 (N_34046,N_32249,N_33243);
or U34047 (N_34047,N_33731,N_33012);
or U34048 (N_34048,N_33223,N_33304);
and U34049 (N_34049,N_33042,N_33781);
and U34050 (N_34050,N_32267,N_32409);
and U34051 (N_34051,N_33208,N_33007);
and U34052 (N_34052,N_32433,N_33506);
and U34053 (N_34053,N_33464,N_32469);
nor U34054 (N_34054,N_32840,N_32752);
nor U34055 (N_34055,N_32025,N_33469);
or U34056 (N_34056,N_33875,N_32571);
or U34057 (N_34057,N_33480,N_33196);
nand U34058 (N_34058,N_33242,N_33559);
nand U34059 (N_34059,N_33239,N_32517);
or U34060 (N_34060,N_33018,N_32337);
or U34061 (N_34061,N_32134,N_33197);
nand U34062 (N_34062,N_32980,N_32911);
nor U34063 (N_34063,N_32554,N_32681);
xor U34064 (N_34064,N_32261,N_33502);
nor U34065 (N_34065,N_33368,N_32692);
nand U34066 (N_34066,N_33770,N_32931);
xor U34067 (N_34067,N_32465,N_32258);
or U34068 (N_34068,N_32493,N_33068);
xnor U34069 (N_34069,N_32510,N_32339);
nor U34070 (N_34070,N_33118,N_33934);
or U34071 (N_34071,N_33008,N_32658);
xor U34072 (N_34072,N_32596,N_33422);
nand U34073 (N_34073,N_33125,N_33862);
and U34074 (N_34074,N_32998,N_33356);
nand U34075 (N_34075,N_33583,N_33590);
and U34076 (N_34076,N_33436,N_32449);
or U34077 (N_34077,N_32519,N_32311);
nand U34078 (N_34078,N_33747,N_32073);
and U34079 (N_34079,N_33358,N_33281);
and U34080 (N_34080,N_33473,N_33124);
nor U34081 (N_34081,N_33619,N_33060);
or U34082 (N_34082,N_32437,N_33056);
or U34083 (N_34083,N_32236,N_33078);
nand U34084 (N_34084,N_33261,N_32853);
nand U34085 (N_34085,N_33740,N_32939);
and U34086 (N_34086,N_32945,N_33966);
nor U34087 (N_34087,N_33161,N_32200);
nor U34088 (N_34088,N_33971,N_33274);
and U34089 (N_34089,N_33280,N_32794);
nor U34090 (N_34090,N_33977,N_33083);
and U34091 (N_34091,N_33105,N_33683);
nand U34092 (N_34092,N_32247,N_33172);
nor U34093 (N_34093,N_32706,N_32112);
and U34094 (N_34094,N_32944,N_32040);
or U34095 (N_34095,N_32222,N_32959);
or U34096 (N_34096,N_32276,N_32460);
or U34097 (N_34097,N_32012,N_32221);
nand U34098 (N_34098,N_33857,N_33230);
nand U34099 (N_34099,N_32826,N_33100);
nand U34100 (N_34100,N_33290,N_33625);
or U34101 (N_34101,N_32499,N_33795);
or U34102 (N_34102,N_33262,N_32987);
or U34103 (N_34103,N_33163,N_32377);
xor U34104 (N_34104,N_32146,N_32640);
nor U34105 (N_34105,N_33753,N_33427);
or U34106 (N_34106,N_33763,N_32144);
or U34107 (N_34107,N_32952,N_32855);
nand U34108 (N_34108,N_33364,N_32780);
xor U34109 (N_34109,N_33757,N_32650);
nor U34110 (N_34110,N_33476,N_32196);
or U34111 (N_34111,N_32463,N_33397);
nand U34112 (N_34112,N_33352,N_32440);
or U34113 (N_34113,N_32342,N_33286);
nor U34114 (N_34114,N_33445,N_32999);
or U34115 (N_34115,N_32180,N_33412);
nand U34116 (N_34116,N_32282,N_32331);
xor U34117 (N_34117,N_33613,N_33079);
nand U34118 (N_34118,N_32751,N_33866);
nor U34119 (N_34119,N_33994,N_32813);
and U34120 (N_34120,N_33727,N_32625);
nor U34121 (N_34121,N_32621,N_32209);
nand U34122 (N_34122,N_32630,N_32006);
or U34123 (N_34123,N_32951,N_32232);
or U34124 (N_34124,N_32070,N_32670);
or U34125 (N_34125,N_33308,N_33481);
and U34126 (N_34126,N_33265,N_33387);
nand U34127 (N_34127,N_33755,N_32926);
or U34128 (N_34128,N_33482,N_32545);
nand U34129 (N_34129,N_33306,N_33858);
or U34130 (N_34130,N_32747,N_33714);
nor U34131 (N_34131,N_33347,N_33188);
or U34132 (N_34132,N_32850,N_33657);
and U34133 (N_34133,N_33895,N_33191);
xnor U34134 (N_34134,N_33179,N_32946);
and U34135 (N_34135,N_32830,N_32714);
or U34136 (N_34136,N_32214,N_33001);
or U34137 (N_34137,N_32487,N_33375);
nor U34138 (N_34138,N_33848,N_32483);
and U34139 (N_34139,N_33718,N_32110);
and U34140 (N_34140,N_32605,N_33303);
and U34141 (N_34141,N_33992,N_33537);
nor U34142 (N_34142,N_32598,N_33094);
and U34143 (N_34143,N_33809,N_33093);
nand U34144 (N_34144,N_32966,N_32489);
and U34145 (N_34145,N_33370,N_33510);
or U34146 (N_34146,N_32528,N_33543);
nor U34147 (N_34147,N_33513,N_33877);
nand U34148 (N_34148,N_33131,N_32065);
nand U34149 (N_34149,N_32682,N_32461);
nor U34150 (N_34150,N_32240,N_32099);
or U34151 (N_34151,N_33392,N_33546);
nand U34152 (N_34152,N_32686,N_32626);
nand U34153 (N_34153,N_33146,N_33253);
and U34154 (N_34154,N_32860,N_33900);
nand U34155 (N_34155,N_32665,N_32928);
and U34156 (N_34156,N_32321,N_33057);
nor U34157 (N_34157,N_32817,N_33915);
or U34158 (N_34158,N_33109,N_33340);
nand U34159 (N_34159,N_33471,N_32120);
nand U34160 (N_34160,N_33844,N_32867);
and U34161 (N_34161,N_32930,N_33067);
nand U34162 (N_34162,N_33701,N_33679);
nand U34163 (N_34163,N_32774,N_33447);
and U34164 (N_34164,N_33522,N_32594);
and U34165 (N_34165,N_33346,N_33704);
and U34166 (N_34166,N_33429,N_32368);
nand U34167 (N_34167,N_33189,N_32674);
nor U34168 (N_34168,N_33493,N_33489);
or U34169 (N_34169,N_32317,N_33601);
xor U34170 (N_34170,N_33573,N_32603);
nor U34171 (N_34171,N_32907,N_32245);
and U34172 (N_34172,N_33115,N_33806);
or U34173 (N_34173,N_32785,N_33616);
nor U34174 (N_34174,N_32845,N_32707);
nand U34175 (N_34175,N_32761,N_33600);
nand U34176 (N_34176,N_33864,N_33497);
nand U34177 (N_34177,N_33821,N_33278);
nand U34178 (N_34178,N_32547,N_32184);
or U34179 (N_34179,N_32917,N_33039);
nand U34180 (N_34180,N_32635,N_32906);
nor U34181 (N_34181,N_33780,N_32264);
and U34182 (N_34182,N_33141,N_32624);
nand U34183 (N_34183,N_32387,N_33802);
nor U34184 (N_34184,N_32161,N_32857);
or U34185 (N_34185,N_33388,N_33377);
and U34186 (N_34186,N_33111,N_33107);
nand U34187 (N_34187,N_32763,N_32565);
nor U34188 (N_34188,N_32434,N_33271);
nand U34189 (N_34189,N_33973,N_32572);
nor U34190 (N_34190,N_32836,N_33720);
or U34191 (N_34191,N_32982,N_32568);
nand U34192 (N_34192,N_32234,N_32283);
nor U34193 (N_34193,N_32173,N_33968);
nand U34194 (N_34194,N_33211,N_33860);
and U34195 (N_34195,N_33080,N_32877);
nor U34196 (N_34196,N_32710,N_33147);
nand U34197 (N_34197,N_33650,N_32858);
or U34198 (N_34198,N_33694,N_32807);
nor U34199 (N_34199,N_33017,N_32022);
nand U34200 (N_34200,N_32008,N_32037);
and U34201 (N_34201,N_33354,N_32275);
and U34202 (N_34202,N_33563,N_32239);
nor U34203 (N_34203,N_33366,N_33050);
or U34204 (N_34204,N_33713,N_32436);
nand U34205 (N_34205,N_33166,N_33769);
xor U34206 (N_34206,N_33453,N_32627);
or U34207 (N_34207,N_33997,N_32213);
nor U34208 (N_34208,N_32150,N_33750);
or U34209 (N_34209,N_32474,N_33046);
or U34210 (N_34210,N_33626,N_33015);
or U34211 (N_34211,N_32032,N_33010);
or U34212 (N_34212,N_32673,N_33437);
nand U34213 (N_34213,N_32767,N_33646);
nor U34214 (N_34214,N_32690,N_33317);
nand U34215 (N_34215,N_33104,N_32125);
nand U34216 (N_34216,N_33468,N_33122);
nor U34217 (N_34217,N_33835,N_32285);
nand U34218 (N_34218,N_32856,N_33120);
and U34219 (N_34219,N_33484,N_32991);
and U34220 (N_34220,N_33962,N_33890);
or U34221 (N_34221,N_33539,N_33527);
and U34222 (N_34222,N_32534,N_33730);
nand U34223 (N_34223,N_32087,N_32582);
nor U34224 (N_34224,N_33993,N_32986);
or U34225 (N_34225,N_32071,N_33981);
or U34226 (N_34226,N_32178,N_33201);
and U34227 (N_34227,N_32511,N_33726);
and U34228 (N_34228,N_32796,N_33246);
nand U34229 (N_34229,N_33210,N_33096);
nand U34230 (N_34230,N_32615,N_32492);
nand U34231 (N_34231,N_33643,N_32663);
nand U34232 (N_34232,N_33918,N_33097);
or U34233 (N_34233,N_32805,N_32689);
nand U34234 (N_34234,N_33833,N_33439);
xor U34235 (N_34235,N_33373,N_33085);
xnor U34236 (N_34236,N_32168,N_32198);
or U34237 (N_34237,N_32391,N_33558);
nand U34238 (N_34238,N_32443,N_32696);
nor U34239 (N_34239,N_32031,N_32897);
and U34240 (N_34240,N_32356,N_32887);
nand U34241 (N_34241,N_33571,N_32229);
nor U34242 (N_34242,N_33221,N_32735);
or U34243 (N_34243,N_33098,N_32581);
nand U34244 (N_34244,N_33855,N_32106);
or U34245 (N_34245,N_33764,N_32369);
nand U34246 (N_34246,N_32109,N_32252);
and U34247 (N_34247,N_33095,N_32126);
or U34248 (N_34248,N_33765,N_32250);
nor U34249 (N_34249,N_33937,N_33719);
and U34250 (N_34250,N_33449,N_32038);
nand U34251 (N_34251,N_33310,N_32558);
and U34252 (N_34252,N_32979,N_32403);
or U34253 (N_34253,N_33156,N_32383);
or U34254 (N_34254,N_33121,N_32098);
nand U34255 (N_34255,N_32371,N_33138);
or U34256 (N_34256,N_33609,N_33779);
or U34257 (N_34257,N_32925,N_32599);
or U34258 (N_34258,N_32298,N_32623);
nor U34259 (N_34259,N_33333,N_32176);
nand U34260 (N_34260,N_33006,N_33697);
nand U34261 (N_34261,N_32651,N_33000);
nor U34262 (N_34262,N_32559,N_33220);
and U34263 (N_34263,N_32684,N_32494);
nor U34264 (N_34264,N_32709,N_32749);
nand U34265 (N_34265,N_32158,N_33778);
nand U34266 (N_34266,N_33542,N_32384);
or U34267 (N_34267,N_32427,N_33487);
nor U34268 (N_34268,N_32400,N_32064);
xnor U34269 (N_34269,N_32241,N_32143);
nand U34270 (N_34270,N_33359,N_33910);
or U34271 (N_34271,N_33393,N_33576);
and U34272 (N_34272,N_33479,N_32014);
or U34273 (N_34273,N_32846,N_33812);
nand U34274 (N_34274,N_33608,N_32808);
and U34275 (N_34275,N_33963,N_32136);
or U34276 (N_34276,N_33294,N_33548);
nand U34277 (N_34277,N_32700,N_33176);
and U34278 (N_34278,N_33801,N_32162);
nor U34279 (N_34279,N_33532,N_32829);
nand U34280 (N_34280,N_32549,N_32701);
nand U34281 (N_34281,N_33030,N_32533);
or U34282 (N_34282,N_33491,N_33160);
or U34283 (N_34283,N_32574,N_32795);
nand U34284 (N_34284,N_33550,N_33224);
nor U34285 (N_34285,N_32981,N_33043);
nand U34286 (N_34286,N_33268,N_33381);
or U34287 (N_34287,N_32290,N_32550);
nor U34288 (N_34288,N_33301,N_33742);
or U34289 (N_34289,N_32938,N_32313);
and U34290 (N_34290,N_32085,N_32183);
and U34291 (N_34291,N_33503,N_33951);
nand U34292 (N_34292,N_32187,N_33034);
nand U34293 (N_34293,N_33520,N_32215);
and U34294 (N_34294,N_33749,N_32733);
and U34295 (N_34295,N_32051,N_33027);
nor U34296 (N_34296,N_32773,N_33020);
nor U34297 (N_34297,N_32307,N_33061);
nand U34298 (N_34298,N_33676,N_32753);
or U34299 (N_34299,N_33045,N_33140);
and U34300 (N_34300,N_33345,N_32348);
and U34301 (N_34301,N_32672,N_33843);
and U34302 (N_34302,N_33361,N_32828);
or U34303 (N_34303,N_33592,N_33565);
and U34304 (N_34304,N_33884,N_32834);
nand U34305 (N_34305,N_32719,N_32140);
or U34306 (N_34306,N_32172,N_33168);
or U34307 (N_34307,N_33715,N_33227);
nand U34308 (N_34308,N_32535,N_32882);
nand U34309 (N_34309,N_32130,N_32688);
or U34310 (N_34310,N_32555,N_32157);
nand U34311 (N_34311,N_33171,N_32026);
nor U34312 (N_34312,N_32491,N_32050);
or U34313 (N_34313,N_33839,N_33582);
and U34314 (N_34314,N_33882,N_32912);
or U34315 (N_34315,N_32797,N_32890);
nor U34316 (N_34316,N_33925,N_33005);
nor U34317 (N_34317,N_33612,N_33671);
and U34318 (N_34318,N_33167,N_32956);
and U34319 (N_34319,N_33233,N_32741);
nand U34320 (N_34320,N_33435,N_33673);
nor U34321 (N_34321,N_32382,N_32152);
nand U34322 (N_34322,N_32057,N_32843);
nor U34323 (N_34323,N_33150,N_32074);
nand U34324 (N_34324,N_33287,N_32978);
nor U34325 (N_34325,N_33617,N_33872);
or U34326 (N_34326,N_32537,N_33837);
nand U34327 (N_34327,N_33421,N_33722);
nor U34328 (N_34328,N_33631,N_32990);
or U34329 (N_34329,N_33316,N_33250);
nor U34330 (N_34330,N_33028,N_32430);
and U34331 (N_34331,N_33929,N_32048);
and U34332 (N_34332,N_33987,N_33645);
or U34333 (N_34333,N_32645,N_32784);
nand U34334 (N_34334,N_32133,N_32647);
or U34335 (N_34335,N_32113,N_33205);
nand U34336 (N_34336,N_33817,N_33832);
xnor U34337 (N_34337,N_33157,N_33399);
xnor U34338 (N_34338,N_32385,N_32045);
nor U34339 (N_34339,N_32776,N_32378);
and U34340 (N_34340,N_33808,N_33228);
nand U34341 (N_34341,N_33475,N_32141);
and U34342 (N_34342,N_32192,N_32224);
nor U34343 (N_34343,N_33568,N_33607);
or U34344 (N_34344,N_33515,N_33674);
nor U34345 (N_34345,N_33212,N_32995);
nand U34346 (N_34346,N_32865,N_33195);
or U34347 (N_34347,N_32913,N_33178);
nand U34348 (N_34348,N_33830,N_33181);
or U34349 (N_34349,N_33825,N_32016);
nor U34350 (N_34350,N_33815,N_32886);
or U34351 (N_34351,N_33062,N_33295);
and U34352 (N_34352,N_33092,N_33614);
and U34353 (N_34353,N_32464,N_32445);
or U34354 (N_34354,N_32948,N_32047);
or U34355 (N_34355,N_32728,N_32167);
nor U34356 (N_34356,N_33751,N_32607);
nor U34357 (N_34357,N_33737,N_32216);
and U34358 (N_34358,N_33457,N_32470);
or U34359 (N_34359,N_33967,N_32595);
or U34360 (N_34360,N_32086,N_33644);
or U34361 (N_34361,N_33184,N_33604);
nor U34362 (N_34362,N_32322,N_32839);
or U34363 (N_34363,N_32854,N_33741);
nand U34364 (N_34364,N_33450,N_33923);
or U34365 (N_34365,N_32438,N_32898);
or U34366 (N_34366,N_32334,N_33661);
and U34367 (N_34367,N_33752,N_33591);
or U34368 (N_34368,N_33385,N_32066);
nor U34369 (N_34369,N_32062,N_33130);
or U34370 (N_34370,N_32578,N_33762);
xnor U34371 (N_34371,N_33709,N_33905);
nor U34372 (N_34372,N_32546,N_32435);
nand U34373 (N_34373,N_33952,N_32636);
nor U34374 (N_34374,N_33868,N_32514);
nand U34375 (N_34375,N_32210,N_33360);
nand U34376 (N_34376,N_33049,N_33022);
or U34377 (N_34377,N_32989,N_33690);
nor U34378 (N_34378,N_32632,N_32823);
nor U34379 (N_34379,N_33116,N_32556);
nand U34380 (N_34380,N_32458,N_32076);
and U34381 (N_34381,N_33894,N_32360);
or U34382 (N_34382,N_33648,N_32820);
or U34383 (N_34383,N_33414,N_33653);
and U34384 (N_34384,N_32611,N_32478);
nand U34385 (N_34385,N_32381,N_32412);
nor U34386 (N_34386,N_33960,N_32965);
or U34387 (N_34387,N_32375,N_33639);
nand U34388 (N_34388,N_33173,N_33424);
and U34389 (N_34389,N_33496,N_33789);
nor U34390 (N_34390,N_32266,N_32811);
nand U34391 (N_34391,N_32802,N_32316);
or U34392 (N_34392,N_33177,N_32359);
and U34393 (N_34393,N_32278,N_32833);
nand U34394 (N_34394,N_33748,N_32347);
and U34395 (N_34395,N_32924,N_32837);
nor U34396 (N_34396,N_32341,N_32128);
nand U34397 (N_34397,N_33428,N_32077);
or U34398 (N_34398,N_32166,N_32212);
or U34399 (N_34399,N_33058,N_33483);
nor U34400 (N_34400,N_33922,N_33207);
nand U34401 (N_34401,N_32251,N_33486);
nand U34402 (N_34402,N_32277,N_32713);
or U34403 (N_34403,N_32799,N_32764);
nand U34404 (N_34404,N_33656,N_33386);
nand U34405 (N_34405,N_33828,N_33598);
and U34406 (N_34406,N_33091,N_33965);
or U34407 (N_34407,N_33859,N_32666);
and U34408 (N_34408,N_33553,N_32693);
or U34409 (N_34409,N_32975,N_32495);
nand U34410 (N_34410,N_32675,N_32035);
nor U34411 (N_34411,N_32677,N_33818);
or U34412 (N_34412,N_33786,N_33193);
or U34413 (N_34413,N_33530,N_33324);
and U34414 (N_34414,N_32254,N_32778);
or U34415 (N_34415,N_32861,N_33685);
nand U34416 (N_34416,N_33512,N_33379);
nor U34417 (N_34417,N_32481,N_33101);
and U34418 (N_34418,N_32668,N_33691);
or U34419 (N_34419,N_32628,N_32185);
xnor U34420 (N_34420,N_32954,N_33746);
nand U34421 (N_34421,N_32081,N_32885);
or U34422 (N_34422,N_33641,N_32521);
and U34423 (N_34423,N_32480,N_33266);
or U34424 (N_34424,N_33723,N_32903);
xnor U34425 (N_34425,N_32659,N_32118);
and U34426 (N_34426,N_32505,N_32332);
nor U34427 (N_34427,N_32792,N_33838);
xor U34428 (N_34428,N_32421,N_32791);
nor U34429 (N_34429,N_32188,N_33696);
or U34430 (N_34430,N_32775,N_32896);
nor U34431 (N_34431,N_32159,N_32899);
nor U34432 (N_34432,N_32575,N_33470);
nor U34433 (N_34433,N_33805,N_33326);
nor U34434 (N_34434,N_32732,N_32407);
and U34435 (N_34435,N_32054,N_33813);
or U34436 (N_34436,N_32553,N_33739);
nor U34437 (N_34437,N_33126,N_32755);
nand U34438 (N_34438,N_33772,N_33309);
nor U34439 (N_34439,N_33052,N_33214);
or U34440 (N_34440,N_33759,N_33716);
or U34441 (N_34441,N_33552,N_32094);
and U34442 (N_34442,N_33190,N_32408);
or U34443 (N_34443,N_33881,N_32186);
nor U34444 (N_34444,N_33182,N_33688);
or U34445 (N_34445,N_33127,N_32415);
nor U34446 (N_34446,N_32524,N_32750);
nor U34447 (N_34447,N_32450,N_33957);
nor U34448 (N_34448,N_32175,N_33972);
nand U34449 (N_34449,N_32541,N_33867);
and U34450 (N_34450,N_33842,N_33892);
nor U34451 (N_34451,N_32639,N_32219);
nor U34452 (N_34452,N_32592,N_32477);
and U34453 (N_34453,N_33288,N_33011);
or U34454 (N_34454,N_32294,N_32910);
nor U34455 (N_34455,N_32312,N_32889);
nor U34456 (N_34456,N_33038,N_32864);
and U34457 (N_34457,N_33819,N_32961);
and U34458 (N_34458,N_33850,N_32069);
or U34459 (N_34459,N_32503,N_33545);
and U34460 (N_34460,N_33311,N_33766);
or U34461 (N_34461,N_32870,N_32123);
or U34462 (N_34462,N_33871,N_32419);
or U34463 (N_34463,N_32358,N_32798);
nand U34464 (N_34464,N_32225,N_32758);
nor U34465 (N_34465,N_33273,N_32042);
nor U34466 (N_34466,N_33279,N_33444);
or U34467 (N_34467,N_32153,N_32793);
nand U34468 (N_34468,N_33672,N_32398);
or U34469 (N_34469,N_32958,N_32013);
and U34470 (N_34470,N_32868,N_32500);
and U34471 (N_34471,N_32679,N_33187);
nand U34472 (N_34472,N_32357,N_32223);
nand U34473 (N_34473,N_32243,N_32844);
nand U34474 (N_34474,N_33245,N_32325);
and U34475 (N_34475,N_32656,N_32302);
nand U34476 (N_34476,N_32740,N_33112);
nand U34477 (N_34477,N_32181,N_32297);
and U34478 (N_34478,N_32079,N_33627);
and U34479 (N_34479,N_33978,N_32467);
and U34480 (N_34480,N_32335,N_32804);
nor U34481 (N_34481,N_32955,N_33441);
or U34482 (N_34482,N_32993,N_33192);
or U34483 (N_34483,N_33396,N_33426);
nand U34484 (N_34484,N_33928,N_32242);
nand U34485 (N_34485,N_33999,N_33845);
and U34486 (N_34486,N_32525,N_33852);
or U34487 (N_34487,N_33363,N_33041);
nor U34488 (N_34488,N_33410,N_32373);
or U34489 (N_34489,N_33423,N_33320);
or U34490 (N_34490,N_33829,N_33357);
and U34491 (N_34491,N_32760,N_32479);
or U34492 (N_34492,N_33632,N_33595);
and U34493 (N_34493,N_32281,N_32648);
nor U34494 (N_34494,N_33870,N_32723);
nor U34495 (N_34495,N_33137,N_33695);
nand U34496 (N_34496,N_32869,N_32617);
or U34497 (N_34497,N_33913,N_32090);
or U34498 (N_34498,N_33216,N_33380);
or U34499 (N_34499,N_32306,N_33970);
or U34500 (N_34500,N_32206,N_32320);
or U34501 (N_34501,N_32148,N_33637);
and U34502 (N_34502,N_32637,N_33088);
nor U34503 (N_34503,N_32315,N_33047);
nor U34504 (N_34504,N_32205,N_32138);
or U34505 (N_34505,N_33785,N_32490);
nand U34506 (N_34506,N_32286,N_32619);
nand U34507 (N_34507,N_33814,N_33323);
nand U34508 (N_34508,N_33432,N_33569);
or U34509 (N_34509,N_32075,N_32475);
nand U34510 (N_34510,N_32333,N_33073);
nand U34511 (N_34511,N_32936,N_32263);
and U34512 (N_34512,N_33135,N_33334);
or U34513 (N_34513,N_33712,N_33175);
nand U34514 (N_34514,N_33040,N_32745);
and U34515 (N_34515,N_32497,N_33796);
nand U34516 (N_34516,N_32455,N_32585);
or U34517 (N_34517,N_33291,N_32697);
nor U34518 (N_34518,N_33562,N_32685);
nor U34519 (N_34519,N_33322,N_33165);
or U34520 (N_34520,N_32366,N_33053);
and U34521 (N_34521,N_33257,N_33931);
nor U34522 (N_34522,N_32273,N_32878);
and U34523 (N_34523,N_33851,N_33807);
and U34524 (N_34524,N_32204,N_33907);
and U34525 (N_34525,N_32721,N_32036);
or U34526 (N_34526,N_32516,N_33466);
nand U34527 (N_34527,N_33700,N_33820);
and U34528 (N_34528,N_33425,N_33081);
or U34529 (N_34529,N_33874,N_33794);
nand U34530 (N_34530,N_32327,N_32532);
nor U34531 (N_34531,N_32034,N_33911);
and U34532 (N_34532,N_32105,N_32768);
nor U34533 (N_34533,N_32114,N_33917);
or U34534 (N_34534,N_32379,N_33132);
nand U34535 (N_34535,N_32388,N_32323);
and U34536 (N_34536,N_33048,N_33580);
nand U34537 (N_34537,N_32699,N_32145);
nor U34538 (N_34538,N_32231,N_33313);
or U34539 (N_34539,N_32631,N_32884);
and U34540 (N_34540,N_33430,N_33792);
or U34541 (N_34541,N_33948,N_32324);
nor U34542 (N_34542,N_33777,N_32743);
nand U34543 (N_34543,N_32259,N_32597);
or U34544 (N_34544,N_32852,N_32248);
and U34545 (N_34545,N_33452,N_33572);
nor U34546 (N_34546,N_32874,N_33054);
or U34547 (N_34547,N_33021,N_32244);
and U34548 (N_34548,N_33706,N_32742);
nor U34549 (N_34549,N_33169,N_33745);
or U34550 (N_34550,N_33465,N_32160);
or U34551 (N_34551,N_33222,N_32888);
nand U34552 (N_34552,N_32257,N_33258);
or U34553 (N_34553,N_33256,N_33810);
nor U34554 (N_34554,N_32919,N_33976);
nor U34555 (N_34555,N_33678,N_33873);
or U34556 (N_34556,N_33754,N_32800);
or U34557 (N_34557,N_32824,N_33974);
nor U34558 (N_34558,N_33947,N_33655);
nand U34559 (N_34559,N_33330,N_32600);
nand U34560 (N_34560,N_33296,N_32270);
or U34561 (N_34561,N_32863,N_33139);
nand U34562 (N_34562,N_32203,N_33025);
or U34563 (N_34563,N_32095,N_33144);
and U34564 (N_34564,N_33117,N_32226);
nand U34565 (N_34565,N_33888,N_32570);
and U34566 (N_34566,N_33721,N_33588);
nand U34567 (N_34567,N_33689,N_33297);
nor U34568 (N_34568,N_32473,N_33633);
or U34569 (N_34569,N_33315,N_33329);
nor U34570 (N_34570,N_32043,N_33578);
or U34571 (N_34571,N_32984,N_33406);
xnor U34572 (N_34572,N_33505,N_32810);
nand U34573 (N_34573,N_33267,N_33897);
and U34574 (N_34574,N_32446,N_33623);
or U34575 (N_34575,N_33524,N_32687);
and U34576 (N_34576,N_32174,N_32111);
xnor U34577 (N_34577,N_32705,N_32646);
or U34578 (N_34578,N_32643,N_33930);
and U34579 (N_34579,N_32527,N_32059);
nand U34580 (N_34580,N_32891,N_32940);
nand U34581 (N_34581,N_33272,N_33402);
nor U34582 (N_34582,N_32488,N_33136);
nor U34583 (N_34583,N_33919,N_32502);
and U34584 (N_34584,N_33415,N_32424);
and U34585 (N_34585,N_33110,N_32873);
and U34586 (N_34586,N_33988,N_32072);
nor U34587 (N_34587,N_33538,N_32002);
and U34588 (N_34588,N_33666,N_32457);
xnor U34589 (N_34589,N_33853,N_33959);
and U34590 (N_34590,N_33799,N_33529);
nor U34591 (N_34591,N_32918,N_32135);
nand U34592 (N_34592,N_32269,N_32314);
nand U34593 (N_34593,N_32256,N_33705);
nor U34594 (N_34594,N_33418,N_32589);
nor U34595 (N_34595,N_33557,N_33991);
or U34596 (N_34596,N_32509,N_33516);
and U34597 (N_34597,N_33912,N_32121);
nand U34598 (N_34598,N_32468,N_33351);
nand U34599 (N_34599,N_32691,N_32061);
xor U34600 (N_34600,N_32921,N_33677);
and U34601 (N_34601,N_32295,N_32872);
nor U34602 (N_34602,N_33490,N_33886);
and U34603 (N_34603,N_32818,N_33394);
and U34604 (N_34604,N_33443,N_33129);
nand U34605 (N_34605,N_33300,N_33949);
nand U34606 (N_34606,N_32579,N_33086);
or U34607 (N_34607,N_32272,N_32336);
and U34608 (N_34608,N_33790,N_33371);
nand U34609 (N_34609,N_33567,N_33621);
and U34610 (N_34610,N_33014,N_32835);
or U34611 (N_34611,N_32551,N_33463);
nand U34612 (N_34612,N_33174,N_32058);
and U34613 (N_34613,N_32744,N_33896);
nor U34614 (N_34614,N_33536,N_33831);
and U34615 (N_34615,N_33328,N_33082);
or U34616 (N_34616,N_32201,N_32523);
and U34617 (N_34617,N_32169,N_32769);
nor U34618 (N_34618,N_32292,N_33787);
or U34619 (N_34619,N_33797,N_33456);
and U34620 (N_34620,N_33634,N_33932);
or U34621 (N_34621,N_33254,N_32608);
xor U34622 (N_34622,N_32195,N_33756);
and U34623 (N_34623,N_33411,N_32217);
nand U34624 (N_34624,N_32716,N_33401);
nand U34625 (N_34625,N_33438,N_33909);
nor U34626 (N_34626,N_33460,N_33555);
nand U34627 (N_34627,N_33498,N_32024);
and U34628 (N_34628,N_32401,N_32237);
or U34629 (N_34629,N_33687,N_33836);
nor U34630 (N_34630,N_32462,N_32208);
nor U34631 (N_34631,N_32350,N_32591);
nor U34632 (N_34632,N_33744,N_32396);
nand U34633 (N_34633,N_32814,N_32593);
or U34634 (N_34634,N_33587,N_33640);
nor U34635 (N_34635,N_33605,N_33292);
nand U34636 (N_34636,N_33255,N_32116);
and U34637 (N_34637,N_33708,N_32738);
xnor U34638 (N_34638,N_32847,N_33840);
xnor U34639 (N_34639,N_33405,N_33283);
nand U34640 (N_34640,N_32049,N_32486);
nor U34641 (N_34641,N_32452,N_32466);
and U34642 (N_34642,N_33180,N_33123);
and U34643 (N_34643,N_32447,N_32235);
nor U34644 (N_34644,N_32905,N_33226);
nand U34645 (N_34645,N_32301,N_32456);
or U34646 (N_34646,N_33409,N_32927);
nand U34647 (N_34647,N_32801,N_32053);
xor U34648 (N_34648,N_33533,N_33349);
nor U34649 (N_34649,N_33089,N_33108);
nor U34650 (N_34650,N_32389,N_33856);
or U34651 (N_34651,N_33004,N_33654);
nand U34652 (N_34652,N_32299,N_33238);
and U34653 (N_34653,N_33164,N_32155);
and U34654 (N_34654,N_32017,N_32088);
or U34655 (N_34655,N_33577,N_33331);
nor U34656 (N_34656,N_32765,N_32132);
nand U34657 (N_34657,N_33090,N_32425);
or U34658 (N_34658,N_33950,N_32506);
nand U34659 (N_34659,N_33589,N_32851);
nand U34660 (N_34660,N_32819,N_32182);
nand U34661 (N_34661,N_33903,N_32046);
nand U34662 (N_34662,N_33684,N_32901);
nand U34663 (N_34663,N_32287,N_33773);
nor U34664 (N_34664,N_33143,N_32363);
xor U34665 (N_34665,N_33348,N_33235);
or U34666 (N_34666,N_33743,N_33927);
nor U34667 (N_34667,N_32825,N_33635);
and U34668 (N_34668,N_33153,N_32762);
nand U34669 (N_34669,N_32923,N_32531);
or U34670 (N_34670,N_32508,N_33343);
nor U34671 (N_34671,N_33561,N_32103);
nor U34672 (N_34672,N_33488,N_32920);
or U34673 (N_34673,N_33440,N_32644);
or U34674 (N_34674,N_32471,N_33847);
and U34675 (N_34675,N_33732,N_33680);
and U34676 (N_34676,N_32432,N_33382);
or U34677 (N_34677,N_32972,N_32177);
or U34678 (N_34678,N_32576,N_33391);
nand U34679 (N_34679,N_32883,N_33738);
nand U34680 (N_34680,N_33072,N_32484);
or U34681 (N_34681,N_33566,N_33955);
nand U34682 (N_34682,N_32501,N_33942);
nor U34683 (N_34683,N_33106,N_32060);
nor U34684 (N_34684,N_32426,N_32428);
or U34685 (N_34685,N_33390,N_33668);
nor U34686 (N_34686,N_32781,N_33816);
or U34687 (N_34687,N_33906,N_33069);
nor U34688 (N_34688,N_33728,N_33521);
nand U34689 (N_34689,N_32983,N_32862);
nor U34690 (N_34690,N_32370,N_33681);
nand U34691 (N_34691,N_32354,N_32055);
nand U34692 (N_34692,N_32164,N_32418);
xor U34693 (N_34693,N_32498,N_33883);
nand U34694 (N_34694,N_33540,N_33051);
or U34695 (N_34695,N_33376,N_32717);
and U34696 (N_34696,N_33325,N_32194);
or U34697 (N_34697,N_32067,N_32393);
nor U34698 (N_34698,N_32416,N_32573);
or U34699 (N_34699,N_33920,N_33158);
nor U34700 (N_34700,N_32916,N_32165);
or U34701 (N_34701,N_32091,N_32590);
and U34702 (N_34702,N_32704,N_33711);
nor U34703 (N_34703,N_33339,N_32996);
nor U34704 (N_34704,N_32725,N_33194);
and U34705 (N_34705,N_33767,N_33252);
nor U34706 (N_34706,N_32859,N_33002);
nor U34707 (N_34707,N_33247,N_32093);
nor U34708 (N_34708,N_32265,N_32513);
nor U34709 (N_34709,N_33155,N_33664);
and U34710 (N_34710,N_32653,N_33019);
nor U34711 (N_34711,N_33282,N_33575);
xnor U34712 (N_34712,N_32260,N_33791);
nor U34713 (N_34713,N_32485,N_33570);
and U34714 (N_34714,N_32137,N_33703);
or U34715 (N_34715,N_32671,N_33518);
and U34716 (N_34716,N_33350,N_33037);
nand U34717 (N_34717,N_32960,N_33642);
nand U34718 (N_34718,N_32649,N_32759);
xor U34719 (N_34719,N_32561,N_32344);
and U34720 (N_34720,N_33241,N_32543);
or U34721 (N_34721,N_32676,N_33063);
nand U34722 (N_34722,N_32655,N_33462);
and U34723 (N_34723,N_32612,N_33455);
or U34724 (N_34724,N_33389,N_33594);
nand U34725 (N_34725,N_33084,N_32193);
or U34726 (N_34726,N_32737,N_33652);
nand U34727 (N_34727,N_32191,N_32557);
and U34728 (N_34728,N_33035,N_32330);
and U34729 (N_34729,N_32848,N_33270);
and U34730 (N_34730,N_32233,N_33549);
nand U34731 (N_34731,N_32015,N_33420);
nor U34732 (N_34732,N_32329,N_33454);
nor U34733 (N_34733,N_33403,N_32892);
xor U34734 (N_34734,N_32771,N_32748);
or U34735 (N_34735,N_32326,N_33827);
nand U34736 (N_34736,N_33975,N_33725);
or U34737 (N_34737,N_32220,N_32448);
nand U34738 (N_34738,N_33603,N_33314);
nor U34739 (N_34739,N_33374,N_33585);
nand U34740 (N_34740,N_33670,N_32604);
nand U34741 (N_34741,N_33055,N_33240);
and U34742 (N_34742,N_33528,N_32092);
or U34743 (N_34743,N_33586,N_32227);
nor U34744 (N_34744,N_32909,N_32255);
nand U34745 (N_34745,N_33758,N_33344);
nor U34746 (N_34746,N_33149,N_32406);
nor U34747 (N_34747,N_32000,N_33638);
or U34748 (N_34748,N_33335,N_33774);
nand U34749 (N_34749,N_33940,N_32789);
nand U34750 (N_34750,N_32394,N_33863);
nor U34751 (N_34751,N_32695,N_33338);
or U34752 (N_34752,N_32618,N_32876);
nand U34753 (N_34753,N_32620,N_32097);
nand U34754 (N_34754,N_32151,N_33263);
and U34755 (N_34755,N_33531,N_32754);
xnor U34756 (N_34756,N_33404,N_33416);
nand U34757 (N_34757,N_33372,N_32003);
or U34758 (N_34758,N_33784,N_33898);
nor U34759 (N_34759,N_33355,N_33926);
nor U34760 (N_34760,N_33507,N_33023);
nand U34761 (N_34761,N_33321,N_32715);
and U34762 (N_34762,N_33148,N_32734);
nor U34763 (N_34763,N_32777,N_33341);
nand U34764 (N_34764,N_33474,N_33823);
nor U34765 (N_34765,N_32935,N_32724);
nand U34766 (N_34766,N_32757,N_32082);
and U34767 (N_34767,N_32922,N_32253);
and U34768 (N_34768,N_33075,N_33921);
and U34769 (N_34769,N_32739,N_32788);
nor U34770 (N_34770,N_32309,N_32803);
or U34771 (N_34771,N_32328,N_32346);
and U34772 (N_34772,N_32967,N_33581);
nand U34773 (N_34773,N_32349,N_32429);
nand U34774 (N_34774,N_32414,N_32271);
or U34775 (N_34775,N_32779,N_33944);
nand U34776 (N_34776,N_33213,N_32881);
or U34777 (N_34777,N_33467,N_32994);
nor U34778 (N_34778,N_32504,N_33342);
or U34779 (N_34779,N_33803,N_32119);
nor U34780 (N_34780,N_32772,N_33945);
or U34781 (N_34781,N_32280,N_33628);
and U34782 (N_34782,N_32352,N_32101);
and U34783 (N_34783,N_33442,N_32894);
nor U34784 (N_34784,N_32096,N_33259);
and U34785 (N_34785,N_33183,N_32973);
nor U34786 (N_34786,N_32142,N_32288);
nand U34787 (N_34787,N_32131,N_33956);
and U34788 (N_34788,N_32932,N_33961);
xor U34789 (N_34789,N_32664,N_32950);
nand U34790 (N_34790,N_33734,N_33509);
or U34791 (N_34791,N_33865,N_32974);
and U34792 (N_34792,N_33693,N_33933);
nor U34793 (N_34793,N_32056,N_32374);
nor U34794 (N_34794,N_32246,N_33804);
or U34795 (N_34795,N_33099,N_32985);
nand U34796 (N_34796,N_33162,N_32340);
nand U34797 (N_34797,N_32660,N_32441);
and U34798 (N_34798,N_32529,N_33980);
nand U34799 (N_34799,N_33016,N_32147);
nand U34800 (N_34800,N_33941,N_33431);
or U34801 (N_34801,N_32661,N_32238);
nor U34802 (N_34802,N_32293,N_32783);
nor U34803 (N_34803,N_33275,N_32351);
nor U34804 (N_34804,N_33119,N_33378);
and U34805 (N_34805,N_32720,N_33876);
or U34806 (N_34806,N_32914,N_32444);
xor U34807 (N_34807,N_32638,N_32362);
or U34808 (N_34808,N_33199,N_33869);
and U34809 (N_34809,N_32577,N_33013);
nor U34810 (N_34810,N_33841,N_33824);
nand U34811 (N_34811,N_33499,N_32310);
and U34812 (N_34812,N_33793,N_32871);
and U34813 (N_34813,N_32018,N_32080);
or U34814 (N_34814,N_32809,N_33551);
or U34815 (N_34815,N_32010,N_33249);
or U34816 (N_34816,N_32367,N_32567);
nor U34817 (N_34817,N_32971,N_33003);
or U34818 (N_34818,N_33651,N_33031);
or U34819 (N_34819,N_33461,N_33026);
nand U34820 (N_34820,N_32633,N_32319);
nor U34821 (N_34821,N_33887,N_33854);
nand U34822 (N_34822,N_33682,N_32969);
or U34823 (N_34823,N_32020,N_33985);
and U34824 (N_34824,N_32727,N_33264);
nor U34825 (N_34825,N_32365,N_32539);
nor U34826 (N_34826,N_33036,N_32305);
and U34827 (N_34827,N_33485,N_33710);
nor U34828 (N_34828,N_32009,N_33861);
nand U34829 (N_34829,N_33954,N_33788);
and U34830 (N_34830,N_32941,N_33229);
nor U34831 (N_34831,N_33276,N_33159);
nor U34832 (N_34832,N_32968,N_33448);
nor U34833 (N_34833,N_33477,N_32454);
nor U34834 (N_34834,N_33152,N_32580);
nand U34835 (N_34835,N_33554,N_32189);
nand U34836 (N_34836,N_32395,N_33251);
and U34837 (N_34837,N_33407,N_32107);
nor U34838 (N_34838,N_32104,N_33660);
and U34839 (N_34839,N_32041,N_33717);
or U34840 (N_34840,N_33982,N_33198);
nand U34841 (N_34841,N_32900,N_32937);
and U34842 (N_34842,N_33504,N_32023);
nand U34843 (N_34843,N_32230,N_32616);
and U34844 (N_34844,N_32915,N_33492);
nor U34845 (N_34845,N_32520,N_32355);
or U34846 (N_34846,N_33771,N_32083);
nor U34847 (N_34847,N_33936,N_33369);
or U34848 (N_34848,N_33990,N_32613);
or U34849 (N_34849,N_33958,N_32832);
nand U34850 (N_34850,N_33946,N_33914);
nor U34851 (N_34851,N_32588,N_33908);
nand U34852 (N_34852,N_32397,N_33724);
or U34853 (N_34853,N_33269,N_32089);
nand U34854 (N_34854,N_33417,N_33044);
or U34855 (N_34855,N_33989,N_33889);
nor U34856 (N_34856,N_33798,N_33629);
or U34857 (N_34857,N_32420,N_33939);
and U34858 (N_34858,N_33151,N_32392);
and U34859 (N_34859,N_32411,N_32654);
nand U34860 (N_34860,N_33074,N_33699);
nor U34861 (N_34861,N_33783,N_32536);
nand U34862 (N_34862,N_32933,N_32821);
and U34863 (N_34863,N_32641,N_33337);
nand U34864 (N_34864,N_33202,N_32030);
or U34865 (N_34865,N_33953,N_32033);
and U34866 (N_34866,N_32822,N_32730);
nand U34867 (N_34867,N_33782,N_32703);
or U34868 (N_34868,N_33142,N_32496);
nor U34869 (N_34869,N_32279,N_32816);
nand U34870 (N_34870,N_32949,N_32343);
xnor U34871 (N_34871,N_33446,N_32364);
or U34872 (N_34872,N_33800,N_32782);
and U34873 (N_34873,N_32806,N_32708);
nand U34874 (N_34874,N_33059,N_33327);
nor U34875 (N_34875,N_32039,N_33362);
or U34876 (N_34876,N_32992,N_33964);
nand U34877 (N_34877,N_33526,N_32552);
nand U34878 (N_34878,N_32812,N_32827);
nand U34879 (N_34879,N_32262,N_32413);
or U34880 (N_34880,N_33353,N_33574);
nand U34881 (N_34881,N_32345,N_32507);
xnor U34882 (N_34882,N_33636,N_32893);
and U34883 (N_34883,N_33204,N_32476);
nand U34884 (N_34884,N_33776,N_32170);
and U34885 (N_34885,N_33707,N_33508);
nand U34886 (N_34886,N_32417,N_33534);
nand U34887 (N_34887,N_32386,N_33620);
nand U34888 (N_34888,N_32694,N_32453);
or U34889 (N_34889,N_32953,N_33186);
nor U34890 (N_34890,N_33289,N_33729);
and U34891 (N_34891,N_33299,N_32291);
and U34892 (N_34892,N_33935,N_33458);
nand U34893 (N_34893,N_32988,N_32318);
or U34894 (N_34894,N_33599,N_32583);
nor U34895 (N_34895,N_32746,N_32902);
nand U34896 (N_34896,N_33986,N_33560);
nand U34897 (N_34897,N_32842,N_33236);
nand U34898 (N_34898,N_32338,N_33413);
or U34899 (N_34899,N_33663,N_33302);
and U34900 (N_34900,N_32004,N_32007);
nand U34901 (N_34901,N_33878,N_33319);
nand U34902 (N_34902,N_32274,N_32402);
and U34903 (N_34903,N_32711,N_33893);
and U34904 (N_34904,N_33336,N_33318);
nor U34905 (N_34905,N_32977,N_33615);
nor U34906 (N_34906,N_32100,N_32199);
nand U34907 (N_34907,N_33332,N_32376);
xnor U34908 (N_34908,N_32005,N_32530);
and U34909 (N_34909,N_33686,N_33983);
nand U34910 (N_34910,N_33408,N_33277);
nand U34911 (N_34911,N_33736,N_32895);
or U34912 (N_34912,N_33365,N_32606);
or U34913 (N_34913,N_32451,N_33451);
nor U34914 (N_34914,N_32027,N_33514);
nor U34915 (N_34915,N_32218,N_33185);
nand U34916 (N_34916,N_33904,N_32815);
or U34917 (N_34917,N_33517,N_32657);
or U34918 (N_34918,N_33692,N_33606);
nor U34919 (N_34919,N_32718,N_32405);
nand U34920 (N_34920,N_33984,N_33667);
nand U34921 (N_34921,N_32542,N_32849);
and U34922 (N_34922,N_32669,N_33611);
or U34923 (N_34923,N_33134,N_32564);
and U34924 (N_34924,N_32731,N_32964);
nor U34925 (N_34925,N_32662,N_33494);
and U34926 (N_34926,N_32841,N_32562);
or U34927 (N_34927,N_32284,N_33525);
xor U34928 (N_34928,N_33434,N_33459);
and U34929 (N_34929,N_32667,N_33501);
or U34930 (N_34930,N_33733,N_33145);
and U34931 (N_34931,N_32947,N_32001);
nand U34932 (N_34932,N_32683,N_33284);
nand U34933 (N_34933,N_33584,N_32068);
and U34934 (N_34934,N_33822,N_33658);
and U34935 (N_34935,N_32866,N_33564);
or U34936 (N_34936,N_33938,N_32163);
and U34937 (N_34937,N_33649,N_32422);
nand U34938 (N_34938,N_32211,N_32908);
or U34939 (N_34939,N_33624,N_33433);
nand U34940 (N_34940,N_33891,N_32680);
nor U34941 (N_34941,N_33596,N_33544);
nand U34942 (N_34942,N_32482,N_33541);
nor U34943 (N_34943,N_32390,N_33901);
and U34944 (N_34944,N_33622,N_32569);
nand U34945 (N_34945,N_33647,N_33998);
nor U34946 (N_34946,N_32602,N_33102);
and U34947 (N_34947,N_32787,N_32548);
nand U34948 (N_34948,N_33305,N_32770);
nand U34949 (N_34949,N_33367,N_32078);
and U34950 (N_34950,N_33761,N_33472);
or U34951 (N_34951,N_33298,N_32459);
nor U34952 (N_34952,N_33849,N_32838);
nor U34953 (N_34953,N_33979,N_33556);
and U34954 (N_34954,N_32702,N_32942);
and U34955 (N_34955,N_33170,N_33511);
or U34956 (N_34956,N_32622,N_33033);
nand U34957 (N_34957,N_33293,N_33307);
nand U34958 (N_34958,N_33662,N_33579);
nand U34959 (N_34959,N_32831,N_32609);
or U34960 (N_34960,N_33547,N_33610);
nor U34961 (N_34961,N_33312,N_33384);
and U34962 (N_34962,N_33285,N_33969);
nand U34963 (N_34963,N_32976,N_33665);
nand U34964 (N_34964,N_32127,N_33248);
or U34965 (N_34965,N_33244,N_32052);
and U34966 (N_34966,N_33032,N_32303);
or U34967 (N_34967,N_33218,N_32021);
and U34968 (N_34968,N_32399,N_32044);
and U34969 (N_34969,N_33024,N_33154);
nor U34970 (N_34970,N_32149,N_33523);
nor U34971 (N_34971,N_32587,N_33232);
nand U34972 (N_34972,N_33128,N_32601);
xnor U34973 (N_34973,N_32268,N_32538);
and U34974 (N_34974,N_33768,N_32179);
and U34975 (N_34975,N_33618,N_32652);
or U34976 (N_34976,N_32423,N_33760);
nor U34977 (N_34977,N_32566,N_32108);
or U34978 (N_34978,N_33076,N_32540);
or U34979 (N_34979,N_33880,N_32139);
nand U34980 (N_34980,N_32117,N_33669);
and U34981 (N_34981,N_32154,N_33217);
and U34982 (N_34982,N_32304,N_32439);
nand U34983 (N_34983,N_33203,N_32712);
nor U34984 (N_34984,N_32970,N_32766);
nor U34985 (N_34985,N_33995,N_32011);
or U34986 (N_34986,N_32722,N_33383);
nor U34987 (N_34987,N_32410,N_33775);
nand U34988 (N_34988,N_32756,N_33519);
or U34989 (N_34989,N_32380,N_33009);
or U34990 (N_34990,N_32736,N_33215);
nor U34991 (N_34991,N_33237,N_32431);
and U34992 (N_34992,N_33225,N_33260);
nor U34993 (N_34993,N_32102,N_32202);
and U34994 (N_34994,N_32190,N_33702);
nand U34995 (N_34995,N_32526,N_32019);
nor U34996 (N_34996,N_32786,N_33400);
nor U34997 (N_34997,N_32171,N_32296);
nor U34998 (N_34998,N_32678,N_33065);
and U34999 (N_34999,N_32642,N_32729);
or U35000 (N_35000,N_32273,N_32820);
nor U35001 (N_35001,N_32386,N_33063);
nand U35002 (N_35002,N_32406,N_33924);
nand U35003 (N_35003,N_32898,N_33809);
nor U35004 (N_35004,N_33461,N_33515);
or U35005 (N_35005,N_33337,N_33380);
nand U35006 (N_35006,N_33302,N_33362);
and U35007 (N_35007,N_32065,N_32513);
and U35008 (N_35008,N_32818,N_32521);
nor U35009 (N_35009,N_33724,N_33898);
or U35010 (N_35010,N_33659,N_33375);
nand U35011 (N_35011,N_33041,N_33276);
and U35012 (N_35012,N_32818,N_33233);
and U35013 (N_35013,N_33043,N_32588);
nand U35014 (N_35014,N_33679,N_33282);
and U35015 (N_35015,N_33697,N_32525);
and U35016 (N_35016,N_32367,N_32788);
nor U35017 (N_35017,N_32489,N_32713);
nand U35018 (N_35018,N_32763,N_33105);
and U35019 (N_35019,N_33000,N_33692);
or U35020 (N_35020,N_32267,N_33588);
or U35021 (N_35021,N_32071,N_32983);
nand U35022 (N_35022,N_32927,N_32279);
and U35023 (N_35023,N_32408,N_33586);
or U35024 (N_35024,N_33196,N_33414);
nand U35025 (N_35025,N_33152,N_32943);
and U35026 (N_35026,N_33010,N_32793);
and U35027 (N_35027,N_32104,N_32410);
nor U35028 (N_35028,N_33695,N_33698);
or U35029 (N_35029,N_32432,N_33086);
or U35030 (N_35030,N_33685,N_32568);
or U35031 (N_35031,N_32010,N_33634);
and U35032 (N_35032,N_33602,N_32547);
nor U35033 (N_35033,N_33072,N_32498);
and U35034 (N_35034,N_33765,N_33323);
nor U35035 (N_35035,N_33875,N_32767);
and U35036 (N_35036,N_33288,N_32393);
nor U35037 (N_35037,N_32369,N_32389);
and U35038 (N_35038,N_32989,N_33045);
or U35039 (N_35039,N_33643,N_33216);
nor U35040 (N_35040,N_33002,N_33100);
nor U35041 (N_35041,N_32504,N_32469);
nand U35042 (N_35042,N_32475,N_33841);
and U35043 (N_35043,N_32271,N_33237);
or U35044 (N_35044,N_33042,N_33522);
nor U35045 (N_35045,N_32218,N_33354);
and U35046 (N_35046,N_33163,N_33992);
and U35047 (N_35047,N_33637,N_32892);
or U35048 (N_35048,N_32032,N_33893);
nand U35049 (N_35049,N_32298,N_33688);
nand U35050 (N_35050,N_32643,N_32052);
or U35051 (N_35051,N_32988,N_32544);
or U35052 (N_35052,N_33691,N_32285);
nand U35053 (N_35053,N_33304,N_33299);
or U35054 (N_35054,N_33248,N_32694);
nor U35055 (N_35055,N_33048,N_32801);
nand U35056 (N_35056,N_32391,N_33595);
and U35057 (N_35057,N_32981,N_32818);
or U35058 (N_35058,N_33628,N_32881);
and U35059 (N_35059,N_33099,N_32451);
or U35060 (N_35060,N_33259,N_32880);
or U35061 (N_35061,N_33710,N_33926);
nand U35062 (N_35062,N_32515,N_32250);
and U35063 (N_35063,N_32961,N_32210);
nor U35064 (N_35064,N_32947,N_32626);
and U35065 (N_35065,N_32825,N_32894);
nor U35066 (N_35066,N_33239,N_32536);
nor U35067 (N_35067,N_33436,N_33446);
nor U35068 (N_35068,N_32628,N_32261);
nor U35069 (N_35069,N_32907,N_33713);
or U35070 (N_35070,N_32326,N_32318);
nand U35071 (N_35071,N_32766,N_32666);
nand U35072 (N_35072,N_32502,N_33215);
and U35073 (N_35073,N_33693,N_33148);
and U35074 (N_35074,N_33932,N_33107);
nor U35075 (N_35075,N_32786,N_32343);
or U35076 (N_35076,N_32655,N_33308);
and U35077 (N_35077,N_32837,N_32891);
and U35078 (N_35078,N_32576,N_33820);
nand U35079 (N_35079,N_33760,N_33701);
nand U35080 (N_35080,N_32325,N_33478);
nand U35081 (N_35081,N_33474,N_32900);
nand U35082 (N_35082,N_32983,N_32433);
or U35083 (N_35083,N_32024,N_32751);
nand U35084 (N_35084,N_33513,N_33173);
nand U35085 (N_35085,N_32172,N_32762);
and U35086 (N_35086,N_33848,N_33593);
or U35087 (N_35087,N_32850,N_32404);
and U35088 (N_35088,N_33009,N_33050);
or U35089 (N_35089,N_32338,N_32019);
and U35090 (N_35090,N_33705,N_33456);
or U35091 (N_35091,N_33538,N_33474);
or U35092 (N_35092,N_32199,N_32175);
and U35093 (N_35093,N_33683,N_33601);
nand U35094 (N_35094,N_32303,N_33937);
nand U35095 (N_35095,N_33005,N_32654);
or U35096 (N_35096,N_32520,N_32682);
and U35097 (N_35097,N_32818,N_33750);
nand U35098 (N_35098,N_33643,N_33548);
and U35099 (N_35099,N_32297,N_32944);
or U35100 (N_35100,N_33154,N_33438);
or U35101 (N_35101,N_33496,N_32650);
or U35102 (N_35102,N_32397,N_32444);
nor U35103 (N_35103,N_33902,N_33928);
nand U35104 (N_35104,N_32947,N_33096);
and U35105 (N_35105,N_32593,N_32647);
nand U35106 (N_35106,N_32985,N_33648);
nor U35107 (N_35107,N_33616,N_32242);
and U35108 (N_35108,N_32087,N_32309);
or U35109 (N_35109,N_32993,N_32665);
xor U35110 (N_35110,N_32181,N_33877);
nand U35111 (N_35111,N_32194,N_32615);
or U35112 (N_35112,N_32474,N_33193);
or U35113 (N_35113,N_32047,N_33374);
or U35114 (N_35114,N_32590,N_32991);
nor U35115 (N_35115,N_33762,N_33964);
or U35116 (N_35116,N_32028,N_32424);
nor U35117 (N_35117,N_33332,N_32612);
nor U35118 (N_35118,N_32779,N_33342);
nor U35119 (N_35119,N_33522,N_32195);
nor U35120 (N_35120,N_33959,N_33902);
xor U35121 (N_35121,N_32940,N_33627);
or U35122 (N_35122,N_33618,N_32450);
xor U35123 (N_35123,N_32913,N_33054);
and U35124 (N_35124,N_32661,N_32183);
and U35125 (N_35125,N_32077,N_33307);
nor U35126 (N_35126,N_33629,N_32244);
and U35127 (N_35127,N_32455,N_33069);
or U35128 (N_35128,N_33624,N_32418);
nor U35129 (N_35129,N_33379,N_32273);
nor U35130 (N_35130,N_33448,N_33495);
or U35131 (N_35131,N_33295,N_32107);
and U35132 (N_35132,N_32320,N_33982);
and U35133 (N_35133,N_33172,N_33271);
nor U35134 (N_35134,N_32313,N_33581);
nor U35135 (N_35135,N_33655,N_33326);
nand U35136 (N_35136,N_33618,N_32575);
or U35137 (N_35137,N_32714,N_32414);
or U35138 (N_35138,N_33110,N_33632);
and U35139 (N_35139,N_33763,N_33978);
or U35140 (N_35140,N_32837,N_32310);
nor U35141 (N_35141,N_32462,N_32366);
or U35142 (N_35142,N_33329,N_32829);
nor U35143 (N_35143,N_32247,N_33535);
nor U35144 (N_35144,N_32713,N_32644);
nor U35145 (N_35145,N_32287,N_32927);
and U35146 (N_35146,N_33709,N_33121);
or U35147 (N_35147,N_33452,N_33094);
nand U35148 (N_35148,N_32975,N_33798);
nand U35149 (N_35149,N_33683,N_33145);
and U35150 (N_35150,N_32434,N_32017);
nor U35151 (N_35151,N_32257,N_33164);
nor U35152 (N_35152,N_33691,N_33057);
nor U35153 (N_35153,N_32004,N_33838);
nand U35154 (N_35154,N_32444,N_33925);
nor U35155 (N_35155,N_32383,N_32883);
or U35156 (N_35156,N_33848,N_33674);
nor U35157 (N_35157,N_32542,N_32360);
nor U35158 (N_35158,N_32984,N_33824);
and U35159 (N_35159,N_33132,N_33043);
nor U35160 (N_35160,N_32813,N_33383);
nand U35161 (N_35161,N_33422,N_32772);
and U35162 (N_35162,N_32518,N_32839);
nor U35163 (N_35163,N_32236,N_33969);
and U35164 (N_35164,N_32671,N_32138);
nand U35165 (N_35165,N_33036,N_33294);
or U35166 (N_35166,N_32154,N_33126);
nor U35167 (N_35167,N_33643,N_32685);
nor U35168 (N_35168,N_32540,N_33618);
nand U35169 (N_35169,N_33212,N_32969);
nand U35170 (N_35170,N_32608,N_32522);
nor U35171 (N_35171,N_33457,N_33539);
and U35172 (N_35172,N_32428,N_32192);
or U35173 (N_35173,N_32738,N_33758);
nand U35174 (N_35174,N_32983,N_33195);
nor U35175 (N_35175,N_32131,N_32487);
and U35176 (N_35176,N_32406,N_32150);
or U35177 (N_35177,N_32178,N_33131);
nand U35178 (N_35178,N_33615,N_32919);
or U35179 (N_35179,N_32593,N_32550);
nor U35180 (N_35180,N_32140,N_33776);
or U35181 (N_35181,N_33845,N_32580);
nor U35182 (N_35182,N_33924,N_33400);
or U35183 (N_35183,N_32638,N_33604);
nor U35184 (N_35184,N_33220,N_33959);
or U35185 (N_35185,N_32580,N_32365);
and U35186 (N_35186,N_33218,N_32105);
xnor U35187 (N_35187,N_32207,N_32357);
or U35188 (N_35188,N_32991,N_33129);
nor U35189 (N_35189,N_32047,N_33774);
or U35190 (N_35190,N_32237,N_33637);
nand U35191 (N_35191,N_32026,N_32850);
nor U35192 (N_35192,N_33556,N_32642);
or U35193 (N_35193,N_33740,N_33887);
or U35194 (N_35194,N_33773,N_33969);
or U35195 (N_35195,N_33328,N_32553);
or U35196 (N_35196,N_33812,N_32926);
xor U35197 (N_35197,N_33300,N_33557);
nor U35198 (N_35198,N_32138,N_32241);
and U35199 (N_35199,N_33534,N_32699);
or U35200 (N_35200,N_32378,N_32857);
or U35201 (N_35201,N_32671,N_33938);
nand U35202 (N_35202,N_33604,N_32091);
and U35203 (N_35203,N_33849,N_32425);
nor U35204 (N_35204,N_33568,N_32732);
nor U35205 (N_35205,N_33252,N_33369);
and U35206 (N_35206,N_33345,N_33670);
nor U35207 (N_35207,N_33151,N_33984);
nor U35208 (N_35208,N_32427,N_33376);
xor U35209 (N_35209,N_32394,N_32002);
nor U35210 (N_35210,N_32713,N_33403);
nor U35211 (N_35211,N_33706,N_33296);
nor U35212 (N_35212,N_33998,N_32070);
nand U35213 (N_35213,N_33286,N_32852);
or U35214 (N_35214,N_32226,N_33094);
nor U35215 (N_35215,N_33010,N_32248);
or U35216 (N_35216,N_32710,N_32836);
nand U35217 (N_35217,N_33034,N_32190);
and U35218 (N_35218,N_32435,N_32323);
nor U35219 (N_35219,N_32489,N_33723);
nor U35220 (N_35220,N_33580,N_33381);
nand U35221 (N_35221,N_32755,N_33342);
and U35222 (N_35222,N_32722,N_33773);
nor U35223 (N_35223,N_32712,N_32907);
xor U35224 (N_35224,N_32634,N_33640);
or U35225 (N_35225,N_32467,N_33428);
or U35226 (N_35226,N_32528,N_32602);
nand U35227 (N_35227,N_32606,N_32178);
or U35228 (N_35228,N_33298,N_32101);
and U35229 (N_35229,N_33719,N_32417);
and U35230 (N_35230,N_32149,N_32385);
nor U35231 (N_35231,N_33445,N_33702);
nand U35232 (N_35232,N_33494,N_32499);
and U35233 (N_35233,N_33194,N_32687);
nor U35234 (N_35234,N_33570,N_32789);
nor U35235 (N_35235,N_32674,N_32641);
or U35236 (N_35236,N_32724,N_33010);
or U35237 (N_35237,N_33023,N_32898);
and U35238 (N_35238,N_32440,N_33587);
and U35239 (N_35239,N_33319,N_33681);
or U35240 (N_35240,N_33923,N_32056);
and U35241 (N_35241,N_33094,N_33969);
or U35242 (N_35242,N_33258,N_33122);
and U35243 (N_35243,N_32284,N_33121);
nor U35244 (N_35244,N_33371,N_32061);
or U35245 (N_35245,N_33664,N_32474);
nand U35246 (N_35246,N_32781,N_32507);
and U35247 (N_35247,N_32031,N_33515);
nand U35248 (N_35248,N_32631,N_33585);
and U35249 (N_35249,N_33800,N_32525);
nand U35250 (N_35250,N_33009,N_32317);
nand U35251 (N_35251,N_32943,N_32764);
and U35252 (N_35252,N_33202,N_33199);
or U35253 (N_35253,N_32391,N_33906);
nand U35254 (N_35254,N_33397,N_33532);
xor U35255 (N_35255,N_33507,N_33146);
or U35256 (N_35256,N_33278,N_33952);
and U35257 (N_35257,N_33735,N_33004);
or U35258 (N_35258,N_32527,N_33862);
and U35259 (N_35259,N_33209,N_32796);
nor U35260 (N_35260,N_32960,N_32751);
nor U35261 (N_35261,N_33575,N_33019);
or U35262 (N_35262,N_32525,N_33505);
nand U35263 (N_35263,N_33225,N_33896);
nand U35264 (N_35264,N_32265,N_33698);
or U35265 (N_35265,N_32457,N_33433);
or U35266 (N_35266,N_33642,N_32493);
and U35267 (N_35267,N_32561,N_33827);
and U35268 (N_35268,N_33178,N_32751);
nand U35269 (N_35269,N_32965,N_32622);
or U35270 (N_35270,N_32561,N_32835);
nand U35271 (N_35271,N_33792,N_32172);
and U35272 (N_35272,N_32086,N_33736);
nand U35273 (N_35273,N_33027,N_32095);
or U35274 (N_35274,N_32837,N_33026);
or U35275 (N_35275,N_32680,N_33347);
nor U35276 (N_35276,N_33486,N_33835);
nor U35277 (N_35277,N_33384,N_32452);
nor U35278 (N_35278,N_33169,N_33544);
nand U35279 (N_35279,N_32125,N_32846);
xor U35280 (N_35280,N_32254,N_32764);
nand U35281 (N_35281,N_33989,N_33659);
nand U35282 (N_35282,N_32063,N_33766);
nor U35283 (N_35283,N_33927,N_32978);
nor U35284 (N_35284,N_33048,N_32096);
nand U35285 (N_35285,N_32219,N_32109);
nor U35286 (N_35286,N_33727,N_33864);
and U35287 (N_35287,N_32513,N_32531);
nand U35288 (N_35288,N_32012,N_33259);
or U35289 (N_35289,N_33382,N_32831);
or U35290 (N_35290,N_33861,N_33365);
and U35291 (N_35291,N_32731,N_33162);
and U35292 (N_35292,N_33803,N_33813);
xor U35293 (N_35293,N_32206,N_33765);
and U35294 (N_35294,N_32374,N_32311);
and U35295 (N_35295,N_32291,N_33599);
nand U35296 (N_35296,N_32501,N_33457);
and U35297 (N_35297,N_32819,N_33128);
nor U35298 (N_35298,N_33812,N_32780);
and U35299 (N_35299,N_32434,N_32643);
or U35300 (N_35300,N_33571,N_33898);
nor U35301 (N_35301,N_33453,N_33995);
nand U35302 (N_35302,N_33718,N_33430);
and U35303 (N_35303,N_32556,N_33743);
and U35304 (N_35304,N_33832,N_33597);
and U35305 (N_35305,N_32395,N_33010);
and U35306 (N_35306,N_33809,N_32146);
nor U35307 (N_35307,N_33357,N_32062);
nor U35308 (N_35308,N_33952,N_33662);
nor U35309 (N_35309,N_32475,N_32224);
or U35310 (N_35310,N_33242,N_32660);
and U35311 (N_35311,N_32000,N_33756);
nor U35312 (N_35312,N_32254,N_32690);
and U35313 (N_35313,N_33944,N_33109);
nor U35314 (N_35314,N_32012,N_33819);
and U35315 (N_35315,N_32266,N_32617);
nand U35316 (N_35316,N_32687,N_32470);
and U35317 (N_35317,N_32600,N_33041);
or U35318 (N_35318,N_32402,N_33776);
nor U35319 (N_35319,N_32337,N_32502);
or U35320 (N_35320,N_33284,N_32035);
or U35321 (N_35321,N_32283,N_33254);
and U35322 (N_35322,N_33919,N_33987);
nand U35323 (N_35323,N_32903,N_32736);
nor U35324 (N_35324,N_33487,N_32622);
or U35325 (N_35325,N_33894,N_32274);
and U35326 (N_35326,N_33027,N_33070);
nor U35327 (N_35327,N_32119,N_33580);
nor U35328 (N_35328,N_33731,N_32665);
nand U35329 (N_35329,N_33909,N_33532);
and U35330 (N_35330,N_33091,N_32199);
and U35331 (N_35331,N_32383,N_32904);
or U35332 (N_35332,N_32927,N_32214);
and U35333 (N_35333,N_33997,N_33898);
nand U35334 (N_35334,N_32803,N_33362);
and U35335 (N_35335,N_32160,N_33889);
and U35336 (N_35336,N_32937,N_32515);
nand U35337 (N_35337,N_32267,N_33950);
nor U35338 (N_35338,N_32335,N_33436);
nor U35339 (N_35339,N_32110,N_32280);
and U35340 (N_35340,N_32430,N_33711);
nand U35341 (N_35341,N_32072,N_33403);
and U35342 (N_35342,N_32226,N_33136);
or U35343 (N_35343,N_32803,N_33440);
or U35344 (N_35344,N_32804,N_33615);
or U35345 (N_35345,N_32728,N_33493);
or U35346 (N_35346,N_32145,N_33301);
or U35347 (N_35347,N_33184,N_32605);
nor U35348 (N_35348,N_33696,N_33846);
or U35349 (N_35349,N_33456,N_32697);
nor U35350 (N_35350,N_33423,N_32420);
xnor U35351 (N_35351,N_32366,N_33537);
nor U35352 (N_35352,N_32399,N_32161);
nor U35353 (N_35353,N_32499,N_32314);
xnor U35354 (N_35354,N_33083,N_33524);
and U35355 (N_35355,N_32188,N_32202);
and U35356 (N_35356,N_32382,N_33576);
nor U35357 (N_35357,N_33990,N_32235);
and U35358 (N_35358,N_32530,N_32618);
nand U35359 (N_35359,N_32805,N_32751);
or U35360 (N_35360,N_32676,N_32313);
nand U35361 (N_35361,N_32989,N_32370);
or U35362 (N_35362,N_33864,N_32536);
and U35363 (N_35363,N_32754,N_33510);
nor U35364 (N_35364,N_33381,N_33029);
and U35365 (N_35365,N_33431,N_33554);
nand U35366 (N_35366,N_33810,N_33087);
and U35367 (N_35367,N_33297,N_33496);
nand U35368 (N_35368,N_32165,N_32253);
and U35369 (N_35369,N_33397,N_33475);
nor U35370 (N_35370,N_33423,N_33395);
or U35371 (N_35371,N_32556,N_33348);
nor U35372 (N_35372,N_33381,N_33518);
and U35373 (N_35373,N_32433,N_33171);
and U35374 (N_35374,N_33967,N_33610);
and U35375 (N_35375,N_33868,N_33603);
nand U35376 (N_35376,N_33877,N_33484);
nand U35377 (N_35377,N_33962,N_32409);
or U35378 (N_35378,N_32932,N_32129);
xor U35379 (N_35379,N_32933,N_32582);
nand U35380 (N_35380,N_32376,N_32211);
or U35381 (N_35381,N_32878,N_32374);
nor U35382 (N_35382,N_33490,N_33385);
nor U35383 (N_35383,N_33242,N_32303);
nand U35384 (N_35384,N_32482,N_33104);
or U35385 (N_35385,N_33162,N_32096);
or U35386 (N_35386,N_32579,N_32453);
and U35387 (N_35387,N_32136,N_32958);
and U35388 (N_35388,N_33509,N_33522);
and U35389 (N_35389,N_33643,N_32726);
or U35390 (N_35390,N_32010,N_33905);
and U35391 (N_35391,N_32676,N_32548);
nor U35392 (N_35392,N_33584,N_32861);
nand U35393 (N_35393,N_33055,N_33381);
and U35394 (N_35394,N_33428,N_33070);
and U35395 (N_35395,N_33027,N_33507);
or U35396 (N_35396,N_33768,N_32691);
nand U35397 (N_35397,N_33709,N_32814);
xor U35398 (N_35398,N_32021,N_32069);
or U35399 (N_35399,N_33367,N_33979);
xor U35400 (N_35400,N_33812,N_33621);
nor U35401 (N_35401,N_33719,N_32897);
nand U35402 (N_35402,N_33088,N_32045);
xnor U35403 (N_35403,N_32766,N_32816);
or U35404 (N_35404,N_32460,N_32431);
xor U35405 (N_35405,N_32990,N_32560);
nand U35406 (N_35406,N_32278,N_33483);
nor U35407 (N_35407,N_33784,N_33516);
nor U35408 (N_35408,N_32016,N_32827);
and U35409 (N_35409,N_32312,N_33324);
or U35410 (N_35410,N_32269,N_33000);
nor U35411 (N_35411,N_33948,N_32051);
nor U35412 (N_35412,N_33744,N_33470);
or U35413 (N_35413,N_32086,N_33215);
or U35414 (N_35414,N_32787,N_32459);
xor U35415 (N_35415,N_32685,N_32351);
nor U35416 (N_35416,N_32268,N_33327);
and U35417 (N_35417,N_32052,N_33256);
and U35418 (N_35418,N_33288,N_32420);
and U35419 (N_35419,N_33389,N_33586);
xor U35420 (N_35420,N_33908,N_32244);
nor U35421 (N_35421,N_32092,N_33766);
or U35422 (N_35422,N_32844,N_33127);
or U35423 (N_35423,N_32197,N_33203);
or U35424 (N_35424,N_33171,N_32695);
and U35425 (N_35425,N_33895,N_32018);
or U35426 (N_35426,N_32886,N_32274);
nand U35427 (N_35427,N_33713,N_33958);
or U35428 (N_35428,N_32760,N_33671);
and U35429 (N_35429,N_32191,N_33766);
nor U35430 (N_35430,N_33160,N_32982);
and U35431 (N_35431,N_32409,N_32238);
nand U35432 (N_35432,N_32266,N_33506);
or U35433 (N_35433,N_33722,N_32884);
or U35434 (N_35434,N_33842,N_33985);
nor U35435 (N_35435,N_33211,N_33294);
nand U35436 (N_35436,N_33785,N_33007);
and U35437 (N_35437,N_33362,N_32596);
nor U35438 (N_35438,N_32823,N_32676);
xor U35439 (N_35439,N_32709,N_33118);
and U35440 (N_35440,N_33609,N_33870);
nand U35441 (N_35441,N_32533,N_33587);
or U35442 (N_35442,N_32627,N_33873);
nand U35443 (N_35443,N_33073,N_33864);
nand U35444 (N_35444,N_32691,N_33035);
and U35445 (N_35445,N_32142,N_33701);
xnor U35446 (N_35446,N_33488,N_32533);
and U35447 (N_35447,N_33134,N_33368);
nor U35448 (N_35448,N_32558,N_33387);
and U35449 (N_35449,N_32687,N_32679);
nand U35450 (N_35450,N_32622,N_32995);
nor U35451 (N_35451,N_32200,N_32172);
or U35452 (N_35452,N_32712,N_32558);
nand U35453 (N_35453,N_32464,N_32476);
or U35454 (N_35454,N_32735,N_32014);
and U35455 (N_35455,N_33304,N_32454);
nand U35456 (N_35456,N_33449,N_33963);
and U35457 (N_35457,N_32938,N_33691);
and U35458 (N_35458,N_32715,N_33138);
and U35459 (N_35459,N_32557,N_32904);
and U35460 (N_35460,N_32269,N_33745);
nor U35461 (N_35461,N_32416,N_33691);
or U35462 (N_35462,N_33425,N_32619);
nand U35463 (N_35463,N_32005,N_33403);
nand U35464 (N_35464,N_33154,N_32858);
and U35465 (N_35465,N_32579,N_33167);
and U35466 (N_35466,N_33634,N_33175);
and U35467 (N_35467,N_32092,N_33687);
nand U35468 (N_35468,N_32046,N_32069);
nand U35469 (N_35469,N_33095,N_33117);
or U35470 (N_35470,N_32096,N_32143);
nand U35471 (N_35471,N_33487,N_32384);
nand U35472 (N_35472,N_33573,N_32667);
nor U35473 (N_35473,N_32730,N_33450);
and U35474 (N_35474,N_33026,N_32125);
xnor U35475 (N_35475,N_32511,N_32412);
and U35476 (N_35476,N_33152,N_33204);
nor U35477 (N_35477,N_33351,N_33607);
and U35478 (N_35478,N_33968,N_32744);
nor U35479 (N_35479,N_33512,N_33088);
nor U35480 (N_35480,N_32286,N_32152);
and U35481 (N_35481,N_32102,N_32333);
and U35482 (N_35482,N_33651,N_32474);
or U35483 (N_35483,N_32943,N_32095);
nor U35484 (N_35484,N_32765,N_33392);
or U35485 (N_35485,N_32301,N_32398);
nand U35486 (N_35486,N_32877,N_32122);
or U35487 (N_35487,N_33377,N_33110);
and U35488 (N_35488,N_33034,N_33157);
nand U35489 (N_35489,N_33262,N_32633);
or U35490 (N_35490,N_33631,N_33661);
nor U35491 (N_35491,N_33317,N_32697);
nor U35492 (N_35492,N_32670,N_33765);
or U35493 (N_35493,N_32227,N_33583);
and U35494 (N_35494,N_32223,N_32260);
or U35495 (N_35495,N_33912,N_32101);
or U35496 (N_35496,N_33127,N_32342);
and U35497 (N_35497,N_33897,N_32385);
xor U35498 (N_35498,N_33318,N_33458);
and U35499 (N_35499,N_33343,N_33962);
and U35500 (N_35500,N_32432,N_32193);
and U35501 (N_35501,N_33493,N_33951);
and U35502 (N_35502,N_33399,N_33798);
and U35503 (N_35503,N_32549,N_33731);
and U35504 (N_35504,N_33824,N_32163);
nor U35505 (N_35505,N_32952,N_33213);
xnor U35506 (N_35506,N_32442,N_32342);
or U35507 (N_35507,N_33942,N_32618);
or U35508 (N_35508,N_32781,N_33853);
nor U35509 (N_35509,N_33997,N_32049);
nand U35510 (N_35510,N_32840,N_32933);
nor U35511 (N_35511,N_32819,N_33614);
or U35512 (N_35512,N_32745,N_33999);
and U35513 (N_35513,N_32088,N_33598);
nor U35514 (N_35514,N_32181,N_32305);
or U35515 (N_35515,N_33942,N_33813);
or U35516 (N_35516,N_33162,N_32292);
or U35517 (N_35517,N_33065,N_33458);
or U35518 (N_35518,N_33960,N_32279);
or U35519 (N_35519,N_32116,N_32445);
nand U35520 (N_35520,N_32315,N_32235);
and U35521 (N_35521,N_32365,N_33407);
nand U35522 (N_35522,N_33308,N_33408);
and U35523 (N_35523,N_32348,N_33296);
nor U35524 (N_35524,N_32902,N_32973);
nor U35525 (N_35525,N_33991,N_33873);
nor U35526 (N_35526,N_32737,N_32324);
nand U35527 (N_35527,N_33116,N_32100);
or U35528 (N_35528,N_33374,N_33313);
or U35529 (N_35529,N_32521,N_33294);
or U35530 (N_35530,N_32434,N_33886);
or U35531 (N_35531,N_33888,N_33358);
and U35532 (N_35532,N_33658,N_32666);
and U35533 (N_35533,N_32369,N_33623);
nand U35534 (N_35534,N_32458,N_32550);
nand U35535 (N_35535,N_32116,N_32737);
and U35536 (N_35536,N_33248,N_33176);
and U35537 (N_35537,N_33281,N_32514);
nand U35538 (N_35538,N_32311,N_32077);
nor U35539 (N_35539,N_32026,N_32128);
or U35540 (N_35540,N_33786,N_32290);
nand U35541 (N_35541,N_32721,N_33335);
or U35542 (N_35542,N_32733,N_32856);
and U35543 (N_35543,N_32634,N_32315);
or U35544 (N_35544,N_32262,N_32625);
nand U35545 (N_35545,N_33798,N_33108);
nor U35546 (N_35546,N_32491,N_32368);
nand U35547 (N_35547,N_33076,N_32465);
or U35548 (N_35548,N_33928,N_33016);
nand U35549 (N_35549,N_33068,N_32564);
and U35550 (N_35550,N_32142,N_32204);
or U35551 (N_35551,N_32291,N_32363);
and U35552 (N_35552,N_33975,N_33928);
and U35553 (N_35553,N_33911,N_33483);
or U35554 (N_35554,N_32162,N_33398);
and U35555 (N_35555,N_32398,N_33897);
nor U35556 (N_35556,N_33622,N_32423);
nor U35557 (N_35557,N_32778,N_32051);
nand U35558 (N_35558,N_32271,N_33581);
nand U35559 (N_35559,N_32425,N_32139);
nor U35560 (N_35560,N_33781,N_33028);
nor U35561 (N_35561,N_33293,N_32684);
and U35562 (N_35562,N_32485,N_32953);
nor U35563 (N_35563,N_33952,N_32066);
nor U35564 (N_35564,N_33104,N_33360);
nand U35565 (N_35565,N_32958,N_33389);
nor U35566 (N_35566,N_33519,N_32885);
xnor U35567 (N_35567,N_33884,N_33646);
nand U35568 (N_35568,N_32306,N_32422);
nand U35569 (N_35569,N_32569,N_32540);
and U35570 (N_35570,N_32937,N_32912);
nand U35571 (N_35571,N_32644,N_33674);
or U35572 (N_35572,N_33080,N_32933);
or U35573 (N_35573,N_32687,N_33866);
or U35574 (N_35574,N_32090,N_33349);
and U35575 (N_35575,N_32104,N_32587);
and U35576 (N_35576,N_32922,N_33214);
nand U35577 (N_35577,N_33731,N_32968);
xnor U35578 (N_35578,N_33834,N_32182);
nand U35579 (N_35579,N_33887,N_32346);
or U35580 (N_35580,N_32731,N_33143);
nor U35581 (N_35581,N_32835,N_33547);
or U35582 (N_35582,N_33891,N_32622);
and U35583 (N_35583,N_32088,N_33324);
or U35584 (N_35584,N_32648,N_32511);
nand U35585 (N_35585,N_33980,N_33987);
nand U35586 (N_35586,N_32003,N_33135);
and U35587 (N_35587,N_33865,N_33551);
or U35588 (N_35588,N_33055,N_33797);
nor U35589 (N_35589,N_32781,N_32934);
nor U35590 (N_35590,N_32866,N_32694);
nor U35591 (N_35591,N_33209,N_32482);
and U35592 (N_35592,N_33876,N_33968);
nor U35593 (N_35593,N_32366,N_33333);
nor U35594 (N_35594,N_32738,N_33453);
nor U35595 (N_35595,N_33645,N_33681);
nor U35596 (N_35596,N_32169,N_32245);
or U35597 (N_35597,N_33595,N_33028);
and U35598 (N_35598,N_32569,N_32642);
or U35599 (N_35599,N_32804,N_33305);
nand U35600 (N_35600,N_32620,N_33439);
and U35601 (N_35601,N_33171,N_32133);
nand U35602 (N_35602,N_33425,N_33516);
nand U35603 (N_35603,N_33460,N_33288);
or U35604 (N_35604,N_33814,N_32987);
and U35605 (N_35605,N_32608,N_32495);
nor U35606 (N_35606,N_33525,N_33447);
or U35607 (N_35607,N_32664,N_33370);
nor U35608 (N_35608,N_33245,N_32431);
and U35609 (N_35609,N_32083,N_33205);
or U35610 (N_35610,N_32303,N_33670);
or U35611 (N_35611,N_33702,N_32269);
nor U35612 (N_35612,N_33806,N_32339);
nand U35613 (N_35613,N_32832,N_32563);
nand U35614 (N_35614,N_32599,N_32744);
or U35615 (N_35615,N_33940,N_32595);
nor U35616 (N_35616,N_32698,N_33943);
nand U35617 (N_35617,N_32824,N_33568);
or U35618 (N_35618,N_32130,N_32577);
and U35619 (N_35619,N_32663,N_33501);
nand U35620 (N_35620,N_32021,N_33118);
and U35621 (N_35621,N_33052,N_32716);
and U35622 (N_35622,N_33173,N_32027);
nor U35623 (N_35623,N_32771,N_33185);
nand U35624 (N_35624,N_33057,N_33196);
nor U35625 (N_35625,N_33771,N_33612);
or U35626 (N_35626,N_33575,N_32610);
nand U35627 (N_35627,N_33426,N_33935);
nor U35628 (N_35628,N_32398,N_33673);
or U35629 (N_35629,N_32224,N_32547);
or U35630 (N_35630,N_32553,N_33782);
or U35631 (N_35631,N_33205,N_32474);
and U35632 (N_35632,N_32959,N_33994);
or U35633 (N_35633,N_33570,N_33659);
nand U35634 (N_35634,N_32114,N_32013);
or U35635 (N_35635,N_32423,N_32854);
nor U35636 (N_35636,N_33537,N_32280);
and U35637 (N_35637,N_32970,N_32770);
nor U35638 (N_35638,N_32524,N_33927);
nor U35639 (N_35639,N_33551,N_32895);
nand U35640 (N_35640,N_32136,N_33820);
nor U35641 (N_35641,N_32017,N_33285);
nor U35642 (N_35642,N_32586,N_32285);
and U35643 (N_35643,N_32143,N_32026);
or U35644 (N_35644,N_32872,N_33369);
and U35645 (N_35645,N_33523,N_32011);
nand U35646 (N_35646,N_33805,N_33538);
xnor U35647 (N_35647,N_32786,N_33168);
nand U35648 (N_35648,N_32577,N_33613);
and U35649 (N_35649,N_33628,N_32690);
nor U35650 (N_35650,N_33717,N_32421);
and U35651 (N_35651,N_33160,N_32876);
nor U35652 (N_35652,N_33378,N_33826);
and U35653 (N_35653,N_33405,N_33642);
nor U35654 (N_35654,N_32081,N_32382);
nand U35655 (N_35655,N_32235,N_32046);
nand U35656 (N_35656,N_32804,N_33469);
and U35657 (N_35657,N_33911,N_32780);
nand U35658 (N_35658,N_32635,N_32129);
nand U35659 (N_35659,N_33873,N_33892);
or U35660 (N_35660,N_32190,N_32918);
nand U35661 (N_35661,N_32216,N_33217);
or U35662 (N_35662,N_32583,N_32303);
nor U35663 (N_35663,N_33934,N_33776);
nand U35664 (N_35664,N_32995,N_32471);
xnor U35665 (N_35665,N_32011,N_32454);
and U35666 (N_35666,N_33408,N_33787);
and U35667 (N_35667,N_33117,N_32486);
nand U35668 (N_35668,N_33693,N_32276);
and U35669 (N_35669,N_33427,N_32875);
or U35670 (N_35670,N_32758,N_33917);
xnor U35671 (N_35671,N_33924,N_33230);
or U35672 (N_35672,N_33257,N_33230);
nor U35673 (N_35673,N_32656,N_32639);
and U35674 (N_35674,N_32180,N_33480);
and U35675 (N_35675,N_32014,N_32537);
nand U35676 (N_35676,N_32462,N_33483);
and U35677 (N_35677,N_33821,N_32623);
nor U35678 (N_35678,N_33956,N_32004);
nor U35679 (N_35679,N_33250,N_32306);
nand U35680 (N_35680,N_33438,N_32228);
or U35681 (N_35681,N_32216,N_33814);
and U35682 (N_35682,N_32242,N_32354);
nand U35683 (N_35683,N_32678,N_32955);
nand U35684 (N_35684,N_33402,N_32966);
nand U35685 (N_35685,N_33274,N_33724);
and U35686 (N_35686,N_33698,N_33094);
nand U35687 (N_35687,N_32374,N_33273);
nand U35688 (N_35688,N_33336,N_33876);
nor U35689 (N_35689,N_32321,N_33601);
nand U35690 (N_35690,N_32441,N_33058);
or U35691 (N_35691,N_33710,N_32242);
nand U35692 (N_35692,N_33182,N_33744);
nor U35693 (N_35693,N_33610,N_32812);
nor U35694 (N_35694,N_32010,N_32443);
nand U35695 (N_35695,N_32425,N_32030);
and U35696 (N_35696,N_32502,N_32748);
or U35697 (N_35697,N_32704,N_33007);
nand U35698 (N_35698,N_33164,N_33166);
and U35699 (N_35699,N_33814,N_32446);
or U35700 (N_35700,N_33672,N_32751);
nand U35701 (N_35701,N_33133,N_32313);
nand U35702 (N_35702,N_33245,N_32380);
nor U35703 (N_35703,N_33526,N_33500);
nor U35704 (N_35704,N_33289,N_33436);
nand U35705 (N_35705,N_33985,N_32832);
nand U35706 (N_35706,N_32117,N_33011);
and U35707 (N_35707,N_33365,N_33709);
and U35708 (N_35708,N_33384,N_33763);
nor U35709 (N_35709,N_32426,N_32165);
xnor U35710 (N_35710,N_33072,N_33993);
and U35711 (N_35711,N_33837,N_32920);
or U35712 (N_35712,N_32381,N_33513);
nor U35713 (N_35713,N_33427,N_32767);
or U35714 (N_35714,N_33792,N_32020);
or U35715 (N_35715,N_33719,N_32151);
nand U35716 (N_35716,N_32156,N_33891);
nand U35717 (N_35717,N_32652,N_33544);
nand U35718 (N_35718,N_32209,N_32850);
and U35719 (N_35719,N_32300,N_33688);
nor U35720 (N_35720,N_33596,N_32243);
or U35721 (N_35721,N_33775,N_33342);
and U35722 (N_35722,N_33108,N_32850);
nor U35723 (N_35723,N_33971,N_32187);
or U35724 (N_35724,N_33786,N_32195);
nand U35725 (N_35725,N_32868,N_32970);
nor U35726 (N_35726,N_32590,N_32864);
and U35727 (N_35727,N_33578,N_32386);
and U35728 (N_35728,N_32280,N_32689);
and U35729 (N_35729,N_32933,N_32447);
nor U35730 (N_35730,N_32380,N_33597);
or U35731 (N_35731,N_32062,N_33630);
or U35732 (N_35732,N_33848,N_32643);
and U35733 (N_35733,N_33740,N_33143);
nor U35734 (N_35734,N_33966,N_33936);
nor U35735 (N_35735,N_33365,N_33588);
nor U35736 (N_35736,N_32379,N_33799);
and U35737 (N_35737,N_32127,N_33305);
nand U35738 (N_35738,N_33702,N_33140);
or U35739 (N_35739,N_32198,N_32713);
nor U35740 (N_35740,N_33684,N_32784);
and U35741 (N_35741,N_32214,N_33650);
and U35742 (N_35742,N_33885,N_32157);
nand U35743 (N_35743,N_33520,N_33014);
nor U35744 (N_35744,N_32856,N_32396);
nand U35745 (N_35745,N_33139,N_32826);
and U35746 (N_35746,N_33226,N_32433);
nor U35747 (N_35747,N_33513,N_33006);
nor U35748 (N_35748,N_32932,N_33117);
and U35749 (N_35749,N_33614,N_32120);
nand U35750 (N_35750,N_33705,N_33033);
or U35751 (N_35751,N_32818,N_33528);
nor U35752 (N_35752,N_32828,N_33328);
or U35753 (N_35753,N_32498,N_33577);
nor U35754 (N_35754,N_32515,N_32246);
nand U35755 (N_35755,N_33199,N_32196);
and U35756 (N_35756,N_33955,N_32570);
and U35757 (N_35757,N_32286,N_32886);
nand U35758 (N_35758,N_32528,N_32140);
nand U35759 (N_35759,N_32359,N_33821);
or U35760 (N_35760,N_33013,N_32218);
and U35761 (N_35761,N_32917,N_33053);
or U35762 (N_35762,N_32593,N_32076);
and U35763 (N_35763,N_33689,N_33047);
and U35764 (N_35764,N_32392,N_32926);
nand U35765 (N_35765,N_32819,N_32373);
nand U35766 (N_35766,N_33388,N_32595);
nand U35767 (N_35767,N_32250,N_33778);
nor U35768 (N_35768,N_33013,N_33268);
nor U35769 (N_35769,N_32722,N_33866);
nand U35770 (N_35770,N_32147,N_32831);
and U35771 (N_35771,N_32528,N_33973);
or U35772 (N_35772,N_32706,N_33746);
or U35773 (N_35773,N_33184,N_33409);
nor U35774 (N_35774,N_33484,N_33058);
and U35775 (N_35775,N_33599,N_33800);
and U35776 (N_35776,N_33450,N_33683);
and U35777 (N_35777,N_32783,N_32020);
nand U35778 (N_35778,N_32986,N_33582);
or U35779 (N_35779,N_33152,N_33406);
xnor U35780 (N_35780,N_32381,N_33567);
or U35781 (N_35781,N_32079,N_32321);
or U35782 (N_35782,N_33981,N_32732);
or U35783 (N_35783,N_32952,N_33074);
and U35784 (N_35784,N_32230,N_33907);
nor U35785 (N_35785,N_33250,N_32596);
and U35786 (N_35786,N_33287,N_32752);
and U35787 (N_35787,N_32440,N_32048);
or U35788 (N_35788,N_33942,N_33472);
nor U35789 (N_35789,N_32317,N_33260);
and U35790 (N_35790,N_33305,N_33333);
or U35791 (N_35791,N_33241,N_32810);
or U35792 (N_35792,N_33809,N_32797);
nor U35793 (N_35793,N_33088,N_32773);
and U35794 (N_35794,N_32689,N_32598);
or U35795 (N_35795,N_33828,N_32758);
nand U35796 (N_35796,N_32682,N_33936);
or U35797 (N_35797,N_32546,N_33795);
or U35798 (N_35798,N_32752,N_32234);
nor U35799 (N_35799,N_33362,N_33360);
nor U35800 (N_35800,N_32130,N_32877);
nand U35801 (N_35801,N_32649,N_33511);
and U35802 (N_35802,N_32968,N_32812);
or U35803 (N_35803,N_33948,N_33254);
nor U35804 (N_35804,N_33996,N_32250);
or U35805 (N_35805,N_32482,N_33190);
or U35806 (N_35806,N_33767,N_33368);
and U35807 (N_35807,N_32658,N_32633);
nor U35808 (N_35808,N_32559,N_32911);
or U35809 (N_35809,N_33970,N_33791);
and U35810 (N_35810,N_33810,N_32268);
nor U35811 (N_35811,N_33363,N_33240);
nand U35812 (N_35812,N_32828,N_32267);
nand U35813 (N_35813,N_33681,N_32382);
or U35814 (N_35814,N_33291,N_33814);
nor U35815 (N_35815,N_32412,N_32249);
nand U35816 (N_35816,N_32037,N_33028);
xnor U35817 (N_35817,N_32714,N_32638);
and U35818 (N_35818,N_32307,N_32753);
nor U35819 (N_35819,N_32477,N_32448);
nor U35820 (N_35820,N_32225,N_32814);
nand U35821 (N_35821,N_33371,N_33694);
nand U35822 (N_35822,N_33017,N_32776);
nor U35823 (N_35823,N_32783,N_33132);
nor U35824 (N_35824,N_32413,N_32044);
or U35825 (N_35825,N_32775,N_33750);
or U35826 (N_35826,N_33885,N_33014);
nor U35827 (N_35827,N_32716,N_32934);
or U35828 (N_35828,N_33071,N_32718);
nor U35829 (N_35829,N_33869,N_32459);
and U35830 (N_35830,N_33826,N_32264);
nor U35831 (N_35831,N_33680,N_33477);
and U35832 (N_35832,N_33597,N_32107);
or U35833 (N_35833,N_32974,N_33643);
nor U35834 (N_35834,N_32507,N_32903);
nand U35835 (N_35835,N_32705,N_32898);
nand U35836 (N_35836,N_33641,N_32633);
and U35837 (N_35837,N_33592,N_32901);
or U35838 (N_35838,N_32592,N_32654);
or U35839 (N_35839,N_32356,N_32280);
and U35840 (N_35840,N_32936,N_32308);
nor U35841 (N_35841,N_33230,N_33311);
and U35842 (N_35842,N_32640,N_33620);
or U35843 (N_35843,N_33227,N_32063);
nor U35844 (N_35844,N_33128,N_33549);
nand U35845 (N_35845,N_32195,N_32172);
or U35846 (N_35846,N_32006,N_33830);
or U35847 (N_35847,N_32236,N_32640);
or U35848 (N_35848,N_33535,N_32515);
nor U35849 (N_35849,N_33505,N_32898);
and U35850 (N_35850,N_32409,N_33793);
nand U35851 (N_35851,N_32728,N_32102);
nand U35852 (N_35852,N_32407,N_33032);
or U35853 (N_35853,N_32439,N_33013);
nor U35854 (N_35854,N_33972,N_32431);
nand U35855 (N_35855,N_32114,N_33959);
or U35856 (N_35856,N_33451,N_33457);
and U35857 (N_35857,N_33624,N_32458);
or U35858 (N_35858,N_33783,N_32376);
nor U35859 (N_35859,N_32071,N_33166);
or U35860 (N_35860,N_32995,N_33226);
or U35861 (N_35861,N_33403,N_32243);
nand U35862 (N_35862,N_32049,N_32719);
nand U35863 (N_35863,N_32030,N_33489);
nor U35864 (N_35864,N_32731,N_33605);
and U35865 (N_35865,N_33213,N_32271);
and U35866 (N_35866,N_32772,N_33523);
nand U35867 (N_35867,N_32331,N_32953);
nor U35868 (N_35868,N_32706,N_32976);
nand U35869 (N_35869,N_33363,N_32431);
nor U35870 (N_35870,N_32554,N_32852);
nor U35871 (N_35871,N_33421,N_32666);
or U35872 (N_35872,N_32628,N_33685);
nor U35873 (N_35873,N_32586,N_32082);
and U35874 (N_35874,N_33774,N_32982);
nand U35875 (N_35875,N_32082,N_32216);
nand U35876 (N_35876,N_32632,N_33711);
and U35877 (N_35877,N_33381,N_32133);
nand U35878 (N_35878,N_32195,N_32166);
nor U35879 (N_35879,N_32298,N_32565);
and U35880 (N_35880,N_33012,N_33172);
nor U35881 (N_35881,N_33856,N_33803);
and U35882 (N_35882,N_32773,N_32738);
and U35883 (N_35883,N_33817,N_32747);
or U35884 (N_35884,N_33925,N_33865);
nand U35885 (N_35885,N_32956,N_32694);
and U35886 (N_35886,N_32030,N_33686);
or U35887 (N_35887,N_32983,N_32088);
and U35888 (N_35888,N_33380,N_32820);
nand U35889 (N_35889,N_33088,N_33176);
and U35890 (N_35890,N_33414,N_33784);
and U35891 (N_35891,N_33110,N_33205);
and U35892 (N_35892,N_33165,N_33981);
nand U35893 (N_35893,N_32546,N_32794);
xor U35894 (N_35894,N_33446,N_33553);
and U35895 (N_35895,N_32578,N_32828);
nand U35896 (N_35896,N_32575,N_32131);
xor U35897 (N_35897,N_32667,N_33506);
or U35898 (N_35898,N_32459,N_32600);
and U35899 (N_35899,N_32175,N_32846);
and U35900 (N_35900,N_33844,N_33893);
or U35901 (N_35901,N_33964,N_32626);
nand U35902 (N_35902,N_32024,N_33823);
and U35903 (N_35903,N_33143,N_32198);
and U35904 (N_35904,N_33362,N_33601);
nand U35905 (N_35905,N_32683,N_33917);
xnor U35906 (N_35906,N_33791,N_32868);
xor U35907 (N_35907,N_32467,N_33655);
and U35908 (N_35908,N_33754,N_32159);
or U35909 (N_35909,N_32813,N_33014);
and U35910 (N_35910,N_32340,N_33973);
nor U35911 (N_35911,N_33799,N_32352);
and U35912 (N_35912,N_32649,N_33896);
nand U35913 (N_35913,N_33234,N_32638);
nand U35914 (N_35914,N_33814,N_33642);
nand U35915 (N_35915,N_33667,N_32890);
and U35916 (N_35916,N_33602,N_33829);
or U35917 (N_35917,N_33654,N_32298);
nand U35918 (N_35918,N_33609,N_32378);
or U35919 (N_35919,N_32597,N_32275);
or U35920 (N_35920,N_33239,N_33514);
nand U35921 (N_35921,N_32302,N_33971);
nor U35922 (N_35922,N_32239,N_33489);
nand U35923 (N_35923,N_32379,N_33164);
and U35924 (N_35924,N_33648,N_33668);
xnor U35925 (N_35925,N_33089,N_32887);
nand U35926 (N_35926,N_32880,N_32199);
nor U35927 (N_35927,N_32308,N_32479);
and U35928 (N_35928,N_33007,N_32495);
nor U35929 (N_35929,N_32037,N_33795);
nand U35930 (N_35930,N_32248,N_32538);
nand U35931 (N_35931,N_33970,N_33102);
and U35932 (N_35932,N_33863,N_33017);
nand U35933 (N_35933,N_32969,N_32477);
and U35934 (N_35934,N_32852,N_32613);
nand U35935 (N_35935,N_32356,N_32558);
or U35936 (N_35936,N_33793,N_32422);
and U35937 (N_35937,N_33479,N_32824);
and U35938 (N_35938,N_33238,N_33657);
and U35939 (N_35939,N_32698,N_32927);
or U35940 (N_35940,N_33598,N_33776);
nor U35941 (N_35941,N_33384,N_32437);
nor U35942 (N_35942,N_33444,N_33852);
and U35943 (N_35943,N_33463,N_32249);
nor U35944 (N_35944,N_32504,N_33355);
and U35945 (N_35945,N_32511,N_32495);
or U35946 (N_35946,N_33778,N_32539);
nor U35947 (N_35947,N_33906,N_33904);
and U35948 (N_35948,N_32809,N_33273);
nand U35949 (N_35949,N_33605,N_33378);
nand U35950 (N_35950,N_32364,N_33199);
nor U35951 (N_35951,N_32225,N_32995);
nor U35952 (N_35952,N_32323,N_33551);
nor U35953 (N_35953,N_33492,N_33139);
nor U35954 (N_35954,N_32032,N_32634);
and U35955 (N_35955,N_33205,N_32033);
nand U35956 (N_35956,N_32512,N_33581);
or U35957 (N_35957,N_32784,N_32855);
nand U35958 (N_35958,N_33338,N_33783);
or U35959 (N_35959,N_32676,N_33892);
and U35960 (N_35960,N_33747,N_32855);
and U35961 (N_35961,N_32848,N_33140);
nand U35962 (N_35962,N_32292,N_32510);
or U35963 (N_35963,N_33071,N_32975);
and U35964 (N_35964,N_33015,N_32641);
or U35965 (N_35965,N_33787,N_33562);
nand U35966 (N_35966,N_32858,N_33360);
and U35967 (N_35967,N_33170,N_33590);
nor U35968 (N_35968,N_33011,N_33576);
nor U35969 (N_35969,N_33240,N_33123);
or U35970 (N_35970,N_32841,N_33311);
nor U35971 (N_35971,N_32941,N_33479);
nand U35972 (N_35972,N_32495,N_32699);
nand U35973 (N_35973,N_32209,N_33725);
or U35974 (N_35974,N_33373,N_33756);
and U35975 (N_35975,N_33679,N_33704);
xnor U35976 (N_35976,N_33135,N_33236);
nor U35977 (N_35977,N_33897,N_33388);
or U35978 (N_35978,N_33052,N_33223);
nand U35979 (N_35979,N_32113,N_33452);
or U35980 (N_35980,N_32178,N_32633);
nor U35981 (N_35981,N_33087,N_32035);
and U35982 (N_35982,N_33309,N_33300);
nand U35983 (N_35983,N_32725,N_32581);
and U35984 (N_35984,N_32108,N_33663);
or U35985 (N_35985,N_33694,N_32329);
and U35986 (N_35986,N_33449,N_33856);
nand U35987 (N_35987,N_33482,N_32590);
nand U35988 (N_35988,N_33511,N_32976);
or U35989 (N_35989,N_33847,N_32912);
xor U35990 (N_35990,N_32362,N_33660);
nand U35991 (N_35991,N_32239,N_32606);
or U35992 (N_35992,N_32065,N_32601);
nor U35993 (N_35993,N_33263,N_32174);
xor U35994 (N_35994,N_33928,N_32734);
nor U35995 (N_35995,N_32560,N_33230);
or U35996 (N_35996,N_33657,N_33000);
and U35997 (N_35997,N_32604,N_33633);
or U35998 (N_35998,N_32657,N_32015);
nand U35999 (N_35999,N_32745,N_32852);
or U36000 (N_36000,N_35204,N_34731);
or U36001 (N_36001,N_35038,N_34658);
and U36002 (N_36002,N_34093,N_35149);
nand U36003 (N_36003,N_35803,N_34025);
xor U36004 (N_36004,N_35647,N_35042);
and U36005 (N_36005,N_35605,N_34035);
nand U36006 (N_36006,N_34006,N_34080);
or U36007 (N_36007,N_34183,N_34337);
nand U36008 (N_36008,N_35078,N_35503);
and U36009 (N_36009,N_34194,N_35944);
and U36010 (N_36010,N_34451,N_34668);
nand U36011 (N_36011,N_35613,N_35339);
and U36012 (N_36012,N_35229,N_35903);
nand U36013 (N_36013,N_35491,N_35215);
nand U36014 (N_36014,N_35840,N_35112);
nor U36015 (N_36015,N_35353,N_35775);
nand U36016 (N_36016,N_34889,N_34079);
nor U36017 (N_36017,N_35879,N_34551);
nor U36018 (N_36018,N_35674,N_34657);
or U36019 (N_36019,N_34594,N_35547);
and U36020 (N_36020,N_34980,N_35401);
and U36021 (N_36021,N_34029,N_35625);
or U36022 (N_36022,N_35332,N_35010);
xor U36023 (N_36023,N_35441,N_34933);
nand U36024 (N_36024,N_35980,N_34923);
nand U36025 (N_36025,N_34009,N_35584);
nor U36026 (N_36026,N_34008,N_34457);
nand U36027 (N_36027,N_34444,N_34972);
nand U36028 (N_36028,N_34791,N_35863);
and U36029 (N_36029,N_35284,N_35272);
nor U36030 (N_36030,N_35178,N_35247);
or U36031 (N_36031,N_34452,N_34569);
nor U36032 (N_36032,N_35323,N_35915);
nor U36033 (N_36033,N_35464,N_35075);
or U36034 (N_36034,N_34467,N_34638);
xnor U36035 (N_36035,N_34756,N_34415);
xor U36036 (N_36036,N_35521,N_35514);
or U36037 (N_36037,N_35437,N_35259);
or U36038 (N_36038,N_35160,N_34475);
or U36039 (N_36039,N_34691,N_34802);
nand U36040 (N_36040,N_35921,N_35893);
nand U36041 (N_36041,N_34436,N_35127);
nor U36042 (N_36042,N_35134,N_35319);
and U36043 (N_36043,N_35322,N_34727);
nor U36044 (N_36044,N_34087,N_34185);
nor U36045 (N_36045,N_34096,N_34995);
nor U36046 (N_36046,N_34970,N_34606);
or U36047 (N_36047,N_35657,N_34860);
or U36048 (N_36048,N_35493,N_35922);
or U36049 (N_36049,N_34201,N_34599);
nand U36050 (N_36050,N_34649,N_35615);
nand U36051 (N_36051,N_34967,N_34073);
nand U36052 (N_36052,N_35796,N_35816);
nand U36053 (N_36053,N_35282,N_34772);
xor U36054 (N_36054,N_35458,N_35295);
and U36055 (N_36055,N_34281,N_35756);
and U36056 (N_36056,N_35805,N_34639);
and U36057 (N_36057,N_35419,N_34764);
and U36058 (N_36058,N_35270,N_35748);
or U36059 (N_36059,N_35049,N_34537);
nand U36060 (N_36060,N_34636,N_35618);
nand U36061 (N_36061,N_34883,N_34242);
nand U36062 (N_36062,N_34767,N_34582);
xnor U36063 (N_36063,N_34674,N_34495);
nor U36064 (N_36064,N_34246,N_34076);
or U36065 (N_36065,N_34485,N_34953);
and U36066 (N_36066,N_35609,N_35036);
nor U36067 (N_36067,N_35450,N_34442);
or U36068 (N_36068,N_34760,N_35594);
and U36069 (N_36069,N_35106,N_35210);
or U36070 (N_36070,N_34884,N_34729);
and U36071 (N_36071,N_34155,N_34742);
nand U36072 (N_36072,N_34497,N_34385);
xor U36073 (N_36073,N_35769,N_35743);
nand U36074 (N_36074,N_35465,N_34612);
xnor U36075 (N_36075,N_35166,N_34125);
nand U36076 (N_36076,N_35612,N_34045);
nand U36077 (N_36077,N_35875,N_34360);
nand U36078 (N_36078,N_34411,N_35601);
nand U36079 (N_36079,N_34382,N_35812);
nor U36080 (N_36080,N_34295,N_34748);
nor U36081 (N_36081,N_34605,N_34325);
and U36082 (N_36082,N_34186,N_34648);
and U36083 (N_36083,N_35826,N_34629);
nand U36084 (N_36084,N_35188,N_35781);
or U36085 (N_36085,N_34854,N_34869);
or U36086 (N_36086,N_34061,N_35302);
or U36087 (N_36087,N_34850,N_35637);
or U36088 (N_36088,N_35161,N_35024);
and U36089 (N_36089,N_35981,N_34853);
nand U36090 (N_36090,N_34321,N_34031);
nand U36091 (N_36091,N_35498,N_35155);
nor U36092 (N_36092,N_35783,N_34575);
and U36093 (N_36093,N_35933,N_35039);
or U36094 (N_36094,N_35866,N_35556);
and U36095 (N_36095,N_34768,N_34574);
and U36096 (N_36096,N_35212,N_35789);
nor U36097 (N_36097,N_35658,N_35909);
or U36098 (N_36098,N_34241,N_34617);
nand U36099 (N_36099,N_34377,N_35835);
or U36100 (N_36100,N_34122,N_35201);
nor U36101 (N_36101,N_35645,N_35545);
nor U36102 (N_36102,N_35105,N_35554);
nor U36103 (N_36103,N_34924,N_35844);
and U36104 (N_36104,N_34642,N_34829);
nand U36105 (N_36105,N_34341,N_35941);
nor U36106 (N_36106,N_35788,N_35813);
and U36107 (N_36107,N_35916,N_34766);
nor U36108 (N_36108,N_34465,N_35052);
and U36109 (N_36109,N_34941,N_35433);
and U36110 (N_36110,N_35258,N_34663);
or U36111 (N_36111,N_34358,N_34693);
nand U36112 (N_36112,N_35607,N_35472);
nor U36113 (N_36113,N_35290,N_34365);
nor U36114 (N_36114,N_35145,N_35018);
nor U36115 (N_36115,N_35585,N_34499);
and U36116 (N_36116,N_35119,N_34438);
nor U36117 (N_36117,N_34506,N_34815);
nand U36118 (N_36118,N_35695,N_35752);
nand U36119 (N_36119,N_34956,N_35574);
nand U36120 (N_36120,N_35340,N_34895);
nor U36121 (N_36121,N_34110,N_34302);
xor U36122 (N_36122,N_35726,N_35715);
nand U36123 (N_36123,N_35670,N_34395);
nand U36124 (N_36124,N_34667,N_35292);
or U36125 (N_36125,N_34255,N_35638);
nand U36126 (N_36126,N_35118,N_35997);
and U36127 (N_36127,N_35734,N_35596);
nor U36128 (N_36128,N_35942,N_35561);
and U36129 (N_36129,N_34330,N_35621);
nand U36130 (N_36130,N_35565,N_34305);
nor U36131 (N_36131,N_35978,N_35964);
and U36132 (N_36132,N_35142,N_34193);
and U36133 (N_36133,N_34548,N_35376);
nand U36134 (N_36134,N_34214,N_35685);
or U36135 (N_36135,N_34244,N_34710);
nand U36136 (N_36136,N_35619,N_34545);
nor U36137 (N_36137,N_34877,N_34412);
nor U36138 (N_36138,N_35883,N_35740);
nand U36139 (N_36139,N_34616,N_34907);
xnor U36140 (N_36140,N_35492,N_35373);
nand U36141 (N_36141,N_34238,N_35254);
or U36142 (N_36142,N_35095,N_35298);
and U36143 (N_36143,N_35570,N_35308);
nor U36144 (N_36144,N_35370,N_34866);
nor U36145 (N_36145,N_35717,N_34051);
nor U36146 (N_36146,N_34205,N_34744);
and U36147 (N_36147,N_35508,N_35611);
and U36148 (N_36148,N_34173,N_34461);
nor U36149 (N_36149,N_35988,N_34531);
or U36150 (N_36150,N_34425,N_34987);
or U36151 (N_36151,N_35531,N_34963);
nand U36152 (N_36152,N_34882,N_34282);
nor U36153 (N_36153,N_35214,N_34627);
or U36154 (N_36154,N_35818,N_35971);
and U36155 (N_36155,N_34213,N_34916);
nand U36156 (N_36156,N_34095,N_34868);
nor U36157 (N_36157,N_35417,N_34216);
and U36158 (N_36158,N_35086,N_35414);
nand U36159 (N_36159,N_34900,N_35771);
or U36160 (N_36160,N_34954,N_34397);
nand U36161 (N_36161,N_35369,N_34345);
or U36162 (N_36162,N_34774,N_35228);
and U36163 (N_36163,N_35143,N_35736);
nor U36164 (N_36164,N_34157,N_34101);
or U36165 (N_36165,N_34023,N_35725);
nand U36166 (N_36166,N_35663,N_34903);
nand U36167 (N_36167,N_34749,N_35868);
nor U36168 (N_36168,N_34979,N_34986);
and U36169 (N_36169,N_35887,N_34273);
and U36170 (N_36170,N_34287,N_34417);
and U36171 (N_36171,N_34588,N_34849);
and U36172 (N_36172,N_34743,N_35713);
or U36173 (N_36173,N_34044,N_35173);
nor U36174 (N_36174,N_35354,N_34250);
and U36175 (N_36175,N_34277,N_35787);
nand U36176 (N_36176,N_34738,N_35268);
nand U36177 (N_36177,N_34806,N_35548);
or U36178 (N_36178,N_34978,N_35785);
nor U36179 (N_36179,N_35129,N_35871);
and U36180 (N_36180,N_34248,N_34820);
and U36181 (N_36181,N_35589,N_35686);
nand U36182 (N_36182,N_34804,N_34554);
nor U36183 (N_36183,N_34245,N_35286);
or U36184 (N_36184,N_34099,N_35749);
nor U36185 (N_36185,N_34137,N_35069);
or U36186 (N_36186,N_34156,N_35230);
and U36187 (N_36187,N_34151,N_35700);
nor U36188 (N_36188,N_35714,N_34602);
or U36189 (N_36189,N_35660,N_34069);
and U36190 (N_36190,N_35635,N_34447);
nor U36191 (N_36191,N_34192,N_34421);
or U36192 (N_36192,N_35123,N_35632);
or U36193 (N_36193,N_35930,N_35819);
nand U36194 (N_36194,N_34346,N_34105);
xnor U36195 (N_36195,N_35375,N_34879);
or U36196 (N_36196,N_35053,N_34567);
or U36197 (N_36197,N_34446,N_34056);
nor U36198 (N_36198,N_35934,N_35085);
and U36199 (N_36199,N_35938,N_34822);
and U36200 (N_36200,N_35037,N_34041);
nand U36201 (N_36201,N_35480,N_35851);
nor U36202 (N_36202,N_34068,N_34565);
nor U36203 (N_36203,N_34534,N_34641);
nor U36204 (N_36204,N_34827,N_34852);
and U36205 (N_36205,N_34206,N_35539);
and U36206 (N_36206,N_34013,N_35343);
or U36207 (N_36207,N_34807,N_34635);
or U36208 (N_36208,N_34038,N_34074);
nand U36209 (N_36209,N_34089,N_34433);
nand U36210 (N_36210,N_34510,N_35683);
or U36211 (N_36211,N_35524,N_34480);
nor U36212 (N_36212,N_34643,N_34523);
nand U36213 (N_36213,N_35378,N_35328);
or U36214 (N_36214,N_34354,N_35359);
nor U36215 (N_36215,N_35677,N_35022);
or U36216 (N_36216,N_34278,N_35336);
nor U36217 (N_36217,N_35741,N_35081);
and U36218 (N_36218,N_34779,N_35864);
or U36219 (N_36219,N_34138,N_34665);
or U36220 (N_36220,N_34524,N_35071);
nor U36221 (N_36221,N_34019,N_35870);
or U36222 (N_36222,N_35445,N_35048);
or U36223 (N_36223,N_34917,N_35967);
nor U36224 (N_36224,N_34855,N_35159);
or U36225 (N_36225,N_35620,N_34857);
nor U36226 (N_36226,N_34703,N_35285);
or U36227 (N_36227,N_35202,N_35832);
or U36228 (N_36228,N_35907,N_34060);
and U36229 (N_36229,N_34655,N_34459);
or U36230 (N_36230,N_34132,N_35935);
nand U36231 (N_36231,N_34613,N_34563);
nand U36232 (N_36232,N_34831,N_35416);
nand U36233 (N_36233,N_35553,N_35684);
nor U36234 (N_36234,N_35076,N_35730);
or U36235 (N_36235,N_34513,N_35368);
or U36236 (N_36236,N_34198,N_34316);
nand U36237 (N_36237,N_35627,N_34429);
and U36238 (N_36238,N_35299,N_34178);
nand U36239 (N_36239,N_35872,N_35062);
nor U36240 (N_36240,N_34946,N_35569);
and U36241 (N_36241,N_35329,N_34862);
or U36242 (N_36242,N_34723,N_35953);
nand U36243 (N_36243,N_35402,N_35301);
nand U36244 (N_36244,N_35562,N_35482);
nor U36245 (N_36245,N_34239,N_35182);
nor U36246 (N_36246,N_35823,N_34410);
or U36247 (N_36247,N_34552,N_35027);
nor U36248 (N_36248,N_34107,N_35096);
or U36249 (N_36249,N_34601,N_35798);
nand U36250 (N_36250,N_35946,N_35624);
nand U36251 (N_36251,N_34596,N_35455);
and U36252 (N_36252,N_35474,N_34189);
or U36253 (N_36253,N_34833,N_34842);
nor U36254 (N_36254,N_34741,N_35197);
and U36255 (N_36255,N_34539,N_34573);
nand U36256 (N_36256,N_34702,N_35296);
and U36257 (N_36257,N_34149,N_35444);
xnor U36258 (N_36258,N_34684,N_34579);
and U36259 (N_36259,N_34293,N_35264);
or U36260 (N_36260,N_35802,N_34726);
and U36261 (N_36261,N_34362,N_34307);
nor U36262 (N_36262,N_35170,N_34159);
or U36263 (N_36263,N_34886,N_34422);
nand U36264 (N_36264,N_34704,N_35033);
and U36265 (N_36265,N_35488,N_35345);
and U36266 (N_36266,N_35747,N_35911);
nand U36267 (N_36267,N_35528,N_34870);
nand U36268 (N_36268,N_34054,N_35512);
or U36269 (N_36269,N_34376,N_34102);
or U36270 (N_36270,N_35557,N_34897);
nand U36271 (N_36271,N_35654,N_34765);
or U36272 (N_36272,N_34816,N_35846);
nand U36273 (N_36273,N_34578,N_35702);
xor U36274 (N_36274,N_34324,N_35446);
or U36275 (N_36275,N_34486,N_34356);
and U36276 (N_36276,N_34477,N_35003);
and U36277 (N_36277,N_34810,N_34180);
or U36278 (N_36278,N_35643,N_34263);
and U36279 (N_36279,N_34709,N_34072);
and U36280 (N_36280,N_34319,N_34094);
or U36281 (N_36281,N_34697,N_35195);
nor U36282 (N_36282,N_35385,N_34176);
nor U36283 (N_36283,N_34310,N_34725);
nor U36284 (N_36284,N_34182,N_34835);
and U36285 (N_36285,N_35337,N_34762);
and U36286 (N_36286,N_35550,N_35833);
or U36287 (N_36287,N_35243,N_35733);
or U36288 (N_36288,N_34312,N_35055);
or U36289 (N_36289,N_34463,N_35758);
nand U36290 (N_36290,N_34919,N_34874);
and U36291 (N_36291,N_35460,N_35927);
nor U36292 (N_36292,N_34040,N_35710);
or U36293 (N_36293,N_35732,N_34247);
and U36294 (N_36294,N_35396,N_34611);
xnor U36295 (N_36295,N_34859,N_34127);
or U36296 (N_36296,N_35600,N_34532);
nor U36297 (N_36297,N_34003,N_35720);
xnor U36298 (N_36298,N_35454,N_34814);
nor U36299 (N_36299,N_34018,N_34067);
and U36300 (N_36300,N_35382,N_35573);
and U36301 (N_36301,N_35659,N_35257);
or U36302 (N_36302,N_35806,N_34934);
nand U36303 (N_36303,N_34808,N_34677);
and U36304 (N_36304,N_34024,N_34938);
nand U36305 (N_36305,N_35393,N_35102);
nor U36306 (N_36306,N_35360,N_35755);
nor U36307 (N_36307,N_35588,N_35463);
nor U36308 (N_36308,N_35772,N_34290);
or U36309 (N_36309,N_34496,N_35793);
nor U36310 (N_36310,N_34650,N_35593);
or U36311 (N_36311,N_34334,N_34374);
and U36312 (N_36312,N_35226,N_35761);
and U36313 (N_36313,N_35869,N_34572);
nor U36314 (N_36314,N_35438,N_35529);
and U36315 (N_36315,N_34195,N_34169);
and U36316 (N_36316,N_34930,N_35716);
nor U36317 (N_36317,N_35398,N_34839);
and U36318 (N_36318,N_35092,N_35485);
nand U36319 (N_36319,N_34587,N_35209);
nor U36320 (N_36320,N_35435,N_34370);
nand U36321 (N_36321,N_35822,N_34114);
or U36322 (N_36322,N_34838,N_35141);
nor U36323 (N_36323,N_35325,N_34873);
and U36324 (N_36324,N_34431,N_34147);
or U36325 (N_36325,N_35121,N_35742);
and U36326 (N_36326,N_35672,N_34867);
and U36327 (N_36327,N_35221,N_35252);
nand U36328 (N_36328,N_35928,N_35087);
or U36329 (N_36329,N_34174,N_34123);
and U36330 (N_36330,N_34799,N_34906);
or U36331 (N_36331,N_34696,N_34542);
nand U36332 (N_36332,N_35361,N_35430);
or U36333 (N_36333,N_34610,N_34407);
nand U36334 (N_36334,N_35206,N_35116);
or U36335 (N_36335,N_35533,N_34538);
nor U36336 (N_36336,N_35384,N_34931);
and U36337 (N_36337,N_34637,N_34179);
or U36338 (N_36338,N_35587,N_35551);
and U36339 (N_36339,N_35825,N_35418);
nor U36340 (N_36340,N_34170,N_35431);
nand U36341 (N_36341,N_35744,N_35780);
and U36342 (N_36342,N_34286,N_34750);
or U36343 (N_36343,N_34973,N_35954);
and U36344 (N_36344,N_34140,N_34490);
or U36345 (N_36345,N_35633,N_34948);
nor U36346 (N_36346,N_34158,N_34303);
or U36347 (N_36347,N_34472,N_34518);
nand U36348 (N_36348,N_35233,N_35504);
nor U36349 (N_36349,N_35023,N_34115);
nor U36350 (N_36350,N_34392,N_35706);
xor U36351 (N_36351,N_35698,N_35745);
or U36352 (N_36352,N_34876,N_35249);
nor U36353 (N_36353,N_34434,N_34878);
nand U36354 (N_36354,N_34199,N_35932);
nand U36355 (N_36355,N_34985,N_34962);
and U36356 (N_36356,N_34836,N_35137);
xor U36357 (N_36357,N_35469,N_35366);
and U36358 (N_36358,N_34759,N_35991);
and U36359 (N_36359,N_35172,N_35673);
nor U36360 (N_36360,N_34445,N_34329);
nor U36361 (N_36361,N_34798,N_35380);
or U36362 (N_36362,N_35865,N_35114);
nor U36363 (N_36363,N_34133,N_34769);
nand U36364 (N_36364,N_34022,N_34468);
or U36365 (N_36365,N_34577,N_35649);
and U36366 (N_36366,N_34350,N_34432);
and U36367 (N_36367,N_34010,N_34543);
or U36368 (N_36368,N_35951,N_34326);
or U36369 (N_36369,N_35581,N_34165);
nor U36370 (N_36370,N_35404,N_35267);
xnor U36371 (N_36371,N_35977,N_34484);
nand U36372 (N_36372,N_34163,N_35111);
and U36373 (N_36373,N_35896,N_34514);
xnor U36374 (N_36374,N_35693,N_34771);
and U36375 (N_36375,N_34315,N_34592);
or U36376 (N_36376,N_35501,N_34982);
nor U36377 (N_36377,N_34783,N_35509);
and U36378 (N_36378,N_35566,N_34556);
nand U36379 (N_36379,N_35827,N_35409);
nor U36380 (N_36380,N_35136,N_35350);
nand U36381 (N_36381,N_34652,N_35175);
nor U36382 (N_36382,N_35255,N_35006);
and U36383 (N_36383,N_35276,N_34983);
nand U36384 (N_36384,N_35293,N_35186);
or U36385 (N_36385,N_35814,N_35540);
nor U36386 (N_36386,N_34904,N_34521);
and U36387 (N_36387,N_35956,N_34653);
and U36388 (N_36388,N_35009,N_35479);
nand U36389 (N_36389,N_34943,N_34586);
nor U36390 (N_36390,N_34818,N_34795);
nand U36391 (N_36391,N_34160,N_35115);
nand U36392 (N_36392,N_34634,N_34671);
nor U36393 (N_36393,N_35211,N_34251);
or U36394 (N_36394,N_34228,N_35807);
or U36395 (N_36395,N_34015,N_34188);
nand U36396 (N_36396,N_35029,N_35728);
nor U36397 (N_36397,N_35975,N_34803);
or U36398 (N_36398,N_34647,N_35628);
or U36399 (N_36399,N_35217,N_34166);
nor U36400 (N_36400,N_35845,N_34793);
and U36401 (N_36401,N_34926,N_34646);
nor U36402 (N_36402,N_34851,N_35013);
nand U36403 (N_36403,N_35348,N_35424);
nor U36404 (N_36404,N_34387,N_34098);
nand U36405 (N_36405,N_35496,N_34112);
and U36406 (N_36406,N_35181,N_34753);
nand U36407 (N_36407,N_34896,N_34581);
nand U36408 (N_36408,N_34722,N_35965);
nor U36409 (N_36409,N_34585,N_35989);
nor U36410 (N_36410,N_35321,N_35709);
or U36411 (N_36411,N_34448,N_34212);
or U36412 (N_36412,N_34498,N_35905);
and U36413 (N_36413,N_34136,N_35442);
and U36414 (N_36414,N_34314,N_34848);
nor U36415 (N_36415,N_35892,N_35064);
nor U36416 (N_36416,N_35044,N_34812);
nand U36417 (N_36417,N_35880,N_35108);
and U36418 (N_36418,N_34714,N_34687);
and U36419 (N_36419,N_34757,N_34561);
nand U36420 (N_36420,N_35766,N_34466);
or U36421 (N_36421,N_34085,N_34530);
nor U36422 (N_36422,N_35364,N_34719);
and U36423 (N_36423,N_34952,N_35180);
and U36424 (N_36424,N_35138,N_34527);
and U36425 (N_36425,N_35598,N_35760);
nand U36426 (N_36426,N_34033,N_35560);
nand U36427 (N_36427,N_34625,N_35487);
and U36428 (N_36428,N_34210,N_35357);
nand U36429 (N_36429,N_34735,N_34824);
and U36430 (N_36430,N_35976,N_35680);
or U36431 (N_36431,N_35821,N_34776);
and U36432 (N_36432,N_34819,N_35241);
nand U36433 (N_36433,N_34327,N_34357);
nor U36434 (N_36434,N_34624,N_35811);
and U36435 (N_36435,N_35139,N_34082);
or U36436 (N_36436,N_34676,N_34823);
nand U36437 (N_36437,N_35028,N_34562);
or U36438 (N_36438,N_34628,N_34232);
nand U36439 (N_36439,N_34109,N_35912);
and U36440 (N_36440,N_35263,N_34294);
and U36441 (N_36441,N_34969,N_35874);
xor U36442 (N_36442,N_35030,N_35784);
nand U36443 (N_36443,N_35603,N_35650);
or U36444 (N_36444,N_35451,N_35171);
nor U36445 (N_36445,N_35985,N_34454);
and U36446 (N_36446,N_35314,N_35676);
or U36447 (N_36447,N_34965,N_35901);
or U36448 (N_36448,N_35099,N_34226);
nor U36449 (N_36449,N_35043,N_34291);
nand U36450 (N_36450,N_35697,N_35996);
nor U36451 (N_36451,N_35926,N_35169);
nor U36452 (N_36452,N_34120,N_34809);
or U36453 (N_36453,N_34017,N_35889);
or U36454 (N_36454,N_35133,N_35117);
or U36455 (N_36455,N_34999,N_34483);
nand U36456 (N_36456,N_34966,N_35379);
and U36457 (N_36457,N_35722,N_34491);
nor U36458 (N_36458,N_34243,N_34414);
and U36459 (N_36459,N_35958,N_35894);
nor U36460 (N_36460,N_35089,N_35227);
nand U36461 (N_36461,N_35347,N_35669);
and U36462 (N_36462,N_35571,N_35391);
nand U36463 (N_36463,N_34104,N_34283);
nor U36464 (N_36464,N_35829,N_35305);
nand U36465 (N_36465,N_34424,N_35436);
or U36466 (N_36466,N_34737,N_35130);
nor U36467 (N_36467,N_34732,N_34191);
or U36468 (N_36468,N_34394,N_35523);
and U36469 (N_36469,N_35936,N_35536);
xor U36470 (N_36470,N_35694,N_35797);
or U36471 (N_36471,N_35499,N_34508);
and U36472 (N_36472,N_34223,N_35843);
or U36473 (N_36473,N_35520,N_35342);
and U36474 (N_36474,N_34111,N_35313);
or U36475 (N_36475,N_35622,N_34754);
or U36476 (N_36476,N_34675,N_35407);
nand U36477 (N_36477,N_35131,N_35895);
or U36478 (N_36478,N_34172,N_35877);
nand U36479 (N_36479,N_34801,N_34746);
nor U36480 (N_36480,N_35176,N_35897);
and U36481 (N_36481,N_34730,N_34705);
nor U36482 (N_36482,N_35261,N_35757);
and U36483 (N_36483,N_34364,N_34998);
or U36484 (N_36484,N_34736,N_34046);
and U36485 (N_36485,N_35815,N_34813);
nor U36486 (N_36486,N_35516,N_35655);
or U36487 (N_36487,N_35665,N_34369);
nor U36488 (N_36488,N_35394,N_35567);
nand U36489 (N_36489,N_35790,N_35886);
nand U36490 (N_36490,N_34240,N_35058);
or U36491 (N_36491,N_34042,N_35462);
xor U36492 (N_36492,N_35098,N_34991);
or U36493 (N_36493,N_35962,N_34168);
nor U36494 (N_36494,N_34280,N_34474);
or U36495 (N_36495,N_35552,N_34817);
nand U36496 (N_36496,N_34786,N_34515);
nor U36497 (N_36497,N_34439,N_35692);
nor U36498 (N_36498,N_35193,N_35671);
xor U36499 (N_36499,N_34048,N_35679);
xnor U36500 (N_36500,N_34547,N_34351);
nand U36501 (N_36501,N_35311,N_35225);
nor U36502 (N_36502,N_34773,N_34419);
and U36503 (N_36503,N_34418,N_34235);
nor U36504 (N_36504,N_35083,N_35770);
or U36505 (N_36505,N_34898,N_35519);
nand U36506 (N_36506,N_35885,N_35990);
nand U36507 (N_36507,N_34141,N_35687);
nand U36508 (N_36508,N_35324,N_34755);
nand U36509 (N_36509,N_34279,N_34215);
or U36510 (N_36510,N_35253,N_35795);
nand U36511 (N_36511,N_34134,N_35801);
nand U36512 (N_36512,N_34590,N_35021);
nand U36513 (N_36513,N_34620,N_35998);
or U36514 (N_36514,N_35580,N_35271);
and U36515 (N_36515,N_34332,N_34028);
and U36516 (N_36516,N_35383,N_35185);
nor U36517 (N_36517,N_35399,N_35973);
or U36518 (N_36518,N_35238,N_34945);
nand U36519 (N_36519,N_35681,N_35856);
or U36520 (N_36520,N_34306,N_35250);
or U36521 (N_36521,N_34175,N_35489);
and U36522 (N_36522,N_34057,N_34470);
nor U36523 (N_36523,N_35810,N_34037);
and U36524 (N_36524,N_34236,N_35050);
nand U36525 (N_36525,N_34284,N_34259);
or U36526 (N_36526,N_35381,N_34950);
or U36527 (N_36527,N_34914,N_34402);
nor U36528 (N_36528,N_35294,N_35273);
nor U36529 (N_36529,N_35363,N_35082);
and U36530 (N_36530,N_35984,N_34656);
and U36531 (N_36531,N_35477,N_34167);
nand U36532 (N_36532,N_34153,N_34086);
and U36533 (N_36533,N_34366,N_34489);
or U36534 (N_36534,N_34386,N_34841);
nor U36535 (N_36535,N_35199,N_35371);
nor U36536 (N_36536,N_34631,N_34942);
nor U36537 (N_36537,N_35242,N_35599);
or U36538 (N_36538,N_34522,N_35992);
nor U36539 (N_36539,N_35779,N_34651);
or U36540 (N_36540,N_34758,N_34113);
and U36541 (N_36541,N_34707,N_34745);
nand U36542 (N_36542,N_34724,N_35857);
nor U36543 (N_36543,N_35739,N_34777);
nand U36544 (N_36544,N_35128,N_34437);
nand U36545 (N_36545,N_34885,N_35318);
nor U36546 (N_36546,N_34274,N_35280);
or U36547 (N_36547,N_34081,N_35326);
and U36548 (N_36548,N_35104,N_35881);
nand U36549 (N_36549,N_35120,N_35675);
or U36550 (N_36550,N_35920,N_35067);
nor U36551 (N_36551,N_34555,N_35586);
nor U36552 (N_36552,N_34309,N_35522);
or U36553 (N_36553,N_34271,N_34164);
and U36554 (N_36554,N_34996,N_34034);
nor U36555 (N_36555,N_35461,N_34682);
and U36556 (N_36556,N_35662,N_35235);
or U36557 (N_36557,N_34420,N_35853);
or U36558 (N_36558,N_34275,N_34712);
nor U36559 (N_36559,N_34152,N_35534);
and U36560 (N_36560,N_34959,N_34103);
nor U36561 (N_36561,N_35011,N_35945);
nor U36562 (N_36562,N_34875,N_34609);
and U36563 (N_36563,N_34359,N_34598);
or U36564 (N_36564,N_35982,N_34352);
nor U36565 (N_36565,N_35731,N_34001);
or U36566 (N_36566,N_35088,N_35473);
nand U36567 (N_36567,N_35244,N_35764);
nor U36568 (N_36568,N_34272,N_35415);
nand U36569 (N_36569,N_34660,N_35817);
nor U36570 (N_36570,N_35542,N_34011);
nor U36571 (N_36571,N_35355,N_34416);
or U36572 (N_36572,N_35091,N_35158);
and U36573 (N_36573,N_34219,N_35765);
or U36574 (N_36574,N_35955,N_35447);
nor U36575 (N_36575,N_34378,N_34221);
and U36576 (N_36576,N_35005,N_35961);
nand U36577 (N_36577,N_34821,N_34560);
nand U36578 (N_36578,N_34528,N_35616);
nand U36579 (N_36579,N_34256,N_35351);
or U36580 (N_36580,N_35162,N_34752);
nor U36581 (N_36581,N_35074,N_34622);
and U36582 (N_36582,N_35763,N_34790);
or U36583 (N_36583,N_35950,N_34899);
nor U36584 (N_36584,N_34728,N_35506);
or U36585 (N_36585,N_34456,N_35315);
or U36586 (N_36586,N_34462,N_35782);
nand U36587 (N_36587,N_35794,N_35146);
nand U36588 (N_36588,N_34559,N_34958);
nor U36589 (N_36589,N_34372,N_35275);
nand U36590 (N_36590,N_35056,N_34672);
or U36591 (N_36591,N_35168,N_34615);
xnor U36592 (N_36592,N_34640,N_34891);
nor U36593 (N_36593,N_34940,N_34285);
nor U36594 (N_36594,N_35093,N_35668);
or U36595 (N_36595,N_34328,N_35014);
nor U36596 (N_36596,N_34217,N_34830);
nor U36597 (N_36597,N_35606,N_34100);
nor U36598 (N_36598,N_35704,N_34005);
nor U36599 (N_36599,N_34910,N_34162);
nand U36600 (N_36600,N_34347,N_35511);
and U36601 (N_36601,N_34526,N_35878);
or U36602 (N_36602,N_35841,N_35831);
or U36603 (N_36603,N_35837,N_34388);
or U36604 (N_36604,N_34570,N_35919);
nor U36605 (N_36605,N_34131,N_35426);
and U36606 (N_36606,N_35641,N_34220);
nand U36607 (N_36607,N_35957,N_34264);
or U36608 (N_36608,N_35631,N_35959);
nand U36609 (N_36609,N_35830,N_34473);
and U36610 (N_36610,N_34678,N_34144);
nand U36611 (N_36611,N_35839,N_35289);
nand U36612 (N_36612,N_34449,N_35644);
and U36613 (N_36613,N_34503,N_34391);
nor U36614 (N_36614,N_35636,N_35163);
and U36615 (N_36615,N_34501,N_35150);
nor U36616 (N_36616,N_35626,N_35634);
and U36617 (N_36617,N_34920,N_34614);
nand U36618 (N_36618,N_34664,N_34846);
nand U36619 (N_36619,N_34988,N_35705);
or U36620 (N_36620,N_34384,N_35327);
nand U36621 (N_36621,N_35617,N_35940);
and U36622 (N_36622,N_34597,N_34856);
nor U36623 (N_36623,N_35054,N_34805);
nor U36624 (N_36624,N_34960,N_34670);
nand U36625 (N_36625,N_35427,N_34488);
and U36626 (N_36626,N_35664,N_35778);
and U36627 (N_36627,N_34070,N_34692);
and U36628 (N_36628,N_35943,N_34064);
or U36629 (N_36629,N_35667,N_34322);
xor U36630 (N_36630,N_34065,N_34355);
or U36631 (N_36631,N_35408,N_34872);
nor U36632 (N_36632,N_35144,N_34481);
or U36633 (N_36633,N_34225,N_34683);
and U36634 (N_36634,N_34413,N_35867);
nand U36635 (N_36635,N_34039,N_35213);
and U36636 (N_36636,N_35576,N_35012);
and U36637 (N_36637,N_35245,N_34700);
or U36638 (N_36638,N_35555,N_34139);
nor U36639 (N_36639,N_35890,N_34440);
nand U36640 (N_36640,N_35240,N_35344);
or U36641 (N_36641,N_34130,N_35691);
and U36642 (N_36642,N_35678,N_35914);
and U36643 (N_36643,N_35300,N_35563);
and U36644 (N_36644,N_34789,N_35507);
nor U36645 (N_36645,N_35157,N_34997);
or U36646 (N_36646,N_35167,N_34108);
and U36647 (N_36647,N_34049,N_34124);
or U36648 (N_36648,N_35754,N_35020);
or U36649 (N_36649,N_34455,N_35929);
and U36650 (N_36650,N_35510,N_34881);
nor U36651 (N_36651,N_34955,N_35639);
nor U36652 (N_36652,N_35820,N_35604);
nor U36653 (N_36653,N_35187,N_34858);
and U36654 (N_36654,N_34536,N_34181);
or U36655 (N_36655,N_34721,N_35952);
nor U36656 (N_36656,N_35986,N_35177);
and U36657 (N_36657,N_34032,N_34549);
nand U36658 (N_36658,N_35884,N_35222);
nand U36659 (N_36659,N_35232,N_34020);
or U36660 (N_36660,N_35579,N_35410);
and U36661 (N_36661,N_35412,N_34014);
or U36662 (N_36662,N_34557,N_34428);
and U36663 (N_36663,N_35640,N_35541);
or U36664 (N_36664,N_34233,N_35559);
xor U36665 (N_36665,N_34381,N_35443);
or U36666 (N_36666,N_35931,N_34084);
and U36667 (N_36667,N_34502,N_34645);
nor U36668 (N_36668,N_35219,N_35727);
or U36669 (N_36669,N_34993,N_35040);
or U36670 (N_36670,N_35791,N_34336);
and U36671 (N_36671,N_34349,N_34929);
nand U36672 (N_36672,N_35824,N_34012);
and U36673 (N_36673,N_35804,N_35148);
or U36674 (N_36674,N_35947,N_34298);
nor U36675 (N_36675,N_34679,N_35471);
nor U36676 (N_36676,N_34913,N_34843);
nor U36677 (N_36677,N_35800,N_35902);
nand U36678 (N_36678,N_35854,N_35004);
or U36679 (N_36679,N_35246,N_35882);
nand U36680 (N_36680,N_35194,N_35910);
nand U36681 (N_36681,N_35428,N_34398);
and U36682 (N_36682,N_35850,N_35046);
nand U36683 (N_36683,N_34864,N_34389);
or U36684 (N_36684,N_35939,N_35505);
nor U36685 (N_36685,N_35400,N_34450);
nand U36686 (N_36686,N_34200,N_35610);
nor U36687 (N_36687,N_35476,N_34021);
and U36688 (N_36688,N_35490,N_34276);
nor U36689 (N_36689,N_35809,N_34202);
nand U36690 (N_36690,N_34690,N_34761);
and U36691 (N_36691,N_35608,N_35937);
nor U36692 (N_36692,N_35218,N_35838);
nor U36693 (N_36693,N_35045,N_35239);
nand U36694 (N_36694,N_35723,N_34142);
nand U36695 (N_36695,N_35031,N_35032);
nor U36696 (N_36696,N_34342,N_35432);
or U36697 (N_36697,N_34659,N_34792);
nor U36698 (N_36698,N_35140,N_34308);
nand U36699 (N_36699,N_34826,N_35497);
nor U36700 (N_36700,N_35223,N_34908);
nor U36701 (N_36701,N_35060,N_34626);
nand U36702 (N_36702,N_34004,N_35690);
nand U36703 (N_36703,N_35746,N_34289);
nor U36704 (N_36704,N_35101,N_34911);
or U36705 (N_36705,N_35494,N_34894);
or U36706 (N_36706,N_34409,N_35558);
and U36707 (N_36707,N_34593,N_34145);
nor U36708 (N_36708,N_35356,N_35568);
and U36709 (N_36709,N_35448,N_34564);
or U36710 (N_36710,N_35572,N_35122);
nor U36711 (N_36711,N_34837,N_35502);
and U36712 (N_36712,N_34845,N_34313);
or U36713 (N_36713,N_35135,N_35459);
nor U36714 (N_36714,N_35303,N_35968);
and U36715 (N_36715,N_34267,N_35651);
and U36716 (N_36716,N_35196,N_35515);
nand U36717 (N_36717,N_35721,N_34661);
nor U36718 (N_36718,N_34740,N_35834);
nor U36719 (N_36719,N_34494,N_35309);
or U36720 (N_36720,N_34915,N_35365);
nor U36721 (N_36721,N_34546,N_35277);
or U36722 (N_36722,N_34964,N_34961);
and U36723 (N_36723,N_35236,N_34343);
nand U36724 (N_36724,N_35154,N_35530);
or U36725 (N_36725,N_34090,N_34126);
nor U36726 (N_36726,N_34148,N_35453);
nand U36727 (N_36727,N_34681,N_34237);
and U36728 (N_36728,N_34512,N_35452);
and U36729 (N_36729,N_35422,N_34887);
or U36730 (N_36730,N_34788,N_34971);
nand U36731 (N_36731,N_35481,N_34493);
or U36732 (N_36732,N_35109,N_34618);
and U36733 (N_36733,N_35179,N_35307);
and U36734 (N_36734,N_35652,N_35972);
or U36735 (N_36735,N_35966,N_35467);
nor U36736 (N_36736,N_34253,N_34224);
and U36737 (N_36737,N_34734,N_35097);
and U36738 (N_36738,N_34204,N_34083);
nand U36739 (N_36739,N_34331,N_35549);
and U36740 (N_36740,N_34000,N_35025);
nand U36741 (N_36741,N_35993,N_35792);
and U36742 (N_36742,N_34595,N_34994);
and U36743 (N_36743,N_34834,N_35405);
or U36744 (N_36744,N_34427,N_34589);
and U36745 (N_36745,N_35513,N_34371);
and U36746 (N_36746,N_34751,N_34763);
nand U36747 (N_36747,N_34566,N_34519);
or U36748 (N_36748,N_35917,N_34423);
and U36749 (N_36749,N_35035,N_34901);
nor U36750 (N_36750,N_35304,N_34252);
nor U36751 (N_36751,N_35701,N_35388);
and U36752 (N_36752,N_34404,N_35189);
nor U36753 (N_36753,N_35047,N_35900);
nor U36754 (N_36754,N_34258,N_35094);
and U36755 (N_36755,N_35429,N_34464);
and U36756 (N_36756,N_34460,N_34135);
nor U36757 (N_36757,N_35862,N_35165);
nand U36758 (N_36758,N_35386,N_34058);
or U36759 (N_36759,N_34507,N_34825);
nor U36760 (N_36760,N_35015,N_35421);
nand U36761 (N_36761,N_35265,N_34249);
nand U36762 (N_36762,N_34301,N_35281);
nor U36763 (N_36763,N_35836,N_35666);
and U36764 (N_36764,N_34405,N_35256);
xor U36765 (N_36765,N_34520,N_35279);
and U36766 (N_36766,N_34207,N_35699);
nor U36767 (N_36767,N_34844,N_34654);
nand U36768 (N_36768,N_35411,N_34928);
and U36769 (N_36769,N_34701,N_35125);
nand U36770 (N_36770,N_34348,N_35016);
nand U36771 (N_36771,N_35362,N_35475);
nor U36772 (N_36772,N_34043,N_34533);
or U36773 (N_36773,N_34863,N_34685);
or U36774 (N_36774,N_35274,N_34426);
nand U36775 (N_36775,N_34716,N_34553);
nand U36776 (N_36776,N_34190,N_35312);
nor U36777 (N_36777,N_34482,N_34540);
or U36778 (N_36778,N_35406,N_35248);
or U36779 (N_36779,N_35440,N_35526);
nand U36780 (N_36780,N_35689,N_34568);
nor U36781 (N_36781,N_34689,N_34871);
nor U36782 (N_36782,N_35859,N_34893);
and U36783 (N_36783,N_35577,N_35861);
nor U36784 (N_36784,N_34211,N_35072);
or U36785 (N_36785,N_35316,N_35059);
and U36786 (N_36786,N_35646,N_34990);
nand U36787 (N_36787,N_35041,N_35237);
nor U36788 (N_36788,N_34161,N_35113);
xor U36789 (N_36789,N_34607,N_35532);
nand U36790 (N_36790,N_34266,N_35392);
and U36791 (N_36791,N_35735,N_35317);
nor U36792 (N_36792,N_34782,N_34951);
nand U36793 (N_36793,N_35466,N_35283);
xor U36794 (N_36794,N_35266,N_34016);
or U36795 (N_36795,N_35629,N_35648);
or U36796 (N_36796,N_35719,N_34623);
nor U36797 (N_36797,N_35151,N_35208);
nand U36798 (N_36798,N_34968,N_34981);
nor U36799 (N_36799,N_35750,N_34698);
nor U36800 (N_36800,N_34396,N_34828);
and U36801 (N_36801,N_35434,N_35852);
or U36802 (N_36802,N_34739,N_34984);
nand U36803 (N_36803,N_35974,N_35183);
and U36804 (N_36804,N_35860,N_35395);
nand U36805 (N_36805,N_35582,N_34695);
nand U36806 (N_36806,N_34230,N_34430);
xnor U36807 (N_36807,N_34921,N_34128);
nor U36808 (N_36808,N_34323,N_34688);
nand U36809 (N_36809,N_34975,N_34304);
and U36810 (N_36810,N_35906,N_35200);
nand U36811 (N_36811,N_35153,N_34666);
and U36812 (N_36812,N_34787,N_34403);
nor U36813 (N_36813,N_34576,N_34909);
or U36814 (N_36814,N_35703,N_35191);
nand U36815 (N_36815,N_34458,N_35876);
and U36816 (N_36816,N_34129,N_34406);
and U36817 (N_36817,N_35583,N_34935);
nand U36818 (N_36818,N_34912,N_35203);
nand U36819 (N_36819,N_34435,N_34106);
nor U36820 (N_36820,N_34121,N_35751);
xor U36821 (N_36821,N_34662,N_35858);
nand U36822 (N_36822,N_34865,N_35899);
nand U36823 (N_36823,N_34055,N_35500);
and U36824 (N_36824,N_35711,N_34150);
or U36825 (N_36825,N_35358,N_34375);
nor U36826 (N_36826,N_35948,N_34932);
nor U36827 (N_36827,N_35124,N_35126);
and U36828 (N_36828,N_34861,N_35855);
or U36829 (N_36829,N_34936,N_34361);
and U36830 (N_36830,N_34775,N_35949);
nor U36831 (N_36831,N_34443,N_35306);
and U36832 (N_36832,N_35103,N_34383);
xnor U36833 (N_36833,N_34300,N_34603);
or U36834 (N_36834,N_35898,N_34203);
and U36835 (N_36835,N_35190,N_35080);
and U36836 (N_36836,N_35423,N_34053);
nor U36837 (N_36837,N_34977,N_34091);
nand U36838 (N_36838,N_35543,N_35591);
and U36839 (N_36839,N_35595,N_34600);
nand U36840 (N_36840,N_35000,N_34373);
nor U36841 (N_36841,N_34143,N_35590);
or U36842 (N_36842,N_34118,N_35963);
or U36843 (N_36843,N_34400,N_34504);
or U36844 (N_36844,N_35420,N_34888);
and U36845 (N_36845,N_35525,N_35320);
or U36846 (N_36846,N_35891,N_35578);
or U36847 (N_36847,N_34957,N_34062);
nand U36848 (N_36848,N_34644,N_34030);
or U36849 (N_36849,N_35372,N_34007);
nand U36850 (N_36850,N_34608,N_35073);
nor U36851 (N_36851,N_34989,N_35969);
nand U36852 (N_36852,N_34720,N_35849);
nor U36853 (N_36853,N_34925,N_34680);
or U36854 (N_36854,N_35808,N_34379);
nor U36855 (N_36855,N_35331,N_35575);
nand U36856 (N_36856,N_35970,N_35708);
nand U36857 (N_36857,N_35068,N_35449);
and U36858 (N_36858,N_34401,N_35753);
and U36859 (N_36859,N_35278,N_34318);
or U36860 (N_36860,N_35224,N_34939);
and U36861 (N_36861,N_35335,N_35367);
or U36862 (N_36862,N_35537,N_34368);
nand U36863 (N_36863,N_35738,N_34847);
nor U36864 (N_36864,N_34116,N_35026);
or U36865 (N_36865,N_34262,N_34227);
or U36866 (N_36866,N_34399,N_35110);
and U36867 (N_36867,N_35925,N_34077);
or U36868 (N_36868,N_34363,N_35960);
and U36869 (N_36869,N_35260,N_35377);
and U36870 (N_36870,N_34478,N_34517);
and U36871 (N_36871,N_35220,N_34949);
and U36872 (N_36872,N_35333,N_35084);
and U36873 (N_36873,N_34171,N_34840);
and U36874 (N_36874,N_34367,N_35777);
nand U36875 (N_36875,N_34353,N_34619);
nand U36876 (N_36876,N_35486,N_34441);
nand U36877 (N_36877,N_34927,N_35478);
and U36878 (N_36878,N_35718,N_35767);
nand U36879 (N_36879,N_35425,N_34380);
nor U36880 (N_36880,N_34583,N_34558);
nor U36881 (N_36881,N_34785,N_35288);
nand U36882 (N_36882,N_35291,N_35174);
nand U36883 (N_36883,N_35538,N_34265);
xor U36884 (N_36884,N_34922,N_34339);
nand U36885 (N_36885,N_35799,N_34027);
nand U36886 (N_36886,N_35908,N_35712);
or U36887 (N_36887,N_34296,N_35070);
nor U36888 (N_36888,N_35983,N_35352);
and U36889 (N_36889,N_35051,N_35107);
or U36890 (N_36890,N_34317,N_34393);
or U36891 (N_36891,N_35592,N_35737);
or U36892 (N_36892,N_34892,N_35413);
nor U36893 (N_36893,N_35987,N_34747);
nand U36894 (N_36894,N_35999,N_34880);
nand U36895 (N_36895,N_35535,N_35602);
nand U36896 (N_36896,N_34097,N_34918);
or U36897 (N_36897,N_34604,N_34784);
and U36898 (N_36898,N_34794,N_34937);
nor U36899 (N_36899,N_35696,N_35231);
xnor U36900 (N_36900,N_35913,N_34699);
nor U36901 (N_36901,N_34047,N_35192);
nor U36902 (N_36902,N_34119,N_35762);
or U36903 (N_36903,N_35847,N_34509);
nor U36904 (N_36904,N_34630,N_34571);
nand U36905 (N_36905,N_34584,N_34669);
or U36906 (N_36906,N_35688,N_35234);
or U36907 (N_36907,N_34633,N_34992);
and U36908 (N_36908,N_35544,N_34075);
nand U36909 (N_36909,N_35527,N_34686);
or U36910 (N_36910,N_35828,N_35653);
nand U36911 (N_36911,N_34026,N_35468);
nand U36912 (N_36912,N_34706,N_34390);
or U36913 (N_36913,N_34036,N_34800);
nand U36914 (N_36914,N_34500,N_34187);
nand U36915 (N_36915,N_34254,N_35063);
nor U36916 (N_36916,N_35403,N_34059);
and U36917 (N_36917,N_34832,N_34197);
or U36918 (N_36918,N_35918,N_35707);
or U36919 (N_36919,N_34591,N_35184);
and U36920 (N_36920,N_34580,N_35630);
nand U36921 (N_36921,N_35390,N_34694);
or U36922 (N_36922,N_35147,N_35842);
and U36923 (N_36923,N_34154,N_34525);
and U36924 (N_36924,N_35786,N_35456);
or U36925 (N_36925,N_34516,N_34338);
and U36926 (N_36926,N_35152,N_35297);
nor U36927 (N_36927,N_35439,N_34292);
or U36928 (N_36928,N_35682,N_34002);
nor U36929 (N_36929,N_34469,N_34270);
nand U36930 (N_36930,N_34718,N_34268);
nor U36931 (N_36931,N_35205,N_35034);
nor U36932 (N_36932,N_35397,N_34050);
nand U36933 (N_36933,N_35614,N_34320);
or U36934 (N_36934,N_34479,N_34770);
nand U36935 (N_36935,N_35729,N_34218);
nor U36936 (N_36936,N_34476,N_34529);
nor U36937 (N_36937,N_34088,N_35776);
nor U36938 (N_36938,N_34052,N_34544);
nand U36939 (N_36939,N_35389,N_34890);
nor U36940 (N_36940,N_35251,N_35546);
or U36941 (N_36941,N_35346,N_35774);
nand U36942 (N_36942,N_35994,N_35207);
nand U36943 (N_36943,N_34117,N_35262);
and U36944 (N_36944,N_35597,N_35995);
nand U36945 (N_36945,N_34711,N_35017);
and U36946 (N_36946,N_34177,N_34078);
nor U36947 (N_36947,N_35066,N_35090);
nor U36948 (N_36948,N_34261,N_34717);
nor U36949 (N_36949,N_35768,N_34453);
or U36950 (N_36950,N_34492,N_34146);
or U36951 (N_36951,N_35065,N_34269);
or U36952 (N_36952,N_35008,N_34229);
and U36953 (N_36953,N_34780,N_35495);
nand U36954 (N_36954,N_35924,N_34811);
nand U36955 (N_36955,N_34632,N_35198);
nand U36956 (N_36956,N_35019,N_34947);
or U36957 (N_36957,N_34335,N_34231);
xor U36958 (N_36958,N_35310,N_35904);
or U36959 (N_36959,N_34260,N_34905);
or U36960 (N_36960,N_35642,N_35341);
nand U36961 (N_36961,N_35077,N_34778);
nand U36962 (N_36962,N_35330,N_34511);
and U36963 (N_36963,N_34297,N_35387);
and U36964 (N_36964,N_35156,N_34344);
nand U36965 (N_36965,N_34621,N_34673);
and U36966 (N_36966,N_34487,N_35457);
nor U36967 (N_36967,N_35100,N_35287);
nor U36968 (N_36968,N_34092,N_35470);
or U36969 (N_36969,N_34063,N_35483);
nand U36970 (N_36970,N_35923,N_35848);
or U36971 (N_36971,N_34976,N_35007);
nor U36972 (N_36972,N_34796,N_35564);
or U36973 (N_36973,N_35773,N_35216);
and U36974 (N_36974,N_35349,N_34902);
and U36975 (N_36975,N_35057,N_34797);
and U36976 (N_36976,N_34257,N_34713);
nand U36977 (N_36977,N_34550,N_35623);
or U36978 (N_36978,N_34071,N_34944);
and U36979 (N_36979,N_35517,N_34184);
nand U36980 (N_36980,N_35374,N_34974);
nor U36981 (N_36981,N_34196,N_34505);
nor U36982 (N_36982,N_34733,N_35888);
or U36983 (N_36983,N_34299,N_34234);
and U36984 (N_36984,N_34715,N_34333);
and U36985 (N_36985,N_34340,N_34208);
and U36986 (N_36986,N_35061,N_35518);
and U36987 (N_36987,N_34288,N_35164);
nor U36988 (N_36988,N_35132,N_34209);
xor U36989 (N_36989,N_35759,N_35002);
nand U36990 (N_36990,N_34066,N_35661);
nor U36991 (N_36991,N_35338,N_34311);
and U36992 (N_36992,N_35079,N_35484);
nand U36993 (N_36993,N_35656,N_35269);
nand U36994 (N_36994,N_35001,N_34222);
or U36995 (N_36995,N_34781,N_34535);
and U36996 (N_36996,N_34471,N_34708);
or U36997 (N_36997,N_35873,N_35724);
xor U36998 (N_36998,N_35979,N_35334);
and U36999 (N_36999,N_34408,N_34541);
or U37000 (N_37000,N_35815,N_34495);
and U37001 (N_37001,N_34009,N_35201);
or U37002 (N_37002,N_34025,N_35355);
or U37003 (N_37003,N_35378,N_34281);
nor U37004 (N_37004,N_35139,N_35818);
nor U37005 (N_37005,N_34917,N_34199);
nand U37006 (N_37006,N_34526,N_34730);
or U37007 (N_37007,N_35668,N_34463);
nor U37008 (N_37008,N_34990,N_35390);
or U37009 (N_37009,N_34395,N_35052);
nand U37010 (N_37010,N_34667,N_34414);
or U37011 (N_37011,N_35890,N_34725);
or U37012 (N_37012,N_34431,N_35113);
or U37013 (N_37013,N_34327,N_35062);
nand U37014 (N_37014,N_35039,N_34675);
or U37015 (N_37015,N_35314,N_34330);
nor U37016 (N_37016,N_35824,N_35803);
and U37017 (N_37017,N_34422,N_35460);
nand U37018 (N_37018,N_35171,N_34975);
and U37019 (N_37019,N_34385,N_34311);
or U37020 (N_37020,N_35665,N_35160);
nor U37021 (N_37021,N_34232,N_34255);
nor U37022 (N_37022,N_35471,N_34196);
or U37023 (N_37023,N_35218,N_34628);
nand U37024 (N_37024,N_34359,N_35679);
nor U37025 (N_37025,N_35556,N_35078);
nor U37026 (N_37026,N_35420,N_34336);
and U37027 (N_37027,N_35839,N_34187);
and U37028 (N_37028,N_34800,N_34347);
or U37029 (N_37029,N_35687,N_35369);
nor U37030 (N_37030,N_34984,N_34978);
and U37031 (N_37031,N_34565,N_35747);
or U37032 (N_37032,N_35657,N_35593);
or U37033 (N_37033,N_35637,N_35368);
nor U37034 (N_37034,N_35442,N_35963);
and U37035 (N_37035,N_34195,N_35556);
or U37036 (N_37036,N_35932,N_34066);
and U37037 (N_37037,N_35416,N_34127);
or U37038 (N_37038,N_35741,N_34421);
nor U37039 (N_37039,N_35555,N_35848);
nor U37040 (N_37040,N_34277,N_34556);
and U37041 (N_37041,N_34451,N_34641);
and U37042 (N_37042,N_34639,N_34923);
nand U37043 (N_37043,N_34837,N_35380);
or U37044 (N_37044,N_34588,N_35703);
nor U37045 (N_37045,N_34408,N_35838);
and U37046 (N_37046,N_35291,N_34008);
and U37047 (N_37047,N_35568,N_35381);
nor U37048 (N_37048,N_34957,N_34098);
nor U37049 (N_37049,N_35288,N_34922);
or U37050 (N_37050,N_35217,N_35100);
nor U37051 (N_37051,N_34377,N_35252);
nand U37052 (N_37052,N_34524,N_34542);
nand U37053 (N_37053,N_35471,N_35578);
and U37054 (N_37054,N_34188,N_35818);
nor U37055 (N_37055,N_34656,N_34657);
nor U37056 (N_37056,N_34288,N_34953);
or U37057 (N_37057,N_35111,N_34005);
and U37058 (N_37058,N_35660,N_34010);
nor U37059 (N_37059,N_34053,N_34553);
nand U37060 (N_37060,N_35270,N_34738);
nand U37061 (N_37061,N_34711,N_35580);
and U37062 (N_37062,N_35586,N_35763);
and U37063 (N_37063,N_35685,N_35305);
nand U37064 (N_37064,N_35041,N_35717);
or U37065 (N_37065,N_34967,N_35589);
nand U37066 (N_37066,N_35782,N_34497);
or U37067 (N_37067,N_34553,N_35126);
nand U37068 (N_37068,N_35398,N_34289);
and U37069 (N_37069,N_35203,N_34702);
or U37070 (N_37070,N_35238,N_35173);
nor U37071 (N_37071,N_35981,N_35875);
nor U37072 (N_37072,N_34833,N_34525);
nor U37073 (N_37073,N_34744,N_35579);
nand U37074 (N_37074,N_35732,N_35175);
nand U37075 (N_37075,N_34180,N_35850);
nor U37076 (N_37076,N_34753,N_35962);
or U37077 (N_37077,N_34004,N_35519);
xor U37078 (N_37078,N_35770,N_35435);
or U37079 (N_37079,N_35117,N_35984);
nand U37080 (N_37080,N_34534,N_35026);
and U37081 (N_37081,N_34649,N_35625);
nor U37082 (N_37082,N_35100,N_34254);
or U37083 (N_37083,N_35739,N_35654);
or U37084 (N_37084,N_34352,N_34942);
nand U37085 (N_37085,N_35882,N_34012);
and U37086 (N_37086,N_35567,N_35357);
nor U37087 (N_37087,N_34297,N_35644);
or U37088 (N_37088,N_34475,N_34549);
nand U37089 (N_37089,N_34800,N_34026);
and U37090 (N_37090,N_35557,N_35815);
nand U37091 (N_37091,N_34638,N_35075);
nor U37092 (N_37092,N_34532,N_34289);
xor U37093 (N_37093,N_34480,N_35934);
and U37094 (N_37094,N_35839,N_34891);
xor U37095 (N_37095,N_34737,N_35685);
and U37096 (N_37096,N_34492,N_35387);
nor U37097 (N_37097,N_35578,N_35945);
nand U37098 (N_37098,N_34380,N_34618);
or U37099 (N_37099,N_34268,N_34141);
nor U37100 (N_37100,N_34338,N_34424);
nor U37101 (N_37101,N_34599,N_35298);
and U37102 (N_37102,N_34338,N_35243);
and U37103 (N_37103,N_34416,N_34266);
or U37104 (N_37104,N_35369,N_34251);
and U37105 (N_37105,N_34081,N_34516);
or U37106 (N_37106,N_34896,N_34675);
nor U37107 (N_37107,N_34011,N_34899);
or U37108 (N_37108,N_34064,N_34896);
nand U37109 (N_37109,N_35072,N_34880);
xnor U37110 (N_37110,N_35737,N_35012);
nor U37111 (N_37111,N_34672,N_35826);
and U37112 (N_37112,N_35805,N_35924);
nor U37113 (N_37113,N_35455,N_34426);
nand U37114 (N_37114,N_35533,N_34260);
nand U37115 (N_37115,N_34360,N_34557);
or U37116 (N_37116,N_35181,N_35965);
nand U37117 (N_37117,N_35364,N_35238);
or U37118 (N_37118,N_34779,N_34935);
nor U37119 (N_37119,N_35076,N_35745);
nand U37120 (N_37120,N_35758,N_35304);
nor U37121 (N_37121,N_35917,N_35730);
and U37122 (N_37122,N_35751,N_35434);
or U37123 (N_37123,N_35410,N_34351);
xnor U37124 (N_37124,N_35918,N_35620);
nor U37125 (N_37125,N_35973,N_34568);
nand U37126 (N_37126,N_35364,N_35409);
nor U37127 (N_37127,N_35266,N_34406);
nor U37128 (N_37128,N_35298,N_35328);
nor U37129 (N_37129,N_34869,N_34913);
or U37130 (N_37130,N_35751,N_35732);
and U37131 (N_37131,N_35646,N_34588);
nor U37132 (N_37132,N_34250,N_34568);
or U37133 (N_37133,N_34710,N_35112);
nor U37134 (N_37134,N_35738,N_35915);
nor U37135 (N_37135,N_35464,N_34213);
and U37136 (N_37136,N_34244,N_35844);
or U37137 (N_37137,N_35156,N_35835);
and U37138 (N_37138,N_34142,N_35956);
and U37139 (N_37139,N_35525,N_34797);
and U37140 (N_37140,N_35848,N_34715);
nand U37141 (N_37141,N_34458,N_35412);
nor U37142 (N_37142,N_35327,N_34771);
nand U37143 (N_37143,N_35325,N_34481);
or U37144 (N_37144,N_34425,N_34338);
or U37145 (N_37145,N_34122,N_34951);
or U37146 (N_37146,N_35966,N_35500);
and U37147 (N_37147,N_34225,N_35135);
xnor U37148 (N_37148,N_34536,N_34563);
nand U37149 (N_37149,N_34966,N_35355);
nor U37150 (N_37150,N_35254,N_35956);
and U37151 (N_37151,N_34822,N_34708);
and U37152 (N_37152,N_35143,N_35929);
nor U37153 (N_37153,N_35271,N_34592);
or U37154 (N_37154,N_35604,N_35463);
nand U37155 (N_37155,N_35990,N_35750);
and U37156 (N_37156,N_34282,N_35550);
and U37157 (N_37157,N_34737,N_34755);
and U37158 (N_37158,N_34661,N_35382);
and U37159 (N_37159,N_35916,N_34960);
or U37160 (N_37160,N_35506,N_35723);
nand U37161 (N_37161,N_34678,N_34006);
and U37162 (N_37162,N_34871,N_35111);
or U37163 (N_37163,N_35948,N_35470);
and U37164 (N_37164,N_34555,N_34160);
nand U37165 (N_37165,N_35626,N_34700);
and U37166 (N_37166,N_35924,N_34359);
and U37167 (N_37167,N_35375,N_34285);
and U37168 (N_37168,N_34497,N_35654);
nor U37169 (N_37169,N_35913,N_35282);
and U37170 (N_37170,N_34927,N_34496);
nand U37171 (N_37171,N_34751,N_35383);
nand U37172 (N_37172,N_35774,N_34863);
nand U37173 (N_37173,N_35974,N_34098);
or U37174 (N_37174,N_35424,N_34330);
nand U37175 (N_37175,N_35595,N_34030);
nand U37176 (N_37176,N_35971,N_35727);
and U37177 (N_37177,N_34746,N_35453);
nand U37178 (N_37178,N_35501,N_34412);
or U37179 (N_37179,N_35060,N_35178);
and U37180 (N_37180,N_34631,N_35171);
nor U37181 (N_37181,N_35823,N_34655);
and U37182 (N_37182,N_34286,N_34749);
nand U37183 (N_37183,N_34338,N_34243);
nor U37184 (N_37184,N_35313,N_35819);
nor U37185 (N_37185,N_34632,N_34910);
nand U37186 (N_37186,N_34258,N_35097);
nand U37187 (N_37187,N_35053,N_34838);
nand U37188 (N_37188,N_34442,N_35938);
nor U37189 (N_37189,N_35586,N_35975);
xor U37190 (N_37190,N_35924,N_35515);
or U37191 (N_37191,N_35626,N_35009);
nor U37192 (N_37192,N_34358,N_35170);
nand U37193 (N_37193,N_35415,N_34192);
or U37194 (N_37194,N_35055,N_34001);
nand U37195 (N_37195,N_35908,N_34037);
nand U37196 (N_37196,N_35945,N_35995);
and U37197 (N_37197,N_34759,N_34878);
and U37198 (N_37198,N_35969,N_35118);
nor U37199 (N_37199,N_34832,N_35027);
or U37200 (N_37200,N_35563,N_35296);
nor U37201 (N_37201,N_34075,N_35865);
xor U37202 (N_37202,N_34049,N_35239);
or U37203 (N_37203,N_34437,N_34527);
nand U37204 (N_37204,N_34403,N_35084);
and U37205 (N_37205,N_34405,N_34055);
xor U37206 (N_37206,N_34344,N_34622);
or U37207 (N_37207,N_34577,N_34434);
nor U37208 (N_37208,N_34728,N_34651);
and U37209 (N_37209,N_34986,N_34779);
and U37210 (N_37210,N_34807,N_34235);
and U37211 (N_37211,N_34211,N_35295);
nor U37212 (N_37212,N_35194,N_35379);
and U37213 (N_37213,N_35616,N_34492);
or U37214 (N_37214,N_34001,N_34700);
or U37215 (N_37215,N_34939,N_35553);
nor U37216 (N_37216,N_34632,N_35813);
or U37217 (N_37217,N_35428,N_34512);
nor U37218 (N_37218,N_35068,N_35698);
and U37219 (N_37219,N_35444,N_35403);
xnor U37220 (N_37220,N_34441,N_35037);
nand U37221 (N_37221,N_35201,N_35242);
and U37222 (N_37222,N_34560,N_35741);
and U37223 (N_37223,N_35075,N_35045);
or U37224 (N_37224,N_34466,N_34796);
nand U37225 (N_37225,N_34967,N_34867);
nand U37226 (N_37226,N_34597,N_34045);
or U37227 (N_37227,N_34675,N_34781);
nand U37228 (N_37228,N_35362,N_34749);
nor U37229 (N_37229,N_35756,N_35982);
nand U37230 (N_37230,N_34573,N_34517);
nand U37231 (N_37231,N_34812,N_35434);
and U37232 (N_37232,N_34797,N_35100);
xor U37233 (N_37233,N_35541,N_35753);
nand U37234 (N_37234,N_34530,N_35660);
or U37235 (N_37235,N_35679,N_34481);
and U37236 (N_37236,N_34544,N_35483);
or U37237 (N_37237,N_34685,N_35496);
nor U37238 (N_37238,N_35283,N_35055);
or U37239 (N_37239,N_34150,N_34159);
and U37240 (N_37240,N_34618,N_34894);
nand U37241 (N_37241,N_34738,N_35088);
or U37242 (N_37242,N_35809,N_35666);
and U37243 (N_37243,N_35418,N_34261);
or U37244 (N_37244,N_35715,N_34575);
or U37245 (N_37245,N_34106,N_34342);
nor U37246 (N_37246,N_34874,N_34540);
or U37247 (N_37247,N_35533,N_34700);
and U37248 (N_37248,N_34528,N_35071);
nor U37249 (N_37249,N_35904,N_34145);
or U37250 (N_37250,N_35306,N_34756);
nor U37251 (N_37251,N_34255,N_34280);
and U37252 (N_37252,N_34726,N_34618);
nor U37253 (N_37253,N_34491,N_34060);
nand U37254 (N_37254,N_35163,N_35619);
or U37255 (N_37255,N_35956,N_35010);
and U37256 (N_37256,N_34743,N_35421);
and U37257 (N_37257,N_34657,N_35225);
and U37258 (N_37258,N_35245,N_35958);
or U37259 (N_37259,N_35878,N_34067);
nand U37260 (N_37260,N_35770,N_34972);
nor U37261 (N_37261,N_35911,N_34480);
nand U37262 (N_37262,N_34919,N_34259);
and U37263 (N_37263,N_35613,N_34686);
and U37264 (N_37264,N_35124,N_35061);
or U37265 (N_37265,N_35091,N_35649);
nor U37266 (N_37266,N_34968,N_34874);
and U37267 (N_37267,N_35752,N_35450);
or U37268 (N_37268,N_34310,N_34637);
nor U37269 (N_37269,N_35248,N_35181);
or U37270 (N_37270,N_34141,N_35376);
or U37271 (N_37271,N_35743,N_34994);
nand U37272 (N_37272,N_35895,N_35320);
nor U37273 (N_37273,N_35602,N_35273);
nor U37274 (N_37274,N_34133,N_35588);
and U37275 (N_37275,N_35621,N_34630);
nand U37276 (N_37276,N_35219,N_34716);
nor U37277 (N_37277,N_35289,N_34398);
nand U37278 (N_37278,N_34623,N_34549);
and U37279 (N_37279,N_35983,N_35940);
nor U37280 (N_37280,N_34080,N_34541);
and U37281 (N_37281,N_35072,N_34669);
nor U37282 (N_37282,N_35814,N_34150);
and U37283 (N_37283,N_35788,N_34819);
nand U37284 (N_37284,N_35124,N_34073);
or U37285 (N_37285,N_35415,N_34985);
nand U37286 (N_37286,N_34840,N_34774);
nor U37287 (N_37287,N_34814,N_35080);
nor U37288 (N_37288,N_35486,N_35104);
or U37289 (N_37289,N_34935,N_34348);
and U37290 (N_37290,N_34311,N_34348);
or U37291 (N_37291,N_34326,N_34199);
and U37292 (N_37292,N_35248,N_34677);
and U37293 (N_37293,N_34680,N_35798);
nand U37294 (N_37294,N_34616,N_34454);
nor U37295 (N_37295,N_35139,N_35123);
and U37296 (N_37296,N_35985,N_35970);
nor U37297 (N_37297,N_35744,N_35400);
nor U37298 (N_37298,N_35530,N_35598);
nand U37299 (N_37299,N_35940,N_34087);
or U37300 (N_37300,N_35504,N_35182);
or U37301 (N_37301,N_34703,N_35197);
nor U37302 (N_37302,N_34773,N_34177);
nand U37303 (N_37303,N_35649,N_35198);
or U37304 (N_37304,N_35531,N_35058);
nand U37305 (N_37305,N_34378,N_34439);
and U37306 (N_37306,N_34971,N_34520);
nor U37307 (N_37307,N_35739,N_34410);
nand U37308 (N_37308,N_35459,N_35245);
and U37309 (N_37309,N_34122,N_35647);
or U37310 (N_37310,N_35124,N_35275);
and U37311 (N_37311,N_34606,N_35556);
and U37312 (N_37312,N_34582,N_34804);
nor U37313 (N_37313,N_35204,N_35900);
nand U37314 (N_37314,N_34051,N_34493);
nand U37315 (N_37315,N_35856,N_34445);
nor U37316 (N_37316,N_35562,N_34220);
xor U37317 (N_37317,N_35209,N_35476);
and U37318 (N_37318,N_35242,N_35583);
and U37319 (N_37319,N_35334,N_34678);
nor U37320 (N_37320,N_35405,N_34681);
or U37321 (N_37321,N_34005,N_34533);
and U37322 (N_37322,N_35767,N_35756);
or U37323 (N_37323,N_34495,N_35997);
or U37324 (N_37324,N_34226,N_34910);
or U37325 (N_37325,N_35556,N_34556);
xnor U37326 (N_37326,N_35139,N_35366);
nor U37327 (N_37327,N_35036,N_34807);
and U37328 (N_37328,N_35342,N_35110);
and U37329 (N_37329,N_35051,N_34496);
nand U37330 (N_37330,N_34744,N_34787);
nor U37331 (N_37331,N_35952,N_35128);
nand U37332 (N_37332,N_34110,N_35106);
and U37333 (N_37333,N_34671,N_34931);
nand U37334 (N_37334,N_34173,N_35585);
or U37335 (N_37335,N_34951,N_35055);
nand U37336 (N_37336,N_35958,N_34861);
nand U37337 (N_37337,N_34095,N_35358);
nor U37338 (N_37338,N_34295,N_34070);
and U37339 (N_37339,N_34202,N_35721);
nand U37340 (N_37340,N_34862,N_35443);
nor U37341 (N_37341,N_34010,N_34057);
nand U37342 (N_37342,N_34789,N_35085);
or U37343 (N_37343,N_35962,N_34357);
xor U37344 (N_37344,N_34890,N_34348);
and U37345 (N_37345,N_35308,N_34048);
nor U37346 (N_37346,N_34846,N_34534);
or U37347 (N_37347,N_34023,N_35751);
nor U37348 (N_37348,N_34834,N_34850);
nand U37349 (N_37349,N_35374,N_34004);
or U37350 (N_37350,N_34695,N_34029);
nand U37351 (N_37351,N_35797,N_34089);
nor U37352 (N_37352,N_34509,N_34911);
and U37353 (N_37353,N_35114,N_35124);
nand U37354 (N_37354,N_35243,N_34986);
nor U37355 (N_37355,N_35978,N_35668);
nor U37356 (N_37356,N_35635,N_34596);
nand U37357 (N_37357,N_34388,N_35889);
or U37358 (N_37358,N_34598,N_35732);
or U37359 (N_37359,N_34332,N_34755);
nor U37360 (N_37360,N_35643,N_35167);
nand U37361 (N_37361,N_35042,N_34477);
or U37362 (N_37362,N_34965,N_34331);
or U37363 (N_37363,N_35220,N_34877);
nor U37364 (N_37364,N_35797,N_35166);
nand U37365 (N_37365,N_34432,N_34623);
nor U37366 (N_37366,N_34286,N_35535);
nor U37367 (N_37367,N_34560,N_35748);
and U37368 (N_37368,N_34418,N_34837);
and U37369 (N_37369,N_35985,N_35944);
and U37370 (N_37370,N_35900,N_34551);
and U37371 (N_37371,N_35905,N_35163);
nor U37372 (N_37372,N_35009,N_34588);
nand U37373 (N_37373,N_34070,N_35328);
nand U37374 (N_37374,N_35967,N_35350);
nand U37375 (N_37375,N_35859,N_35607);
nand U37376 (N_37376,N_34501,N_34069);
nand U37377 (N_37377,N_35483,N_34302);
or U37378 (N_37378,N_35663,N_34978);
or U37379 (N_37379,N_34271,N_34894);
nor U37380 (N_37380,N_35733,N_35700);
and U37381 (N_37381,N_35916,N_35837);
or U37382 (N_37382,N_34913,N_34148);
nor U37383 (N_37383,N_35545,N_35893);
nand U37384 (N_37384,N_34435,N_35512);
nor U37385 (N_37385,N_35760,N_34260);
nor U37386 (N_37386,N_35514,N_34108);
and U37387 (N_37387,N_34992,N_34401);
or U37388 (N_37388,N_34194,N_34028);
nor U37389 (N_37389,N_35413,N_35693);
nand U37390 (N_37390,N_34108,N_35896);
or U37391 (N_37391,N_34367,N_35686);
or U37392 (N_37392,N_35720,N_34207);
xnor U37393 (N_37393,N_35691,N_34237);
and U37394 (N_37394,N_35528,N_34882);
or U37395 (N_37395,N_34990,N_34322);
or U37396 (N_37396,N_34430,N_34113);
and U37397 (N_37397,N_34311,N_34790);
or U37398 (N_37398,N_35319,N_35595);
or U37399 (N_37399,N_34413,N_35913);
nand U37400 (N_37400,N_35168,N_34465);
and U37401 (N_37401,N_35080,N_34306);
or U37402 (N_37402,N_35258,N_34689);
and U37403 (N_37403,N_34188,N_35047);
nand U37404 (N_37404,N_35323,N_35177);
nand U37405 (N_37405,N_35144,N_35675);
or U37406 (N_37406,N_35307,N_34414);
or U37407 (N_37407,N_34308,N_35715);
nand U37408 (N_37408,N_35252,N_35818);
and U37409 (N_37409,N_34222,N_35850);
nor U37410 (N_37410,N_34998,N_34217);
and U37411 (N_37411,N_35035,N_35934);
nand U37412 (N_37412,N_34662,N_35638);
or U37413 (N_37413,N_35603,N_35805);
and U37414 (N_37414,N_34328,N_35908);
nand U37415 (N_37415,N_35217,N_34678);
and U37416 (N_37416,N_35944,N_35720);
or U37417 (N_37417,N_35011,N_35565);
nand U37418 (N_37418,N_34906,N_34110);
nor U37419 (N_37419,N_34979,N_34072);
or U37420 (N_37420,N_34778,N_34009);
or U37421 (N_37421,N_34937,N_35801);
nand U37422 (N_37422,N_34927,N_35374);
nor U37423 (N_37423,N_35279,N_35854);
nand U37424 (N_37424,N_35208,N_35287);
nor U37425 (N_37425,N_34195,N_35763);
and U37426 (N_37426,N_35864,N_35075);
nor U37427 (N_37427,N_34951,N_35451);
nand U37428 (N_37428,N_34670,N_34095);
or U37429 (N_37429,N_35719,N_34206);
or U37430 (N_37430,N_35270,N_35136);
nand U37431 (N_37431,N_34879,N_35897);
and U37432 (N_37432,N_35156,N_34072);
nand U37433 (N_37433,N_35349,N_35180);
or U37434 (N_37434,N_35016,N_35061);
nor U37435 (N_37435,N_34772,N_35465);
and U37436 (N_37436,N_34006,N_35223);
and U37437 (N_37437,N_34781,N_35891);
nor U37438 (N_37438,N_35953,N_34875);
nand U37439 (N_37439,N_34359,N_35816);
or U37440 (N_37440,N_34565,N_34648);
nand U37441 (N_37441,N_34491,N_34020);
nand U37442 (N_37442,N_35786,N_35136);
nor U37443 (N_37443,N_34902,N_34891);
or U37444 (N_37444,N_35292,N_34557);
nor U37445 (N_37445,N_35591,N_34562);
or U37446 (N_37446,N_34307,N_34239);
and U37447 (N_37447,N_35411,N_34438);
nor U37448 (N_37448,N_35150,N_34743);
and U37449 (N_37449,N_35596,N_35741);
or U37450 (N_37450,N_35636,N_34413);
nand U37451 (N_37451,N_35334,N_34924);
or U37452 (N_37452,N_34866,N_34985);
and U37453 (N_37453,N_35329,N_35664);
or U37454 (N_37454,N_34876,N_34605);
nand U37455 (N_37455,N_35964,N_35997);
nand U37456 (N_37456,N_34201,N_34606);
nor U37457 (N_37457,N_34212,N_34865);
nor U37458 (N_37458,N_34753,N_34715);
nand U37459 (N_37459,N_35884,N_35578);
nand U37460 (N_37460,N_35280,N_34740);
xor U37461 (N_37461,N_35896,N_34390);
nand U37462 (N_37462,N_34725,N_34912);
nand U37463 (N_37463,N_35813,N_35620);
nand U37464 (N_37464,N_34755,N_34889);
nand U37465 (N_37465,N_34335,N_35475);
or U37466 (N_37466,N_35488,N_34077);
nor U37467 (N_37467,N_34377,N_34422);
or U37468 (N_37468,N_34437,N_34416);
or U37469 (N_37469,N_35920,N_34585);
nand U37470 (N_37470,N_35902,N_35766);
or U37471 (N_37471,N_35822,N_35188);
nand U37472 (N_37472,N_34336,N_34463);
and U37473 (N_37473,N_35145,N_35851);
or U37474 (N_37474,N_35275,N_35882);
nand U37475 (N_37475,N_35867,N_35345);
nand U37476 (N_37476,N_34359,N_35631);
nor U37477 (N_37477,N_34797,N_35516);
nor U37478 (N_37478,N_35417,N_35223);
and U37479 (N_37479,N_35234,N_35369);
or U37480 (N_37480,N_35348,N_35462);
or U37481 (N_37481,N_34385,N_34252);
and U37482 (N_37482,N_34672,N_35296);
nor U37483 (N_37483,N_35424,N_35258);
nand U37484 (N_37484,N_35896,N_34578);
nor U37485 (N_37485,N_34304,N_35363);
nor U37486 (N_37486,N_35850,N_34593);
or U37487 (N_37487,N_34354,N_35541);
nor U37488 (N_37488,N_34228,N_34799);
nand U37489 (N_37489,N_34401,N_35825);
or U37490 (N_37490,N_34141,N_35431);
or U37491 (N_37491,N_34872,N_34067);
and U37492 (N_37492,N_34325,N_35210);
and U37493 (N_37493,N_35169,N_35949);
or U37494 (N_37494,N_35645,N_35808);
nand U37495 (N_37495,N_34876,N_35458);
and U37496 (N_37496,N_35845,N_35170);
nand U37497 (N_37497,N_34476,N_34614);
and U37498 (N_37498,N_35215,N_35641);
and U37499 (N_37499,N_35758,N_34743);
nor U37500 (N_37500,N_35255,N_34240);
or U37501 (N_37501,N_35018,N_35190);
nand U37502 (N_37502,N_34150,N_35058);
or U37503 (N_37503,N_34352,N_35342);
nor U37504 (N_37504,N_34603,N_35532);
nand U37505 (N_37505,N_34699,N_34432);
nand U37506 (N_37506,N_35241,N_34573);
and U37507 (N_37507,N_35394,N_35107);
nand U37508 (N_37508,N_35243,N_35607);
nand U37509 (N_37509,N_34347,N_34617);
xnor U37510 (N_37510,N_35345,N_35565);
and U37511 (N_37511,N_35441,N_34521);
nand U37512 (N_37512,N_34934,N_35420);
or U37513 (N_37513,N_34768,N_35996);
nand U37514 (N_37514,N_34511,N_34080);
nor U37515 (N_37515,N_34121,N_34884);
nor U37516 (N_37516,N_34794,N_34273);
nor U37517 (N_37517,N_34391,N_34325);
or U37518 (N_37518,N_35364,N_35463);
xor U37519 (N_37519,N_34988,N_35425);
nor U37520 (N_37520,N_34856,N_34890);
and U37521 (N_37521,N_35313,N_35372);
nor U37522 (N_37522,N_34850,N_35631);
or U37523 (N_37523,N_34193,N_34001);
nand U37524 (N_37524,N_34387,N_35195);
and U37525 (N_37525,N_34240,N_34581);
nor U37526 (N_37526,N_35085,N_34955);
or U37527 (N_37527,N_34744,N_35707);
nand U37528 (N_37528,N_35330,N_34327);
nor U37529 (N_37529,N_35522,N_35519);
nand U37530 (N_37530,N_34397,N_35281);
or U37531 (N_37531,N_35083,N_34720);
nand U37532 (N_37532,N_35603,N_35661);
nand U37533 (N_37533,N_35630,N_34467);
or U37534 (N_37534,N_34812,N_35292);
or U37535 (N_37535,N_35531,N_34052);
and U37536 (N_37536,N_35042,N_34977);
and U37537 (N_37537,N_34162,N_34499);
nand U37538 (N_37538,N_35562,N_35950);
and U37539 (N_37539,N_35082,N_35717);
nor U37540 (N_37540,N_34545,N_34022);
and U37541 (N_37541,N_35033,N_34396);
nand U37542 (N_37542,N_34591,N_35375);
or U37543 (N_37543,N_34257,N_34403);
nor U37544 (N_37544,N_34052,N_35833);
nand U37545 (N_37545,N_35716,N_35141);
nand U37546 (N_37546,N_35892,N_34502);
nor U37547 (N_37547,N_34529,N_35157);
or U37548 (N_37548,N_34318,N_34805);
nand U37549 (N_37549,N_34593,N_34318);
nor U37550 (N_37550,N_35492,N_34075);
nor U37551 (N_37551,N_34703,N_35887);
nor U37552 (N_37552,N_35069,N_35262);
nor U37553 (N_37553,N_34849,N_34863);
or U37554 (N_37554,N_35149,N_34268);
nor U37555 (N_37555,N_35182,N_35272);
or U37556 (N_37556,N_35324,N_35269);
nand U37557 (N_37557,N_34220,N_35309);
or U37558 (N_37558,N_35815,N_34419);
nor U37559 (N_37559,N_34236,N_35323);
and U37560 (N_37560,N_35167,N_34206);
and U37561 (N_37561,N_34065,N_35775);
or U37562 (N_37562,N_34044,N_35921);
and U37563 (N_37563,N_34372,N_34907);
nand U37564 (N_37564,N_35105,N_35476);
nor U37565 (N_37565,N_34999,N_34346);
nand U37566 (N_37566,N_35806,N_35965);
and U37567 (N_37567,N_35668,N_34971);
nand U37568 (N_37568,N_34579,N_34432);
xor U37569 (N_37569,N_34505,N_34084);
nor U37570 (N_37570,N_35876,N_34885);
nor U37571 (N_37571,N_35130,N_35948);
and U37572 (N_37572,N_35530,N_35473);
or U37573 (N_37573,N_34408,N_34974);
nand U37574 (N_37574,N_35222,N_35033);
nand U37575 (N_37575,N_35326,N_35088);
or U37576 (N_37576,N_35312,N_34575);
nor U37577 (N_37577,N_34684,N_34808);
or U37578 (N_37578,N_35319,N_34862);
nand U37579 (N_37579,N_35007,N_34200);
nor U37580 (N_37580,N_34941,N_34059);
or U37581 (N_37581,N_35749,N_34095);
or U37582 (N_37582,N_35947,N_35497);
and U37583 (N_37583,N_34508,N_35087);
or U37584 (N_37584,N_35943,N_34407);
or U37585 (N_37585,N_34798,N_35201);
and U37586 (N_37586,N_34207,N_35271);
or U37587 (N_37587,N_34266,N_35373);
nand U37588 (N_37588,N_34973,N_34202);
nor U37589 (N_37589,N_34406,N_35115);
nor U37590 (N_37590,N_34223,N_34692);
or U37591 (N_37591,N_34322,N_35278);
xnor U37592 (N_37592,N_35369,N_35729);
nor U37593 (N_37593,N_35812,N_34465);
or U37594 (N_37594,N_35551,N_34893);
or U37595 (N_37595,N_35437,N_35866);
nor U37596 (N_37596,N_35093,N_35177);
nor U37597 (N_37597,N_35511,N_35833);
or U37598 (N_37598,N_35188,N_34047);
xnor U37599 (N_37599,N_35907,N_35241);
nand U37600 (N_37600,N_35214,N_34575);
and U37601 (N_37601,N_35258,N_35218);
nand U37602 (N_37602,N_35522,N_34247);
nor U37603 (N_37603,N_34840,N_34755);
or U37604 (N_37604,N_34298,N_35360);
and U37605 (N_37605,N_35282,N_35454);
and U37606 (N_37606,N_35645,N_35906);
nand U37607 (N_37607,N_35977,N_34724);
and U37608 (N_37608,N_35641,N_35841);
nand U37609 (N_37609,N_35662,N_35467);
nand U37610 (N_37610,N_35658,N_34693);
and U37611 (N_37611,N_35517,N_35487);
nor U37612 (N_37612,N_34947,N_35247);
nand U37613 (N_37613,N_34342,N_34156);
nand U37614 (N_37614,N_35053,N_34989);
nor U37615 (N_37615,N_34497,N_34675);
nand U37616 (N_37616,N_35673,N_34927);
nand U37617 (N_37617,N_35608,N_35375);
and U37618 (N_37618,N_34836,N_34299);
nand U37619 (N_37619,N_34737,N_35686);
nor U37620 (N_37620,N_34878,N_34108);
nand U37621 (N_37621,N_34828,N_35569);
nor U37622 (N_37622,N_35657,N_35097);
or U37623 (N_37623,N_34971,N_34699);
and U37624 (N_37624,N_35241,N_35314);
nand U37625 (N_37625,N_34605,N_35996);
or U37626 (N_37626,N_35481,N_34131);
nand U37627 (N_37627,N_35470,N_34974);
nand U37628 (N_37628,N_35669,N_34890);
and U37629 (N_37629,N_34676,N_35700);
nand U37630 (N_37630,N_34023,N_35453);
nor U37631 (N_37631,N_35244,N_34506);
or U37632 (N_37632,N_34797,N_34736);
or U37633 (N_37633,N_35093,N_34692);
or U37634 (N_37634,N_35515,N_34284);
or U37635 (N_37635,N_34478,N_35168);
nor U37636 (N_37636,N_34899,N_35459);
nand U37637 (N_37637,N_35943,N_35836);
nor U37638 (N_37638,N_35989,N_35931);
nand U37639 (N_37639,N_34043,N_35952);
nor U37640 (N_37640,N_35700,N_35653);
nor U37641 (N_37641,N_34857,N_35080);
xor U37642 (N_37642,N_34048,N_35429);
nand U37643 (N_37643,N_35110,N_35073);
nand U37644 (N_37644,N_34960,N_35522);
nor U37645 (N_37645,N_35544,N_35764);
or U37646 (N_37646,N_35289,N_35397);
nor U37647 (N_37647,N_35796,N_34781);
and U37648 (N_37648,N_34915,N_35861);
or U37649 (N_37649,N_35237,N_34673);
and U37650 (N_37650,N_35393,N_35292);
and U37651 (N_37651,N_35615,N_35374);
nand U37652 (N_37652,N_34762,N_34401);
nor U37653 (N_37653,N_35044,N_34950);
nand U37654 (N_37654,N_34412,N_34958);
nor U37655 (N_37655,N_35891,N_34055);
nand U37656 (N_37656,N_35779,N_34987);
nor U37657 (N_37657,N_35327,N_34281);
nand U37658 (N_37658,N_35289,N_34408);
and U37659 (N_37659,N_35737,N_35904);
nor U37660 (N_37660,N_34311,N_35387);
nor U37661 (N_37661,N_34018,N_35271);
nand U37662 (N_37662,N_35987,N_35940);
and U37663 (N_37663,N_34060,N_35868);
nand U37664 (N_37664,N_35582,N_34771);
and U37665 (N_37665,N_34315,N_34231);
nand U37666 (N_37666,N_35425,N_35520);
nand U37667 (N_37667,N_35830,N_35236);
nor U37668 (N_37668,N_35673,N_35003);
or U37669 (N_37669,N_35332,N_35883);
nand U37670 (N_37670,N_34981,N_34506);
nand U37671 (N_37671,N_35892,N_34032);
nor U37672 (N_37672,N_34523,N_35641);
nor U37673 (N_37673,N_34333,N_35908);
or U37674 (N_37674,N_34878,N_35611);
or U37675 (N_37675,N_34692,N_34914);
and U37676 (N_37676,N_35313,N_34529);
and U37677 (N_37677,N_34350,N_34904);
or U37678 (N_37678,N_35090,N_34411);
nor U37679 (N_37679,N_34459,N_35317);
nand U37680 (N_37680,N_34874,N_34501);
and U37681 (N_37681,N_35655,N_35115);
and U37682 (N_37682,N_34288,N_35492);
nand U37683 (N_37683,N_34282,N_34727);
and U37684 (N_37684,N_35211,N_35812);
and U37685 (N_37685,N_35713,N_34564);
and U37686 (N_37686,N_34880,N_35355);
and U37687 (N_37687,N_34672,N_35579);
nand U37688 (N_37688,N_35831,N_34239);
or U37689 (N_37689,N_34102,N_34798);
and U37690 (N_37690,N_34754,N_34750);
or U37691 (N_37691,N_34739,N_34738);
nand U37692 (N_37692,N_35310,N_34362);
nor U37693 (N_37693,N_34844,N_35873);
nor U37694 (N_37694,N_34612,N_35777);
nor U37695 (N_37695,N_35674,N_35266);
or U37696 (N_37696,N_34429,N_35924);
or U37697 (N_37697,N_35663,N_35483);
nand U37698 (N_37698,N_35450,N_34315);
nor U37699 (N_37699,N_35373,N_35058);
nand U37700 (N_37700,N_34596,N_35441);
nand U37701 (N_37701,N_35271,N_35515);
xor U37702 (N_37702,N_34288,N_35412);
nand U37703 (N_37703,N_34648,N_34028);
nand U37704 (N_37704,N_35776,N_35676);
nand U37705 (N_37705,N_35225,N_35785);
or U37706 (N_37706,N_35960,N_35297);
nor U37707 (N_37707,N_35418,N_35938);
or U37708 (N_37708,N_34718,N_34008);
and U37709 (N_37709,N_35324,N_35006);
nor U37710 (N_37710,N_35835,N_35856);
or U37711 (N_37711,N_35679,N_34205);
nor U37712 (N_37712,N_35673,N_35372);
nand U37713 (N_37713,N_34128,N_34021);
nor U37714 (N_37714,N_35667,N_35747);
nand U37715 (N_37715,N_35813,N_35499);
nand U37716 (N_37716,N_34290,N_34354);
and U37717 (N_37717,N_35496,N_34303);
nor U37718 (N_37718,N_35234,N_35847);
nor U37719 (N_37719,N_35570,N_34589);
nand U37720 (N_37720,N_35451,N_34867);
nor U37721 (N_37721,N_34188,N_35770);
or U37722 (N_37722,N_35308,N_35378);
or U37723 (N_37723,N_34953,N_35509);
or U37724 (N_37724,N_34748,N_34536);
nor U37725 (N_37725,N_34158,N_35760);
nand U37726 (N_37726,N_35298,N_34478);
or U37727 (N_37727,N_35451,N_35958);
and U37728 (N_37728,N_34182,N_35745);
and U37729 (N_37729,N_35750,N_35982);
or U37730 (N_37730,N_34360,N_35265);
and U37731 (N_37731,N_34961,N_35408);
and U37732 (N_37732,N_35127,N_35061);
nor U37733 (N_37733,N_35924,N_35102);
or U37734 (N_37734,N_35345,N_35006);
nor U37735 (N_37735,N_34172,N_35036);
nand U37736 (N_37736,N_35737,N_35620);
and U37737 (N_37737,N_34380,N_34543);
nor U37738 (N_37738,N_34604,N_35230);
or U37739 (N_37739,N_35179,N_35829);
nand U37740 (N_37740,N_34040,N_34873);
and U37741 (N_37741,N_35653,N_35591);
or U37742 (N_37742,N_34849,N_35081);
nor U37743 (N_37743,N_35157,N_35990);
nand U37744 (N_37744,N_35845,N_35087);
nor U37745 (N_37745,N_34564,N_35445);
or U37746 (N_37746,N_34566,N_35238);
nor U37747 (N_37747,N_34422,N_35432);
and U37748 (N_37748,N_35344,N_35586);
and U37749 (N_37749,N_35552,N_35114);
or U37750 (N_37750,N_35609,N_35111);
nor U37751 (N_37751,N_35110,N_34833);
nand U37752 (N_37752,N_34212,N_34611);
nand U37753 (N_37753,N_35836,N_35558);
nor U37754 (N_37754,N_35710,N_35828);
nand U37755 (N_37755,N_34516,N_34097);
and U37756 (N_37756,N_35043,N_35084);
nand U37757 (N_37757,N_34201,N_35894);
and U37758 (N_37758,N_35097,N_34864);
nand U37759 (N_37759,N_34771,N_34529);
or U37760 (N_37760,N_34237,N_34188);
or U37761 (N_37761,N_34910,N_34830);
and U37762 (N_37762,N_34488,N_35289);
nand U37763 (N_37763,N_34112,N_35318);
nor U37764 (N_37764,N_34151,N_35942);
and U37765 (N_37765,N_34561,N_34898);
xor U37766 (N_37766,N_34499,N_35639);
nand U37767 (N_37767,N_35004,N_34021);
nand U37768 (N_37768,N_34700,N_35251);
nand U37769 (N_37769,N_35296,N_35467);
nand U37770 (N_37770,N_35168,N_35415);
nand U37771 (N_37771,N_34518,N_35913);
or U37772 (N_37772,N_34266,N_34849);
nand U37773 (N_37773,N_35686,N_34266);
nand U37774 (N_37774,N_35727,N_34412);
or U37775 (N_37775,N_34466,N_34995);
nor U37776 (N_37776,N_34608,N_35308);
or U37777 (N_37777,N_34375,N_34235);
nand U37778 (N_37778,N_34152,N_35686);
and U37779 (N_37779,N_34951,N_35703);
or U37780 (N_37780,N_35522,N_35097);
or U37781 (N_37781,N_34129,N_35235);
or U37782 (N_37782,N_34046,N_34799);
nor U37783 (N_37783,N_34665,N_35142);
nand U37784 (N_37784,N_34431,N_35508);
nand U37785 (N_37785,N_34628,N_35557);
and U37786 (N_37786,N_34543,N_35028);
and U37787 (N_37787,N_34133,N_35428);
or U37788 (N_37788,N_34608,N_35852);
nor U37789 (N_37789,N_35417,N_35221);
nand U37790 (N_37790,N_34709,N_35838);
nand U37791 (N_37791,N_34936,N_35036);
nand U37792 (N_37792,N_35523,N_35724);
nand U37793 (N_37793,N_34300,N_35007);
and U37794 (N_37794,N_35691,N_34806);
nor U37795 (N_37795,N_34243,N_34014);
or U37796 (N_37796,N_34503,N_35213);
nand U37797 (N_37797,N_35363,N_34335);
or U37798 (N_37798,N_35028,N_34440);
or U37799 (N_37799,N_34361,N_34387);
or U37800 (N_37800,N_35703,N_34031);
and U37801 (N_37801,N_35492,N_35891);
nor U37802 (N_37802,N_35295,N_34480);
or U37803 (N_37803,N_34005,N_35267);
nand U37804 (N_37804,N_34888,N_35281);
or U37805 (N_37805,N_35325,N_35777);
nand U37806 (N_37806,N_35779,N_34823);
nand U37807 (N_37807,N_35227,N_34430);
nand U37808 (N_37808,N_35169,N_34870);
or U37809 (N_37809,N_35704,N_35761);
nand U37810 (N_37810,N_34272,N_35510);
nor U37811 (N_37811,N_34292,N_34080);
nor U37812 (N_37812,N_35266,N_34395);
nor U37813 (N_37813,N_34266,N_34025);
nor U37814 (N_37814,N_34216,N_35028);
or U37815 (N_37815,N_34471,N_35419);
or U37816 (N_37816,N_34223,N_34941);
nor U37817 (N_37817,N_34409,N_35543);
nand U37818 (N_37818,N_35782,N_34465);
xnor U37819 (N_37819,N_35454,N_34479);
and U37820 (N_37820,N_35110,N_34973);
and U37821 (N_37821,N_34896,N_35458);
nor U37822 (N_37822,N_35481,N_34024);
or U37823 (N_37823,N_34562,N_34740);
or U37824 (N_37824,N_35551,N_34682);
and U37825 (N_37825,N_34278,N_35264);
or U37826 (N_37826,N_34182,N_34232);
or U37827 (N_37827,N_35010,N_35022);
nor U37828 (N_37828,N_34620,N_34249);
nor U37829 (N_37829,N_34150,N_35118);
nand U37830 (N_37830,N_34206,N_34860);
nand U37831 (N_37831,N_34866,N_34642);
or U37832 (N_37832,N_34900,N_34314);
nand U37833 (N_37833,N_34455,N_34066);
nor U37834 (N_37834,N_35992,N_34255);
and U37835 (N_37835,N_34274,N_35627);
nand U37836 (N_37836,N_35418,N_35471);
or U37837 (N_37837,N_34919,N_34320);
or U37838 (N_37838,N_35604,N_35435);
and U37839 (N_37839,N_35472,N_34959);
or U37840 (N_37840,N_34151,N_35753);
or U37841 (N_37841,N_34995,N_34204);
and U37842 (N_37842,N_34850,N_35760);
nor U37843 (N_37843,N_35199,N_34221);
nand U37844 (N_37844,N_34552,N_35951);
or U37845 (N_37845,N_34270,N_35628);
nand U37846 (N_37846,N_34389,N_35602);
nor U37847 (N_37847,N_35834,N_34264);
or U37848 (N_37848,N_35129,N_34069);
and U37849 (N_37849,N_35350,N_34964);
and U37850 (N_37850,N_34685,N_34610);
nor U37851 (N_37851,N_34011,N_35178);
and U37852 (N_37852,N_34019,N_34390);
or U37853 (N_37853,N_35676,N_35388);
xnor U37854 (N_37854,N_34302,N_35788);
or U37855 (N_37855,N_34018,N_34680);
nor U37856 (N_37856,N_34072,N_35707);
or U37857 (N_37857,N_34449,N_34096);
and U37858 (N_37858,N_35926,N_34893);
nor U37859 (N_37859,N_34826,N_35642);
nand U37860 (N_37860,N_35851,N_34445);
nor U37861 (N_37861,N_34018,N_35843);
or U37862 (N_37862,N_34608,N_34368);
nor U37863 (N_37863,N_35007,N_35080);
nand U37864 (N_37864,N_34287,N_35535);
nor U37865 (N_37865,N_34569,N_35760);
nand U37866 (N_37866,N_35053,N_34663);
and U37867 (N_37867,N_35445,N_35062);
nor U37868 (N_37868,N_35957,N_35140);
and U37869 (N_37869,N_35680,N_35654);
nand U37870 (N_37870,N_34403,N_35237);
or U37871 (N_37871,N_35305,N_34849);
or U37872 (N_37872,N_34316,N_35267);
nor U37873 (N_37873,N_35056,N_35585);
or U37874 (N_37874,N_35970,N_34392);
nor U37875 (N_37875,N_35962,N_34853);
nor U37876 (N_37876,N_35558,N_34820);
nor U37877 (N_37877,N_34653,N_35962);
nand U37878 (N_37878,N_35961,N_34127);
nand U37879 (N_37879,N_34924,N_35202);
or U37880 (N_37880,N_35325,N_34412);
and U37881 (N_37881,N_34988,N_34581);
or U37882 (N_37882,N_34046,N_34649);
and U37883 (N_37883,N_34982,N_35161);
nand U37884 (N_37884,N_35666,N_35232);
nor U37885 (N_37885,N_34356,N_34366);
and U37886 (N_37886,N_35073,N_34079);
and U37887 (N_37887,N_34844,N_35945);
and U37888 (N_37888,N_35641,N_34805);
nor U37889 (N_37889,N_35240,N_35602);
nor U37890 (N_37890,N_35773,N_35206);
nand U37891 (N_37891,N_34804,N_35244);
and U37892 (N_37892,N_35229,N_34176);
or U37893 (N_37893,N_35061,N_35631);
and U37894 (N_37894,N_35549,N_34996);
or U37895 (N_37895,N_34753,N_35410);
nand U37896 (N_37896,N_35029,N_35982);
and U37897 (N_37897,N_35807,N_35492);
and U37898 (N_37898,N_34447,N_35608);
and U37899 (N_37899,N_35989,N_35050);
nand U37900 (N_37900,N_35493,N_34862);
or U37901 (N_37901,N_35046,N_35841);
nor U37902 (N_37902,N_35672,N_35483);
and U37903 (N_37903,N_35084,N_35218);
nor U37904 (N_37904,N_35802,N_35997);
and U37905 (N_37905,N_35203,N_34289);
or U37906 (N_37906,N_35171,N_35878);
nor U37907 (N_37907,N_34830,N_35460);
nor U37908 (N_37908,N_34025,N_35414);
nor U37909 (N_37909,N_34581,N_35126);
or U37910 (N_37910,N_35790,N_34120);
nor U37911 (N_37911,N_35617,N_35001);
nand U37912 (N_37912,N_35253,N_35179);
nand U37913 (N_37913,N_34156,N_35964);
nor U37914 (N_37914,N_35087,N_34979);
and U37915 (N_37915,N_34566,N_35256);
nand U37916 (N_37916,N_35780,N_35335);
nand U37917 (N_37917,N_34915,N_34722);
nand U37918 (N_37918,N_35943,N_35580);
xor U37919 (N_37919,N_35062,N_34062);
nor U37920 (N_37920,N_34637,N_35026);
or U37921 (N_37921,N_35690,N_35728);
or U37922 (N_37922,N_34821,N_34637);
and U37923 (N_37923,N_35594,N_34203);
nor U37924 (N_37924,N_34939,N_34343);
and U37925 (N_37925,N_35498,N_34525);
or U37926 (N_37926,N_35999,N_34913);
and U37927 (N_37927,N_35423,N_35341);
xnor U37928 (N_37928,N_34358,N_34441);
or U37929 (N_37929,N_34684,N_34799);
and U37930 (N_37930,N_34237,N_34769);
nor U37931 (N_37931,N_35912,N_35228);
or U37932 (N_37932,N_35705,N_34269);
nand U37933 (N_37933,N_35899,N_34088);
or U37934 (N_37934,N_34832,N_35968);
nand U37935 (N_37935,N_34914,N_35686);
and U37936 (N_37936,N_35765,N_35837);
nor U37937 (N_37937,N_35646,N_34320);
or U37938 (N_37938,N_34320,N_34975);
nor U37939 (N_37939,N_34003,N_35736);
nor U37940 (N_37940,N_35971,N_35242);
nand U37941 (N_37941,N_34879,N_35765);
nand U37942 (N_37942,N_34199,N_35160);
nor U37943 (N_37943,N_35050,N_35249);
nor U37944 (N_37944,N_35074,N_34262);
nand U37945 (N_37945,N_34971,N_34675);
nand U37946 (N_37946,N_34940,N_35969);
and U37947 (N_37947,N_34419,N_34042);
or U37948 (N_37948,N_35221,N_35814);
and U37949 (N_37949,N_34885,N_35831);
or U37950 (N_37950,N_34190,N_34466);
xor U37951 (N_37951,N_35173,N_34949);
and U37952 (N_37952,N_35826,N_34418);
xnor U37953 (N_37953,N_34032,N_35657);
nor U37954 (N_37954,N_35766,N_34357);
nor U37955 (N_37955,N_34525,N_35463);
nor U37956 (N_37956,N_35213,N_35747);
nand U37957 (N_37957,N_34088,N_35499);
nand U37958 (N_37958,N_35040,N_35449);
nor U37959 (N_37959,N_34757,N_34812);
xor U37960 (N_37960,N_35322,N_35830);
and U37961 (N_37961,N_34425,N_35990);
nand U37962 (N_37962,N_34860,N_34461);
nor U37963 (N_37963,N_34533,N_35616);
or U37964 (N_37964,N_35197,N_35375);
or U37965 (N_37965,N_35253,N_34752);
and U37966 (N_37966,N_34569,N_35305);
or U37967 (N_37967,N_35047,N_34526);
or U37968 (N_37968,N_34931,N_34758);
or U37969 (N_37969,N_34312,N_35702);
nor U37970 (N_37970,N_34458,N_34972);
or U37971 (N_37971,N_35573,N_35865);
xor U37972 (N_37972,N_35032,N_35393);
or U37973 (N_37973,N_35298,N_35297);
or U37974 (N_37974,N_34533,N_34354);
or U37975 (N_37975,N_34983,N_35994);
nor U37976 (N_37976,N_34793,N_35236);
nor U37977 (N_37977,N_35410,N_35034);
nand U37978 (N_37978,N_35156,N_35548);
nand U37979 (N_37979,N_35709,N_34608);
or U37980 (N_37980,N_34290,N_34512);
nor U37981 (N_37981,N_35761,N_35536);
or U37982 (N_37982,N_34127,N_35677);
nand U37983 (N_37983,N_35256,N_34813);
nor U37984 (N_37984,N_35636,N_35071);
or U37985 (N_37985,N_34378,N_35025);
nor U37986 (N_37986,N_35052,N_35776);
or U37987 (N_37987,N_34336,N_35861);
and U37988 (N_37988,N_35866,N_35550);
and U37989 (N_37989,N_34019,N_35458);
and U37990 (N_37990,N_34927,N_35916);
nand U37991 (N_37991,N_35229,N_35389);
or U37992 (N_37992,N_34061,N_34760);
xor U37993 (N_37993,N_35767,N_35790);
and U37994 (N_37994,N_35149,N_34086);
nor U37995 (N_37995,N_34922,N_34734);
and U37996 (N_37996,N_35112,N_34040);
and U37997 (N_37997,N_34632,N_34937);
nor U37998 (N_37998,N_35703,N_34537);
or U37999 (N_37999,N_35961,N_34118);
or U38000 (N_38000,N_37589,N_37663);
nor U38001 (N_38001,N_36304,N_37688);
nand U38002 (N_38002,N_37930,N_36853);
nand U38003 (N_38003,N_37281,N_37186);
or U38004 (N_38004,N_37945,N_36081);
or U38005 (N_38005,N_36651,N_36328);
or U38006 (N_38006,N_36367,N_37680);
nor U38007 (N_38007,N_37320,N_36250);
nand U38008 (N_38008,N_37564,N_37559);
nor U38009 (N_38009,N_36720,N_36243);
or U38010 (N_38010,N_37443,N_37062);
and U38011 (N_38011,N_37334,N_37814);
nand U38012 (N_38012,N_37361,N_36575);
nand U38013 (N_38013,N_37227,N_37393);
nand U38014 (N_38014,N_36798,N_37793);
nor U38015 (N_38015,N_37053,N_37411);
nor U38016 (N_38016,N_36525,N_36880);
and U38017 (N_38017,N_37436,N_36169);
nand U38018 (N_38018,N_36240,N_37604);
xor U38019 (N_38019,N_36141,N_36646);
or U38020 (N_38020,N_37236,N_37901);
or U38021 (N_38021,N_36282,N_36697);
nor U38022 (N_38022,N_37545,N_36685);
nand U38023 (N_38023,N_37843,N_37075);
nand U38024 (N_38024,N_36285,N_37746);
nor U38025 (N_38025,N_37728,N_37040);
or U38026 (N_38026,N_37175,N_36036);
and U38027 (N_38027,N_36186,N_36184);
nor U38028 (N_38028,N_37685,N_36069);
nor U38029 (N_38029,N_36345,N_36579);
and U38030 (N_38030,N_36013,N_37494);
nor U38031 (N_38031,N_36356,N_36007);
nor U38032 (N_38032,N_37890,N_36123);
and U38033 (N_38033,N_37992,N_37629);
and U38034 (N_38034,N_36956,N_36978);
nor U38035 (N_38035,N_36666,N_37765);
nand U38036 (N_38036,N_36911,N_36902);
or U38037 (N_38037,N_36124,N_37584);
and U38038 (N_38038,N_37250,N_37855);
nor U38039 (N_38039,N_36607,N_37705);
nor U38040 (N_38040,N_36025,N_36842);
nand U38041 (N_38041,N_36516,N_37557);
nor U38042 (N_38042,N_36675,N_37838);
or U38043 (N_38043,N_36619,N_36783);
and U38044 (N_38044,N_37234,N_36212);
and U38045 (N_38045,N_36887,N_37834);
xor U38046 (N_38046,N_37318,N_37998);
or U38047 (N_38047,N_37370,N_36095);
or U38048 (N_38048,N_37521,N_36699);
and U38049 (N_38049,N_37201,N_36787);
nor U38050 (N_38050,N_36636,N_36227);
and U38051 (N_38051,N_37285,N_36496);
nor U38052 (N_38052,N_36475,N_36102);
or U38053 (N_38053,N_36335,N_36654);
nor U38054 (N_38054,N_36079,N_36959);
nand U38055 (N_38055,N_36406,N_36620);
nor U38056 (N_38056,N_36316,N_36108);
and U38057 (N_38057,N_36991,N_37060);
nor U38058 (N_38058,N_37081,N_37755);
nand U38059 (N_38059,N_36032,N_36995);
nor U38060 (N_38060,N_36612,N_37230);
and U38061 (N_38061,N_36520,N_37734);
nor U38062 (N_38062,N_37172,N_36495);
nor U38063 (N_38063,N_37546,N_37110);
nand U38064 (N_38064,N_37007,N_37089);
xor U38065 (N_38065,N_36837,N_36490);
xnor U38066 (N_38066,N_37377,N_37129);
and U38067 (N_38067,N_37555,N_36979);
or U38068 (N_38068,N_37136,N_37104);
and U38069 (N_38069,N_36633,N_37255);
nand U38070 (N_38070,N_36364,N_37983);
and U38071 (N_38071,N_36056,N_37469);
xor U38072 (N_38072,N_37977,N_36093);
or U38073 (N_38073,N_36080,N_37033);
nand U38074 (N_38074,N_36778,N_36001);
nor U38075 (N_38075,N_37074,N_37079);
and U38076 (N_38076,N_36353,N_36306);
nand U38077 (N_38077,N_37824,N_36347);
nor U38078 (N_38078,N_36738,N_36663);
or U38079 (N_38079,N_37517,N_36550);
or U38080 (N_38080,N_36524,N_36363);
nand U38081 (N_38081,N_36258,N_37309);
or U38082 (N_38082,N_37094,N_36688);
or U38083 (N_38083,N_37923,N_37528);
nor U38084 (N_38084,N_36867,N_36270);
and U38085 (N_38085,N_36561,N_37384);
or U38086 (N_38086,N_37023,N_36760);
nand U38087 (N_38087,N_36052,N_36324);
nand U38088 (N_38088,N_36439,N_37775);
and U38089 (N_38089,N_36091,N_36393);
or U38090 (N_38090,N_37390,N_36936);
or U38091 (N_38091,N_37940,N_36856);
nor U38092 (N_38092,N_36661,N_37468);
nand U38093 (N_38093,N_37723,N_37841);
nor U38094 (N_38094,N_37386,N_36313);
and U38095 (N_38095,N_37541,N_36779);
and U38096 (N_38096,N_36728,N_37988);
nor U38097 (N_38097,N_36850,N_37866);
nand U38098 (N_38098,N_36368,N_37100);
and U38099 (N_38099,N_37064,N_37102);
nand U38100 (N_38100,N_37140,N_36724);
nor U38101 (N_38101,N_37433,N_37976);
nor U38102 (N_38102,N_37424,N_36875);
and U38103 (N_38103,N_37985,N_37605);
nor U38104 (N_38104,N_37753,N_36327);
nand U38105 (N_38105,N_36523,N_36017);
nand U38106 (N_38106,N_37303,N_37679);
or U38107 (N_38107,N_37562,N_37877);
nor U38108 (N_38108,N_36209,N_37482);
nand U38109 (N_38109,N_36061,N_37566);
nand U38110 (N_38110,N_36544,N_36121);
nand U38111 (N_38111,N_36385,N_36522);
nor U38112 (N_38112,N_36411,N_36404);
nand U38113 (N_38113,N_37238,N_37830);
nand U38114 (N_38114,N_36729,N_36952);
or U38115 (N_38115,N_36592,N_36461);
nor U38116 (N_38116,N_37353,N_37054);
nor U38117 (N_38117,N_36326,N_36541);
nor U38118 (N_38118,N_37633,N_37774);
and U38119 (N_38119,N_37360,N_37844);
nor U38120 (N_38120,N_37152,N_37720);
or U38121 (N_38121,N_36564,N_37550);
nor U38122 (N_38122,N_36008,N_37966);
or U38123 (N_38123,N_36866,N_36676);
or U38124 (N_38124,N_37766,N_36259);
and U38125 (N_38125,N_36279,N_37187);
nand U38126 (N_38126,N_37256,N_36932);
or U38127 (N_38127,N_36921,N_37453);
and U38128 (N_38128,N_36819,N_36252);
and U38129 (N_38129,N_36031,N_36801);
or U38130 (N_38130,N_37741,N_36648);
nor U38131 (N_38131,N_37308,N_37167);
or U38132 (N_38132,N_36230,N_37724);
nor U38133 (N_38133,N_36482,N_37665);
nor U38134 (N_38134,N_37455,N_36931);
or U38135 (N_38135,N_37055,N_37061);
or U38136 (N_38136,N_36832,N_37692);
nor U38137 (N_38137,N_36774,N_36777);
nor U38138 (N_38138,N_36623,N_37896);
nor U38139 (N_38139,N_37748,N_36092);
and U38140 (N_38140,N_36305,N_36397);
and U38141 (N_38141,N_37533,N_36148);
and U38142 (N_38142,N_36621,N_37592);
nand U38143 (N_38143,N_37942,N_37925);
or U38144 (N_38144,N_37614,N_37088);
or U38145 (N_38145,N_37972,N_36785);
nand U38146 (N_38146,N_36613,N_37237);
nor U38147 (N_38147,N_36381,N_37931);
nor U38148 (N_38148,N_36300,N_37233);
nand U38149 (N_38149,N_36907,N_37403);
nand U38150 (N_38150,N_36929,N_37625);
nand U38151 (N_38151,N_37943,N_36048);
nor U38152 (N_38152,N_37590,N_37247);
or U38153 (N_38153,N_36752,N_37000);
nor U38154 (N_38154,N_36540,N_36749);
nor U38155 (N_38155,N_37861,N_37707);
or U38156 (N_38156,N_37691,N_36357);
nor U38157 (N_38157,N_37941,N_37702);
and U38158 (N_38158,N_36140,N_37908);
nor U38159 (N_38159,N_36692,N_36903);
and U38160 (N_38160,N_37730,N_36387);
nor U38161 (N_38161,N_37619,N_36582);
or U38162 (N_38162,N_36926,N_36042);
nand U38163 (N_38163,N_37512,N_37177);
and U38164 (N_38164,N_36493,N_37388);
and U38165 (N_38165,N_37179,N_36156);
nor U38166 (N_38166,N_37761,N_36735);
and U38167 (N_38167,N_37822,N_37875);
or U38168 (N_38168,N_36830,N_36764);
and U38169 (N_38169,N_36040,N_37495);
and U38170 (N_38170,N_36310,N_37463);
nor U38171 (N_38171,N_36810,N_37769);
or U38172 (N_38172,N_36770,N_36910);
nor U38173 (N_38173,N_37103,N_37457);
and U38174 (N_38174,N_37410,N_36375);
nor U38175 (N_38175,N_37211,N_36792);
or U38176 (N_38176,N_36154,N_37056);
or U38177 (N_38177,N_37727,N_36580);
and U38178 (N_38178,N_36268,N_37488);
or U38179 (N_38179,N_36436,N_37960);
nor U38180 (N_38180,N_37603,N_37314);
nor U38181 (N_38181,N_36394,N_36665);
or U38182 (N_38182,N_37899,N_37666);
nor U38183 (N_38183,N_37754,N_36768);
nand U38184 (N_38184,N_37485,N_37645);
nor U38185 (N_38185,N_37818,N_36177);
and U38186 (N_38186,N_36292,N_36740);
nor U38187 (N_38187,N_36362,N_36103);
and U38188 (N_38188,N_36918,N_36873);
nor U38189 (N_38189,N_37714,N_37354);
nand U38190 (N_38190,N_37624,N_36839);
nor U38191 (N_38191,N_36147,N_36222);
nor U38192 (N_38192,N_37504,N_37507);
nand U38193 (N_38193,N_36137,N_36742);
and U38194 (N_38194,N_37395,N_37848);
or U38195 (N_38195,N_36788,N_37194);
or U38196 (N_38196,N_36396,N_36349);
nand U38197 (N_38197,N_37525,N_37904);
and U38198 (N_38198,N_37639,N_36275);
nor U38199 (N_38199,N_37704,N_36727);
nor U38200 (N_38200,N_36281,N_37419);
and U38201 (N_38201,N_36127,N_37535);
and U38202 (N_38202,N_37965,N_36553);
and U38203 (N_38203,N_37228,N_36504);
or U38204 (N_38204,N_36710,N_36456);
and U38205 (N_38205,N_37414,N_37523);
nand U38206 (N_38206,N_36595,N_37750);
nand U38207 (N_38207,N_37339,N_36078);
and U38208 (N_38208,N_37682,N_36446);
nor U38209 (N_38209,N_37034,N_36199);
nor U38210 (N_38210,N_37917,N_37014);
xnor U38211 (N_38211,N_37291,N_37997);
nor U38212 (N_38212,N_36448,N_37646);
nor U38213 (N_38213,N_37460,N_36552);
nand U38214 (N_38214,N_36732,N_37602);
nor U38215 (N_38215,N_36000,N_36346);
and U38216 (N_38216,N_36440,N_37563);
or U38217 (N_38217,N_36129,N_36500);
nand U38218 (N_38218,N_36467,N_37371);
or U38219 (N_38219,N_37322,N_37542);
xnor U38220 (N_38220,N_37212,N_37251);
nor U38221 (N_38221,N_36046,N_36262);
or U38222 (N_38222,N_37153,N_36371);
or U38223 (N_38223,N_36437,N_36115);
and U38224 (N_38224,N_37658,N_36445);
nor U38225 (N_38225,N_36958,N_36369);
or U38226 (N_38226,N_37782,N_37405);
nor U38227 (N_38227,N_36064,N_36034);
or U38228 (N_38228,N_36805,N_37017);
nand U38229 (N_38229,N_37929,N_37437);
and U38230 (N_38230,N_37618,N_37560);
or U38231 (N_38231,N_37305,N_37743);
nand U38232 (N_38232,N_37125,N_36981);
nor U38233 (N_38233,N_36014,N_37058);
nor U38234 (N_38234,N_37148,N_37332);
and U38235 (N_38235,N_37781,N_36506);
nor U38236 (N_38236,N_37697,N_36847);
nand U38237 (N_38237,N_36898,N_37547);
nor U38238 (N_38238,N_36861,N_36751);
and U38239 (N_38239,N_36869,N_37514);
nor U38240 (N_38240,N_36529,N_37127);
or U38241 (N_38241,N_37406,N_36090);
nand U38242 (N_38242,N_36965,N_36024);
and U38243 (N_38243,N_36970,N_36374);
or U38244 (N_38244,N_37587,N_36038);
xor U38245 (N_38245,N_36457,N_36094);
and U38246 (N_38246,N_37135,N_36757);
nor U38247 (N_38247,N_37576,N_37464);
and U38248 (N_38248,N_37372,N_37572);
or U38249 (N_38249,N_36941,N_37345);
nor U38250 (N_38250,N_36984,N_36722);
nand U38251 (N_38251,N_36100,N_37188);
or U38252 (N_38252,N_37948,N_37116);
xnor U38253 (N_38253,N_37107,N_37001);
and U38254 (N_38254,N_36293,N_37969);
or U38255 (N_38255,N_37610,N_37570);
nor U38256 (N_38256,N_36597,N_37134);
nand U38257 (N_38257,N_36355,N_36639);
nand U38258 (N_38258,N_36200,N_36844);
and U38259 (N_38259,N_37239,N_36105);
or U38260 (N_38260,N_37190,N_37245);
nor U38261 (N_38261,N_37120,N_37816);
nand U38262 (N_38262,N_37577,N_37317);
nor U38263 (N_38263,N_37181,N_36016);
nand U38264 (N_38264,N_37163,N_37779);
nand U38265 (N_38265,N_37496,N_37657);
nand U38266 (N_38266,N_36672,N_37902);
nor U38267 (N_38267,N_36492,N_36015);
nor U38268 (N_38268,N_37235,N_37751);
and U38269 (N_38269,N_37197,N_36963);
nor U38270 (N_38270,N_36705,N_36291);
xnor U38271 (N_38271,N_37579,N_36269);
nor U38272 (N_38272,N_36241,N_37312);
nand U38273 (N_38273,N_37086,N_37527);
and U38274 (N_38274,N_36365,N_36423);
nor U38275 (N_38275,N_36530,N_36332);
and U38276 (N_38276,N_37072,N_36643);
nor U38277 (N_38277,N_36674,N_36754);
nor U38278 (N_38278,N_36973,N_37293);
or U38279 (N_38279,N_37615,N_37809);
xnor U38280 (N_38280,N_36338,N_36152);
and U38281 (N_38281,N_37850,N_36739);
and U38282 (N_38282,N_37404,N_37800);
or U38283 (N_38283,N_37262,N_37826);
nor U38284 (N_38284,N_36974,N_36473);
and U38285 (N_38285,N_36517,N_37348);
and U38286 (N_38286,N_36569,N_37078);
or U38287 (N_38287,N_37003,N_36756);
nand U38288 (N_38288,N_37659,N_37683);
nand U38289 (N_38289,N_36149,N_36950);
and U38290 (N_38290,N_36260,N_36410);
and U38291 (N_38291,N_37939,N_37823);
and U38292 (N_38292,N_36334,N_36657);
or U38293 (N_38293,N_36168,N_37807);
nand U38294 (N_38294,N_37763,N_37336);
nand U38295 (N_38295,N_37365,N_36287);
and U38296 (N_38296,N_37880,N_37927);
nor U38297 (N_38297,N_37738,N_37068);
or U38298 (N_38298,N_37280,N_37158);
xor U38299 (N_38299,N_36426,N_36689);
or U38300 (N_38300,N_36167,N_37726);
nor U38301 (N_38301,N_36226,N_37654);
nor U38302 (N_38302,N_36750,N_37069);
nor U38303 (N_38303,N_37733,N_37051);
nand U38304 (N_38304,N_36939,N_37422);
nor U38305 (N_38305,N_37634,N_36930);
or U38306 (N_38306,N_37096,N_36398);
xnor U38307 (N_38307,N_36714,N_37092);
nor U38308 (N_38308,N_36700,N_36403);
xor U38309 (N_38309,N_36745,N_36784);
nand U38310 (N_38310,N_37794,N_36173);
or U38311 (N_38311,N_37366,N_37480);
nand U38312 (N_38312,N_36645,N_37027);
or U38313 (N_38313,N_37400,N_37952);
nand U38314 (N_38314,N_37612,N_36693);
and U38315 (N_38315,N_37044,N_37222);
and U38316 (N_38316,N_37347,N_36295);
nand U38317 (N_38317,N_37747,N_36055);
or U38318 (N_38318,N_37947,N_37038);
nand U38319 (N_38319,N_36348,N_37041);
nand U38320 (N_38320,N_37621,N_36631);
or U38321 (N_38321,N_36706,N_36023);
and U38322 (N_38322,N_37173,N_37483);
and U38323 (N_38323,N_36872,N_37381);
and U38324 (N_38324,N_36987,N_37343);
nor U38325 (N_38325,N_37505,N_37519);
nand U38326 (N_38326,N_36659,N_36433);
nor U38327 (N_38327,N_37133,N_37744);
or U38328 (N_38328,N_36992,N_36715);
nor U38329 (N_38329,N_37984,N_37694);
and U38330 (N_38330,N_37828,N_36874);
and U38331 (N_38331,N_36668,N_37740);
and U38332 (N_38332,N_37304,N_37138);
nand U38333 (N_38333,N_36145,N_37288);
and U38334 (N_38334,N_37195,N_37835);
nor U38335 (N_38335,N_36189,N_36808);
nand U38336 (N_38336,N_37427,N_36174);
or U38337 (N_38337,N_37350,N_37164);
or U38338 (N_38338,N_37836,N_37777);
nand U38339 (N_38339,N_37795,N_36855);
nor U38340 (N_38340,N_37508,N_37856);
or U38341 (N_38341,N_36486,N_37891);
nor U38342 (N_38342,N_37315,N_37106);
nand U38343 (N_38343,N_37953,N_37306);
nor U38344 (N_38344,N_36547,N_36736);
nand U38345 (N_38345,N_37813,N_36953);
nor U38346 (N_38346,N_36134,N_37821);
and U38347 (N_38347,N_36204,N_36421);
nor U38348 (N_38348,N_37429,N_37653);
nand U38349 (N_38349,N_37892,N_37271);
nor U38350 (N_38350,N_36565,N_37652);
nor U38351 (N_38351,N_37289,N_36841);
nor U38352 (N_38352,N_36944,N_36994);
or U38353 (N_38353,N_37417,N_36075);
nor U38354 (N_38354,N_37674,N_37854);
nor U38355 (N_38355,N_36976,N_37906);
or U38356 (N_38356,N_37582,N_37771);
nor U38357 (N_38357,N_36201,N_36532);
nor U38358 (N_38358,N_36548,N_37099);
nand U38359 (N_38359,N_37989,N_37471);
nor U38360 (N_38360,N_36614,N_36908);
nand U38361 (N_38361,N_36806,N_37554);
and U38362 (N_38362,N_36585,N_36864);
nand U38363 (N_38363,N_36261,N_36286);
and U38364 (N_38364,N_36388,N_36558);
and U38365 (N_38365,N_36109,N_37911);
or U38366 (N_38366,N_36247,N_36505);
or U38367 (N_38367,N_36202,N_37080);
and U38368 (N_38368,N_37524,N_36884);
or U38369 (N_38369,N_37817,N_37510);
nand U38370 (N_38370,N_36343,N_37790);
and U38371 (N_38371,N_37796,N_36341);
or U38372 (N_38372,N_36155,N_37246);
and U38373 (N_38373,N_37392,N_37708);
and U38374 (N_38374,N_37415,N_37752);
nor U38375 (N_38375,N_36588,N_36846);
and U38376 (N_38376,N_37839,N_37851);
nor U38377 (N_38377,N_36242,N_37588);
and U38378 (N_38378,N_36962,N_36231);
nor U38379 (N_38379,N_37520,N_37955);
and U38380 (N_38380,N_37673,N_36463);
or U38381 (N_38381,N_37253,N_37178);
nor U38382 (N_38382,N_36917,N_36143);
nand U38383 (N_38383,N_36961,N_37018);
xnor U38384 (N_38384,N_37274,N_37160);
and U38385 (N_38385,N_36626,N_36744);
or U38386 (N_38386,N_36319,N_37016);
nand U38387 (N_38387,N_36004,N_36883);
nor U38388 (N_38388,N_36998,N_37651);
nand U38389 (N_38389,N_36586,N_36681);
nor U38390 (N_38390,N_37376,N_36707);
and U38391 (N_38391,N_36629,N_37413);
and U38392 (N_38392,N_36488,N_37544);
nor U38393 (N_38393,N_36765,N_37569);
nand U38394 (N_38394,N_36063,N_37394);
nand U38395 (N_38395,N_36333,N_36458);
nor U38396 (N_38396,N_37265,N_36807);
nand U38397 (N_38397,N_37349,N_36190);
nor U38398 (N_38398,N_37076,N_36136);
nand U38399 (N_38399,N_36361,N_36820);
nor U38400 (N_38400,N_36288,N_36667);
or U38401 (N_38401,N_36342,N_37159);
nor U38402 (N_38402,N_36593,N_37565);
and U38403 (N_38403,N_36429,N_37640);
nor U38404 (N_38404,N_36704,N_36142);
and U38405 (N_38405,N_36957,N_37995);
and U38406 (N_38406,N_36132,N_37380);
or U38407 (N_38407,N_36811,N_37805);
xor U38408 (N_38408,N_37273,N_36825);
and U38409 (N_38409,N_37540,N_37325);
or U38410 (N_38410,N_37888,N_36759);
xor U38411 (N_38411,N_37558,N_37863);
or U38412 (N_38412,N_36465,N_36924);
nor U38413 (N_38413,N_37206,N_37351);
nand U38414 (N_38414,N_37876,N_36723);
nand U38415 (N_38415,N_37170,N_37489);
or U38416 (N_38416,N_36376,N_36382);
nand U38417 (N_38417,N_37829,N_37290);
nor U38418 (N_38418,N_36664,N_37184);
or U38419 (N_38419,N_37719,N_36562);
and U38420 (N_38420,N_37101,N_36871);
and U38421 (N_38421,N_36859,N_37887);
or U38422 (N_38422,N_36472,N_37898);
and U38423 (N_38423,N_36178,N_36721);
nand U38424 (N_38424,N_37176,N_37529);
nand U38425 (N_38425,N_37865,N_36237);
or U38426 (N_38426,N_37077,N_37287);
nor U38427 (N_38427,N_37113,N_36405);
nor U38428 (N_38428,N_36669,N_36144);
xnor U38429 (N_38429,N_37174,N_36717);
nor U38430 (N_38430,N_37874,N_36975);
or U38431 (N_38431,N_36464,N_36238);
nor U38432 (N_38432,N_36097,N_37169);
nand U38433 (N_38433,N_37762,N_37905);
nand U38434 (N_38434,N_37025,N_37442);
and U38435 (N_38435,N_36373,N_37950);
nand U38436 (N_38436,N_37295,N_37012);
nor U38437 (N_38437,N_37951,N_37214);
or U38438 (N_38438,N_36746,N_37499);
nand U38439 (N_38439,N_37567,N_37690);
nor U38440 (N_38440,N_36021,N_36459);
nand U38441 (N_38441,N_37431,N_36302);
nand U38442 (N_38442,N_36223,N_36428);
nand U38443 (N_38443,N_37141,N_36159);
nor U38444 (N_38444,N_36826,N_37241);
nor U38445 (N_38445,N_36407,N_37581);
and U38446 (N_38446,N_37678,N_36818);
and U38447 (N_38447,N_37391,N_36315);
nor U38448 (N_38448,N_36814,N_36430);
nor U38449 (N_38449,N_37215,N_36563);
or U38450 (N_38450,N_36686,N_36366);
nor U38451 (N_38451,N_37049,N_36219);
or U38452 (N_38452,N_36698,N_37401);
nor U38453 (N_38453,N_36590,N_36782);
nand U38454 (N_38454,N_36249,N_36863);
or U38455 (N_38455,N_36893,N_37297);
and U38456 (N_38456,N_37418,N_36390);
nor U38457 (N_38457,N_36307,N_36424);
nand U38458 (N_38458,N_36892,N_36925);
nor U38459 (N_38459,N_36919,N_36849);
or U38460 (N_38460,N_36794,N_36330);
nor U38461 (N_38461,N_37448,N_36946);
nand U38462 (N_38462,N_36126,N_37321);
nor U38463 (N_38463,N_36019,N_36531);
nor U38464 (N_38464,N_36833,N_37979);
or U38465 (N_38465,N_36567,N_36114);
nor U38466 (N_38466,N_37548,N_37398);
and U38467 (N_38467,N_36519,N_37956);
nor U38468 (N_38468,N_37537,N_36125);
nand U38469 (N_38469,N_37845,N_37664);
nand U38470 (N_38470,N_36581,N_36890);
nand U38471 (N_38471,N_36006,N_36821);
nor U38472 (N_38472,N_36761,N_36678);
and U38473 (N_38473,N_37032,N_37119);
nand U38474 (N_38474,N_36197,N_37689);
nand U38475 (N_38475,N_37737,N_37909);
and U38476 (N_38476,N_36422,N_36412);
nand U38477 (N_38477,N_37675,N_37229);
nor U38478 (N_38478,N_36401,N_36053);
or U38479 (N_38479,N_36606,N_36089);
nor U38480 (N_38480,N_37873,N_37725);
and U38481 (N_38481,N_37242,N_37301);
and U38482 (N_38482,N_36916,N_36217);
nor U38483 (N_38483,N_37208,N_36927);
nand U38484 (N_38484,N_36662,N_36860);
nand U38485 (N_38485,N_36543,N_36474);
nor U38486 (N_38486,N_36196,N_37593);
nor U38487 (N_38487,N_37871,N_37819);
nand U38488 (N_38488,N_36836,N_36769);
or U38489 (N_38489,N_37676,N_36650);
nor U38490 (N_38490,N_36290,N_37200);
nand U38491 (N_38491,N_36848,N_37860);
nor U38492 (N_38492,N_37698,N_36680);
and U38493 (N_38493,N_37412,N_37473);
nor U38494 (N_38494,N_37772,N_36914);
nand U38495 (N_38495,N_36901,N_37907);
and U38496 (N_38496,N_37611,N_37447);
nand U38497 (N_38497,N_36526,N_37421);
nand U38498 (N_38498,N_36767,N_37470);
or U38499 (N_38499,N_37859,N_37601);
nor U38500 (N_38500,N_37893,N_36577);
nand U38501 (N_38501,N_36044,N_36796);
and U38502 (N_38502,N_36635,N_37922);
nor U38503 (N_38503,N_37492,N_36726);
or U38504 (N_38504,N_37827,N_37713);
nor U38505 (N_38505,N_36298,N_36703);
or U38506 (N_38506,N_36072,N_36022);
and U38507 (N_38507,N_37010,N_36413);
nor U38508 (N_38508,N_37812,N_37359);
xor U38509 (N_38509,N_36730,N_37783);
nor U38510 (N_38510,N_36028,N_37538);
xor U38511 (N_38511,N_36267,N_36501);
or U38512 (N_38512,N_36487,N_37571);
nor U38513 (N_38513,N_36166,N_37935);
nor U38514 (N_38514,N_37833,N_36762);
or U38515 (N_38515,N_37070,N_36617);
and U38516 (N_38516,N_36857,N_36600);
and U38517 (N_38517,N_37849,N_36207);
or U38518 (N_38518,N_37884,N_36185);
nand U38519 (N_38519,N_36104,N_36059);
or U38520 (N_38520,N_36949,N_36176);
nand U38521 (N_38521,N_37626,N_36203);
nor U38522 (N_38522,N_37193,N_37606);
nand U38523 (N_38523,N_36570,N_37420);
or U38524 (N_38524,N_37858,N_36660);
and U38525 (N_38525,N_36537,N_37937);
or U38526 (N_38526,N_36557,N_36303);
nor U38527 (N_38527,N_37655,N_36491);
nor U38528 (N_38528,N_36747,N_36862);
nor U38529 (N_38529,N_36737,N_37944);
nand U38530 (N_38530,N_37852,N_36881);
nand U38531 (N_38531,N_36748,N_37369);
and U38532 (N_38532,N_37091,N_37362);
nand U38533 (N_38533,N_36120,N_36160);
nand U38534 (N_38534,N_37973,N_37310);
and U38535 (N_38535,N_36886,N_37402);
and U38536 (N_38536,N_36510,N_36711);
or U38537 (N_38537,N_36966,N_37378);
and U38538 (N_38538,N_37693,N_36434);
or U38539 (N_38539,N_37531,N_37971);
nand U38540 (N_38540,N_37272,N_37283);
nand U38541 (N_38541,N_37085,N_37205);
or U38542 (N_38542,N_37881,N_37311);
nand U38543 (N_38543,N_36476,N_37477);
nor U38544 (N_38544,N_36503,N_36058);
nor U38545 (N_38545,N_37047,N_36823);
and U38546 (N_38546,N_37991,N_37598);
and U38547 (N_38547,N_37710,N_36283);
nor U38548 (N_38548,N_36119,N_36683);
nand U38549 (N_38549,N_36462,N_37963);
or U38550 (N_38550,N_36899,N_36943);
nand U38551 (N_38551,N_37648,N_37696);
nand U38552 (N_38552,N_36509,N_37112);
or U38553 (N_38553,N_36455,N_36937);
nand U38554 (N_38554,N_37426,N_37474);
and U38555 (N_38555,N_36624,N_36576);
nor U38556 (N_38556,N_36566,N_36183);
or U38557 (N_38557,N_36071,N_37065);
or U38558 (N_38558,N_36266,N_36047);
and U38559 (N_38559,N_37028,N_36980);
nor U38560 (N_38560,N_36640,N_37885);
nor U38561 (N_38561,N_37526,N_37623);
and U38562 (N_38562,N_36583,N_37389);
nand U38563 (N_38563,N_36870,N_36477);
or U38564 (N_38564,N_37093,N_37223);
nand U38565 (N_38565,N_36983,N_37649);
nor U38566 (N_38566,N_36793,N_36851);
or U38567 (N_38567,N_36573,N_36632);
or U38568 (N_38568,N_37776,N_37650);
or U38569 (N_38569,N_37660,N_36340);
or U38570 (N_38570,N_37687,N_37915);
nor U38571 (N_38571,N_36400,N_37756);
and U38572 (N_38572,N_37073,N_37760);
nand U38573 (N_38573,N_36386,N_36608);
nand U38574 (N_38574,N_36498,N_36947);
nor U38575 (N_38575,N_37721,N_36215);
nor U38576 (N_38576,N_37472,N_36027);
or U38577 (N_38577,N_37043,N_37192);
nor U38578 (N_38578,N_37607,N_37142);
nand U38579 (N_38579,N_36112,N_37316);
nand U38580 (N_38580,N_37637,N_37050);
or U38581 (N_38581,N_37168,N_36809);
and U38582 (N_38582,N_37982,N_37344);
or U38583 (N_38583,N_37831,N_36020);
nand U38584 (N_38584,N_36276,N_36904);
nor U38585 (N_38585,N_37082,N_36896);
nand U38586 (N_38586,N_37166,N_36891);
nand U38587 (N_38587,N_36653,N_36098);
or U38588 (N_38588,N_36301,N_36272);
and U38589 (N_38589,N_37785,N_37278);
or U38590 (N_38590,N_37661,N_36494);
and U38591 (N_38591,N_37502,N_36905);
or U38592 (N_38592,N_36011,N_36776);
and U38593 (N_38593,N_37578,N_36070);
or U38594 (N_38594,N_36030,N_36277);
nand U38595 (N_38595,N_37889,N_37806);
or U38596 (N_38596,N_37342,N_37154);
nor U38597 (N_38597,N_36451,N_37742);
and U38598 (N_38598,N_36171,N_36271);
xnor U38599 (N_38599,N_37030,N_37244);
and U38600 (N_38600,N_36951,N_36244);
nor U38601 (N_38601,N_37684,N_36996);
or U38602 (N_38602,N_37778,N_36344);
and U38603 (N_38603,N_36392,N_37263);
and U38604 (N_38604,N_36205,N_37481);
nor U38605 (N_38605,N_36066,N_37008);
or U38606 (N_38606,N_37118,N_37869);
or U38607 (N_38607,N_36615,N_36453);
nand U38608 (N_38608,N_37276,N_36789);
and U38609 (N_38609,N_36049,N_37981);
nand U38610 (N_38610,N_37294,N_37994);
or U38611 (N_38611,N_36838,N_36803);
and U38612 (N_38612,N_37919,N_37042);
and U38613 (N_38613,N_36352,N_37225);
nand U38614 (N_38614,N_37631,N_36191);
and U38615 (N_38615,N_37045,N_37387);
nand U38616 (N_38616,N_37467,N_37949);
and U38617 (N_38617,N_37185,N_36713);
and U38618 (N_38618,N_36425,N_37961);
nor U38619 (N_38619,N_37996,N_36515);
nand U38620 (N_38620,N_36214,N_36444);
or U38621 (N_38621,N_36435,N_37798);
or U38622 (N_38622,N_37924,N_37335);
or U38623 (N_38623,N_37552,N_36449);
nand U38624 (N_38624,N_36559,N_37518);
and U38625 (N_38625,N_37539,N_37617);
or U38626 (N_38626,N_37264,N_37671);
nor U38627 (N_38627,N_37011,N_37792);
nand U38628 (N_38628,N_36677,N_36988);
nor U38629 (N_38629,N_37260,N_36797);
nand U38630 (N_38630,N_36802,N_36225);
or U38631 (N_38631,N_37019,N_37423);
or U38632 (N_38632,N_36795,N_36033);
nor U38633 (N_38633,N_36719,N_37484);
and U38634 (N_38634,N_37218,N_37451);
nor U38635 (N_38635,N_37867,N_36466);
nand U38636 (N_38636,N_37270,N_36229);
nor U38637 (N_38637,N_36454,N_37717);
and U38638 (N_38638,N_37493,N_36945);
and U38639 (N_38639,N_37232,N_36195);
and U38640 (N_38640,N_37331,N_36452);
nand U38641 (N_38641,N_36265,N_36960);
nor U38642 (N_38642,N_37458,N_36415);
nor U38643 (N_38643,N_36321,N_37644);
nand U38644 (N_38644,N_36471,N_36065);
nor U38645 (N_38645,N_36766,N_36206);
or U38646 (N_38646,N_36741,N_36647);
and U38647 (N_38647,N_36035,N_37114);
nand U38648 (N_38648,N_37580,N_37221);
or U38649 (N_38649,N_36935,N_37978);
or U38650 (N_38650,N_37151,N_37627);
nor U38651 (N_38651,N_36997,N_37990);
or U38652 (N_38652,N_36299,N_37147);
and U38653 (N_38653,N_37319,N_37853);
and U38654 (N_38654,N_36968,N_36743);
or U38655 (N_38655,N_36989,N_36151);
nor U38656 (N_38656,N_37248,N_37910);
or U38657 (N_38657,N_37912,N_37459);
or U38658 (N_38658,N_37435,N_36731);
and U38659 (N_38659,N_37324,N_36443);
nand U38660 (N_38660,N_37432,N_36772);
nor U38661 (N_38661,N_36161,N_36799);
and U38662 (N_38662,N_36218,N_37475);
nand U38663 (N_38663,N_37445,N_36117);
nor U38664 (N_38664,N_36734,N_36311);
nor U38665 (N_38665,N_36618,N_37217);
and U38666 (N_38666,N_37700,N_36470);
or U38667 (N_38667,N_36383,N_36489);
nor U38668 (N_38668,N_36555,N_37846);
and U38669 (N_38669,N_37677,N_36478);
or U38670 (N_38670,N_36781,N_36483);
or U38671 (N_38671,N_37355,N_36211);
nor U38672 (N_38672,N_37416,N_37641);
and U38673 (N_38673,N_36535,N_36419);
nor U38674 (N_38674,N_37895,N_36554);
nand U38675 (N_38675,N_37358,N_37063);
or U38676 (N_38676,N_36533,N_36331);
nand U38677 (N_38677,N_36248,N_37780);
nor U38678 (N_38678,N_37699,N_36556);
nand U38679 (N_38679,N_37804,N_37408);
xor U38680 (N_38680,N_36395,N_36447);
and U38681 (N_38681,N_36228,N_37379);
and U38682 (N_38682,N_36877,N_37959);
nand U38683 (N_38683,N_37139,N_36427);
and U38684 (N_38684,N_37026,N_36096);
nand U38685 (N_38685,N_37837,N_37962);
nor U38686 (N_38686,N_37269,N_37202);
nor U38687 (N_38687,N_37553,N_36915);
and U38688 (N_38688,N_36118,N_37701);
nor U38689 (N_38689,N_36928,N_37231);
nand U38690 (N_38690,N_37568,N_37487);
and U38691 (N_38691,N_36208,N_36077);
nor U38692 (N_38692,N_37757,N_36026);
or U38693 (N_38693,N_37428,N_37357);
and U38694 (N_38694,N_36273,N_37522);
and U38695 (N_38695,N_36673,N_37130);
xor U38696 (N_38696,N_37254,N_36043);
nand U38697 (N_38697,N_36018,N_36709);
or U38698 (N_38698,N_36131,N_36432);
nor U38699 (N_38699,N_36644,N_36193);
nor U38700 (N_38700,N_37759,N_37450);
nor U38701 (N_38701,N_36441,N_37111);
or U38702 (N_38702,N_37328,N_37006);
or U38703 (N_38703,N_36591,N_36906);
and U38704 (N_38704,N_37333,N_36182);
nand U38705 (N_38705,N_36786,N_37466);
or U38706 (N_38706,N_36878,N_37409);
or U38707 (N_38707,N_36399,N_36753);
nand U38708 (N_38708,N_37681,N_36895);
or U38709 (N_38709,N_36083,N_36670);
nor U38710 (N_38710,N_37338,N_37476);
nand U38711 (N_38711,N_37670,N_36948);
nor U38712 (N_38712,N_37878,N_36885);
or U38713 (N_38713,N_36312,N_36900);
and U38714 (N_38714,N_36468,N_37444);
and U38715 (N_38715,N_37052,N_37886);
or U38716 (N_38716,N_36284,N_37551);
or U38717 (N_38717,N_37037,N_37842);
or U38718 (N_38718,N_36634,N_37918);
or U38719 (N_38719,N_37286,N_37199);
and U38720 (N_38720,N_36993,N_37196);
nand U38721 (N_38721,N_37146,N_37036);
and U38722 (N_38722,N_37132,N_36236);
nor U38723 (N_38723,N_37832,N_37597);
and U38724 (N_38724,N_36009,N_36010);
or U38725 (N_38725,N_36187,N_37936);
and U38726 (N_38726,N_37642,N_36220);
nand U38727 (N_38727,N_36057,N_36153);
nor U38728 (N_38728,N_36508,N_37216);
or U38729 (N_38729,N_37573,N_37503);
nor U38730 (N_38730,N_36414,N_36696);
nor U38731 (N_38731,N_37259,N_36822);
nand U38732 (N_38732,N_37628,N_36627);
or U38733 (N_38733,N_36628,N_36840);
and U38734 (N_38734,N_36599,N_36460);
or U38735 (N_38735,N_36546,N_36923);
xor U38736 (N_38736,N_37933,N_36868);
and U38737 (N_38737,N_36074,N_36763);
and U38738 (N_38738,N_37430,N_36245);
or U38739 (N_38739,N_37620,N_37543);
nand U38740 (N_38740,N_36545,N_36684);
and U38741 (N_38741,N_37802,N_37585);
nand U38742 (N_38742,N_37084,N_36113);
nor U38743 (N_38743,N_37669,N_37329);
nor U38744 (N_38744,N_36339,N_37957);
or U38745 (N_38745,N_36971,N_37249);
or U38746 (N_38746,N_37788,N_36507);
and U38747 (N_38747,N_37509,N_37374);
and U38748 (N_38748,N_36602,N_36322);
nor U38749 (N_38749,N_37009,N_36812);
or U38750 (N_38750,N_36005,N_37109);
and U38751 (N_38751,N_37530,N_36264);
nor U38752 (N_38752,N_36450,N_37022);
nor U38753 (N_38753,N_37946,N_37020);
nand U38754 (N_38754,N_36480,N_36157);
or U38755 (N_38755,N_36351,N_37213);
and U38756 (N_38756,N_37695,N_37300);
and U38757 (N_38757,N_36251,N_36671);
nand U38758 (N_38758,N_36076,N_37862);
nor U38759 (N_38759,N_37449,N_37596);
nor U38760 (N_38760,N_37095,N_36589);
nand U38761 (N_38761,N_36835,N_37261);
nand U38762 (N_38762,N_36106,N_36986);
nor U38763 (N_38763,N_37257,N_36354);
nor U38764 (N_38764,N_36256,N_36146);
nand U38765 (N_38765,N_36972,N_37591);
nand U38766 (N_38766,N_36320,N_37667);
and U38767 (N_38767,N_37145,N_37980);
nand U38768 (N_38768,N_37586,N_37712);
nor U38769 (N_38769,N_37534,N_37438);
nand U38770 (N_38770,N_37958,N_36107);
or U38771 (N_38771,N_36638,N_36420);
and U38772 (N_38772,N_37736,N_37549);
nand U38773 (N_38773,N_37057,N_36130);
or U38774 (N_38774,N_37556,N_36518);
nor U38775 (N_38775,N_37024,N_37968);
nor U38776 (N_38776,N_37439,N_37108);
and U38777 (N_38777,N_37974,N_37609);
nor U38778 (N_38778,N_36955,N_37296);
and U38779 (N_38779,N_36712,N_36539);
and U38780 (N_38780,N_37090,N_36158);
nor U38781 (N_38781,N_37815,N_36969);
nand U38782 (N_38782,N_36170,N_37716);
nand U38783 (N_38783,N_37128,N_37299);
xor U38784 (N_38784,N_37307,N_36954);
or U38785 (N_38785,N_37913,N_36637);
or U38786 (N_38786,N_36834,N_37486);
nor U38787 (N_38787,N_36188,N_37773);
or U38788 (N_38788,N_37180,N_36967);
nand U38789 (N_38789,N_37647,N_37616);
nor U38790 (N_38790,N_36417,N_36641);
nand U38791 (N_38791,N_37921,N_37498);
nand U38792 (N_38792,N_36831,N_36484);
or U38793 (N_38793,N_37126,N_37872);
nand U38794 (N_38794,N_36502,N_36309);
xnor U38795 (N_38795,N_36790,N_37975);
or U38796 (N_38796,N_36922,N_36865);
and U38797 (N_38797,N_36656,N_37599);
or U38798 (N_38798,N_37396,N_36725);
nand U38799 (N_38799,N_37462,N_37015);
and U38800 (N_38800,N_36181,N_36234);
or U38801 (N_38801,N_36442,N_37268);
nor U38802 (N_38802,N_36701,N_36274);
or U38803 (N_38803,N_36702,N_37382);
or U38804 (N_38804,N_37425,N_37059);
or U38805 (N_38805,N_37686,N_37282);
nor U38806 (N_38806,N_36358,N_37258);
or U38807 (N_38807,N_36073,N_37441);
or U38808 (N_38808,N_37461,N_37226);
nand U38809 (N_38809,N_36813,N_36210);
xnor U38810 (N_38810,N_37346,N_37938);
nand U38811 (N_38811,N_36511,N_37954);
nand U38812 (N_38812,N_37123,N_36598);
or U38813 (N_38813,N_37868,N_37204);
nand U38814 (N_38814,N_37934,N_36037);
or U38815 (N_38815,N_37302,N_37900);
and U38816 (N_38816,N_37764,N_36977);
nor U38817 (N_38817,N_36192,N_36012);
and U38818 (N_38818,N_37367,N_37986);
nand U38819 (N_38819,N_37284,N_36894);
nand U38820 (N_38820,N_37722,N_36499);
xnor U38821 (N_38821,N_36616,N_37879);
or U38822 (N_38822,N_36536,N_36050);
nor U38823 (N_38823,N_36999,N_37745);
nor U38824 (N_38824,N_37224,N_37672);
nor U38825 (N_38825,N_36318,N_36278);
or U38826 (N_38826,N_37575,N_36879);
nor U38827 (N_38827,N_37243,N_36775);
or U38828 (N_38828,N_37662,N_37266);
nor U38829 (N_38829,N_37718,N_37252);
nand U38830 (N_38830,N_36408,N_36521);
nand U38831 (N_38831,N_37375,N_36135);
nor U38832 (N_38832,N_36067,N_36854);
or U38833 (N_38833,N_36690,N_37031);
nand U38834 (N_38834,N_37021,N_37967);
and U38835 (N_38835,N_37002,N_37883);
nand U38836 (N_38836,N_37013,N_36596);
or U38837 (N_38837,N_37600,N_36897);
or U38838 (N_38838,N_37005,N_37364);
nand U38839 (N_38839,N_37456,N_37330);
and U38840 (N_38840,N_37277,N_36594);
and U38841 (N_38841,N_37668,N_37046);
or U38842 (N_38842,N_36329,N_37399);
nor U38843 (N_38843,N_36111,N_36733);
nor U38844 (N_38844,N_36086,N_37137);
and U38845 (N_38845,N_36221,N_36370);
and U38846 (N_38846,N_37811,N_36815);
and U38847 (N_38847,N_36128,N_36845);
or U38848 (N_38848,N_37156,N_36560);
nand U38849 (N_38849,N_37870,N_37635);
or U38850 (N_38850,N_37157,N_37434);
xor U38851 (N_38851,N_36101,N_36658);
and U38852 (N_38852,N_36888,N_37632);
nor U38853 (N_38853,N_37643,N_37066);
or U38854 (N_38854,N_37739,N_36163);
or U38855 (N_38855,N_36087,N_37926);
nor U38856 (N_38856,N_36534,N_37117);
or U38857 (N_38857,N_36964,N_36695);
or U38858 (N_38858,N_37155,N_37121);
or U38859 (N_38859,N_36325,N_36239);
or U38860 (N_38860,N_36062,N_36527);
or U38861 (N_38861,N_37516,N_36263);
or U38862 (N_38862,N_36933,N_36694);
nand U38863 (N_38863,N_37327,N_37326);
nand U38864 (N_38864,N_36990,N_37786);
nor U38865 (N_38865,N_36336,N_36224);
nor U38866 (N_38866,N_37731,N_37098);
and U38867 (N_38867,N_36985,N_37115);
nand U38868 (N_38868,N_37916,N_36481);
nor U38869 (N_38869,N_37993,N_37506);
xor U38870 (N_38870,N_36314,N_36655);
or U38871 (N_38871,N_37048,N_37511);
or U38872 (N_38872,N_37964,N_37706);
and U38873 (N_38873,N_37035,N_37656);
and U38874 (N_38874,N_36568,N_36175);
and U38875 (N_38875,N_36758,N_36549);
and U38876 (N_38876,N_36858,N_37711);
and U38877 (N_38877,N_36041,N_37165);
nand U38878 (N_38878,N_37914,N_36172);
and U38879 (N_38879,N_36054,N_37171);
xor U38880 (N_38880,N_37267,N_36133);
nand U38881 (N_38881,N_37465,N_37363);
nand U38882 (N_38882,N_37801,N_37373);
and U38883 (N_38883,N_37143,N_37131);
nand U38884 (N_38884,N_36604,N_36716);
nor U38885 (N_38885,N_37500,N_36391);
and U38886 (N_38886,N_36180,N_37847);
nand U38887 (N_38887,N_36232,N_36337);
or U38888 (N_38888,N_37613,N_36800);
xor U38889 (N_38889,N_37189,N_36652);
or U38890 (N_38890,N_36198,N_36682);
and U38891 (N_38891,N_36691,N_37729);
xor U38892 (N_38892,N_36150,N_37341);
or U38893 (N_38893,N_36828,N_36164);
and U38894 (N_38894,N_36317,N_36389);
or U38895 (N_38895,N_37150,N_36122);
nand U38896 (N_38896,N_36572,N_36882);
and U38897 (N_38897,N_37513,N_36082);
or U38898 (N_38898,N_36817,N_36791);
and U38899 (N_38899,N_37161,N_37279);
and U38900 (N_38900,N_37219,N_37122);
or U38901 (N_38901,N_37897,N_37920);
nor U38902 (N_38902,N_36360,N_36538);
nor U38903 (N_38903,N_36982,N_37292);
and U38904 (N_38904,N_37987,N_36718);
nand U38905 (N_38905,N_36216,N_36045);
or U38906 (N_38906,N_37446,N_37337);
nor U38907 (N_38907,N_36708,N_36827);
nor U38908 (N_38908,N_37203,N_36773);
nand U38909 (N_38909,N_36642,N_36574);
or U38910 (N_38910,N_36942,N_36469);
and U38911 (N_38911,N_37894,N_37162);
nand U38912 (N_38912,N_37970,N_37191);
or U38913 (N_38913,N_37182,N_36485);
nor U38914 (N_38914,N_36940,N_36416);
nor U38915 (N_38915,N_36584,N_36431);
or U38916 (N_38916,N_36497,N_36029);
nand U38917 (N_38917,N_36542,N_36162);
nor U38918 (N_38918,N_37630,N_36289);
and U38919 (N_38919,N_37105,N_36780);
nand U38920 (N_38920,N_37087,N_37857);
and U38921 (N_38921,N_36528,N_37240);
nor U38922 (N_38922,N_36611,N_37275);
nand U38923 (N_38923,N_37220,N_36039);
and U38924 (N_38924,N_36912,N_36003);
nand U38925 (N_38925,N_36934,N_37594);
nor U38926 (N_38926,N_37803,N_37352);
and U38927 (N_38927,N_37097,N_36909);
and U38928 (N_38928,N_36308,N_36068);
nor U38929 (N_38929,N_37799,N_36920);
or U38930 (N_38930,N_37932,N_37383);
or U38931 (N_38931,N_36372,N_37715);
and U38932 (N_38932,N_37784,N_36514);
nor U38933 (N_38933,N_36084,N_36213);
nand U38934 (N_38934,N_37999,N_36051);
or U38935 (N_38935,N_37622,N_36687);
or U38936 (N_38936,N_37536,N_36649);
or U38937 (N_38937,N_36418,N_36255);
nand U38938 (N_38938,N_36194,N_36233);
and U38939 (N_38939,N_36138,N_36876);
nor U38940 (N_38940,N_36139,N_37210);
nand U38941 (N_38941,N_36771,N_36246);
or U38942 (N_38942,N_36438,N_36294);
and U38943 (N_38943,N_36110,N_36350);
and U38944 (N_38944,N_37758,N_37583);
or U38945 (N_38945,N_36297,N_37183);
nand U38946 (N_38946,N_37071,N_37497);
nor U38947 (N_38947,N_37928,N_37368);
nor U38948 (N_38948,N_37004,N_36512);
and U38949 (N_38949,N_36257,N_36409);
nor U38950 (N_38950,N_37083,N_36622);
or U38951 (N_38951,N_37903,N_37515);
or U38952 (N_38952,N_36601,N_37882);
and U38953 (N_38953,N_36913,N_36938);
and U38954 (N_38954,N_36610,N_37209);
or U38955 (N_38955,N_37825,N_37207);
and U38956 (N_38956,N_37124,N_37767);
and U38957 (N_38957,N_37149,N_37789);
and U38958 (N_38958,N_37067,N_37491);
and U38959 (N_38959,N_36551,N_36587);
and U38960 (N_38960,N_36088,N_36843);
nand U38961 (N_38961,N_37636,N_36513);
nand U38962 (N_38962,N_37808,N_37532);
and U38963 (N_38963,N_37768,N_36630);
nor U38964 (N_38964,N_37313,N_37029);
nor U38965 (N_38965,N_37864,N_36323);
nand U38966 (N_38966,N_37820,N_36179);
or U38967 (N_38967,N_37840,N_37709);
or U38968 (N_38968,N_36359,N_37608);
and U38969 (N_38969,N_37440,N_36889);
and U38970 (N_38970,N_36116,N_37340);
nor U38971 (N_38971,N_37323,N_37561);
nand U38972 (N_38972,N_37385,N_37501);
nor U38973 (N_38973,N_37298,N_36479);
nand U38974 (N_38974,N_37810,N_37595);
nor U38975 (N_38975,N_36085,N_37490);
nor U38976 (N_38976,N_37638,N_36099);
nor U38977 (N_38977,N_37198,N_37797);
nand U38978 (N_38978,N_37703,N_37574);
or U38979 (N_38979,N_36609,N_36402);
nor U38980 (N_38980,N_36378,N_37787);
or U38981 (N_38981,N_36578,N_36235);
or U38982 (N_38982,N_37791,N_36605);
and U38983 (N_38983,N_37479,N_36002);
nor U38984 (N_38984,N_37478,N_37407);
and U38985 (N_38985,N_36296,N_36280);
and U38986 (N_38986,N_36571,N_36816);
nor U38987 (N_38987,N_36824,N_36165);
and U38988 (N_38988,N_36852,N_37749);
and U38989 (N_38989,N_37770,N_37039);
nand U38990 (N_38990,N_36379,N_36384);
and U38991 (N_38991,N_37356,N_36380);
nand U38992 (N_38992,N_36625,N_37452);
nor U38993 (N_38993,N_36603,N_37397);
or U38994 (N_38994,N_37454,N_37735);
or U38995 (N_38995,N_36254,N_36755);
nor U38996 (N_38996,N_36253,N_36377);
and U38997 (N_38997,N_36060,N_37732);
nand U38998 (N_38998,N_36679,N_36804);
nor U38999 (N_38999,N_36829,N_37144);
or U39000 (N_39000,N_36241,N_36105);
or U39001 (N_39001,N_36708,N_37047);
and U39002 (N_39002,N_36924,N_36826);
nor U39003 (N_39003,N_36345,N_37727);
xor U39004 (N_39004,N_37323,N_36126);
or U39005 (N_39005,N_36632,N_36037);
or U39006 (N_39006,N_36272,N_37181);
nand U39007 (N_39007,N_36246,N_37603);
and U39008 (N_39008,N_37057,N_36406);
and U39009 (N_39009,N_37358,N_36539);
nor U39010 (N_39010,N_37888,N_36042);
nand U39011 (N_39011,N_36465,N_37870);
or U39012 (N_39012,N_36788,N_36487);
and U39013 (N_39013,N_36809,N_36595);
nor U39014 (N_39014,N_36228,N_36216);
nor U39015 (N_39015,N_37016,N_36476);
nor U39016 (N_39016,N_36574,N_36262);
nand U39017 (N_39017,N_36147,N_37633);
and U39018 (N_39018,N_37619,N_36149);
nand U39019 (N_39019,N_36889,N_36175);
nand U39020 (N_39020,N_37339,N_37812);
nor U39021 (N_39021,N_36711,N_36507);
nand U39022 (N_39022,N_37953,N_37244);
nor U39023 (N_39023,N_37448,N_36251);
and U39024 (N_39024,N_37181,N_37495);
or U39025 (N_39025,N_36228,N_37237);
and U39026 (N_39026,N_37112,N_37867);
or U39027 (N_39027,N_37589,N_37281);
or U39028 (N_39028,N_36687,N_37348);
and U39029 (N_39029,N_36088,N_37726);
and U39030 (N_39030,N_36049,N_36327);
or U39031 (N_39031,N_36669,N_37342);
or U39032 (N_39032,N_37599,N_37135);
nand U39033 (N_39033,N_36595,N_37704);
nor U39034 (N_39034,N_37807,N_37908);
nor U39035 (N_39035,N_36015,N_36150);
or U39036 (N_39036,N_37022,N_37338);
nand U39037 (N_39037,N_37118,N_36347);
and U39038 (N_39038,N_36461,N_37646);
or U39039 (N_39039,N_36685,N_37660);
or U39040 (N_39040,N_36125,N_36328);
or U39041 (N_39041,N_37540,N_36821);
nand U39042 (N_39042,N_36325,N_36675);
and U39043 (N_39043,N_36693,N_37500);
and U39044 (N_39044,N_37462,N_36855);
or U39045 (N_39045,N_37798,N_37986);
or U39046 (N_39046,N_36157,N_37610);
and U39047 (N_39047,N_36049,N_36211);
and U39048 (N_39048,N_36511,N_37351);
nand U39049 (N_39049,N_37873,N_36194);
nand U39050 (N_39050,N_36531,N_37932);
and U39051 (N_39051,N_37659,N_37442);
and U39052 (N_39052,N_36674,N_37968);
and U39053 (N_39053,N_36691,N_37779);
and U39054 (N_39054,N_36989,N_37489);
nor U39055 (N_39055,N_37429,N_37846);
nand U39056 (N_39056,N_37635,N_36351);
nor U39057 (N_39057,N_36991,N_37607);
or U39058 (N_39058,N_36834,N_37378);
nor U39059 (N_39059,N_37107,N_37647);
or U39060 (N_39060,N_37560,N_37156);
and U39061 (N_39061,N_36567,N_36192);
nor U39062 (N_39062,N_36313,N_37505);
nand U39063 (N_39063,N_36040,N_36678);
or U39064 (N_39064,N_37734,N_37744);
nor U39065 (N_39065,N_37928,N_37641);
and U39066 (N_39066,N_37568,N_36463);
or U39067 (N_39067,N_37254,N_36520);
nor U39068 (N_39068,N_36110,N_37582);
nand U39069 (N_39069,N_36655,N_36620);
and U39070 (N_39070,N_37674,N_36826);
nand U39071 (N_39071,N_37379,N_36833);
and U39072 (N_39072,N_37075,N_36533);
and U39073 (N_39073,N_36233,N_36835);
nor U39074 (N_39074,N_37908,N_36137);
or U39075 (N_39075,N_36721,N_36794);
nand U39076 (N_39076,N_37800,N_37848);
and U39077 (N_39077,N_37409,N_37104);
and U39078 (N_39078,N_37541,N_37872);
nand U39079 (N_39079,N_36957,N_36969);
nand U39080 (N_39080,N_37881,N_36929);
nor U39081 (N_39081,N_36782,N_37384);
nand U39082 (N_39082,N_37515,N_37630);
xnor U39083 (N_39083,N_36862,N_36433);
nand U39084 (N_39084,N_37280,N_36499);
nand U39085 (N_39085,N_37488,N_36994);
or U39086 (N_39086,N_37894,N_37793);
or U39087 (N_39087,N_36503,N_36904);
nor U39088 (N_39088,N_36353,N_37033);
or U39089 (N_39089,N_37954,N_37794);
xor U39090 (N_39090,N_36247,N_36176);
nor U39091 (N_39091,N_37453,N_37362);
nand U39092 (N_39092,N_36264,N_37328);
or U39093 (N_39093,N_36565,N_36318);
nand U39094 (N_39094,N_37130,N_36393);
or U39095 (N_39095,N_36645,N_36917);
nor U39096 (N_39096,N_36479,N_37651);
nor U39097 (N_39097,N_36070,N_37221);
and U39098 (N_39098,N_36960,N_37019);
and U39099 (N_39099,N_36840,N_36561);
or U39100 (N_39100,N_37430,N_37439);
nand U39101 (N_39101,N_36995,N_36008);
nand U39102 (N_39102,N_37366,N_36936);
and U39103 (N_39103,N_36982,N_36524);
nor U39104 (N_39104,N_36738,N_37253);
nand U39105 (N_39105,N_36968,N_36593);
and U39106 (N_39106,N_37666,N_36583);
nor U39107 (N_39107,N_36880,N_37258);
xor U39108 (N_39108,N_36590,N_36767);
and U39109 (N_39109,N_37322,N_36346);
nor U39110 (N_39110,N_37648,N_36167);
nand U39111 (N_39111,N_36617,N_36535);
nand U39112 (N_39112,N_36387,N_36103);
nand U39113 (N_39113,N_37385,N_36185);
and U39114 (N_39114,N_37258,N_37614);
or U39115 (N_39115,N_36015,N_36187);
nor U39116 (N_39116,N_37035,N_37653);
and U39117 (N_39117,N_37292,N_36959);
nand U39118 (N_39118,N_37343,N_36484);
nor U39119 (N_39119,N_36692,N_37794);
and U39120 (N_39120,N_36029,N_37071);
nand U39121 (N_39121,N_37170,N_37681);
nand U39122 (N_39122,N_36488,N_36574);
and U39123 (N_39123,N_36800,N_37140);
and U39124 (N_39124,N_36847,N_37656);
or U39125 (N_39125,N_36692,N_36450);
or U39126 (N_39126,N_37347,N_37944);
and U39127 (N_39127,N_36613,N_36810);
or U39128 (N_39128,N_36071,N_37615);
and U39129 (N_39129,N_37668,N_36974);
nor U39130 (N_39130,N_36120,N_37885);
and U39131 (N_39131,N_37351,N_36084);
nor U39132 (N_39132,N_36159,N_36772);
nand U39133 (N_39133,N_36539,N_37379);
nand U39134 (N_39134,N_36084,N_36162);
and U39135 (N_39135,N_37056,N_36768);
or U39136 (N_39136,N_37662,N_36921);
nor U39137 (N_39137,N_37093,N_36361);
or U39138 (N_39138,N_36791,N_36849);
and U39139 (N_39139,N_37956,N_36751);
nor U39140 (N_39140,N_36664,N_36632);
nand U39141 (N_39141,N_37261,N_36877);
or U39142 (N_39142,N_36068,N_36965);
or U39143 (N_39143,N_36226,N_36803);
nand U39144 (N_39144,N_37210,N_36869);
or U39145 (N_39145,N_37576,N_37313);
nand U39146 (N_39146,N_37678,N_36540);
nand U39147 (N_39147,N_36770,N_37917);
nor U39148 (N_39148,N_36873,N_37906);
and U39149 (N_39149,N_36925,N_37794);
nand U39150 (N_39150,N_37684,N_37509);
and U39151 (N_39151,N_37430,N_37914);
nand U39152 (N_39152,N_36718,N_37438);
nand U39153 (N_39153,N_37501,N_36149);
or U39154 (N_39154,N_37031,N_36948);
or U39155 (N_39155,N_36881,N_36648);
and U39156 (N_39156,N_36570,N_36930);
and U39157 (N_39157,N_37509,N_37123);
nor U39158 (N_39158,N_36691,N_36422);
nand U39159 (N_39159,N_37247,N_36252);
or U39160 (N_39160,N_36827,N_37896);
nor U39161 (N_39161,N_36449,N_36286);
and U39162 (N_39162,N_36197,N_37842);
nand U39163 (N_39163,N_37910,N_37155);
or U39164 (N_39164,N_37387,N_36038);
nor U39165 (N_39165,N_37226,N_37258);
nand U39166 (N_39166,N_37720,N_36654);
and U39167 (N_39167,N_36742,N_36146);
or U39168 (N_39168,N_37963,N_36360);
xnor U39169 (N_39169,N_36863,N_37624);
or U39170 (N_39170,N_37339,N_36806);
nand U39171 (N_39171,N_36832,N_37695);
and U39172 (N_39172,N_37639,N_37992);
xor U39173 (N_39173,N_36379,N_37563);
or U39174 (N_39174,N_37458,N_37336);
and U39175 (N_39175,N_37548,N_36146);
nand U39176 (N_39176,N_36615,N_37881);
and U39177 (N_39177,N_37970,N_36636);
nor U39178 (N_39178,N_37824,N_37572);
and U39179 (N_39179,N_36506,N_37976);
and U39180 (N_39180,N_37059,N_37907);
nor U39181 (N_39181,N_36790,N_37763);
nand U39182 (N_39182,N_37930,N_36784);
nand U39183 (N_39183,N_36576,N_37341);
nand U39184 (N_39184,N_36878,N_37160);
nor U39185 (N_39185,N_37191,N_37603);
and U39186 (N_39186,N_37623,N_36804);
nor U39187 (N_39187,N_36128,N_37716);
or U39188 (N_39188,N_37050,N_36050);
or U39189 (N_39189,N_37820,N_37256);
nor U39190 (N_39190,N_37098,N_37693);
and U39191 (N_39191,N_36008,N_36997);
nand U39192 (N_39192,N_37663,N_37151);
nand U39193 (N_39193,N_36226,N_37206);
xnor U39194 (N_39194,N_36335,N_36126);
and U39195 (N_39195,N_37741,N_36455);
or U39196 (N_39196,N_37890,N_36829);
nand U39197 (N_39197,N_36028,N_37151);
or U39198 (N_39198,N_37385,N_36577);
nor U39199 (N_39199,N_37190,N_37244);
nor U39200 (N_39200,N_36997,N_36689);
and U39201 (N_39201,N_37808,N_36654);
and U39202 (N_39202,N_36363,N_36953);
or U39203 (N_39203,N_36393,N_37436);
and U39204 (N_39204,N_36037,N_37092);
or U39205 (N_39205,N_37667,N_36596);
nor U39206 (N_39206,N_37417,N_36925);
nor U39207 (N_39207,N_36834,N_37795);
nor U39208 (N_39208,N_36933,N_36474);
and U39209 (N_39209,N_36005,N_37830);
nor U39210 (N_39210,N_36784,N_37081);
and U39211 (N_39211,N_37813,N_36672);
and U39212 (N_39212,N_37144,N_36007);
nor U39213 (N_39213,N_36906,N_37431);
and U39214 (N_39214,N_37009,N_36627);
and U39215 (N_39215,N_36197,N_36958);
or U39216 (N_39216,N_37533,N_37408);
nand U39217 (N_39217,N_36908,N_36134);
nor U39218 (N_39218,N_37987,N_37086);
nand U39219 (N_39219,N_37707,N_37148);
and U39220 (N_39220,N_36883,N_37476);
or U39221 (N_39221,N_37529,N_36697);
and U39222 (N_39222,N_37485,N_36589);
and U39223 (N_39223,N_37672,N_36261);
nand U39224 (N_39224,N_37076,N_36462);
and U39225 (N_39225,N_37877,N_37675);
nand U39226 (N_39226,N_36554,N_36710);
nand U39227 (N_39227,N_37670,N_36779);
or U39228 (N_39228,N_37445,N_37731);
nand U39229 (N_39229,N_36338,N_36253);
nand U39230 (N_39230,N_36305,N_37386);
nand U39231 (N_39231,N_37012,N_36566);
and U39232 (N_39232,N_36733,N_37190);
or U39233 (N_39233,N_37383,N_37169);
or U39234 (N_39234,N_37754,N_36271);
and U39235 (N_39235,N_36798,N_36300);
nand U39236 (N_39236,N_36378,N_36621);
and U39237 (N_39237,N_36502,N_36185);
nor U39238 (N_39238,N_36889,N_37166);
and U39239 (N_39239,N_37387,N_37013);
nand U39240 (N_39240,N_36508,N_36332);
nand U39241 (N_39241,N_36494,N_37782);
or U39242 (N_39242,N_36798,N_37474);
xor U39243 (N_39243,N_36311,N_37485);
and U39244 (N_39244,N_36642,N_36149);
and U39245 (N_39245,N_37443,N_37786);
nand U39246 (N_39246,N_37097,N_36728);
or U39247 (N_39247,N_36184,N_36680);
and U39248 (N_39248,N_37860,N_36837);
and U39249 (N_39249,N_36607,N_36433);
nor U39250 (N_39250,N_36089,N_37357);
and U39251 (N_39251,N_37773,N_37639);
and U39252 (N_39252,N_37167,N_37674);
nor U39253 (N_39253,N_37252,N_36562);
and U39254 (N_39254,N_37036,N_37517);
nor U39255 (N_39255,N_37017,N_37429);
and U39256 (N_39256,N_36329,N_37860);
nor U39257 (N_39257,N_36445,N_36184);
or U39258 (N_39258,N_37928,N_36693);
and U39259 (N_39259,N_37335,N_36540);
or U39260 (N_39260,N_37062,N_36444);
or U39261 (N_39261,N_37047,N_37311);
nand U39262 (N_39262,N_37431,N_36619);
nor U39263 (N_39263,N_36019,N_36171);
nand U39264 (N_39264,N_36425,N_36289);
nand U39265 (N_39265,N_36187,N_37622);
or U39266 (N_39266,N_36586,N_36876);
nand U39267 (N_39267,N_37394,N_37156);
and U39268 (N_39268,N_37468,N_36217);
nand U39269 (N_39269,N_37373,N_36626);
or U39270 (N_39270,N_36181,N_36201);
and U39271 (N_39271,N_36812,N_36324);
or U39272 (N_39272,N_36616,N_36667);
and U39273 (N_39273,N_36469,N_36980);
and U39274 (N_39274,N_36383,N_37167);
and U39275 (N_39275,N_36254,N_37235);
nor U39276 (N_39276,N_37726,N_37739);
and U39277 (N_39277,N_36512,N_36427);
or U39278 (N_39278,N_36588,N_37352);
and U39279 (N_39279,N_36347,N_36114);
nor U39280 (N_39280,N_36641,N_37978);
nor U39281 (N_39281,N_36764,N_37153);
nand U39282 (N_39282,N_37659,N_37369);
nor U39283 (N_39283,N_37993,N_36334);
nor U39284 (N_39284,N_37864,N_37066);
nand U39285 (N_39285,N_37380,N_37034);
nor U39286 (N_39286,N_36706,N_36122);
nand U39287 (N_39287,N_37767,N_36779);
and U39288 (N_39288,N_36375,N_37960);
and U39289 (N_39289,N_37243,N_36025);
and U39290 (N_39290,N_37103,N_37598);
xnor U39291 (N_39291,N_37397,N_37407);
nand U39292 (N_39292,N_36655,N_36247);
nand U39293 (N_39293,N_37140,N_36066);
nor U39294 (N_39294,N_37396,N_37951);
or U39295 (N_39295,N_36697,N_37874);
and U39296 (N_39296,N_37402,N_37898);
or U39297 (N_39297,N_37612,N_37622);
nand U39298 (N_39298,N_37496,N_36233);
nor U39299 (N_39299,N_36472,N_37580);
nand U39300 (N_39300,N_37814,N_37194);
nand U39301 (N_39301,N_37689,N_37514);
and U39302 (N_39302,N_36952,N_37069);
nand U39303 (N_39303,N_37821,N_36552);
and U39304 (N_39304,N_36035,N_36482);
or U39305 (N_39305,N_36617,N_36975);
nand U39306 (N_39306,N_36182,N_37646);
or U39307 (N_39307,N_36696,N_37541);
nand U39308 (N_39308,N_37235,N_37284);
nand U39309 (N_39309,N_36596,N_36388);
or U39310 (N_39310,N_36573,N_36340);
nand U39311 (N_39311,N_37349,N_36295);
and U39312 (N_39312,N_36804,N_37930);
or U39313 (N_39313,N_37266,N_37808);
or U39314 (N_39314,N_36065,N_37422);
and U39315 (N_39315,N_36920,N_36756);
nor U39316 (N_39316,N_37779,N_36816);
nand U39317 (N_39317,N_36510,N_37424);
and U39318 (N_39318,N_36514,N_37662);
nor U39319 (N_39319,N_36507,N_36655);
or U39320 (N_39320,N_37332,N_37902);
or U39321 (N_39321,N_37632,N_37524);
or U39322 (N_39322,N_36916,N_36485);
xnor U39323 (N_39323,N_37623,N_37744);
nand U39324 (N_39324,N_36658,N_37909);
nand U39325 (N_39325,N_36677,N_36199);
nor U39326 (N_39326,N_36402,N_36510);
and U39327 (N_39327,N_37665,N_36243);
or U39328 (N_39328,N_37412,N_37918);
nor U39329 (N_39329,N_37703,N_36149);
nor U39330 (N_39330,N_37857,N_36866);
nand U39331 (N_39331,N_37568,N_37126);
nor U39332 (N_39332,N_36185,N_37186);
or U39333 (N_39333,N_36619,N_37700);
nand U39334 (N_39334,N_36596,N_37956);
or U39335 (N_39335,N_37117,N_37393);
and U39336 (N_39336,N_37019,N_36856);
xor U39337 (N_39337,N_37587,N_37910);
and U39338 (N_39338,N_36523,N_37172);
and U39339 (N_39339,N_37530,N_37842);
nor U39340 (N_39340,N_36553,N_36989);
nand U39341 (N_39341,N_37242,N_36634);
nor U39342 (N_39342,N_37838,N_37351);
or U39343 (N_39343,N_36268,N_37752);
nor U39344 (N_39344,N_36624,N_36931);
and U39345 (N_39345,N_37429,N_37002);
nor U39346 (N_39346,N_36345,N_37233);
and U39347 (N_39347,N_36708,N_37898);
nor U39348 (N_39348,N_37942,N_36657);
and U39349 (N_39349,N_36020,N_36417);
nand U39350 (N_39350,N_36289,N_37533);
nand U39351 (N_39351,N_37088,N_36876);
nand U39352 (N_39352,N_37597,N_36882);
and U39353 (N_39353,N_37197,N_37547);
nand U39354 (N_39354,N_36977,N_36495);
and U39355 (N_39355,N_37767,N_37650);
or U39356 (N_39356,N_36660,N_37967);
and U39357 (N_39357,N_36836,N_36261);
nand U39358 (N_39358,N_37405,N_37374);
and U39359 (N_39359,N_37792,N_37037);
and U39360 (N_39360,N_36679,N_37914);
or U39361 (N_39361,N_37091,N_37142);
nand U39362 (N_39362,N_37269,N_37983);
or U39363 (N_39363,N_37478,N_37042);
or U39364 (N_39364,N_37532,N_36631);
nor U39365 (N_39365,N_36765,N_36689);
nand U39366 (N_39366,N_37042,N_36825);
or U39367 (N_39367,N_37611,N_37595);
nor U39368 (N_39368,N_37138,N_37869);
nand U39369 (N_39369,N_37303,N_36491);
and U39370 (N_39370,N_36663,N_37980);
or U39371 (N_39371,N_37282,N_36808);
nand U39372 (N_39372,N_36076,N_37184);
and U39373 (N_39373,N_37221,N_37378);
nor U39374 (N_39374,N_37096,N_37851);
and U39375 (N_39375,N_36822,N_36232);
nor U39376 (N_39376,N_36170,N_37115);
and U39377 (N_39377,N_37594,N_36508);
or U39378 (N_39378,N_36658,N_36628);
nor U39379 (N_39379,N_36306,N_36529);
and U39380 (N_39380,N_37722,N_36256);
nor U39381 (N_39381,N_36531,N_36821);
nand U39382 (N_39382,N_37710,N_37371);
nand U39383 (N_39383,N_36993,N_37081);
nor U39384 (N_39384,N_36570,N_37784);
nand U39385 (N_39385,N_36533,N_36269);
nand U39386 (N_39386,N_37154,N_37232);
nand U39387 (N_39387,N_36367,N_37687);
xnor U39388 (N_39388,N_37836,N_36278);
and U39389 (N_39389,N_36396,N_37619);
and U39390 (N_39390,N_37878,N_36978);
nor U39391 (N_39391,N_37206,N_37777);
nor U39392 (N_39392,N_37312,N_37752);
nand U39393 (N_39393,N_37542,N_37316);
xnor U39394 (N_39394,N_37806,N_36000);
nand U39395 (N_39395,N_37712,N_37795);
nand U39396 (N_39396,N_37423,N_36453);
nor U39397 (N_39397,N_37362,N_37018);
nand U39398 (N_39398,N_36874,N_36595);
nand U39399 (N_39399,N_37699,N_37609);
and U39400 (N_39400,N_36687,N_36410);
nand U39401 (N_39401,N_37180,N_36043);
and U39402 (N_39402,N_37418,N_37894);
nand U39403 (N_39403,N_37066,N_37299);
and U39404 (N_39404,N_37246,N_36886);
nand U39405 (N_39405,N_37811,N_37434);
or U39406 (N_39406,N_37919,N_36552);
or U39407 (N_39407,N_37390,N_36439);
nand U39408 (N_39408,N_36149,N_37536);
nor U39409 (N_39409,N_37228,N_36714);
or U39410 (N_39410,N_37118,N_36500);
nand U39411 (N_39411,N_36998,N_36443);
nand U39412 (N_39412,N_37535,N_37228);
and U39413 (N_39413,N_37519,N_36451);
or U39414 (N_39414,N_37970,N_37105);
or U39415 (N_39415,N_37794,N_37905);
nor U39416 (N_39416,N_37348,N_36622);
and U39417 (N_39417,N_36263,N_36307);
nor U39418 (N_39418,N_36555,N_36589);
or U39419 (N_39419,N_36346,N_37445);
nor U39420 (N_39420,N_37666,N_36838);
or U39421 (N_39421,N_36992,N_36274);
nand U39422 (N_39422,N_36745,N_36958);
and U39423 (N_39423,N_36483,N_37675);
or U39424 (N_39424,N_37966,N_37646);
and U39425 (N_39425,N_36082,N_36224);
nor U39426 (N_39426,N_36730,N_36009);
and U39427 (N_39427,N_36316,N_36968);
and U39428 (N_39428,N_36635,N_36104);
or U39429 (N_39429,N_36756,N_36871);
nand U39430 (N_39430,N_37314,N_37531);
nor U39431 (N_39431,N_36360,N_36428);
and U39432 (N_39432,N_36623,N_37579);
and U39433 (N_39433,N_36172,N_37290);
and U39434 (N_39434,N_37166,N_37199);
nor U39435 (N_39435,N_37403,N_36303);
or U39436 (N_39436,N_36298,N_37259);
nor U39437 (N_39437,N_36628,N_37748);
or U39438 (N_39438,N_37935,N_36697);
and U39439 (N_39439,N_37740,N_37187);
or U39440 (N_39440,N_37109,N_37579);
nand U39441 (N_39441,N_36341,N_37565);
nor U39442 (N_39442,N_37816,N_37631);
nand U39443 (N_39443,N_37510,N_36655);
nor U39444 (N_39444,N_36580,N_36127);
nor U39445 (N_39445,N_36729,N_36846);
and U39446 (N_39446,N_36165,N_37464);
nor U39447 (N_39447,N_37516,N_36503);
and U39448 (N_39448,N_36213,N_37243);
or U39449 (N_39449,N_37609,N_37863);
or U39450 (N_39450,N_37267,N_37472);
and U39451 (N_39451,N_36187,N_37368);
and U39452 (N_39452,N_36430,N_37760);
nor U39453 (N_39453,N_36208,N_36715);
and U39454 (N_39454,N_36193,N_36803);
or U39455 (N_39455,N_36284,N_37764);
and U39456 (N_39456,N_36814,N_36279);
and U39457 (N_39457,N_36237,N_36658);
or U39458 (N_39458,N_36751,N_37058);
and U39459 (N_39459,N_36496,N_37930);
and U39460 (N_39460,N_36562,N_37621);
or U39461 (N_39461,N_36368,N_37181);
nor U39462 (N_39462,N_37567,N_36516);
and U39463 (N_39463,N_36644,N_36883);
nor U39464 (N_39464,N_37433,N_37144);
nor U39465 (N_39465,N_36985,N_36650);
nor U39466 (N_39466,N_36096,N_37204);
nor U39467 (N_39467,N_36187,N_36099);
nand U39468 (N_39468,N_37160,N_36471);
or U39469 (N_39469,N_37403,N_36689);
xor U39470 (N_39470,N_37329,N_36700);
nor U39471 (N_39471,N_36070,N_36638);
and U39472 (N_39472,N_36281,N_36352);
or U39473 (N_39473,N_37066,N_36112);
and U39474 (N_39474,N_36904,N_36393);
or U39475 (N_39475,N_37826,N_36206);
nand U39476 (N_39476,N_36349,N_36162);
nand U39477 (N_39477,N_37016,N_36965);
and U39478 (N_39478,N_36921,N_37347);
nand U39479 (N_39479,N_36912,N_36352);
nand U39480 (N_39480,N_36315,N_37203);
or U39481 (N_39481,N_36697,N_37880);
or U39482 (N_39482,N_36042,N_37688);
and U39483 (N_39483,N_36266,N_36079);
nand U39484 (N_39484,N_36433,N_36803);
nand U39485 (N_39485,N_37051,N_37413);
nor U39486 (N_39486,N_36667,N_37589);
nor U39487 (N_39487,N_36609,N_36798);
or U39488 (N_39488,N_36067,N_37295);
nand U39489 (N_39489,N_37878,N_37089);
and U39490 (N_39490,N_37144,N_36767);
or U39491 (N_39491,N_37688,N_36678);
and U39492 (N_39492,N_36680,N_37537);
or U39493 (N_39493,N_37231,N_37080);
and U39494 (N_39494,N_36530,N_36545);
and U39495 (N_39495,N_36115,N_37237);
xnor U39496 (N_39496,N_36609,N_36007);
and U39497 (N_39497,N_37534,N_37571);
nor U39498 (N_39498,N_36104,N_37853);
nand U39499 (N_39499,N_37443,N_37216);
and U39500 (N_39500,N_37143,N_36727);
nor U39501 (N_39501,N_36467,N_37059);
or U39502 (N_39502,N_37865,N_37018);
xor U39503 (N_39503,N_36914,N_36035);
and U39504 (N_39504,N_37058,N_36889);
or U39505 (N_39505,N_36221,N_37037);
nand U39506 (N_39506,N_37106,N_37710);
and U39507 (N_39507,N_36787,N_37154);
nor U39508 (N_39508,N_36116,N_37880);
and U39509 (N_39509,N_37204,N_36342);
nor U39510 (N_39510,N_36924,N_37903);
and U39511 (N_39511,N_37929,N_37886);
and U39512 (N_39512,N_36272,N_37956);
nand U39513 (N_39513,N_37115,N_37732);
and U39514 (N_39514,N_37505,N_37692);
and U39515 (N_39515,N_36777,N_36446);
or U39516 (N_39516,N_36693,N_36473);
and U39517 (N_39517,N_37861,N_37408);
nor U39518 (N_39518,N_36375,N_37367);
nor U39519 (N_39519,N_37458,N_36147);
and U39520 (N_39520,N_36450,N_37745);
or U39521 (N_39521,N_37628,N_37982);
nor U39522 (N_39522,N_37016,N_36386);
and U39523 (N_39523,N_36405,N_36653);
nor U39524 (N_39524,N_36386,N_36882);
nand U39525 (N_39525,N_36283,N_37326);
or U39526 (N_39526,N_36226,N_37905);
or U39527 (N_39527,N_37850,N_36824);
nor U39528 (N_39528,N_36571,N_36375);
nand U39529 (N_39529,N_36660,N_36620);
or U39530 (N_39530,N_36880,N_36576);
and U39531 (N_39531,N_36023,N_36327);
nor U39532 (N_39532,N_37258,N_37266);
or U39533 (N_39533,N_36923,N_36088);
nand U39534 (N_39534,N_37934,N_36263);
xor U39535 (N_39535,N_37143,N_37325);
nor U39536 (N_39536,N_36985,N_36415);
or U39537 (N_39537,N_36597,N_37120);
nor U39538 (N_39538,N_36184,N_37920);
nor U39539 (N_39539,N_36118,N_36466);
nor U39540 (N_39540,N_37328,N_37213);
nor U39541 (N_39541,N_37394,N_37235);
or U39542 (N_39542,N_36068,N_37067);
and U39543 (N_39543,N_36178,N_36101);
nor U39544 (N_39544,N_36263,N_37203);
nand U39545 (N_39545,N_36094,N_36114);
nand U39546 (N_39546,N_36537,N_37333);
nand U39547 (N_39547,N_37311,N_37050);
nor U39548 (N_39548,N_36305,N_37216);
nand U39549 (N_39549,N_37279,N_37600);
and U39550 (N_39550,N_36488,N_37721);
or U39551 (N_39551,N_37253,N_37452);
or U39552 (N_39552,N_36084,N_36508);
or U39553 (N_39553,N_37241,N_36672);
nand U39554 (N_39554,N_36793,N_36634);
nand U39555 (N_39555,N_37497,N_36995);
or U39556 (N_39556,N_36969,N_36753);
xnor U39557 (N_39557,N_37584,N_36713);
and U39558 (N_39558,N_36147,N_36865);
or U39559 (N_39559,N_37528,N_36224);
nor U39560 (N_39560,N_36849,N_36954);
nor U39561 (N_39561,N_37400,N_37589);
and U39562 (N_39562,N_36632,N_37533);
nor U39563 (N_39563,N_37408,N_37856);
or U39564 (N_39564,N_37518,N_36800);
nand U39565 (N_39565,N_37562,N_37017);
nor U39566 (N_39566,N_36075,N_37137);
or U39567 (N_39567,N_36820,N_37356);
nand U39568 (N_39568,N_37497,N_36234);
or U39569 (N_39569,N_37579,N_37587);
nand U39570 (N_39570,N_36768,N_37029);
nand U39571 (N_39571,N_36420,N_37752);
nor U39572 (N_39572,N_37206,N_36612);
and U39573 (N_39573,N_36457,N_36454);
nor U39574 (N_39574,N_36477,N_36433);
or U39575 (N_39575,N_37075,N_36384);
nor U39576 (N_39576,N_37765,N_36633);
and U39577 (N_39577,N_36430,N_36580);
or U39578 (N_39578,N_37939,N_36429);
or U39579 (N_39579,N_37236,N_37074);
nor U39580 (N_39580,N_36029,N_37775);
nand U39581 (N_39581,N_36895,N_37578);
nor U39582 (N_39582,N_37826,N_36534);
nor U39583 (N_39583,N_36225,N_36404);
and U39584 (N_39584,N_37260,N_36036);
nor U39585 (N_39585,N_37071,N_36591);
nor U39586 (N_39586,N_37756,N_37904);
or U39587 (N_39587,N_36999,N_36457);
nand U39588 (N_39588,N_36923,N_37925);
or U39589 (N_39589,N_37053,N_37319);
or U39590 (N_39590,N_36766,N_36019);
nand U39591 (N_39591,N_36973,N_36463);
and U39592 (N_39592,N_36592,N_36521);
or U39593 (N_39593,N_37456,N_37153);
and U39594 (N_39594,N_36876,N_37485);
or U39595 (N_39595,N_37476,N_36113);
or U39596 (N_39596,N_37366,N_36942);
or U39597 (N_39597,N_36995,N_36218);
and U39598 (N_39598,N_37171,N_37076);
nor U39599 (N_39599,N_36191,N_36447);
nand U39600 (N_39600,N_37766,N_37044);
nor U39601 (N_39601,N_36103,N_37403);
or U39602 (N_39602,N_36280,N_36928);
and U39603 (N_39603,N_36712,N_36180);
nand U39604 (N_39604,N_36291,N_37518);
nor U39605 (N_39605,N_36610,N_36690);
xor U39606 (N_39606,N_37608,N_36271);
or U39607 (N_39607,N_36248,N_36784);
and U39608 (N_39608,N_36828,N_36625);
and U39609 (N_39609,N_37987,N_36059);
or U39610 (N_39610,N_37548,N_36262);
and U39611 (N_39611,N_36259,N_36987);
nand U39612 (N_39612,N_36688,N_37377);
nand U39613 (N_39613,N_37743,N_36898);
and U39614 (N_39614,N_36221,N_37604);
or U39615 (N_39615,N_37690,N_37909);
and U39616 (N_39616,N_36354,N_37983);
or U39617 (N_39617,N_37199,N_37116);
and U39618 (N_39618,N_36823,N_36029);
nand U39619 (N_39619,N_36252,N_37128);
and U39620 (N_39620,N_37342,N_37126);
nand U39621 (N_39621,N_36038,N_36733);
or U39622 (N_39622,N_37713,N_36695);
nand U39623 (N_39623,N_37202,N_37592);
nor U39624 (N_39624,N_36917,N_36952);
xor U39625 (N_39625,N_36533,N_37680);
and U39626 (N_39626,N_36345,N_36819);
nor U39627 (N_39627,N_36288,N_37030);
nand U39628 (N_39628,N_36430,N_36120);
and U39629 (N_39629,N_37419,N_36078);
nand U39630 (N_39630,N_37163,N_37599);
xnor U39631 (N_39631,N_36454,N_36556);
or U39632 (N_39632,N_36013,N_37288);
or U39633 (N_39633,N_36834,N_37662);
or U39634 (N_39634,N_37558,N_37212);
or U39635 (N_39635,N_37638,N_37086);
and U39636 (N_39636,N_37440,N_36541);
nor U39637 (N_39637,N_37614,N_36406);
or U39638 (N_39638,N_37933,N_36878);
or U39639 (N_39639,N_37557,N_36032);
and U39640 (N_39640,N_36591,N_37241);
nand U39641 (N_39641,N_37960,N_36319);
nand U39642 (N_39642,N_37453,N_37162);
and U39643 (N_39643,N_37426,N_36762);
or U39644 (N_39644,N_36004,N_36249);
or U39645 (N_39645,N_37748,N_36319);
and U39646 (N_39646,N_36141,N_36622);
nand U39647 (N_39647,N_37607,N_37829);
xor U39648 (N_39648,N_37689,N_37982);
nor U39649 (N_39649,N_37919,N_36913);
or U39650 (N_39650,N_36524,N_37676);
nor U39651 (N_39651,N_37493,N_37829);
or U39652 (N_39652,N_37422,N_36596);
nor U39653 (N_39653,N_36246,N_37279);
and U39654 (N_39654,N_36006,N_37276);
nand U39655 (N_39655,N_37299,N_36987);
nand U39656 (N_39656,N_36298,N_36805);
nor U39657 (N_39657,N_36871,N_36873);
nand U39658 (N_39658,N_36213,N_36432);
or U39659 (N_39659,N_37705,N_37456);
and U39660 (N_39660,N_37942,N_37414);
or U39661 (N_39661,N_37592,N_36899);
or U39662 (N_39662,N_36370,N_36771);
and U39663 (N_39663,N_36038,N_36153);
nor U39664 (N_39664,N_37531,N_37097);
and U39665 (N_39665,N_37765,N_37241);
or U39666 (N_39666,N_37577,N_37314);
and U39667 (N_39667,N_36304,N_36831);
nand U39668 (N_39668,N_37494,N_36589);
nor U39669 (N_39669,N_37204,N_37929);
nor U39670 (N_39670,N_36661,N_36671);
nor U39671 (N_39671,N_36187,N_37129);
or U39672 (N_39672,N_37606,N_36091);
nor U39673 (N_39673,N_37439,N_36247);
nand U39674 (N_39674,N_37499,N_36159);
and U39675 (N_39675,N_37702,N_37073);
or U39676 (N_39676,N_36973,N_37218);
and U39677 (N_39677,N_37159,N_37557);
and U39678 (N_39678,N_36886,N_36121);
or U39679 (N_39679,N_37596,N_36078);
or U39680 (N_39680,N_36743,N_36869);
nand U39681 (N_39681,N_36816,N_37290);
or U39682 (N_39682,N_37923,N_36807);
or U39683 (N_39683,N_36680,N_36797);
nand U39684 (N_39684,N_37341,N_37717);
nor U39685 (N_39685,N_37179,N_37185);
nor U39686 (N_39686,N_37515,N_36440);
and U39687 (N_39687,N_36228,N_37322);
nand U39688 (N_39688,N_36156,N_36222);
nor U39689 (N_39689,N_37049,N_36838);
nor U39690 (N_39690,N_37701,N_36572);
and U39691 (N_39691,N_37001,N_37763);
or U39692 (N_39692,N_36369,N_36789);
nand U39693 (N_39693,N_36385,N_36457);
and U39694 (N_39694,N_37665,N_36456);
nor U39695 (N_39695,N_36660,N_36427);
and U39696 (N_39696,N_37632,N_37514);
or U39697 (N_39697,N_37713,N_37587);
and U39698 (N_39698,N_36293,N_36001);
or U39699 (N_39699,N_36350,N_36791);
or U39700 (N_39700,N_36601,N_37294);
nor U39701 (N_39701,N_37593,N_37646);
and U39702 (N_39702,N_37076,N_37229);
and U39703 (N_39703,N_36578,N_37574);
or U39704 (N_39704,N_37702,N_36498);
nor U39705 (N_39705,N_36049,N_36292);
or U39706 (N_39706,N_36913,N_37371);
or U39707 (N_39707,N_37311,N_37646);
or U39708 (N_39708,N_37399,N_36738);
and U39709 (N_39709,N_36151,N_37741);
or U39710 (N_39710,N_36158,N_37786);
or U39711 (N_39711,N_37880,N_37548);
nor U39712 (N_39712,N_36059,N_37907);
and U39713 (N_39713,N_37081,N_36276);
and U39714 (N_39714,N_36180,N_37024);
nor U39715 (N_39715,N_36554,N_37832);
xor U39716 (N_39716,N_37454,N_37889);
or U39717 (N_39717,N_36059,N_37644);
and U39718 (N_39718,N_37849,N_37013);
nor U39719 (N_39719,N_36862,N_37848);
nor U39720 (N_39720,N_37605,N_36983);
nor U39721 (N_39721,N_37238,N_37521);
nor U39722 (N_39722,N_36800,N_37175);
nor U39723 (N_39723,N_37697,N_37360);
or U39724 (N_39724,N_37153,N_36055);
or U39725 (N_39725,N_36585,N_36167);
nand U39726 (N_39726,N_36874,N_36917);
nor U39727 (N_39727,N_36168,N_36911);
nor U39728 (N_39728,N_36748,N_36172);
nand U39729 (N_39729,N_37875,N_37162);
nand U39730 (N_39730,N_37250,N_37032);
nand U39731 (N_39731,N_37958,N_37481);
and U39732 (N_39732,N_37844,N_36998);
nand U39733 (N_39733,N_36168,N_37671);
or U39734 (N_39734,N_37430,N_36596);
and U39735 (N_39735,N_37803,N_36428);
and U39736 (N_39736,N_36388,N_36646);
or U39737 (N_39737,N_36512,N_37792);
or U39738 (N_39738,N_36810,N_37089);
or U39739 (N_39739,N_36430,N_37791);
or U39740 (N_39740,N_36710,N_36096);
nor U39741 (N_39741,N_36741,N_36062);
or U39742 (N_39742,N_37429,N_37853);
nand U39743 (N_39743,N_36140,N_36026);
and U39744 (N_39744,N_37373,N_37883);
and U39745 (N_39745,N_37312,N_36999);
nor U39746 (N_39746,N_36236,N_37750);
nand U39747 (N_39747,N_37120,N_37277);
or U39748 (N_39748,N_36938,N_37957);
and U39749 (N_39749,N_37832,N_36486);
nand U39750 (N_39750,N_36931,N_37473);
and U39751 (N_39751,N_36861,N_36680);
nand U39752 (N_39752,N_36992,N_36239);
nor U39753 (N_39753,N_36335,N_36393);
and U39754 (N_39754,N_37055,N_37962);
nand U39755 (N_39755,N_36983,N_37637);
and U39756 (N_39756,N_37300,N_36956);
nor U39757 (N_39757,N_37312,N_36932);
and U39758 (N_39758,N_37736,N_37244);
nand U39759 (N_39759,N_36082,N_36088);
nand U39760 (N_39760,N_37392,N_37129);
nand U39761 (N_39761,N_36807,N_37295);
nand U39762 (N_39762,N_36205,N_37673);
nand U39763 (N_39763,N_36650,N_37025);
or U39764 (N_39764,N_37889,N_37625);
or U39765 (N_39765,N_36805,N_36331);
nor U39766 (N_39766,N_37229,N_37889);
and U39767 (N_39767,N_37654,N_37822);
nor U39768 (N_39768,N_36504,N_36396);
nand U39769 (N_39769,N_37799,N_37984);
or U39770 (N_39770,N_36602,N_36255);
or U39771 (N_39771,N_36346,N_36874);
and U39772 (N_39772,N_37319,N_36787);
nand U39773 (N_39773,N_37521,N_37260);
and U39774 (N_39774,N_36764,N_36332);
and U39775 (N_39775,N_36293,N_36198);
and U39776 (N_39776,N_36606,N_37019);
nand U39777 (N_39777,N_37712,N_37176);
nor U39778 (N_39778,N_37856,N_37672);
nand U39779 (N_39779,N_36775,N_36684);
nand U39780 (N_39780,N_37507,N_37902);
or U39781 (N_39781,N_36217,N_37414);
nand U39782 (N_39782,N_36106,N_36013);
nand U39783 (N_39783,N_36419,N_36347);
xnor U39784 (N_39784,N_37945,N_37079);
nor U39785 (N_39785,N_37165,N_37470);
and U39786 (N_39786,N_36611,N_36118);
xnor U39787 (N_39787,N_36225,N_36094);
nor U39788 (N_39788,N_37808,N_36228);
nand U39789 (N_39789,N_37060,N_37626);
nor U39790 (N_39790,N_36611,N_37783);
nor U39791 (N_39791,N_36762,N_36459);
or U39792 (N_39792,N_37979,N_37503);
nand U39793 (N_39793,N_37702,N_36456);
or U39794 (N_39794,N_37862,N_36306);
nor U39795 (N_39795,N_37242,N_36562);
and U39796 (N_39796,N_37756,N_36177);
and U39797 (N_39797,N_36035,N_37165);
and U39798 (N_39798,N_37637,N_36839);
xor U39799 (N_39799,N_36688,N_36562);
and U39800 (N_39800,N_37277,N_36244);
nand U39801 (N_39801,N_37602,N_36917);
and U39802 (N_39802,N_37415,N_36284);
nor U39803 (N_39803,N_37600,N_36539);
nor U39804 (N_39804,N_37547,N_36326);
nand U39805 (N_39805,N_36886,N_37979);
nor U39806 (N_39806,N_36909,N_36736);
and U39807 (N_39807,N_37900,N_36456);
or U39808 (N_39808,N_36876,N_37728);
nor U39809 (N_39809,N_36151,N_37221);
or U39810 (N_39810,N_36464,N_37605);
nor U39811 (N_39811,N_37882,N_36784);
nand U39812 (N_39812,N_37982,N_36583);
and U39813 (N_39813,N_37278,N_36391);
nand U39814 (N_39814,N_37379,N_37894);
nor U39815 (N_39815,N_37195,N_37627);
and U39816 (N_39816,N_36154,N_37562);
and U39817 (N_39817,N_36773,N_36091);
and U39818 (N_39818,N_37942,N_36953);
and U39819 (N_39819,N_36555,N_36833);
or U39820 (N_39820,N_37206,N_36238);
and U39821 (N_39821,N_36657,N_36481);
nand U39822 (N_39822,N_37876,N_37642);
nor U39823 (N_39823,N_36391,N_36137);
nor U39824 (N_39824,N_36274,N_36727);
or U39825 (N_39825,N_37968,N_37135);
nand U39826 (N_39826,N_36627,N_37354);
or U39827 (N_39827,N_36184,N_37424);
or U39828 (N_39828,N_37082,N_36643);
nand U39829 (N_39829,N_36784,N_37677);
or U39830 (N_39830,N_36947,N_37627);
and U39831 (N_39831,N_36365,N_36701);
nand U39832 (N_39832,N_37385,N_37927);
nand U39833 (N_39833,N_37776,N_36272);
nand U39834 (N_39834,N_37512,N_37872);
nor U39835 (N_39835,N_36032,N_36663);
nand U39836 (N_39836,N_37312,N_36488);
or U39837 (N_39837,N_36230,N_37975);
or U39838 (N_39838,N_37302,N_37763);
or U39839 (N_39839,N_37038,N_36945);
nor U39840 (N_39840,N_36166,N_36099);
nand U39841 (N_39841,N_36887,N_36464);
nor U39842 (N_39842,N_36958,N_36586);
nand U39843 (N_39843,N_36483,N_37968);
or U39844 (N_39844,N_36363,N_37567);
nand U39845 (N_39845,N_37052,N_36482);
nand U39846 (N_39846,N_37159,N_37600);
nor U39847 (N_39847,N_37394,N_37180);
nor U39848 (N_39848,N_36807,N_37060);
and U39849 (N_39849,N_37624,N_36061);
or U39850 (N_39850,N_37640,N_37908);
and U39851 (N_39851,N_36622,N_37447);
xor U39852 (N_39852,N_36400,N_37355);
nand U39853 (N_39853,N_37851,N_37350);
or U39854 (N_39854,N_37039,N_37918);
nor U39855 (N_39855,N_36162,N_37796);
nor U39856 (N_39856,N_36839,N_37551);
or U39857 (N_39857,N_36185,N_36595);
nand U39858 (N_39858,N_37499,N_36032);
or U39859 (N_39859,N_37072,N_37389);
nor U39860 (N_39860,N_36939,N_36740);
nand U39861 (N_39861,N_37312,N_36870);
nand U39862 (N_39862,N_37459,N_37610);
nand U39863 (N_39863,N_36982,N_37888);
and U39864 (N_39864,N_37681,N_36625);
nand U39865 (N_39865,N_36072,N_37363);
and U39866 (N_39866,N_37939,N_36141);
nor U39867 (N_39867,N_36521,N_37884);
or U39868 (N_39868,N_36919,N_36954);
nand U39869 (N_39869,N_37148,N_37636);
or U39870 (N_39870,N_37200,N_36716);
and U39871 (N_39871,N_37191,N_37881);
nor U39872 (N_39872,N_37102,N_37204);
and U39873 (N_39873,N_37137,N_36396);
nand U39874 (N_39874,N_37910,N_37613);
nand U39875 (N_39875,N_37903,N_37686);
xor U39876 (N_39876,N_37797,N_36294);
and U39877 (N_39877,N_37589,N_37391);
nor U39878 (N_39878,N_37900,N_37980);
nand U39879 (N_39879,N_36997,N_36558);
and U39880 (N_39880,N_37488,N_37844);
nand U39881 (N_39881,N_37093,N_36944);
nor U39882 (N_39882,N_37895,N_37997);
or U39883 (N_39883,N_36543,N_36533);
nand U39884 (N_39884,N_36920,N_36129);
nor U39885 (N_39885,N_37625,N_36703);
and U39886 (N_39886,N_37308,N_36188);
nand U39887 (N_39887,N_36264,N_37375);
nor U39888 (N_39888,N_36748,N_36396);
and U39889 (N_39889,N_37007,N_37026);
and U39890 (N_39890,N_36735,N_37816);
and U39891 (N_39891,N_36999,N_37489);
or U39892 (N_39892,N_36463,N_37227);
or U39893 (N_39893,N_36342,N_37059);
and U39894 (N_39894,N_36847,N_37822);
and U39895 (N_39895,N_36885,N_36288);
nand U39896 (N_39896,N_36990,N_37147);
nor U39897 (N_39897,N_37644,N_37107);
nor U39898 (N_39898,N_36957,N_36494);
nand U39899 (N_39899,N_36645,N_37329);
and U39900 (N_39900,N_36349,N_36531);
nor U39901 (N_39901,N_36238,N_36211);
or U39902 (N_39902,N_36043,N_36585);
or U39903 (N_39903,N_37124,N_37901);
xor U39904 (N_39904,N_36749,N_36983);
nand U39905 (N_39905,N_37512,N_36436);
nor U39906 (N_39906,N_37071,N_37957);
nand U39907 (N_39907,N_37264,N_36056);
nand U39908 (N_39908,N_36392,N_36741);
or U39909 (N_39909,N_37835,N_37327);
or U39910 (N_39910,N_36254,N_37806);
and U39911 (N_39911,N_37485,N_37183);
nand U39912 (N_39912,N_36500,N_37594);
and U39913 (N_39913,N_36249,N_37759);
and U39914 (N_39914,N_36302,N_36025);
nand U39915 (N_39915,N_37798,N_36913);
nand U39916 (N_39916,N_36216,N_36032);
nor U39917 (N_39917,N_37087,N_36523);
and U39918 (N_39918,N_37772,N_37620);
and U39919 (N_39919,N_37370,N_37532);
and U39920 (N_39920,N_36547,N_36681);
nor U39921 (N_39921,N_37883,N_36639);
nor U39922 (N_39922,N_36271,N_36275);
nor U39923 (N_39923,N_37371,N_36783);
nand U39924 (N_39924,N_36203,N_37394);
and U39925 (N_39925,N_37114,N_36160);
and U39926 (N_39926,N_37157,N_36085);
or U39927 (N_39927,N_37762,N_36929);
nand U39928 (N_39928,N_37858,N_37834);
nand U39929 (N_39929,N_37311,N_36388);
and U39930 (N_39930,N_37266,N_36522);
and U39931 (N_39931,N_37932,N_36855);
and U39932 (N_39932,N_37457,N_36593);
xor U39933 (N_39933,N_36731,N_37876);
and U39934 (N_39934,N_37268,N_36471);
or U39935 (N_39935,N_36767,N_37630);
or U39936 (N_39936,N_36849,N_37946);
or U39937 (N_39937,N_36468,N_36496);
and U39938 (N_39938,N_37941,N_37114);
nand U39939 (N_39939,N_37090,N_36398);
nand U39940 (N_39940,N_36594,N_36425);
and U39941 (N_39941,N_37827,N_37778);
nand U39942 (N_39942,N_36172,N_37547);
nand U39943 (N_39943,N_36048,N_36470);
nand U39944 (N_39944,N_36537,N_36291);
nor U39945 (N_39945,N_36896,N_37816);
or U39946 (N_39946,N_36184,N_37778);
or U39947 (N_39947,N_37127,N_36058);
nor U39948 (N_39948,N_37649,N_37908);
and U39949 (N_39949,N_36359,N_37074);
nand U39950 (N_39950,N_37337,N_37008);
nand U39951 (N_39951,N_37659,N_36678);
nor U39952 (N_39952,N_36672,N_36358);
nor U39953 (N_39953,N_36150,N_37597);
nor U39954 (N_39954,N_37322,N_37663);
nor U39955 (N_39955,N_37763,N_37570);
nand U39956 (N_39956,N_37809,N_36595);
and U39957 (N_39957,N_36246,N_36046);
and U39958 (N_39958,N_37408,N_36493);
or U39959 (N_39959,N_37196,N_36001);
nand U39960 (N_39960,N_36582,N_37734);
nor U39961 (N_39961,N_37755,N_37153);
nor U39962 (N_39962,N_36855,N_37351);
xor U39963 (N_39963,N_36761,N_37645);
nand U39964 (N_39964,N_36101,N_37194);
and U39965 (N_39965,N_37043,N_36633);
and U39966 (N_39966,N_36065,N_37870);
xnor U39967 (N_39967,N_37440,N_36665);
and U39968 (N_39968,N_36106,N_36392);
nor U39969 (N_39969,N_37043,N_37223);
or U39970 (N_39970,N_37002,N_36871);
nand U39971 (N_39971,N_37438,N_36658);
and U39972 (N_39972,N_37049,N_37454);
nand U39973 (N_39973,N_36278,N_36016);
nand U39974 (N_39974,N_36310,N_36661);
and U39975 (N_39975,N_37433,N_37944);
and U39976 (N_39976,N_36465,N_36390);
nand U39977 (N_39977,N_36604,N_37788);
nor U39978 (N_39978,N_37034,N_36205);
or U39979 (N_39979,N_37011,N_36425);
nor U39980 (N_39980,N_37827,N_37384);
nand U39981 (N_39981,N_37566,N_37676);
and U39982 (N_39982,N_37933,N_37953);
nand U39983 (N_39983,N_37107,N_36346);
nand U39984 (N_39984,N_37887,N_36971);
nor U39985 (N_39985,N_37244,N_36807);
and U39986 (N_39986,N_36511,N_36913);
or U39987 (N_39987,N_36769,N_37611);
or U39988 (N_39988,N_37671,N_36593);
nand U39989 (N_39989,N_36034,N_37567);
nand U39990 (N_39990,N_37101,N_37658);
nand U39991 (N_39991,N_37149,N_36705);
nand U39992 (N_39992,N_37553,N_36650);
or U39993 (N_39993,N_36272,N_37543);
or U39994 (N_39994,N_37729,N_37442);
and U39995 (N_39995,N_37447,N_36608);
nor U39996 (N_39996,N_36095,N_37273);
nor U39997 (N_39997,N_37575,N_37310);
xor U39998 (N_39998,N_37248,N_37016);
nor U39999 (N_39999,N_37808,N_37286);
and U40000 (N_40000,N_38969,N_38824);
nand U40001 (N_40001,N_38121,N_38482);
and U40002 (N_40002,N_39200,N_38361);
and U40003 (N_40003,N_39593,N_38263);
xnor U40004 (N_40004,N_38949,N_39681);
or U40005 (N_40005,N_38841,N_38382);
or U40006 (N_40006,N_38289,N_38698);
and U40007 (N_40007,N_38722,N_38139);
nand U40008 (N_40008,N_38916,N_39847);
xor U40009 (N_40009,N_38055,N_39603);
nand U40010 (N_40010,N_38486,N_39547);
nand U40011 (N_40011,N_38491,N_38025);
nor U40012 (N_40012,N_39737,N_38012);
and U40013 (N_40013,N_38011,N_39504);
nor U40014 (N_40014,N_39123,N_38913);
nand U40015 (N_40015,N_39598,N_38353);
nor U40016 (N_40016,N_39389,N_39570);
nor U40017 (N_40017,N_38048,N_39410);
or U40018 (N_40018,N_39060,N_38475);
and U40019 (N_40019,N_38907,N_38216);
and U40020 (N_40020,N_39280,N_39127);
nor U40021 (N_40021,N_39174,N_38926);
nor U40022 (N_40022,N_39205,N_39134);
nand U40023 (N_40023,N_39740,N_38256);
and U40024 (N_40024,N_38032,N_38168);
or U40025 (N_40025,N_39006,N_38746);
nor U40026 (N_40026,N_39054,N_39886);
and U40027 (N_40027,N_39961,N_39351);
and U40028 (N_40028,N_38999,N_38845);
nand U40029 (N_40029,N_38508,N_38606);
or U40030 (N_40030,N_38861,N_39822);
and U40031 (N_40031,N_38073,N_38511);
and U40032 (N_40032,N_38792,N_38914);
and U40033 (N_40033,N_39744,N_38943);
and U40034 (N_40034,N_39275,N_38325);
or U40035 (N_40035,N_38148,N_38649);
nor U40036 (N_40036,N_38854,N_39602);
nor U40037 (N_40037,N_38478,N_38112);
xor U40038 (N_40038,N_38909,N_39771);
and U40039 (N_40039,N_38173,N_39187);
and U40040 (N_40040,N_39114,N_38529);
or U40041 (N_40041,N_39942,N_39459);
or U40042 (N_40042,N_39573,N_39214);
or U40043 (N_40043,N_39755,N_38822);
and U40044 (N_40044,N_38596,N_38858);
nand U40045 (N_40045,N_39180,N_39609);
and U40046 (N_40046,N_38806,N_39201);
nand U40047 (N_40047,N_39369,N_39909);
and U40048 (N_40048,N_38740,N_38417);
nand U40049 (N_40049,N_39465,N_38928);
nor U40050 (N_40050,N_39703,N_38947);
or U40051 (N_40051,N_38349,N_39050);
nor U40052 (N_40052,N_39367,N_38401);
nand U40053 (N_40053,N_38128,N_39904);
nor U40054 (N_40054,N_38471,N_38844);
nor U40055 (N_40055,N_39199,N_39937);
nor U40056 (N_40056,N_38652,N_38117);
and U40057 (N_40057,N_38391,N_38126);
xor U40058 (N_40058,N_39754,N_38747);
or U40059 (N_40059,N_39005,N_39568);
nor U40060 (N_40060,N_38262,N_38019);
nor U40061 (N_40061,N_39955,N_39823);
or U40062 (N_40062,N_39505,N_38572);
or U40063 (N_40063,N_39648,N_39320);
or U40064 (N_40064,N_38591,N_38451);
or U40065 (N_40065,N_39748,N_38005);
nor U40066 (N_40066,N_39153,N_39322);
or U40067 (N_40067,N_38118,N_39594);
nand U40068 (N_40068,N_38889,N_39009);
and U40069 (N_40069,N_38489,N_38975);
nand U40070 (N_40070,N_39846,N_39219);
nor U40071 (N_40071,N_38415,N_38389);
nand U40072 (N_40072,N_38338,N_38782);
nand U40073 (N_40073,N_39232,N_39697);
nor U40074 (N_40074,N_39251,N_38155);
nor U40075 (N_40075,N_38929,N_38265);
and U40076 (N_40076,N_38908,N_38487);
nand U40077 (N_40077,N_38376,N_39494);
nand U40078 (N_40078,N_38773,N_38789);
or U40079 (N_40079,N_39430,N_39715);
nand U40080 (N_40080,N_39419,N_39233);
or U40081 (N_40081,N_38984,N_39622);
nor U40082 (N_40082,N_39665,N_39943);
or U40083 (N_40083,N_39802,N_39049);
and U40084 (N_40084,N_38692,N_39302);
nor U40085 (N_40085,N_38464,N_39796);
xor U40086 (N_40086,N_38468,N_39628);
nand U40087 (N_40087,N_39575,N_39963);
nand U40088 (N_40088,N_38093,N_39061);
nand U40089 (N_40089,N_39976,N_38754);
nand U40090 (N_40090,N_38250,N_38729);
or U40091 (N_40091,N_39217,N_38702);
nor U40092 (N_40092,N_38170,N_38114);
and U40093 (N_40093,N_38257,N_39297);
nand U40094 (N_40094,N_38452,N_38835);
or U40095 (N_40095,N_39495,N_39024);
or U40096 (N_40096,N_38871,N_39076);
and U40097 (N_40097,N_39989,N_38197);
nor U40098 (N_40098,N_39376,N_38420);
nand U40099 (N_40099,N_39818,N_39307);
or U40100 (N_40100,N_38020,N_39089);
nand U40101 (N_40101,N_38049,N_38588);
nand U40102 (N_40102,N_38558,N_39877);
nor U40103 (N_40103,N_39295,N_38672);
or U40104 (N_40104,N_39861,N_39361);
or U40105 (N_40105,N_38052,N_38661);
and U40106 (N_40106,N_38879,N_38608);
nor U40107 (N_40107,N_38067,N_39707);
nand U40108 (N_40108,N_38815,N_38795);
nor U40109 (N_40109,N_38527,N_39285);
or U40110 (N_40110,N_38569,N_38665);
nand U40111 (N_40111,N_38676,N_38666);
nand U40112 (N_40112,N_38431,N_39212);
or U40113 (N_40113,N_38528,N_38053);
nor U40114 (N_40114,N_38850,N_38274);
nor U40115 (N_40115,N_38832,N_39651);
nand U40116 (N_40116,N_39002,N_39436);
nor U40117 (N_40117,N_39552,N_39468);
nor U40118 (N_40118,N_39265,N_38291);
or U40119 (N_40119,N_38490,N_39309);
or U40120 (N_40120,N_39451,N_38057);
or U40121 (N_40121,N_39031,N_38954);
nand U40122 (N_40122,N_38033,N_39709);
or U40123 (N_40123,N_39305,N_39919);
nand U40124 (N_40124,N_38247,N_39438);
or U40125 (N_40125,N_38959,N_38674);
or U40126 (N_40126,N_39348,N_38517);
xor U40127 (N_40127,N_39638,N_39752);
nor U40128 (N_40128,N_39023,N_39028);
or U40129 (N_40129,N_38883,N_38074);
or U40130 (N_40130,N_39927,N_38650);
or U40131 (N_40131,N_39433,N_39968);
nor U40132 (N_40132,N_39655,N_38812);
nand U40133 (N_40133,N_38612,N_38022);
and U40134 (N_40134,N_38671,N_38158);
nor U40135 (N_40135,N_38171,N_39340);
nand U40136 (N_40136,N_38253,N_38640);
and U40137 (N_40137,N_38326,N_38316);
nor U40138 (N_40138,N_39081,N_39642);
and U40139 (N_40139,N_38739,N_38357);
nor U40140 (N_40140,N_38736,N_39167);
nor U40141 (N_40141,N_39188,N_38419);
nand U40142 (N_40142,N_38026,N_38085);
nand U40143 (N_40143,N_39728,N_38394);
nor U40144 (N_40144,N_39907,N_39313);
nand U40145 (N_40145,N_39824,N_39267);
and U40146 (N_40146,N_38570,N_39700);
nand U40147 (N_40147,N_39645,N_38664);
and U40148 (N_40148,N_39284,N_38154);
nand U40149 (N_40149,N_38064,N_39776);
nand U40150 (N_40150,N_38258,N_39033);
or U40151 (N_40151,N_39413,N_38921);
and U40152 (N_40152,N_39162,N_39420);
nor U40153 (N_40153,N_39170,N_38567);
nor U40154 (N_40154,N_39514,N_39101);
or U40155 (N_40155,N_39166,N_38878);
nor U40156 (N_40156,N_39473,N_38534);
nand U40157 (N_40157,N_39241,N_39213);
and U40158 (N_40158,N_39222,N_39027);
nor U40159 (N_40159,N_38393,N_38427);
and U40160 (N_40160,N_39334,N_38646);
nand U40161 (N_40161,N_39580,N_39917);
nor U40162 (N_40162,N_39992,N_38068);
and U40163 (N_40163,N_39960,N_38494);
nand U40164 (N_40164,N_38436,N_39062);
or U40165 (N_40165,N_39795,N_39261);
nor U40166 (N_40166,N_39844,N_38399);
nand U40167 (N_40167,N_39287,N_38227);
nand U40168 (N_40168,N_39887,N_39503);
nand U40169 (N_40169,N_39319,N_38450);
nand U40170 (N_40170,N_39312,N_39202);
nor U40171 (N_40171,N_38737,N_38181);
and U40172 (N_40172,N_38461,N_38360);
or U40173 (N_40173,N_38138,N_39442);
nor U40174 (N_40174,N_39996,N_38079);
or U40175 (N_40175,N_38960,N_38767);
or U40176 (N_40176,N_39781,N_38220);
or U40177 (N_40177,N_38149,N_38412);
nor U40178 (N_40178,N_38404,N_39765);
nor U40179 (N_40179,N_38002,N_39513);
and U40180 (N_40180,N_38849,N_39331);
nand U40181 (N_40181,N_39146,N_38243);
or U40182 (N_40182,N_38586,N_39726);
nor U40183 (N_40183,N_38018,N_38367);
and U40184 (N_40184,N_38091,N_38329);
nand U40185 (N_40185,N_38900,N_38565);
and U40186 (N_40186,N_39646,N_39160);
and U40187 (N_40187,N_38398,N_38087);
or U40188 (N_40188,N_39093,N_38245);
nor U40189 (N_40189,N_39018,N_39059);
or U40190 (N_40190,N_39132,N_38381);
or U40191 (N_40191,N_39627,N_38651);
or U40192 (N_40192,N_38364,N_39116);
or U40193 (N_40193,N_39432,N_39685);
nor U40194 (N_40194,N_39292,N_39673);
nand U40195 (N_40195,N_39536,N_39444);
or U40196 (N_40196,N_39591,N_38560);
or U40197 (N_40197,N_38614,N_39911);
nor U40198 (N_40198,N_39945,N_39038);
nor U40199 (N_40199,N_39656,N_39522);
or U40200 (N_40200,N_38551,N_39281);
nand U40201 (N_40201,N_39032,N_39527);
nand U40202 (N_40202,N_39113,N_39183);
nand U40203 (N_40203,N_39982,N_38140);
nor U40204 (N_40204,N_39938,N_38995);
nor U40205 (N_40205,N_39778,N_39242);
and U40206 (N_40206,N_38352,N_39194);
nand U40207 (N_40207,N_39617,N_39094);
and U40208 (N_40208,N_39901,N_39492);
or U40209 (N_40209,N_38753,N_39896);
or U40210 (N_40210,N_38449,N_38413);
nand U40211 (N_40211,N_39549,N_39868);
or U40212 (N_40212,N_38609,N_38297);
nor U40213 (N_40213,N_39429,N_38579);
nand U40214 (N_40214,N_38115,N_38716);
and U40215 (N_40215,N_38153,N_38617);
and U40216 (N_40216,N_39667,N_38638);
or U40217 (N_40217,N_38749,N_38484);
and U40218 (N_40218,N_38083,N_39130);
nand U40219 (N_40219,N_39831,N_38628);
nor U40220 (N_40220,N_38056,N_39110);
and U40221 (N_40221,N_38331,N_38231);
or U40222 (N_40222,N_38081,N_38276);
nor U40223 (N_40223,N_39924,N_39077);
nor U40224 (N_40224,N_39891,N_38496);
nand U40225 (N_40225,N_39865,N_38834);
nand U40226 (N_40226,N_39608,N_39355);
and U40227 (N_40227,N_39954,N_39375);
or U40228 (N_40228,N_38899,N_38385);
nand U40229 (N_40229,N_38189,N_38448);
or U40230 (N_40230,N_38620,N_39838);
or U40231 (N_40231,N_39317,N_38632);
nor U40232 (N_40232,N_39586,N_38629);
nand U40233 (N_40233,N_38945,N_39025);
nand U40234 (N_40234,N_38028,N_39720);
and U40235 (N_40235,N_38513,N_39888);
nor U40236 (N_40236,N_38800,N_38814);
and U40237 (N_40237,N_39131,N_39449);
and U40238 (N_40238,N_38619,N_38965);
nand U40239 (N_40239,N_39425,N_39812);
nand U40240 (N_40240,N_39143,N_38555);
or U40241 (N_40241,N_39724,N_39158);
nand U40242 (N_40242,N_39860,N_39182);
nor U40243 (N_40243,N_39582,N_39121);
nand U40244 (N_40244,N_39540,N_39095);
or U40245 (N_40245,N_38964,N_38136);
nor U40246 (N_40246,N_38974,N_38784);
nor U40247 (N_40247,N_39652,N_39446);
or U40248 (N_40248,N_38212,N_39806);
nor U40249 (N_40249,N_38470,N_38318);
and U40250 (N_40250,N_38686,N_38510);
nand U40251 (N_40251,N_39706,N_38356);
and U40252 (N_40252,N_39329,N_38141);
nor U40253 (N_40253,N_38681,N_39934);
and U40254 (N_40254,N_38595,N_39756);
nor U40255 (N_40255,N_38147,N_38347);
and U40256 (N_40256,N_38346,N_39064);
and U40257 (N_40257,N_38285,N_38700);
nor U40258 (N_40258,N_39784,N_38472);
nand U40259 (N_40259,N_39829,N_38823);
nand U40260 (N_40260,N_39820,N_39149);
nor U40261 (N_40261,N_38282,N_39854);
nand U40262 (N_40262,N_39493,N_39995);
nand U40263 (N_40263,N_39004,N_38842);
or U40264 (N_40264,N_39262,N_39288);
xnor U40265 (N_40265,N_38497,N_39350);
or U40266 (N_40266,N_39843,N_38460);
or U40267 (N_40267,N_38456,N_38980);
and U40268 (N_40268,N_39852,N_38167);
and U40269 (N_40269,N_39816,N_39920);
or U40270 (N_40270,N_38807,N_39620);
nor U40271 (N_40271,N_39014,N_38601);
or U40272 (N_40272,N_38295,N_38890);
and U40273 (N_40273,N_38695,N_38599);
nor U40274 (N_40274,N_39516,N_38124);
nor U40275 (N_40275,N_38175,N_38868);
or U40276 (N_40276,N_38034,N_39734);
nand U40277 (N_40277,N_38457,N_38594);
and U40278 (N_40278,N_38611,N_38576);
nor U40279 (N_40279,N_38582,N_39303);
nor U40280 (N_40280,N_39308,N_38424);
and U40281 (N_40281,N_38341,N_38384);
or U40282 (N_40282,N_39408,N_39533);
nand U40283 (N_40283,N_39129,N_39358);
and U40284 (N_40284,N_39629,N_39104);
or U40285 (N_40285,N_38687,N_38694);
nor U40286 (N_40286,N_38712,N_38137);
or U40287 (N_40287,N_39330,N_38309);
or U40288 (N_40288,N_38647,N_38793);
nand U40289 (N_40289,N_38645,N_39346);
and U40290 (N_40290,N_38375,N_38195);
or U40291 (N_40291,N_39086,N_39423);
nor U40292 (N_40292,N_39612,N_38226);
nand U40293 (N_40293,N_39624,N_39326);
nand U40294 (N_40294,N_39531,N_38962);
or U40295 (N_40295,N_39647,N_39769);
and U40296 (N_40296,N_39067,N_38312);
or U40297 (N_40297,N_38771,N_38013);
or U40298 (N_40298,N_38493,N_39417);
and U40299 (N_40299,N_38799,N_38886);
nand U40300 (N_40300,N_38780,N_39405);
and U40301 (N_40301,N_38354,N_39633);
and U40302 (N_40302,N_39529,N_38634);
nand U40303 (N_40303,N_39984,N_39133);
and U40304 (N_40304,N_38116,N_38271);
or U40305 (N_40305,N_38077,N_39507);
or U40306 (N_40306,N_39487,N_39368);
and U40307 (N_40307,N_39008,N_38429);
nand U40308 (N_40308,N_39892,N_38607);
nor U40309 (N_40309,N_38229,N_39699);
or U40310 (N_40310,N_38092,N_39867);
nor U40311 (N_40311,N_38242,N_38506);
xnor U40312 (N_40312,N_38821,N_38481);
or U40313 (N_40313,N_38304,N_38339);
or U40314 (N_40314,N_38235,N_39075);
and U40315 (N_40315,N_38993,N_38000);
xnor U40316 (N_40316,N_39532,N_38462);
nor U40317 (N_40317,N_38030,N_39597);
and U40318 (N_40318,N_39112,N_38830);
and U40319 (N_40319,N_38183,N_38761);
or U40320 (N_40320,N_38725,N_38217);
nor U40321 (N_40321,N_38987,N_39866);
nor U40322 (N_40322,N_38006,N_39282);
or U40323 (N_40323,N_38330,N_39056);
nor U40324 (N_40324,N_39352,N_39443);
and U40325 (N_40325,N_39454,N_39988);
and U40326 (N_40326,N_38473,N_38322);
and U40327 (N_40327,N_39286,N_38583);
xor U40328 (N_40328,N_39338,N_39566);
or U40329 (N_40329,N_38630,N_38531);
and U40330 (N_40330,N_39767,N_39936);
or U40331 (N_40331,N_39238,N_38730);
and U40332 (N_40332,N_38985,N_39256);
nor U40333 (N_40333,N_39569,N_39415);
nor U40334 (N_40334,N_38798,N_38514);
and U40335 (N_40335,N_38548,N_39467);
or U40336 (N_40336,N_38266,N_39336);
or U40337 (N_40337,N_38060,N_38015);
nor U40338 (N_40338,N_39387,N_39498);
and U40339 (N_40339,N_39677,N_38445);
nand U40340 (N_40340,N_39366,N_38580);
or U40341 (N_40341,N_39929,N_38224);
nor U40342 (N_40342,N_38161,N_38163);
or U40343 (N_40343,N_39154,N_38058);
and U40344 (N_40344,N_38305,N_39916);
xor U40345 (N_40345,N_38303,N_39951);
and U40346 (N_40346,N_39759,N_38996);
and U40347 (N_40347,N_38742,N_39364);
nor U40348 (N_40348,N_38281,N_39424);
nor U40349 (N_40349,N_38904,N_39175);
nand U40350 (N_40350,N_38221,N_38122);
nor U40351 (N_40351,N_39395,N_38935);
nor U40352 (N_40352,N_38192,N_39821);
and U40353 (N_40353,N_39559,N_38775);
nand U40354 (N_40354,N_38751,N_39718);
nand U40355 (N_40355,N_39216,N_38293);
or U40356 (N_40356,N_38703,N_38788);
or U40357 (N_40357,N_39614,N_39777);
nand U40358 (N_40358,N_38443,N_39453);
nor U40359 (N_40359,N_38240,N_38371);
nor U40360 (N_40360,N_38976,N_38094);
nand U40361 (N_40361,N_39741,N_38867);
and U40362 (N_40362,N_38707,N_38539);
nor U40363 (N_40363,N_39485,N_38622);
or U40364 (N_40364,N_38961,N_38816);
and U40365 (N_40365,N_38956,N_38008);
and U40366 (N_40366,N_39875,N_38499);
nor U40367 (N_40367,N_39779,N_38639);
and U40368 (N_40368,N_38853,N_39774);
nand U40369 (N_40369,N_38683,N_38922);
or U40370 (N_40370,N_39046,N_39998);
nand U40371 (N_40371,N_38210,N_38724);
and U40372 (N_40372,N_38833,N_39897);
and U40373 (N_40373,N_38106,N_38562);
nor U40374 (N_40374,N_39546,N_39007);
nor U40375 (N_40375,N_39825,N_39991);
nand U40376 (N_40376,N_38104,N_39710);
xor U40377 (N_40377,N_39020,N_38102);
and U40378 (N_40378,N_38791,N_39595);
and U40379 (N_40379,N_38159,N_39688);
nor U40380 (N_40380,N_38306,N_39657);
nand U40381 (N_40381,N_39925,N_39750);
nand U40382 (N_40382,N_39611,N_38244);
or U40383 (N_40383,N_39626,N_38923);
and U40384 (N_40384,N_39965,N_39065);
nor U40385 (N_40385,N_38837,N_39817);
or U40386 (N_40386,N_39043,N_38589);
nor U40387 (N_40387,N_39768,N_39128);
or U40388 (N_40388,N_39363,N_38642);
and U40389 (N_40389,N_39422,N_38095);
and U40390 (N_40390,N_39203,N_39833);
or U40391 (N_40391,N_38874,N_38089);
and U40392 (N_40392,N_39138,N_38100);
nand U40393 (N_40393,N_38260,N_39660);
and U40394 (N_40394,N_39906,N_39870);
or U40395 (N_40395,N_38119,N_39797);
nand U40396 (N_40396,N_39905,N_39252);
nand U40397 (N_40397,N_39902,N_38556);
or U40398 (N_40398,N_39551,N_39773);
nand U40399 (N_40399,N_38504,N_39809);
or U40400 (N_40400,N_38906,N_39360);
nand U40401 (N_40401,N_39583,N_39702);
nand U40402 (N_40402,N_39509,N_39794);
nand U40403 (N_40403,N_38469,N_38069);
nor U40404 (N_40404,N_39402,N_38332);
and U40405 (N_40405,N_39713,N_39915);
and U40406 (N_40406,N_38054,N_39592);
nor U40407 (N_40407,N_38172,N_39291);
and U40408 (N_40408,N_38787,N_38180);
nand U40409 (N_40409,N_39962,N_39607);
or U40410 (N_40410,N_38454,N_38587);
nor U40411 (N_40411,N_38455,N_38414);
and U40412 (N_40412,N_38463,N_38178);
nor U40413 (N_40413,N_39235,N_39761);
nor U40414 (N_40414,N_39599,N_39445);
nand U40415 (N_40415,N_38040,N_38007);
nor U40416 (N_40416,N_39084,N_38270);
and U40417 (N_40417,N_38395,N_39135);
and U40418 (N_40418,N_39173,N_39140);
xor U40419 (N_40419,N_39930,N_38203);
and U40420 (N_40420,N_39482,N_38523);
nand U40421 (N_40421,N_38765,N_39071);
and U40422 (N_40422,N_39933,N_39881);
nor U40423 (N_40423,N_38208,N_38533);
or U40424 (N_40424,N_38726,N_38828);
nor U40425 (N_40425,N_39457,N_38768);
and U40426 (N_40426,N_38045,N_39474);
and U40427 (N_40427,N_38659,N_38946);
xnor U40428 (N_40428,N_38035,N_38750);
nand U40429 (N_40429,N_39021,N_38453);
nand U40430 (N_40430,N_38826,N_38623);
or U40431 (N_40431,N_39452,N_38425);
and U40432 (N_40432,N_38160,N_39489);
nand U40433 (N_40433,N_38038,N_38062);
or U40434 (N_40434,N_38774,N_39659);
nor U40435 (N_40435,N_38134,N_38363);
and U40436 (N_40436,N_39841,N_38763);
or U40437 (N_40437,N_39356,N_39786);
nor U40438 (N_40438,N_39808,N_39680);
nand U40439 (N_40439,N_39725,N_38706);
or U40440 (N_40440,N_39729,N_39108);
and U40441 (N_40441,N_39386,N_39082);
and U40442 (N_40442,N_39192,N_38930);
and U40443 (N_40443,N_39016,N_38809);
nor U40444 (N_40444,N_39119,N_39392);
or U40445 (N_40445,N_39126,N_38135);
nand U40446 (N_40446,N_39010,N_38108);
nand U40447 (N_40447,N_38758,N_38031);
nor U40448 (N_40448,N_39039,N_38574);
nand U40449 (N_40449,N_39380,N_38994);
or U40450 (N_40450,N_38741,N_38836);
or U40451 (N_40451,N_38934,N_39115);
nand U40452 (N_40452,N_38537,N_38519);
and U40453 (N_40453,N_39189,N_38526);
and U40454 (N_40454,N_39675,N_39944);
nand U40455 (N_40455,N_39751,N_38225);
and U40456 (N_40456,N_39542,N_39159);
nor U40457 (N_40457,N_38552,N_39990);
nor U40458 (N_40458,N_39840,N_39971);
or U40459 (N_40459,N_38447,N_39246);
or U40460 (N_40460,N_39105,N_39974);
and U40461 (N_40461,N_38880,N_39550);
or U40462 (N_40462,N_39362,N_39826);
or U40463 (N_40463,N_39506,N_38564);
or U40464 (N_40464,N_38898,N_39686);
or U40465 (N_40465,N_38997,N_39800);
xnor U40466 (N_40466,N_38027,N_38711);
xnor U40467 (N_40467,N_39895,N_39198);
or U40468 (N_40468,N_39749,N_39264);
nor U40469 (N_40469,N_39828,N_39001);
nand U40470 (N_40470,N_38669,N_39880);
nand U40471 (N_40471,N_38400,N_38315);
and U40472 (N_40472,N_39382,N_39562);
and U40473 (N_40473,N_39785,N_38046);
nor U40474 (N_40474,N_38423,N_39663);
or U40475 (N_40475,N_38972,N_39102);
and U40476 (N_40476,N_39874,N_38190);
nand U40477 (N_40477,N_39339,N_39541);
nor U40478 (N_40478,N_39544,N_39577);
and U40479 (N_40479,N_38545,N_38014);
nand U40480 (N_40480,N_38697,N_39088);
or U40481 (N_40481,N_38314,N_39560);
or U40482 (N_40482,N_39947,N_39179);
nand U40483 (N_40483,N_39558,N_38182);
nand U40484 (N_40484,N_38076,N_38635);
nor U40485 (N_40485,N_39618,N_39240);
or U40486 (N_40486,N_39239,N_38931);
or U40487 (N_40487,N_39083,N_39578);
nand U40488 (N_40488,N_39178,N_39206);
or U40489 (N_40489,N_38887,N_39882);
nand U40490 (N_40490,N_39528,N_38718);
nor U40491 (N_40491,N_39388,N_38543);
nand U40492 (N_40492,N_38123,N_39191);
nand U40493 (N_40493,N_39122,N_39714);
nand U40494 (N_40494,N_38233,N_39952);
xnor U40495 (N_40495,N_39230,N_39775);
and U40496 (N_40496,N_39848,N_39690);
or U40497 (N_40497,N_39359,N_38870);
nand U40498 (N_40498,N_38897,N_39928);
nand U40499 (N_40499,N_38319,N_38001);
and U40500 (N_40500,N_38405,N_39842);
nor U40501 (N_40501,N_39914,N_38201);
and U40502 (N_40502,N_39407,N_39664);
nor U40503 (N_40503,N_39394,N_39353);
and U40504 (N_40504,N_39365,N_39670);
nand U40505 (N_40505,N_38327,N_39790);
nand U40506 (N_40506,N_38259,N_39401);
nand U40507 (N_40507,N_39946,N_39456);
nand U40508 (N_40508,N_38086,N_39538);
and U40509 (N_40509,N_38408,N_38133);
or U40510 (N_40510,N_38783,N_39899);
or U40511 (N_40511,N_38299,N_39152);
nand U40512 (N_40512,N_39565,N_39502);
nor U40513 (N_40513,N_39856,N_38905);
or U40514 (N_40514,N_38036,N_39118);
nor U40515 (N_40515,N_38892,N_39385);
nand U40516 (N_40516,N_39488,N_39753);
nand U40517 (N_40517,N_39588,N_39763);
nand U40518 (N_40518,N_38684,N_39883);
nor U40519 (N_40519,N_39501,N_39783);
or U40520 (N_40520,N_39209,N_38685);
nor U40521 (N_40521,N_38578,N_39687);
xnor U40522 (N_40522,N_39328,N_39448);
nor U40523 (N_40523,N_39545,N_38021);
and U40524 (N_40524,N_38351,N_39377);
nand U40525 (N_40525,N_38177,N_38760);
nand U40526 (N_40526,N_39236,N_38105);
nand U40527 (N_40527,N_39440,N_38553);
nand U40528 (N_40528,N_38550,N_39383);
and U40529 (N_40529,N_38287,N_38495);
nor U40530 (N_40530,N_39409,N_39472);
or U40531 (N_40531,N_39548,N_39782);
or U40532 (N_40532,N_39641,N_39871);
or U40533 (N_40533,N_39211,N_39539);
and U40534 (N_40534,N_38938,N_38549);
and U40535 (N_40535,N_38597,N_39147);
nand U40536 (N_40536,N_38915,N_38912);
and U40537 (N_40537,N_39636,N_39237);
nor U40538 (N_40538,N_39691,N_39643);
or U40539 (N_40539,N_39078,N_38621);
or U40540 (N_40540,N_39747,N_38082);
or U40541 (N_40541,N_39063,N_38010);
and U40542 (N_40542,N_39512,N_39975);
xor U40543 (N_40543,N_39898,N_38196);
or U40544 (N_40544,N_39730,N_39414);
or U40545 (N_40545,N_38680,N_39908);
nand U40546 (N_40546,N_39803,N_39469);
and U40547 (N_40547,N_38708,N_38663);
nor U40548 (N_40548,N_38717,N_38734);
nand U40549 (N_40549,N_39980,N_38411);
and U40550 (N_40550,N_38705,N_38416);
and U40551 (N_40551,N_39913,N_38857);
or U40552 (N_40552,N_39567,N_38967);
nand U40553 (N_40553,N_39839,N_38267);
nor U40554 (N_40554,N_39258,N_38166);
nor U40555 (N_40555,N_39333,N_39835);
or U40556 (N_40556,N_38380,N_38328);
nor U40557 (N_40557,N_38097,N_39900);
and U40558 (N_40558,N_39787,N_38542);
or U40559 (N_40559,N_38080,N_38186);
and U40560 (N_40560,N_39111,N_39682);
nor U40561 (N_40561,N_38350,N_38075);
or U40562 (N_40562,N_39052,N_39496);
and U40563 (N_40563,N_38043,N_39259);
and U40564 (N_40564,N_38598,N_39606);
or U40565 (N_40565,N_39226,N_38653);
nand U40566 (N_40566,N_39431,N_39210);
and U40567 (N_40567,N_39231,N_39486);
and U40568 (N_40568,N_38983,N_39969);
or U40569 (N_40569,N_39117,N_38313);
nand U40570 (N_40570,N_39653,N_38268);
nand U40571 (N_40571,N_38693,N_39249);
nor U40572 (N_40572,N_38864,N_38234);
nor U40573 (N_40573,N_38230,N_39635);
or U40574 (N_40574,N_38273,N_39462);
and U40575 (N_40575,N_38343,N_39483);
nand U40576 (N_40576,N_39799,N_38869);
nand U40577 (N_40577,N_38362,N_38344);
and U40578 (N_40578,N_38368,N_39374);
nand U40579 (N_40579,N_38566,N_38648);
nor U40580 (N_40580,N_39296,N_39649);
and U40581 (N_40581,N_38403,N_39862);
and U40582 (N_40582,N_39450,N_39863);
and U40583 (N_40583,N_39106,N_38678);
and U40584 (N_40584,N_39683,N_38113);
and U40585 (N_40585,N_39074,N_39396);
nor U40586 (N_40586,N_38625,N_38875);
or U40587 (N_40587,N_39096,N_38039);
nand U40588 (N_40588,N_38492,N_39255);
nor U40589 (N_40589,N_38373,N_38745);
nand U40590 (N_40590,N_39745,N_39712);
nor U40591 (N_40591,N_38099,N_38146);
or U40592 (N_40592,N_38320,N_38715);
and U40593 (N_40593,N_38779,N_39525);
nand U40594 (N_40594,N_38441,N_38223);
or U40595 (N_40595,N_38334,N_38948);
nor U40596 (N_40596,N_39590,N_39640);
nand U40597 (N_40597,N_38605,N_39970);
nor U40598 (N_40598,N_38103,N_39274);
and U40599 (N_40599,N_38571,N_39398);
and U40600 (N_40600,N_38321,N_39716);
or U40601 (N_40601,N_39403,N_38446);
nor U40602 (N_40602,N_39632,N_38396);
nand U40603 (N_40603,N_38902,N_38882);
nor U40604 (N_40604,N_38125,N_38500);
nor U40605 (N_40605,N_38667,N_38422);
nand U40606 (N_40606,N_39674,N_38776);
nand U40607 (N_40607,N_38557,N_39515);
or U40608 (N_40608,N_38286,N_39379);
and U40609 (N_40609,N_39391,N_39137);
nor U40610 (N_40610,N_39220,N_39658);
nor U40611 (N_40611,N_39957,N_39141);
and U40612 (N_40612,N_38406,N_38061);
nand U40613 (N_40613,N_38090,N_38988);
and U40614 (N_40614,N_39694,N_39080);
nor U40615 (N_40615,N_39306,N_38919);
nor U40616 (N_40616,N_39819,N_38627);
or U40617 (N_40617,N_38577,N_38236);
and U40618 (N_40618,N_39918,N_38377);
and U40619 (N_40619,N_39807,N_39257);
nor U40620 (N_40620,N_39072,N_39994);
or U40621 (N_40621,N_39412,N_39526);
nor U40622 (N_40622,N_39543,N_39851);
and U40623 (N_40623,N_39956,N_38637);
and U40624 (N_40624,N_39186,N_39148);
and U40625 (N_40625,N_39579,N_39036);
nand U40626 (N_40626,N_38246,N_38143);
or U40627 (N_40627,N_38215,N_39644);
nand U40628 (N_40628,N_38335,N_38059);
xnor U40629 (N_40629,N_39341,N_39354);
or U40630 (N_40630,N_39051,N_39125);
or U40631 (N_40631,N_39248,N_38785);
nand U40632 (N_40632,N_38254,N_38337);
or U40633 (N_40633,N_39810,N_38222);
and U40634 (N_40634,N_38942,N_38184);
nand U40635 (N_40635,N_38714,N_39695);
and U40636 (N_40636,N_38498,N_38770);
nand U40637 (N_40637,N_39983,N_39793);
and U40638 (N_40638,N_38616,N_39972);
and U40639 (N_40639,N_39103,N_39434);
or U40640 (N_40640,N_38856,N_39857);
nor U40641 (N_40641,N_38848,N_38434);
and U40642 (N_40642,N_38721,N_39204);
nor U40643 (N_40643,N_39458,N_39177);
and U40644 (N_40644,N_39742,N_38164);
or U40645 (N_40645,N_38937,N_39335);
nand U40646 (N_40646,N_39223,N_39510);
or U40647 (N_40647,N_38825,N_38624);
nand U40648 (N_40648,N_38016,N_38209);
nand U40649 (N_40649,N_38421,N_38509);
nand U40650 (N_40650,N_39518,N_39195);
nor U40651 (N_40651,N_38072,N_39894);
nor U40652 (N_40652,N_39878,N_38838);
or U40653 (N_40653,N_38439,N_39073);
or U40654 (N_40654,N_38759,N_38801);
and U40655 (N_40655,N_38355,N_38888);
or U40656 (N_40656,N_39184,N_38851);
or U40657 (N_40657,N_39163,N_38813);
nor U40658 (N_40658,N_38986,N_38275);
and U40659 (N_40659,N_38568,N_38877);
nor U40660 (N_40660,N_38269,N_38071);
nor U40661 (N_40661,N_38797,N_38392);
nand U40662 (N_40662,N_38107,N_38162);
nand U40663 (N_40663,N_39476,N_39349);
or U40664 (N_40664,N_38710,N_39689);
nand U40665 (N_40665,N_38430,N_38743);
nand U40666 (N_40666,N_38530,N_39227);
nor U40667 (N_40667,N_39610,N_39441);
nor U40668 (N_40668,N_38872,N_38536);
xor U40669 (N_40669,N_38374,N_39679);
and U40670 (N_40670,N_38786,N_38713);
nand U40671 (N_40671,N_38541,N_39661);
and U40672 (N_40672,N_39225,N_39370);
nor U40673 (N_40673,N_39939,N_38280);
nand U40674 (N_40674,N_39311,N_39301);
or U40675 (N_40675,N_39853,N_39428);
or U40676 (N_40676,N_39738,N_39022);
or U40677 (N_40677,N_39427,N_39940);
and U40678 (N_40678,N_39357,N_38593);
nand U40679 (N_40679,N_39966,N_39439);
nand U40680 (N_40680,N_39400,N_39711);
xnor U40681 (N_40681,N_39884,N_39953);
nor U40682 (N_40682,N_39780,N_38302);
and U40683 (N_40683,N_38188,N_39979);
nor U40684 (N_40684,N_39299,N_39029);
nand U40685 (N_40685,N_38843,N_38507);
nor U40686 (N_40686,N_39669,N_39986);
and U40687 (N_40687,N_38677,N_39554);
nor U40688 (N_40688,N_38044,N_38829);
nor U40689 (N_40689,N_38958,N_39693);
and U40690 (N_40690,N_39950,N_39373);
or U40691 (N_40691,N_39384,N_38009);
nand U40692 (N_40692,N_39318,N_39662);
and U40693 (N_40693,N_38479,N_38410);
and U40694 (N_40694,N_38088,N_38581);
or U40695 (N_40695,N_38881,N_39012);
nand U40696 (N_40696,N_39830,N_38604);
nor U40697 (N_40697,N_39157,N_38723);
or U40698 (N_40698,N_38592,N_38643);
or U40699 (N_40699,N_39654,N_38925);
nor U40700 (N_40700,N_39727,N_38185);
and U40701 (N_40701,N_38600,N_38433);
and U40702 (N_40702,N_38884,N_39371);
or U40703 (N_40703,N_39298,N_39722);
nor U40704 (N_40704,N_39732,N_39491);
nor U40705 (N_40705,N_39704,N_39764);
and U40706 (N_40706,N_39404,N_38699);
and U40707 (N_40707,N_39421,N_38109);
or U40708 (N_40708,N_38369,N_38174);
and U40709 (N_40709,N_38757,N_38602);
nand U40710 (N_40710,N_38041,N_39789);
or U40711 (N_40711,N_39193,N_39684);
nand U40712 (N_40712,N_39247,N_38781);
nand U40713 (N_40713,N_38893,N_39321);
nand U40714 (N_40714,N_38924,N_39109);
nand U40715 (N_40715,N_38156,N_38911);
nor U40716 (N_40716,N_38037,N_39092);
nand U40717 (N_40717,N_38819,N_38501);
or U40718 (N_40718,N_39987,N_38839);
or U40719 (N_40719,N_39270,N_39721);
or U40720 (N_40720,N_38670,N_38691);
and U40721 (N_40721,N_38193,N_38252);
or U40722 (N_40722,N_38859,N_38989);
nand U40723 (N_40723,N_38386,N_39276);
xnor U40724 (N_40724,N_39068,N_38251);
nand U40725 (N_40725,N_39042,N_39479);
nand U40726 (N_40726,N_38294,N_38748);
nand U40727 (N_40727,N_38024,N_38891);
nand U40728 (N_40728,N_38966,N_39523);
nand U40729 (N_40729,N_38977,N_38078);
and U40730 (N_40730,N_39026,N_39827);
or U40731 (N_40731,N_38435,N_38918);
or U40732 (N_40732,N_39136,N_38426);
or U40733 (N_40733,N_39964,N_39574);
and U40734 (N_40734,N_39263,N_39941);
or U40735 (N_40735,N_39099,N_38324);
or U40736 (N_40736,N_39030,N_39418);
and U40737 (N_40737,N_39723,N_38769);
nor U40738 (N_40738,N_39912,N_38978);
and U40739 (N_40739,N_39698,N_39142);
nor U40740 (N_40740,N_39150,N_38644);
nand U40741 (N_40741,N_39534,N_39798);
nand U40742 (N_40742,N_38547,N_39310);
or U40743 (N_40743,N_39692,N_38145);
or U40744 (N_40744,N_39098,N_39079);
and U40745 (N_40745,N_38204,N_38827);
nor U40746 (N_40746,N_39973,N_38483);
or U40747 (N_40747,N_38518,N_38805);
nor U40748 (N_40748,N_38176,N_38179);
or U40749 (N_40749,N_38719,N_39480);
or U40750 (N_40750,N_39215,N_38290);
and U40751 (N_40751,N_39766,N_39254);
nand U40752 (N_40752,N_39273,N_39228);
or U40753 (N_40753,N_39760,N_38277);
nand U40754 (N_40754,N_38029,N_39165);
and U40755 (N_40755,N_38804,N_38333);
nor U40756 (N_40756,N_39762,N_39958);
or U40757 (N_40757,N_39572,N_38733);
nand U40758 (N_40758,N_38348,N_39197);
nand U40759 (N_40759,N_38520,N_39268);
and U40760 (N_40760,N_39057,N_38852);
nor U40761 (N_40761,N_38296,N_38979);
nand U40762 (N_40762,N_38660,N_39323);
nand U40763 (N_40763,N_39168,N_38017);
or U40764 (N_40764,N_39041,N_38794);
or U40765 (N_40765,N_39563,N_38228);
and U40766 (N_40766,N_39037,N_39045);
or U40767 (N_40767,N_38144,N_39234);
nor U40768 (N_40768,N_38480,N_39805);
nand U40769 (N_40769,N_38584,N_39124);
nor U40770 (N_40770,N_38573,N_38437);
or U40771 (N_40771,N_39455,N_39345);
nand U40772 (N_40772,N_38308,N_39561);
and U40773 (N_40773,N_38428,N_39985);
nor U40774 (N_40774,N_39207,N_38727);
and U40775 (N_40775,N_39616,N_39977);
or U40776 (N_40776,N_39623,N_39813);
and U40777 (N_40777,N_38546,N_39708);
nor U40778 (N_40778,N_38885,N_38110);
and U40779 (N_40779,N_39347,N_38679);
nand U40780 (N_40780,N_39733,N_38292);
nor U40781 (N_40781,N_39100,N_38610);
nand U40782 (N_40782,N_38973,N_39978);
and U40783 (N_40783,N_38311,N_39601);
and U40784 (N_40784,N_38633,N_38811);
and U40785 (N_40785,N_39343,N_38248);
or U40786 (N_40786,N_39926,N_38772);
or U40787 (N_40787,N_39229,N_38950);
and U40788 (N_40788,N_38590,N_38120);
nand U40789 (N_40789,N_39497,N_38790);
or U40790 (N_40790,N_38895,N_39085);
nor U40791 (N_40791,N_39600,N_39058);
nor U40792 (N_40792,N_38264,N_38365);
or U40793 (N_40793,N_39269,N_39717);
or U40794 (N_40794,N_38432,N_38944);
and U40795 (N_40795,N_38084,N_39873);
and U40796 (N_40796,N_38070,N_38142);
nand U40797 (N_40797,N_38239,N_38358);
nor U40798 (N_40798,N_39294,N_39260);
nand U40799 (N_40799,N_39290,N_38709);
nand U40800 (N_40800,N_39922,N_38505);
nor U40801 (N_40801,N_39378,N_39315);
or U40802 (N_40802,N_38957,N_39277);
nor U40803 (N_40803,N_38990,N_39224);
nor U40804 (N_40804,N_38283,N_38205);
nand U40805 (N_40805,N_39272,N_38340);
or U40806 (N_40806,N_39564,N_39120);
and U40807 (N_40807,N_38129,N_38165);
nand U40808 (N_40808,N_38388,N_38300);
or U40809 (N_40809,N_39500,N_39139);
nand U40810 (N_40810,N_38538,N_38766);
and U40811 (N_40811,N_39701,N_38673);
nand U40812 (N_40812,N_39872,N_38525);
nand U40813 (N_40813,N_39993,N_39537);
nand U40814 (N_40814,N_39519,N_38846);
nand U40815 (N_40815,N_38876,N_39475);
or U40816 (N_40816,N_38284,N_39399);
nor U40817 (N_40817,N_39948,N_39304);
or U40818 (N_40818,N_39447,N_38796);
and U40819 (N_40819,N_39325,N_39571);
xor U40820 (N_40820,N_38255,N_39293);
or U40821 (N_40821,N_38418,N_39406);
nor U40822 (N_40822,N_39013,N_38963);
nand U40823 (N_40823,N_38238,N_39499);
nor U40824 (N_40824,N_38618,N_38535);
and U40825 (N_40825,N_38310,N_39164);
and U40826 (N_40826,N_38301,N_38379);
nor U40827 (N_40827,N_39949,N_38458);
nor U40828 (N_40828,N_39156,N_39801);
or U40829 (N_40829,N_38953,N_38873);
nand U40830 (N_40830,N_39731,N_39011);
and U40831 (N_40831,N_38219,N_38096);
or U40832 (N_40832,N_38998,N_39524);
or U40833 (N_40833,N_38860,N_39196);
nor U40834 (N_40834,N_38955,N_39864);
nor U40835 (N_40835,N_38563,N_39017);
nor U40836 (N_40836,N_38372,N_39171);
or U40837 (N_40837,N_38554,N_39736);
or U40838 (N_40838,N_38532,N_38981);
or U40839 (N_40839,N_38626,N_38755);
nor U40840 (N_40840,N_39155,N_39271);
nand U40841 (N_40841,N_39672,N_39837);
or U40842 (N_40842,N_38261,N_38752);
nor U40843 (N_40843,N_38003,N_38862);
and U40844 (N_40844,N_38279,N_39517);
nor U40845 (N_40845,N_38762,N_39832);
and U40846 (N_40846,N_39596,N_38098);
and U40847 (N_40847,N_39997,N_39278);
xor U40848 (N_40848,N_39735,N_39845);
and U40849 (N_40849,N_38004,N_38488);
and U40850 (N_40850,N_39889,N_38951);
or U40851 (N_40851,N_38968,N_39055);
and U40852 (N_40852,N_39381,N_38323);
or U40853 (N_40853,N_39161,N_39604);
nand U40854 (N_40854,N_39743,N_38982);
and U40855 (N_40855,N_38051,N_39804);
and U40856 (N_40856,N_38764,N_39921);
nand U40857 (N_40857,N_38522,N_39337);
nor U40858 (N_40858,N_39151,N_38130);
and U40859 (N_40859,N_39676,N_39250);
xor U40860 (N_40860,N_38901,N_38336);
nor U40861 (N_40861,N_39416,N_39477);
or U40862 (N_40862,N_39520,N_39245);
nand U40863 (N_40863,N_39097,N_38438);
nor U40864 (N_40864,N_38151,N_39461);
and U40865 (N_40865,N_38810,N_38199);
and U40866 (N_40866,N_39858,N_38689);
nand U40867 (N_40867,N_38409,N_38910);
or U40868 (N_40868,N_39244,N_38150);
nor U40869 (N_40869,N_39555,N_39218);
nor U40870 (N_40870,N_39530,N_39460);
or U40871 (N_40871,N_39834,N_39019);
nor U40872 (N_40872,N_39876,N_38200);
and U40873 (N_40873,N_38249,N_39893);
and U40874 (N_40874,N_39144,N_38521);
and U40875 (N_40875,N_39190,N_39811);
or U40876 (N_40876,N_39739,N_39393);
nand U40877 (N_40877,N_38127,N_39671);
or U40878 (N_40878,N_39324,N_38467);
or U40879 (N_40879,N_38191,N_39266);
nand U40880 (N_40880,N_38540,N_38202);
nand U40881 (N_40881,N_39719,N_38920);
and U40882 (N_40882,N_39463,N_38970);
or U40883 (N_40883,N_39070,N_39869);
or U40884 (N_40884,N_38214,N_39634);
nor U40885 (N_40885,N_39705,N_39490);
nor U40886 (N_40886,N_39931,N_38383);
nor U40887 (N_40887,N_38390,N_39553);
or U40888 (N_40888,N_39625,N_39176);
nor U40889 (N_40889,N_39253,N_39044);
or U40890 (N_40890,N_38831,N_38992);
and U40891 (N_40891,N_39015,N_38307);
or U40892 (N_40892,N_38675,N_39300);
or U40893 (N_40893,N_39048,N_39426);
and U40894 (N_40894,N_38132,N_39435);
and U40895 (N_40895,N_39619,N_38559);
and U40896 (N_40896,N_38206,N_38512);
xor U40897 (N_40897,N_39576,N_38198);
or U40898 (N_40898,N_38657,N_39581);
or U40899 (N_40899,N_39040,N_38288);
or U40900 (N_40900,N_39836,N_38896);
and U40901 (N_40901,N_39621,N_38840);
nand U40902 (N_40902,N_39788,N_38613);
or U40903 (N_40903,N_38941,N_38863);
nand U40904 (N_40904,N_38631,N_39589);
xnor U40905 (N_40905,N_38152,N_38575);
and U40906 (N_40906,N_38818,N_38387);
nor U40907 (N_40907,N_39791,N_39757);
or U40908 (N_40908,N_39639,N_38866);
nand U40909 (N_40909,N_38731,N_38459);
xnor U40910 (N_40910,N_39283,N_38298);
and U40911 (N_40911,N_39859,N_38561);
nand U40912 (N_40912,N_39316,N_38218);
and U40913 (N_40913,N_39584,N_39034);
nand U40914 (N_40914,N_38524,N_38194);
nor U40915 (N_40915,N_38023,N_38047);
nand U40916 (N_40916,N_39631,N_38688);
or U40917 (N_40917,N_38933,N_38917);
or U40918 (N_40918,N_39464,N_39650);
nor U40919 (N_40919,N_38370,N_38655);
nor U40920 (N_40920,N_38728,N_39557);
nand U40921 (N_40921,N_38662,N_38777);
nand U40922 (N_40922,N_39047,N_38756);
or U40923 (N_40923,N_38378,N_38397);
nand U40924 (N_40924,N_39981,N_39814);
and U40925 (N_40925,N_38971,N_39185);
or U40926 (N_40926,N_38808,N_38207);
and U40927 (N_40927,N_38585,N_38169);
nor U40928 (N_40928,N_39000,N_38442);
and U40929 (N_40929,N_38732,N_38803);
or U40930 (N_40930,N_39090,N_39587);
nor U40931 (N_40931,N_39390,N_39556);
or U40932 (N_40932,N_39792,N_39087);
or U40933 (N_40933,N_38066,N_39437);
or U40934 (N_40934,N_39850,N_38237);
nor U40935 (N_40935,N_38502,N_38847);
and U40936 (N_40936,N_38940,N_39066);
or U40937 (N_40937,N_38682,N_38359);
or U40938 (N_40938,N_38735,N_39511);
or U40939 (N_40939,N_39091,N_38317);
nand U40940 (N_40940,N_38211,N_38187);
or U40941 (N_40941,N_39959,N_39508);
and U40942 (N_40942,N_39332,N_38241);
and U40943 (N_40943,N_39342,N_39107);
and U40944 (N_40944,N_39411,N_38927);
or U40945 (N_40945,N_38690,N_39999);
and U40946 (N_40946,N_39314,N_38440);
nand U40947 (N_40947,N_38131,N_38503);
nand U40948 (N_40948,N_39481,N_39003);
nand U40949 (N_40949,N_38516,N_39289);
nand U40950 (N_40950,N_39478,N_39903);
and U40951 (N_40951,N_38704,N_39466);
and U40952 (N_40952,N_39885,N_38063);
and U40953 (N_40953,N_39344,N_39208);
nand U40954 (N_40954,N_39169,N_38477);
nand U40955 (N_40955,N_39470,N_39327);
nor U40956 (N_40956,N_39855,N_39471);
and U40957 (N_40957,N_39279,N_38641);
nor U40958 (N_40958,N_38345,N_38444);
nor U40959 (N_40959,N_38050,N_39666);
or U40960 (N_40960,N_39035,N_38738);
nand U40961 (N_40961,N_38272,N_38042);
and U40962 (N_40962,N_39923,N_39484);
and U40963 (N_40963,N_38952,N_39585);
xnor U40964 (N_40964,N_38865,N_39935);
nand U40965 (N_40965,N_38407,N_39615);
or U40966 (N_40966,N_38939,N_38991);
nand U40967 (N_40967,N_38465,N_38157);
xor U40968 (N_40968,N_38932,N_38278);
or U40969 (N_40969,N_38342,N_38802);
nand U40970 (N_40970,N_39221,N_39668);
nand U40971 (N_40971,N_38744,N_39849);
or U40972 (N_40972,N_38817,N_39772);
nand U40973 (N_40973,N_38696,N_38515);
nand U40974 (N_40974,N_39243,N_38720);
or U40975 (N_40975,N_38101,N_38485);
or U40976 (N_40976,N_38936,N_39053);
and U40977 (N_40977,N_38232,N_38903);
xor U40978 (N_40978,N_39932,N_38668);
nand U40979 (N_40979,N_39967,N_38402);
or U40980 (N_40980,N_39637,N_38855);
nor U40981 (N_40981,N_39758,N_38474);
or U40982 (N_40982,N_38615,N_39397);
and U40983 (N_40983,N_39746,N_39770);
and U40984 (N_40984,N_38778,N_38366);
and U40985 (N_40985,N_39605,N_39069);
nand U40986 (N_40986,N_38894,N_39172);
or U40987 (N_40987,N_38213,N_39372);
and U40988 (N_40988,N_38466,N_38603);
nor U40989 (N_40989,N_38820,N_39181);
nand U40990 (N_40990,N_39145,N_39521);
nor U40991 (N_40991,N_38656,N_39613);
and U40992 (N_40992,N_39696,N_38654);
and U40993 (N_40993,N_38658,N_39879);
nand U40994 (N_40994,N_39815,N_38065);
or U40995 (N_40995,N_38701,N_39630);
or U40996 (N_40996,N_39910,N_39535);
nand U40997 (N_40997,N_38636,N_38476);
and U40998 (N_40998,N_38111,N_39890);
nand U40999 (N_40999,N_39678,N_38544);
nor U41000 (N_41000,N_38327,N_38261);
nor U41001 (N_41001,N_38732,N_39766);
and U41002 (N_41002,N_38341,N_38296);
and U41003 (N_41003,N_38169,N_38497);
or U41004 (N_41004,N_38196,N_39978);
nand U41005 (N_41005,N_39079,N_38112);
or U41006 (N_41006,N_39210,N_38480);
nand U41007 (N_41007,N_38698,N_38597);
nand U41008 (N_41008,N_39324,N_39201);
and U41009 (N_41009,N_38562,N_39350);
nor U41010 (N_41010,N_38173,N_38211);
and U41011 (N_41011,N_39908,N_38349);
nor U41012 (N_41012,N_39160,N_39020);
or U41013 (N_41013,N_38303,N_39411);
and U41014 (N_41014,N_38826,N_38769);
and U41015 (N_41015,N_39924,N_38951);
and U41016 (N_41016,N_38719,N_38579);
nor U41017 (N_41017,N_38150,N_39296);
nand U41018 (N_41018,N_39777,N_39980);
and U41019 (N_41019,N_38310,N_39580);
nor U41020 (N_41020,N_38238,N_38656);
and U41021 (N_41021,N_39970,N_39188);
nand U41022 (N_41022,N_38525,N_39805);
or U41023 (N_41023,N_39391,N_39447);
or U41024 (N_41024,N_39151,N_39417);
and U41025 (N_41025,N_38770,N_39061);
or U41026 (N_41026,N_39494,N_38623);
and U41027 (N_41027,N_39068,N_39637);
or U41028 (N_41028,N_39846,N_39732);
xnor U41029 (N_41029,N_38296,N_38434);
and U41030 (N_41030,N_39519,N_39761);
nor U41031 (N_41031,N_38535,N_38183);
nand U41032 (N_41032,N_39139,N_39728);
and U41033 (N_41033,N_38876,N_39092);
or U41034 (N_41034,N_39854,N_38900);
nor U41035 (N_41035,N_38820,N_39437);
or U41036 (N_41036,N_38611,N_38444);
nor U41037 (N_41037,N_38258,N_39304);
or U41038 (N_41038,N_38101,N_38528);
nand U41039 (N_41039,N_39201,N_38180);
and U41040 (N_41040,N_38050,N_39806);
and U41041 (N_41041,N_39640,N_39752);
and U41042 (N_41042,N_39527,N_38118);
and U41043 (N_41043,N_39868,N_38674);
or U41044 (N_41044,N_38153,N_39669);
nor U41045 (N_41045,N_39065,N_39604);
or U41046 (N_41046,N_38424,N_38776);
nand U41047 (N_41047,N_38006,N_39090);
or U41048 (N_41048,N_38569,N_38791);
or U41049 (N_41049,N_39507,N_38841);
and U41050 (N_41050,N_38747,N_39279);
nor U41051 (N_41051,N_38880,N_39807);
and U41052 (N_41052,N_39533,N_39768);
or U41053 (N_41053,N_39831,N_38126);
nor U41054 (N_41054,N_39475,N_39881);
or U41055 (N_41055,N_39560,N_38765);
xor U41056 (N_41056,N_38562,N_39885);
nor U41057 (N_41057,N_38649,N_38857);
and U41058 (N_41058,N_39790,N_39510);
and U41059 (N_41059,N_39044,N_38468);
and U41060 (N_41060,N_38547,N_38259);
or U41061 (N_41061,N_38973,N_39957);
nand U41062 (N_41062,N_38957,N_38169);
nand U41063 (N_41063,N_39158,N_38578);
or U41064 (N_41064,N_38747,N_39668);
nand U41065 (N_41065,N_38982,N_39498);
and U41066 (N_41066,N_38169,N_38609);
or U41067 (N_41067,N_38961,N_39335);
nand U41068 (N_41068,N_39042,N_38719);
or U41069 (N_41069,N_38958,N_38689);
nand U41070 (N_41070,N_39174,N_38089);
and U41071 (N_41071,N_39985,N_39453);
and U41072 (N_41072,N_39125,N_38967);
nand U41073 (N_41073,N_39584,N_39267);
or U41074 (N_41074,N_38528,N_38009);
or U41075 (N_41075,N_39501,N_39475);
nand U41076 (N_41076,N_38757,N_38905);
and U41077 (N_41077,N_39577,N_38736);
and U41078 (N_41078,N_38848,N_39009);
nor U41079 (N_41079,N_38523,N_39742);
and U41080 (N_41080,N_39221,N_39501);
and U41081 (N_41081,N_38236,N_38050);
nor U41082 (N_41082,N_39687,N_38967);
nand U41083 (N_41083,N_39326,N_38517);
or U41084 (N_41084,N_39094,N_38422);
and U41085 (N_41085,N_38306,N_38871);
and U41086 (N_41086,N_39990,N_39127);
and U41087 (N_41087,N_39142,N_39559);
or U41088 (N_41088,N_38909,N_39774);
nor U41089 (N_41089,N_39637,N_39581);
and U41090 (N_41090,N_38183,N_39923);
or U41091 (N_41091,N_39434,N_39415);
nand U41092 (N_41092,N_38979,N_39770);
and U41093 (N_41093,N_38253,N_38368);
or U41094 (N_41094,N_39932,N_38521);
or U41095 (N_41095,N_39250,N_39215);
or U41096 (N_41096,N_38323,N_39495);
or U41097 (N_41097,N_39128,N_38725);
nand U41098 (N_41098,N_39580,N_38654);
nor U41099 (N_41099,N_39267,N_39183);
or U41100 (N_41100,N_38039,N_39946);
or U41101 (N_41101,N_39392,N_39743);
nand U41102 (N_41102,N_39936,N_38384);
or U41103 (N_41103,N_38764,N_39577);
and U41104 (N_41104,N_38632,N_39547);
nand U41105 (N_41105,N_39793,N_38148);
and U41106 (N_41106,N_38223,N_38940);
nand U41107 (N_41107,N_38636,N_39651);
or U41108 (N_41108,N_38868,N_39287);
and U41109 (N_41109,N_38422,N_39287);
or U41110 (N_41110,N_38156,N_38408);
nand U41111 (N_41111,N_39479,N_38628);
nor U41112 (N_41112,N_39392,N_38789);
nand U41113 (N_41113,N_39826,N_39321);
nand U41114 (N_41114,N_38930,N_39743);
nand U41115 (N_41115,N_38322,N_38740);
and U41116 (N_41116,N_39405,N_38215);
nor U41117 (N_41117,N_38972,N_38065);
and U41118 (N_41118,N_38449,N_38094);
nand U41119 (N_41119,N_38385,N_39945);
and U41120 (N_41120,N_38437,N_38984);
or U41121 (N_41121,N_39062,N_38584);
and U41122 (N_41122,N_38839,N_39439);
nor U41123 (N_41123,N_38497,N_38104);
nor U41124 (N_41124,N_39247,N_38561);
or U41125 (N_41125,N_39957,N_38465);
nor U41126 (N_41126,N_39311,N_38545);
xnor U41127 (N_41127,N_39194,N_39665);
and U41128 (N_41128,N_38280,N_39795);
and U41129 (N_41129,N_39916,N_39292);
nor U41130 (N_41130,N_39144,N_38906);
nand U41131 (N_41131,N_38469,N_38478);
nor U41132 (N_41132,N_39269,N_39460);
or U41133 (N_41133,N_38772,N_38841);
nand U41134 (N_41134,N_38771,N_39746);
or U41135 (N_41135,N_38257,N_39089);
and U41136 (N_41136,N_39997,N_38352);
and U41137 (N_41137,N_39817,N_39646);
and U41138 (N_41138,N_39920,N_38495);
nor U41139 (N_41139,N_39688,N_38493);
and U41140 (N_41140,N_38766,N_39914);
and U41141 (N_41141,N_39780,N_39739);
and U41142 (N_41142,N_39471,N_38346);
nor U41143 (N_41143,N_38650,N_38368);
or U41144 (N_41144,N_39451,N_38234);
nor U41145 (N_41145,N_39410,N_38368);
nor U41146 (N_41146,N_38213,N_38061);
nand U41147 (N_41147,N_39071,N_38321);
nor U41148 (N_41148,N_39773,N_39565);
nand U41149 (N_41149,N_38159,N_39134);
and U41150 (N_41150,N_39750,N_39172);
and U41151 (N_41151,N_38417,N_38379);
nor U41152 (N_41152,N_39999,N_38637);
nand U41153 (N_41153,N_38880,N_39913);
nor U41154 (N_41154,N_38689,N_39489);
and U41155 (N_41155,N_38335,N_39203);
and U41156 (N_41156,N_39749,N_38739);
nand U41157 (N_41157,N_38141,N_38381);
and U41158 (N_41158,N_38536,N_39956);
nand U41159 (N_41159,N_38327,N_38082);
nor U41160 (N_41160,N_38449,N_38740);
and U41161 (N_41161,N_38686,N_39384);
or U41162 (N_41162,N_38467,N_39697);
or U41163 (N_41163,N_38345,N_38475);
nand U41164 (N_41164,N_39326,N_39773);
nand U41165 (N_41165,N_38674,N_39663);
nor U41166 (N_41166,N_38464,N_39045);
nor U41167 (N_41167,N_39590,N_39146);
nor U41168 (N_41168,N_38726,N_39501);
nand U41169 (N_41169,N_38580,N_38297);
or U41170 (N_41170,N_38265,N_38650);
nor U41171 (N_41171,N_38887,N_39205);
and U41172 (N_41172,N_39354,N_39665);
nand U41173 (N_41173,N_39436,N_39167);
or U41174 (N_41174,N_38481,N_39478);
nand U41175 (N_41175,N_39938,N_38243);
nor U41176 (N_41176,N_38587,N_39213);
or U41177 (N_41177,N_39774,N_38211);
and U41178 (N_41178,N_39323,N_38136);
nor U41179 (N_41179,N_38747,N_39581);
nand U41180 (N_41180,N_38170,N_39239);
or U41181 (N_41181,N_39225,N_39348);
nand U41182 (N_41182,N_39091,N_39570);
or U41183 (N_41183,N_38146,N_39599);
or U41184 (N_41184,N_39885,N_38638);
nand U41185 (N_41185,N_39143,N_39111);
nand U41186 (N_41186,N_38457,N_38320);
nor U41187 (N_41187,N_39677,N_38546);
nand U41188 (N_41188,N_38842,N_38297);
nor U41189 (N_41189,N_39977,N_38052);
or U41190 (N_41190,N_38542,N_39342);
and U41191 (N_41191,N_38039,N_38785);
or U41192 (N_41192,N_39755,N_38884);
nor U41193 (N_41193,N_38002,N_38718);
nand U41194 (N_41194,N_39103,N_38619);
or U41195 (N_41195,N_39502,N_38730);
nor U41196 (N_41196,N_38508,N_38963);
and U41197 (N_41197,N_39849,N_38441);
nand U41198 (N_41198,N_39733,N_38184);
nor U41199 (N_41199,N_38791,N_38773);
nand U41200 (N_41200,N_39529,N_39103);
and U41201 (N_41201,N_38833,N_38247);
nor U41202 (N_41202,N_38960,N_38701);
and U41203 (N_41203,N_39888,N_39661);
nand U41204 (N_41204,N_38651,N_38637);
or U41205 (N_41205,N_39597,N_39020);
nor U41206 (N_41206,N_38974,N_39606);
and U41207 (N_41207,N_39945,N_38396);
nor U41208 (N_41208,N_39936,N_38026);
or U41209 (N_41209,N_39956,N_39270);
nand U41210 (N_41210,N_38677,N_39546);
and U41211 (N_41211,N_38545,N_39519);
nor U41212 (N_41212,N_38729,N_38499);
and U41213 (N_41213,N_38064,N_38042);
or U41214 (N_41214,N_39279,N_39541);
nand U41215 (N_41215,N_38477,N_39461);
xor U41216 (N_41216,N_39984,N_38735);
nand U41217 (N_41217,N_39645,N_38834);
nor U41218 (N_41218,N_39138,N_38989);
nand U41219 (N_41219,N_39789,N_38738);
or U41220 (N_41220,N_39624,N_39422);
nor U41221 (N_41221,N_39857,N_38921);
nand U41222 (N_41222,N_39221,N_39613);
xnor U41223 (N_41223,N_39686,N_38922);
nand U41224 (N_41224,N_39954,N_38922);
and U41225 (N_41225,N_38214,N_38679);
nand U41226 (N_41226,N_38171,N_39234);
nand U41227 (N_41227,N_38179,N_38587);
nand U41228 (N_41228,N_39457,N_39133);
or U41229 (N_41229,N_38866,N_39197);
and U41230 (N_41230,N_38649,N_38655);
and U41231 (N_41231,N_39781,N_38858);
or U41232 (N_41232,N_39394,N_38890);
xnor U41233 (N_41233,N_38338,N_39028);
nand U41234 (N_41234,N_38380,N_39113);
nand U41235 (N_41235,N_38845,N_38355);
nand U41236 (N_41236,N_38024,N_39365);
or U41237 (N_41237,N_39356,N_38449);
nand U41238 (N_41238,N_38032,N_39657);
and U41239 (N_41239,N_38569,N_39848);
nor U41240 (N_41240,N_39684,N_38034);
and U41241 (N_41241,N_38607,N_39284);
or U41242 (N_41242,N_39962,N_39388);
or U41243 (N_41243,N_38073,N_39240);
or U41244 (N_41244,N_39684,N_39879);
xnor U41245 (N_41245,N_39073,N_39902);
nor U41246 (N_41246,N_38992,N_39742);
or U41247 (N_41247,N_39093,N_39500);
nor U41248 (N_41248,N_39104,N_39673);
or U41249 (N_41249,N_39055,N_38663);
nor U41250 (N_41250,N_38188,N_38433);
and U41251 (N_41251,N_39879,N_38599);
nand U41252 (N_41252,N_38593,N_39653);
nor U41253 (N_41253,N_38237,N_38954);
nor U41254 (N_41254,N_38150,N_39598);
nor U41255 (N_41255,N_39910,N_38034);
or U41256 (N_41256,N_39853,N_39712);
or U41257 (N_41257,N_38327,N_39434);
nand U41258 (N_41258,N_38460,N_39381);
and U41259 (N_41259,N_39300,N_39393);
or U41260 (N_41260,N_39950,N_38118);
or U41261 (N_41261,N_38338,N_39676);
nand U41262 (N_41262,N_38784,N_38789);
nand U41263 (N_41263,N_39655,N_38678);
nand U41264 (N_41264,N_38532,N_39092);
or U41265 (N_41265,N_39757,N_39086);
nor U41266 (N_41266,N_38486,N_38107);
nand U41267 (N_41267,N_39753,N_39172);
nor U41268 (N_41268,N_38996,N_38972);
nor U41269 (N_41269,N_39066,N_38572);
or U41270 (N_41270,N_38083,N_38453);
and U41271 (N_41271,N_38764,N_39446);
and U41272 (N_41272,N_39569,N_39262);
nand U41273 (N_41273,N_39868,N_38450);
and U41274 (N_41274,N_38855,N_39599);
nand U41275 (N_41275,N_39391,N_39756);
and U41276 (N_41276,N_39401,N_39088);
and U41277 (N_41277,N_38132,N_38255);
nor U41278 (N_41278,N_39727,N_39829);
or U41279 (N_41279,N_39587,N_39803);
nor U41280 (N_41280,N_38332,N_39274);
xnor U41281 (N_41281,N_39140,N_39378);
nor U41282 (N_41282,N_38295,N_39519);
nor U41283 (N_41283,N_38439,N_39345);
nand U41284 (N_41284,N_38595,N_39105);
nor U41285 (N_41285,N_39182,N_38328);
nor U41286 (N_41286,N_38446,N_38697);
or U41287 (N_41287,N_39361,N_38181);
nand U41288 (N_41288,N_39627,N_39359);
and U41289 (N_41289,N_39879,N_39581);
or U41290 (N_41290,N_39697,N_38962);
nand U41291 (N_41291,N_38667,N_39787);
and U41292 (N_41292,N_39839,N_38276);
or U41293 (N_41293,N_39426,N_39934);
and U41294 (N_41294,N_39079,N_39040);
nor U41295 (N_41295,N_38498,N_39262);
nor U41296 (N_41296,N_39243,N_38226);
nand U41297 (N_41297,N_38103,N_38985);
nand U41298 (N_41298,N_39319,N_39285);
nand U41299 (N_41299,N_38150,N_39309);
nand U41300 (N_41300,N_38198,N_38395);
nand U41301 (N_41301,N_38122,N_39308);
or U41302 (N_41302,N_38097,N_39712);
nor U41303 (N_41303,N_39995,N_39666);
or U41304 (N_41304,N_38459,N_39725);
nand U41305 (N_41305,N_38551,N_38466);
nor U41306 (N_41306,N_39923,N_38054);
or U41307 (N_41307,N_39420,N_39400);
or U41308 (N_41308,N_39647,N_38838);
nor U41309 (N_41309,N_38171,N_38226);
nor U41310 (N_41310,N_38401,N_38664);
nor U41311 (N_41311,N_39360,N_38678);
or U41312 (N_41312,N_39505,N_38679);
nor U41313 (N_41313,N_39136,N_39091);
nor U41314 (N_41314,N_38608,N_38600);
nor U41315 (N_41315,N_39522,N_38736);
and U41316 (N_41316,N_39000,N_38678);
nand U41317 (N_41317,N_38767,N_38907);
nor U41318 (N_41318,N_38408,N_39915);
or U41319 (N_41319,N_39646,N_39316);
nand U41320 (N_41320,N_39922,N_39865);
nand U41321 (N_41321,N_38818,N_38951);
and U41322 (N_41322,N_39512,N_38240);
nor U41323 (N_41323,N_39833,N_38738);
nand U41324 (N_41324,N_38099,N_38919);
and U41325 (N_41325,N_38300,N_38077);
or U41326 (N_41326,N_39437,N_39030);
and U41327 (N_41327,N_39547,N_38785);
and U41328 (N_41328,N_39320,N_39788);
nor U41329 (N_41329,N_38566,N_39691);
and U41330 (N_41330,N_39867,N_39487);
or U41331 (N_41331,N_39338,N_39403);
nor U41332 (N_41332,N_38314,N_38763);
or U41333 (N_41333,N_39663,N_39879);
or U41334 (N_41334,N_39520,N_38508);
nor U41335 (N_41335,N_38496,N_39835);
nor U41336 (N_41336,N_39385,N_39557);
or U41337 (N_41337,N_38239,N_38312);
nand U41338 (N_41338,N_39004,N_39615);
and U41339 (N_41339,N_38748,N_39028);
nor U41340 (N_41340,N_38497,N_39019);
or U41341 (N_41341,N_39136,N_39529);
nand U41342 (N_41342,N_39447,N_38362);
nand U41343 (N_41343,N_38545,N_39580);
nor U41344 (N_41344,N_39181,N_39804);
and U41345 (N_41345,N_38259,N_39475);
nand U41346 (N_41346,N_38899,N_38048);
and U41347 (N_41347,N_39717,N_38194);
and U41348 (N_41348,N_38759,N_38050);
and U41349 (N_41349,N_38718,N_38314);
nand U41350 (N_41350,N_38851,N_38683);
or U41351 (N_41351,N_38553,N_38250);
or U41352 (N_41352,N_38204,N_38963);
and U41353 (N_41353,N_38454,N_39876);
nor U41354 (N_41354,N_38754,N_38023);
or U41355 (N_41355,N_38655,N_38265);
or U41356 (N_41356,N_39919,N_38066);
nand U41357 (N_41357,N_38728,N_39679);
nor U41358 (N_41358,N_38529,N_39368);
or U41359 (N_41359,N_38929,N_38864);
or U41360 (N_41360,N_39544,N_39139);
or U41361 (N_41361,N_39375,N_39892);
and U41362 (N_41362,N_38890,N_38693);
and U41363 (N_41363,N_38978,N_38814);
and U41364 (N_41364,N_39580,N_39108);
or U41365 (N_41365,N_39291,N_39473);
nand U41366 (N_41366,N_39084,N_38505);
and U41367 (N_41367,N_38895,N_38772);
nand U41368 (N_41368,N_38626,N_38117);
and U41369 (N_41369,N_38420,N_39047);
nand U41370 (N_41370,N_39463,N_38879);
nor U41371 (N_41371,N_38350,N_38325);
nand U41372 (N_41372,N_38971,N_39174);
and U41373 (N_41373,N_38637,N_38863);
and U41374 (N_41374,N_38893,N_39154);
nor U41375 (N_41375,N_38664,N_38896);
and U41376 (N_41376,N_38274,N_38712);
and U41377 (N_41377,N_39736,N_39790);
nand U41378 (N_41378,N_39861,N_38410);
nand U41379 (N_41379,N_39902,N_39820);
and U41380 (N_41380,N_39934,N_38481);
and U41381 (N_41381,N_39856,N_38430);
nand U41382 (N_41382,N_39863,N_39908);
xnor U41383 (N_41383,N_38995,N_38124);
or U41384 (N_41384,N_39678,N_39475);
and U41385 (N_41385,N_38378,N_39445);
xor U41386 (N_41386,N_39847,N_39945);
and U41387 (N_41387,N_39747,N_38547);
or U41388 (N_41388,N_39630,N_39608);
and U41389 (N_41389,N_38547,N_39789);
and U41390 (N_41390,N_39901,N_38660);
nand U41391 (N_41391,N_39342,N_39263);
nor U41392 (N_41392,N_38957,N_38551);
nor U41393 (N_41393,N_38861,N_39884);
or U41394 (N_41394,N_39211,N_38526);
xnor U41395 (N_41395,N_38742,N_38385);
or U41396 (N_41396,N_39165,N_39811);
nor U41397 (N_41397,N_38097,N_39560);
nand U41398 (N_41398,N_39473,N_39873);
nand U41399 (N_41399,N_38102,N_39422);
nand U41400 (N_41400,N_38411,N_38170);
or U41401 (N_41401,N_38659,N_39328);
and U41402 (N_41402,N_39758,N_38090);
and U41403 (N_41403,N_39334,N_39300);
nand U41404 (N_41404,N_39795,N_39315);
nor U41405 (N_41405,N_38009,N_38342);
and U41406 (N_41406,N_39264,N_38070);
nor U41407 (N_41407,N_39928,N_39253);
and U41408 (N_41408,N_39483,N_39839);
nor U41409 (N_41409,N_38457,N_38494);
and U41410 (N_41410,N_39360,N_38276);
and U41411 (N_41411,N_38508,N_38997);
or U41412 (N_41412,N_38359,N_39316);
nand U41413 (N_41413,N_38718,N_39460);
or U41414 (N_41414,N_39737,N_39173);
nor U41415 (N_41415,N_38826,N_38342);
or U41416 (N_41416,N_38267,N_39997);
and U41417 (N_41417,N_38484,N_38760);
or U41418 (N_41418,N_38093,N_39479);
or U41419 (N_41419,N_38321,N_39510);
nand U41420 (N_41420,N_38939,N_38927);
nand U41421 (N_41421,N_38439,N_38412);
nor U41422 (N_41422,N_38460,N_39256);
nand U41423 (N_41423,N_39162,N_39764);
nor U41424 (N_41424,N_39050,N_38168);
nand U41425 (N_41425,N_38569,N_39593);
nand U41426 (N_41426,N_39755,N_38857);
or U41427 (N_41427,N_39121,N_39894);
or U41428 (N_41428,N_38514,N_38343);
nor U41429 (N_41429,N_38686,N_39126);
nand U41430 (N_41430,N_39107,N_39740);
nor U41431 (N_41431,N_38824,N_39899);
and U41432 (N_41432,N_39174,N_39532);
nor U41433 (N_41433,N_38399,N_39209);
nor U41434 (N_41434,N_38953,N_39383);
nand U41435 (N_41435,N_39462,N_39294);
and U41436 (N_41436,N_38639,N_39622);
nor U41437 (N_41437,N_39062,N_38288);
xor U41438 (N_41438,N_38914,N_39576);
or U41439 (N_41439,N_38747,N_38004);
nor U41440 (N_41440,N_39935,N_38997);
and U41441 (N_41441,N_39316,N_39683);
or U41442 (N_41442,N_38794,N_39269);
and U41443 (N_41443,N_38191,N_39757);
nand U41444 (N_41444,N_39153,N_38638);
and U41445 (N_41445,N_39121,N_39262);
and U41446 (N_41446,N_39489,N_39536);
and U41447 (N_41447,N_38635,N_39826);
or U41448 (N_41448,N_39661,N_38789);
or U41449 (N_41449,N_38861,N_38066);
nor U41450 (N_41450,N_38941,N_38848);
and U41451 (N_41451,N_38867,N_39818);
nor U41452 (N_41452,N_38736,N_38201);
nand U41453 (N_41453,N_38635,N_38662);
nor U41454 (N_41454,N_38470,N_38127);
nor U41455 (N_41455,N_39985,N_38553);
nand U41456 (N_41456,N_38439,N_38327);
nand U41457 (N_41457,N_39961,N_38480);
and U41458 (N_41458,N_39954,N_38422);
nand U41459 (N_41459,N_39940,N_38466);
or U41460 (N_41460,N_38407,N_38114);
nor U41461 (N_41461,N_39709,N_39011);
nand U41462 (N_41462,N_39069,N_38823);
and U41463 (N_41463,N_39328,N_38137);
or U41464 (N_41464,N_39603,N_39676);
and U41465 (N_41465,N_38959,N_39399);
or U41466 (N_41466,N_39923,N_38016);
or U41467 (N_41467,N_38029,N_38489);
nand U41468 (N_41468,N_38759,N_39682);
or U41469 (N_41469,N_38668,N_38358);
nor U41470 (N_41470,N_39065,N_38061);
and U41471 (N_41471,N_39597,N_39094);
or U41472 (N_41472,N_38958,N_39147);
nand U41473 (N_41473,N_38028,N_38783);
or U41474 (N_41474,N_39683,N_38253);
and U41475 (N_41475,N_39547,N_38641);
nor U41476 (N_41476,N_38900,N_39091);
or U41477 (N_41477,N_39730,N_38876);
or U41478 (N_41478,N_38000,N_38967);
or U41479 (N_41479,N_38541,N_39217);
nand U41480 (N_41480,N_39028,N_38358);
nand U41481 (N_41481,N_38096,N_38869);
nor U41482 (N_41482,N_39628,N_38154);
nand U41483 (N_41483,N_39423,N_38970);
nor U41484 (N_41484,N_38831,N_39553);
and U41485 (N_41485,N_38433,N_39341);
nand U41486 (N_41486,N_38925,N_38001);
or U41487 (N_41487,N_39008,N_39999);
nor U41488 (N_41488,N_38676,N_39363);
or U41489 (N_41489,N_39324,N_39177);
nor U41490 (N_41490,N_39169,N_38656);
nand U41491 (N_41491,N_38104,N_38630);
nand U41492 (N_41492,N_38104,N_39985);
nand U41493 (N_41493,N_39273,N_38363);
nor U41494 (N_41494,N_39120,N_39670);
and U41495 (N_41495,N_38034,N_38621);
and U41496 (N_41496,N_38094,N_38501);
or U41497 (N_41497,N_39567,N_38991);
nand U41498 (N_41498,N_39055,N_38134);
nand U41499 (N_41499,N_39669,N_39664);
or U41500 (N_41500,N_38575,N_39904);
and U41501 (N_41501,N_39485,N_39247);
and U41502 (N_41502,N_39418,N_38038);
or U41503 (N_41503,N_38663,N_38781);
nor U41504 (N_41504,N_39040,N_38599);
xor U41505 (N_41505,N_38973,N_38133);
nor U41506 (N_41506,N_39981,N_38243);
or U41507 (N_41507,N_39768,N_39594);
xor U41508 (N_41508,N_38498,N_39064);
nand U41509 (N_41509,N_39864,N_39179);
and U41510 (N_41510,N_38519,N_38523);
nor U41511 (N_41511,N_39519,N_38168);
or U41512 (N_41512,N_39120,N_38618);
nand U41513 (N_41513,N_39385,N_39591);
nand U41514 (N_41514,N_39664,N_39478);
nand U41515 (N_41515,N_39673,N_39679);
nand U41516 (N_41516,N_39015,N_39384);
nor U41517 (N_41517,N_38646,N_39108);
nand U41518 (N_41518,N_39089,N_39756);
nand U41519 (N_41519,N_39908,N_38999);
or U41520 (N_41520,N_39351,N_38498);
or U41521 (N_41521,N_38612,N_38980);
or U41522 (N_41522,N_38711,N_38953);
and U41523 (N_41523,N_38938,N_38844);
nor U41524 (N_41524,N_38320,N_39551);
or U41525 (N_41525,N_39940,N_39273);
or U41526 (N_41526,N_39369,N_38872);
and U41527 (N_41527,N_38600,N_39766);
nor U41528 (N_41528,N_39903,N_38877);
nor U41529 (N_41529,N_38271,N_38528);
nand U41530 (N_41530,N_38338,N_39960);
or U41531 (N_41531,N_39773,N_38876);
xor U41532 (N_41532,N_39297,N_38190);
nand U41533 (N_41533,N_39470,N_39225);
and U41534 (N_41534,N_39207,N_38946);
and U41535 (N_41535,N_38040,N_39469);
nor U41536 (N_41536,N_38059,N_39536);
nand U41537 (N_41537,N_39792,N_39359);
and U41538 (N_41538,N_38716,N_38743);
and U41539 (N_41539,N_39047,N_38026);
nor U41540 (N_41540,N_39598,N_38192);
xor U41541 (N_41541,N_38833,N_39220);
or U41542 (N_41542,N_39804,N_38350);
nand U41543 (N_41543,N_39783,N_38636);
nor U41544 (N_41544,N_38111,N_38171);
and U41545 (N_41545,N_38755,N_38386);
nor U41546 (N_41546,N_39573,N_39471);
nand U41547 (N_41547,N_38415,N_38135);
and U41548 (N_41548,N_38383,N_39197);
or U41549 (N_41549,N_38037,N_39919);
or U41550 (N_41550,N_39399,N_38305);
nor U41551 (N_41551,N_38568,N_39008);
nor U41552 (N_41552,N_39805,N_39034);
and U41553 (N_41553,N_38304,N_38705);
nor U41554 (N_41554,N_38413,N_38143);
nor U41555 (N_41555,N_38000,N_38985);
nor U41556 (N_41556,N_38723,N_39746);
and U41557 (N_41557,N_38899,N_38178);
and U41558 (N_41558,N_39606,N_38144);
nor U41559 (N_41559,N_38806,N_38726);
and U41560 (N_41560,N_39704,N_39452);
and U41561 (N_41561,N_39514,N_39835);
and U41562 (N_41562,N_39637,N_39797);
and U41563 (N_41563,N_38775,N_39314);
and U41564 (N_41564,N_39276,N_38347);
or U41565 (N_41565,N_39585,N_39879);
nand U41566 (N_41566,N_38942,N_39441);
nand U41567 (N_41567,N_38030,N_39170);
or U41568 (N_41568,N_38450,N_39035);
nand U41569 (N_41569,N_38291,N_38292);
or U41570 (N_41570,N_38861,N_38493);
and U41571 (N_41571,N_39474,N_39967);
or U41572 (N_41572,N_39152,N_39908);
or U41573 (N_41573,N_39575,N_39209);
nand U41574 (N_41574,N_39221,N_38697);
nor U41575 (N_41575,N_39749,N_38659);
nand U41576 (N_41576,N_38640,N_39664);
nand U41577 (N_41577,N_38035,N_38921);
xnor U41578 (N_41578,N_38675,N_39659);
nand U41579 (N_41579,N_38005,N_39043);
and U41580 (N_41580,N_39130,N_38708);
or U41581 (N_41581,N_39695,N_38067);
nor U41582 (N_41582,N_39744,N_38910);
nor U41583 (N_41583,N_39383,N_39869);
and U41584 (N_41584,N_39936,N_39967);
and U41585 (N_41585,N_38301,N_38721);
nand U41586 (N_41586,N_38713,N_39419);
nor U41587 (N_41587,N_38900,N_38808);
or U41588 (N_41588,N_38206,N_38102);
nand U41589 (N_41589,N_38145,N_39682);
nand U41590 (N_41590,N_38719,N_39216);
nor U41591 (N_41591,N_38033,N_38438);
and U41592 (N_41592,N_38789,N_38192);
nor U41593 (N_41593,N_38335,N_38886);
nand U41594 (N_41594,N_39372,N_38088);
and U41595 (N_41595,N_39762,N_39678);
nor U41596 (N_41596,N_38220,N_38826);
nor U41597 (N_41597,N_39188,N_38189);
xnor U41598 (N_41598,N_39471,N_39160);
and U41599 (N_41599,N_38407,N_39272);
or U41600 (N_41600,N_39983,N_38224);
or U41601 (N_41601,N_39489,N_38147);
or U41602 (N_41602,N_39655,N_38646);
or U41603 (N_41603,N_39824,N_39008);
nor U41604 (N_41604,N_38059,N_39878);
nand U41605 (N_41605,N_39810,N_38415);
and U41606 (N_41606,N_39928,N_38227);
and U41607 (N_41607,N_38850,N_39894);
or U41608 (N_41608,N_38643,N_39221);
nand U41609 (N_41609,N_39474,N_38622);
and U41610 (N_41610,N_39268,N_38872);
and U41611 (N_41611,N_38588,N_39945);
nand U41612 (N_41612,N_38812,N_38919);
and U41613 (N_41613,N_38867,N_39068);
and U41614 (N_41614,N_38978,N_39843);
nand U41615 (N_41615,N_39036,N_38840);
or U41616 (N_41616,N_38464,N_39580);
and U41617 (N_41617,N_39870,N_38807);
nand U41618 (N_41618,N_38502,N_39835);
or U41619 (N_41619,N_39946,N_39730);
nand U41620 (N_41620,N_38862,N_39336);
and U41621 (N_41621,N_38980,N_38631);
nand U41622 (N_41622,N_38884,N_38678);
and U41623 (N_41623,N_38076,N_38937);
nor U41624 (N_41624,N_39880,N_38502);
or U41625 (N_41625,N_39268,N_38651);
nor U41626 (N_41626,N_39289,N_39265);
nand U41627 (N_41627,N_38410,N_39420);
nand U41628 (N_41628,N_39028,N_39480);
and U41629 (N_41629,N_38558,N_38564);
and U41630 (N_41630,N_39434,N_39263);
and U41631 (N_41631,N_38195,N_39874);
and U41632 (N_41632,N_39594,N_38221);
or U41633 (N_41633,N_39492,N_39702);
or U41634 (N_41634,N_38630,N_38022);
nand U41635 (N_41635,N_38615,N_39676);
nand U41636 (N_41636,N_39397,N_39282);
nor U41637 (N_41637,N_39448,N_39071);
nor U41638 (N_41638,N_39448,N_39879);
or U41639 (N_41639,N_39238,N_39229);
or U41640 (N_41640,N_38934,N_39906);
nand U41641 (N_41641,N_38092,N_39741);
and U41642 (N_41642,N_39670,N_39263);
and U41643 (N_41643,N_39030,N_38664);
nand U41644 (N_41644,N_38569,N_38646);
nand U41645 (N_41645,N_38663,N_38339);
or U41646 (N_41646,N_38409,N_38826);
and U41647 (N_41647,N_38874,N_39681);
and U41648 (N_41648,N_38918,N_39011);
and U41649 (N_41649,N_39718,N_39861);
nor U41650 (N_41650,N_38880,N_38577);
nor U41651 (N_41651,N_38425,N_38083);
nor U41652 (N_41652,N_38239,N_39136);
nor U41653 (N_41653,N_39692,N_38416);
nand U41654 (N_41654,N_39338,N_38501);
nor U41655 (N_41655,N_39636,N_38817);
and U41656 (N_41656,N_39881,N_39391);
or U41657 (N_41657,N_38107,N_38981);
nand U41658 (N_41658,N_39420,N_39138);
or U41659 (N_41659,N_39153,N_39297);
xnor U41660 (N_41660,N_39832,N_38892);
and U41661 (N_41661,N_39804,N_38388);
nor U41662 (N_41662,N_38633,N_39802);
or U41663 (N_41663,N_38095,N_39765);
nor U41664 (N_41664,N_39420,N_38702);
or U41665 (N_41665,N_39445,N_38747);
nand U41666 (N_41666,N_38314,N_38165);
nand U41667 (N_41667,N_39086,N_39306);
and U41668 (N_41668,N_39997,N_39098);
or U41669 (N_41669,N_39585,N_38301);
and U41670 (N_41670,N_39138,N_39647);
or U41671 (N_41671,N_38707,N_39261);
nand U41672 (N_41672,N_38516,N_39834);
and U41673 (N_41673,N_38271,N_39256);
nand U41674 (N_41674,N_38960,N_39492);
nand U41675 (N_41675,N_38507,N_39186);
and U41676 (N_41676,N_38500,N_39984);
nor U41677 (N_41677,N_39055,N_38996);
and U41678 (N_41678,N_39640,N_39418);
nor U41679 (N_41679,N_38689,N_39368);
nor U41680 (N_41680,N_38111,N_39358);
xor U41681 (N_41681,N_39565,N_39450);
nor U41682 (N_41682,N_39808,N_39219);
xor U41683 (N_41683,N_39530,N_38124);
or U41684 (N_41684,N_38134,N_38000);
nand U41685 (N_41685,N_38010,N_39615);
nand U41686 (N_41686,N_39280,N_38576);
or U41687 (N_41687,N_38430,N_39983);
nand U41688 (N_41688,N_38077,N_38455);
and U41689 (N_41689,N_39661,N_39880);
and U41690 (N_41690,N_38054,N_38710);
nand U41691 (N_41691,N_39037,N_39254);
and U41692 (N_41692,N_39721,N_39630);
or U41693 (N_41693,N_39102,N_38001);
or U41694 (N_41694,N_39407,N_38560);
and U41695 (N_41695,N_39325,N_38490);
and U41696 (N_41696,N_39938,N_38113);
and U41697 (N_41697,N_38369,N_38700);
or U41698 (N_41698,N_38154,N_39452);
nand U41699 (N_41699,N_39256,N_39829);
nand U41700 (N_41700,N_38354,N_39188);
and U41701 (N_41701,N_39535,N_39439);
or U41702 (N_41702,N_39776,N_39315);
nor U41703 (N_41703,N_39663,N_38462);
xor U41704 (N_41704,N_38039,N_39626);
and U41705 (N_41705,N_38221,N_38015);
nor U41706 (N_41706,N_38050,N_38010);
nor U41707 (N_41707,N_39672,N_39039);
and U41708 (N_41708,N_38945,N_39732);
xor U41709 (N_41709,N_38479,N_38905);
nor U41710 (N_41710,N_39748,N_38464);
or U41711 (N_41711,N_39009,N_39451);
and U41712 (N_41712,N_39844,N_38924);
xnor U41713 (N_41713,N_39541,N_38755);
nand U41714 (N_41714,N_38008,N_38537);
nand U41715 (N_41715,N_38564,N_38460);
or U41716 (N_41716,N_39561,N_39202);
nor U41717 (N_41717,N_38396,N_38343);
xor U41718 (N_41718,N_39188,N_38143);
or U41719 (N_41719,N_39727,N_38664);
and U41720 (N_41720,N_38674,N_38776);
nand U41721 (N_41721,N_38301,N_38123);
nand U41722 (N_41722,N_39138,N_39664);
nor U41723 (N_41723,N_39143,N_39333);
or U41724 (N_41724,N_39033,N_38804);
or U41725 (N_41725,N_38701,N_39650);
or U41726 (N_41726,N_38275,N_38444);
nand U41727 (N_41727,N_39953,N_39443);
and U41728 (N_41728,N_38453,N_38615);
or U41729 (N_41729,N_38459,N_39739);
nor U41730 (N_41730,N_38954,N_39883);
and U41731 (N_41731,N_38947,N_38108);
nor U41732 (N_41732,N_39647,N_39638);
nor U41733 (N_41733,N_38331,N_38991);
nand U41734 (N_41734,N_39945,N_39966);
and U41735 (N_41735,N_38570,N_39560);
and U41736 (N_41736,N_38099,N_38743);
nand U41737 (N_41737,N_38392,N_38423);
nor U41738 (N_41738,N_39486,N_39031);
or U41739 (N_41739,N_39241,N_39707);
or U41740 (N_41740,N_38295,N_39445);
nor U41741 (N_41741,N_38388,N_39603);
and U41742 (N_41742,N_39704,N_38853);
or U41743 (N_41743,N_38367,N_38042);
or U41744 (N_41744,N_39852,N_39864);
or U41745 (N_41745,N_38167,N_38120);
nor U41746 (N_41746,N_38770,N_38097);
nor U41747 (N_41747,N_38044,N_39010);
nand U41748 (N_41748,N_39259,N_39923);
and U41749 (N_41749,N_38945,N_39590);
nand U41750 (N_41750,N_38619,N_39352);
nor U41751 (N_41751,N_39597,N_39919);
nor U41752 (N_41752,N_38336,N_38572);
nand U41753 (N_41753,N_38976,N_38694);
and U41754 (N_41754,N_39002,N_38984);
nor U41755 (N_41755,N_39403,N_38117);
nand U41756 (N_41756,N_39769,N_38623);
nor U41757 (N_41757,N_39488,N_38308);
or U41758 (N_41758,N_39108,N_38551);
and U41759 (N_41759,N_38577,N_39336);
and U41760 (N_41760,N_38198,N_38889);
nor U41761 (N_41761,N_39202,N_38894);
and U41762 (N_41762,N_38585,N_38594);
or U41763 (N_41763,N_39729,N_38535);
or U41764 (N_41764,N_39693,N_39455);
or U41765 (N_41765,N_38752,N_39438);
and U41766 (N_41766,N_39809,N_39312);
nor U41767 (N_41767,N_38014,N_39795);
or U41768 (N_41768,N_38381,N_38807);
nand U41769 (N_41769,N_39058,N_39560);
or U41770 (N_41770,N_39938,N_39827);
or U41771 (N_41771,N_38866,N_39658);
nand U41772 (N_41772,N_38063,N_38404);
nor U41773 (N_41773,N_39752,N_39040);
and U41774 (N_41774,N_38271,N_38199);
nand U41775 (N_41775,N_39899,N_39969);
or U41776 (N_41776,N_39946,N_38529);
and U41777 (N_41777,N_38877,N_38883);
or U41778 (N_41778,N_38803,N_39151);
and U41779 (N_41779,N_39131,N_38068);
and U41780 (N_41780,N_39071,N_39711);
nand U41781 (N_41781,N_38915,N_39672);
nor U41782 (N_41782,N_38142,N_38913);
or U41783 (N_41783,N_39740,N_38792);
nor U41784 (N_41784,N_39720,N_39226);
nor U41785 (N_41785,N_38118,N_39377);
nor U41786 (N_41786,N_39996,N_38891);
xnor U41787 (N_41787,N_38171,N_38675);
nand U41788 (N_41788,N_38297,N_39146);
nor U41789 (N_41789,N_39817,N_38070);
nor U41790 (N_41790,N_38253,N_38975);
and U41791 (N_41791,N_38040,N_39191);
nor U41792 (N_41792,N_38336,N_39732);
or U41793 (N_41793,N_38911,N_39142);
nand U41794 (N_41794,N_38815,N_38298);
nand U41795 (N_41795,N_38865,N_39588);
or U41796 (N_41796,N_39868,N_39246);
nand U41797 (N_41797,N_39251,N_38880);
and U41798 (N_41798,N_38571,N_39087);
nand U41799 (N_41799,N_38491,N_38542);
and U41800 (N_41800,N_39288,N_38598);
or U41801 (N_41801,N_38069,N_38559);
nor U41802 (N_41802,N_38193,N_39723);
nand U41803 (N_41803,N_39483,N_38677);
nor U41804 (N_41804,N_39964,N_38863);
or U41805 (N_41805,N_39545,N_38048);
and U41806 (N_41806,N_38198,N_39449);
nor U41807 (N_41807,N_39636,N_38235);
nor U41808 (N_41808,N_38096,N_38387);
xor U41809 (N_41809,N_38424,N_38463);
nand U41810 (N_41810,N_38119,N_38109);
or U41811 (N_41811,N_39378,N_39367);
or U41812 (N_41812,N_39131,N_39754);
nand U41813 (N_41813,N_38358,N_39751);
nor U41814 (N_41814,N_39239,N_39566);
and U41815 (N_41815,N_38287,N_38391);
nand U41816 (N_41816,N_38779,N_39931);
or U41817 (N_41817,N_38709,N_39442);
nor U41818 (N_41818,N_39544,N_39239);
or U41819 (N_41819,N_39852,N_39645);
and U41820 (N_41820,N_39772,N_39624);
or U41821 (N_41821,N_38311,N_38673);
nand U41822 (N_41822,N_39270,N_39525);
or U41823 (N_41823,N_38774,N_38380);
or U41824 (N_41824,N_39511,N_38545);
nor U41825 (N_41825,N_39957,N_39296);
nand U41826 (N_41826,N_39680,N_39087);
or U41827 (N_41827,N_38188,N_38161);
nand U41828 (N_41828,N_38511,N_38060);
nor U41829 (N_41829,N_39318,N_38968);
nand U41830 (N_41830,N_38358,N_39173);
nor U41831 (N_41831,N_39593,N_38913);
nand U41832 (N_41832,N_38654,N_39703);
nor U41833 (N_41833,N_39201,N_38167);
and U41834 (N_41834,N_38076,N_39834);
nand U41835 (N_41835,N_39892,N_39282);
nor U41836 (N_41836,N_39232,N_38247);
nor U41837 (N_41837,N_38925,N_39411);
nand U41838 (N_41838,N_38769,N_39136);
nor U41839 (N_41839,N_38391,N_38388);
nand U41840 (N_41840,N_39176,N_38631);
nand U41841 (N_41841,N_38719,N_38301);
nor U41842 (N_41842,N_39933,N_39020);
and U41843 (N_41843,N_39956,N_38012);
nor U41844 (N_41844,N_38383,N_38425);
nor U41845 (N_41845,N_38062,N_39122);
nor U41846 (N_41846,N_39800,N_38287);
or U41847 (N_41847,N_39406,N_38811);
or U41848 (N_41848,N_38525,N_38780);
nand U41849 (N_41849,N_39426,N_38289);
nand U41850 (N_41850,N_39343,N_38840);
and U41851 (N_41851,N_38019,N_38037);
nand U41852 (N_41852,N_39557,N_39353);
or U41853 (N_41853,N_39206,N_38607);
and U41854 (N_41854,N_39225,N_39946);
and U41855 (N_41855,N_38318,N_39213);
and U41856 (N_41856,N_39276,N_38066);
and U41857 (N_41857,N_38274,N_39245);
nor U41858 (N_41858,N_39435,N_39276);
nand U41859 (N_41859,N_39889,N_39576);
xor U41860 (N_41860,N_38242,N_38191);
and U41861 (N_41861,N_39774,N_38226);
or U41862 (N_41862,N_38483,N_38698);
or U41863 (N_41863,N_38674,N_38870);
nand U41864 (N_41864,N_38842,N_38968);
and U41865 (N_41865,N_39405,N_38034);
and U41866 (N_41866,N_39045,N_38122);
and U41867 (N_41867,N_38773,N_39642);
nand U41868 (N_41868,N_39499,N_38602);
nand U41869 (N_41869,N_39930,N_38133);
or U41870 (N_41870,N_39667,N_39822);
and U41871 (N_41871,N_38028,N_38532);
nor U41872 (N_41872,N_39889,N_39036);
or U41873 (N_41873,N_38924,N_38875);
or U41874 (N_41874,N_38955,N_39892);
or U41875 (N_41875,N_38477,N_38873);
and U41876 (N_41876,N_38451,N_38609);
or U41877 (N_41877,N_39660,N_38736);
nand U41878 (N_41878,N_39223,N_38338);
nor U41879 (N_41879,N_38188,N_38318);
or U41880 (N_41880,N_38264,N_38639);
or U41881 (N_41881,N_39929,N_39243);
or U41882 (N_41882,N_38995,N_38661);
nor U41883 (N_41883,N_38834,N_39637);
and U41884 (N_41884,N_39296,N_39598);
or U41885 (N_41885,N_39262,N_39350);
nor U41886 (N_41886,N_38951,N_38568);
or U41887 (N_41887,N_38451,N_39227);
and U41888 (N_41888,N_38811,N_39363);
xor U41889 (N_41889,N_39378,N_38812);
or U41890 (N_41890,N_38927,N_38546);
nand U41891 (N_41891,N_38332,N_39682);
nand U41892 (N_41892,N_39456,N_38086);
and U41893 (N_41893,N_39264,N_39947);
and U41894 (N_41894,N_38123,N_38464);
nor U41895 (N_41895,N_38150,N_38830);
nand U41896 (N_41896,N_38795,N_39136);
nand U41897 (N_41897,N_39395,N_39434);
and U41898 (N_41898,N_38279,N_38135);
xor U41899 (N_41899,N_38621,N_39292);
nand U41900 (N_41900,N_38991,N_38321);
or U41901 (N_41901,N_38554,N_39178);
nor U41902 (N_41902,N_38881,N_39510);
and U41903 (N_41903,N_39908,N_39391);
and U41904 (N_41904,N_39142,N_39720);
nor U41905 (N_41905,N_38291,N_38274);
or U41906 (N_41906,N_39278,N_38086);
nand U41907 (N_41907,N_39198,N_39281);
nor U41908 (N_41908,N_38762,N_38924);
or U41909 (N_41909,N_39028,N_39405);
or U41910 (N_41910,N_39666,N_39348);
nand U41911 (N_41911,N_39796,N_39153);
or U41912 (N_41912,N_38082,N_39523);
nor U41913 (N_41913,N_39178,N_38051);
nor U41914 (N_41914,N_38654,N_39604);
and U41915 (N_41915,N_38591,N_38618);
or U41916 (N_41916,N_38943,N_39401);
and U41917 (N_41917,N_38525,N_38017);
and U41918 (N_41918,N_38381,N_39402);
nand U41919 (N_41919,N_39445,N_38951);
nor U41920 (N_41920,N_38790,N_38039);
or U41921 (N_41921,N_38294,N_38161);
and U41922 (N_41922,N_39860,N_38682);
nor U41923 (N_41923,N_39426,N_39452);
and U41924 (N_41924,N_39456,N_39171);
nand U41925 (N_41925,N_38761,N_39247);
and U41926 (N_41926,N_38876,N_38501);
nor U41927 (N_41927,N_38618,N_38901);
or U41928 (N_41928,N_39591,N_39078);
nand U41929 (N_41929,N_38790,N_39057);
nor U41930 (N_41930,N_39787,N_39941);
nor U41931 (N_41931,N_39118,N_39055);
or U41932 (N_41932,N_39964,N_38315);
and U41933 (N_41933,N_38571,N_38679);
nand U41934 (N_41934,N_38064,N_38328);
and U41935 (N_41935,N_39647,N_39762);
nand U41936 (N_41936,N_38829,N_38000);
and U41937 (N_41937,N_39018,N_39860);
nor U41938 (N_41938,N_38776,N_39183);
nand U41939 (N_41939,N_38758,N_39722);
and U41940 (N_41940,N_39272,N_39068);
or U41941 (N_41941,N_38922,N_38562);
and U41942 (N_41942,N_38652,N_38573);
nor U41943 (N_41943,N_39495,N_38411);
or U41944 (N_41944,N_38395,N_38299);
and U41945 (N_41945,N_38967,N_39051);
nor U41946 (N_41946,N_39850,N_38698);
or U41947 (N_41947,N_39139,N_39750);
nand U41948 (N_41948,N_38547,N_39720);
nand U41949 (N_41949,N_39005,N_39355);
or U41950 (N_41950,N_39772,N_38712);
or U41951 (N_41951,N_38714,N_39981);
nor U41952 (N_41952,N_38381,N_39918);
or U41953 (N_41953,N_38030,N_39290);
nor U41954 (N_41954,N_38400,N_39550);
nor U41955 (N_41955,N_38153,N_38955);
or U41956 (N_41956,N_38154,N_39349);
nor U41957 (N_41957,N_39046,N_39744);
or U41958 (N_41958,N_38450,N_38772);
nand U41959 (N_41959,N_39364,N_38868);
nor U41960 (N_41960,N_38975,N_38089);
or U41961 (N_41961,N_38221,N_39932);
nand U41962 (N_41962,N_38512,N_39876);
and U41963 (N_41963,N_39542,N_38448);
nand U41964 (N_41964,N_38932,N_39151);
nor U41965 (N_41965,N_39319,N_38301);
or U41966 (N_41966,N_39957,N_39122);
and U41967 (N_41967,N_38253,N_38472);
nand U41968 (N_41968,N_38859,N_38589);
nor U41969 (N_41969,N_38930,N_38972);
nand U41970 (N_41970,N_38919,N_38954);
nor U41971 (N_41971,N_38144,N_38107);
and U41972 (N_41972,N_39145,N_38775);
nand U41973 (N_41973,N_39764,N_39371);
or U41974 (N_41974,N_39688,N_38418);
or U41975 (N_41975,N_39933,N_39265);
or U41976 (N_41976,N_39657,N_38688);
or U41977 (N_41977,N_39372,N_39512);
nand U41978 (N_41978,N_38866,N_38145);
or U41979 (N_41979,N_39775,N_38433);
nor U41980 (N_41980,N_39863,N_38582);
or U41981 (N_41981,N_38279,N_38858);
and U41982 (N_41982,N_39384,N_39667);
nor U41983 (N_41983,N_39843,N_38095);
nand U41984 (N_41984,N_39056,N_39691);
nor U41985 (N_41985,N_38606,N_39117);
or U41986 (N_41986,N_39240,N_38158);
nor U41987 (N_41987,N_39397,N_38816);
nand U41988 (N_41988,N_39226,N_39234);
and U41989 (N_41989,N_39952,N_38320);
or U41990 (N_41990,N_39136,N_39476);
and U41991 (N_41991,N_39556,N_38214);
nand U41992 (N_41992,N_38371,N_39083);
and U41993 (N_41993,N_39251,N_39980);
nor U41994 (N_41994,N_39992,N_39981);
nor U41995 (N_41995,N_38737,N_39155);
nand U41996 (N_41996,N_38712,N_39302);
and U41997 (N_41997,N_39882,N_39660);
or U41998 (N_41998,N_39801,N_39552);
or U41999 (N_41999,N_39662,N_39049);
nor U42000 (N_42000,N_40647,N_41400);
nand U42001 (N_42001,N_40001,N_40015);
nor U42002 (N_42002,N_41008,N_40207);
nor U42003 (N_42003,N_41371,N_40652);
nor U42004 (N_42004,N_41203,N_40136);
nor U42005 (N_42005,N_41897,N_40351);
or U42006 (N_42006,N_40567,N_41399);
or U42007 (N_42007,N_40365,N_41157);
nor U42008 (N_42008,N_41092,N_40154);
nor U42009 (N_42009,N_41293,N_40887);
or U42010 (N_42010,N_41802,N_41971);
and U42011 (N_42011,N_41094,N_40788);
nor U42012 (N_42012,N_40186,N_41450);
nand U42013 (N_42013,N_41103,N_41583);
nor U42014 (N_42014,N_41539,N_40398);
nor U42015 (N_42015,N_41719,N_40522);
xnor U42016 (N_42016,N_40843,N_40609);
nor U42017 (N_42017,N_40328,N_40244);
or U42018 (N_42018,N_40124,N_41618);
nor U42019 (N_42019,N_41771,N_40461);
and U42020 (N_42020,N_41975,N_41240);
nor U42021 (N_42021,N_40452,N_40261);
or U42022 (N_42022,N_41022,N_40920);
or U42023 (N_42023,N_41273,N_41494);
and U42024 (N_42024,N_40013,N_40911);
nor U42025 (N_42025,N_40455,N_41788);
and U42026 (N_42026,N_41844,N_41243);
or U42027 (N_42027,N_41491,N_40610);
or U42028 (N_42028,N_41853,N_41924);
or U42029 (N_42029,N_40664,N_40739);
or U42030 (N_42030,N_41019,N_40504);
nand U42031 (N_42031,N_40801,N_41267);
or U42032 (N_42032,N_41635,N_41080);
or U42033 (N_42033,N_40336,N_41960);
and U42034 (N_42034,N_41790,N_41229);
nand U42035 (N_42035,N_40368,N_40113);
or U42036 (N_42036,N_40440,N_40982);
or U42037 (N_42037,N_40663,N_40648);
or U42038 (N_42038,N_41508,N_41449);
nor U42039 (N_42039,N_41529,N_41965);
nor U42040 (N_42040,N_41624,N_41416);
nand U42041 (N_42041,N_40688,N_40490);
or U42042 (N_42042,N_41239,N_41585);
nand U42043 (N_42043,N_40571,N_40890);
and U42044 (N_42044,N_41190,N_41928);
or U42045 (N_42045,N_40088,N_41630);
nand U42046 (N_42046,N_40587,N_40027);
nor U42047 (N_42047,N_40685,N_41470);
and U42048 (N_42048,N_40471,N_41434);
and U42049 (N_42049,N_41230,N_40293);
nor U42050 (N_42050,N_40391,N_40709);
or U42051 (N_42051,N_40594,N_40119);
nand U42052 (N_42052,N_40856,N_40242);
and U42053 (N_42053,N_41672,N_41794);
nor U42054 (N_42054,N_40271,N_40860);
or U42055 (N_42055,N_40921,N_41525);
nand U42056 (N_42056,N_40120,N_40450);
nand U42057 (N_42057,N_40620,N_40466);
and U42058 (N_42058,N_41165,N_40807);
nand U42059 (N_42059,N_40183,N_41860);
and U42060 (N_42060,N_40806,N_40770);
nor U42061 (N_42061,N_40575,N_41173);
nand U42062 (N_42062,N_40515,N_40332);
nor U42063 (N_42063,N_41763,N_40977);
and U42064 (N_42064,N_40809,N_41934);
or U42065 (N_42065,N_40416,N_40393);
and U42066 (N_42066,N_40605,N_41455);
nor U42067 (N_42067,N_40396,N_40048);
or U42068 (N_42068,N_41615,N_41476);
nor U42069 (N_42069,N_41251,N_40697);
nor U42070 (N_42070,N_40202,N_40347);
nand U42071 (N_42071,N_40895,N_41791);
and U42072 (N_42072,N_41957,N_41872);
nand U42073 (N_42073,N_41256,N_40803);
and U42074 (N_42074,N_40769,N_41502);
nand U42075 (N_42075,N_41647,N_40341);
and U42076 (N_42076,N_40129,N_40392);
nor U42077 (N_42077,N_41246,N_40475);
and U42078 (N_42078,N_40681,N_41797);
xor U42079 (N_42079,N_41706,N_41424);
nor U42080 (N_42080,N_41111,N_40296);
nand U42081 (N_42081,N_41048,N_41822);
or U42082 (N_42082,N_41033,N_41687);
nand U42083 (N_42083,N_40908,N_41845);
nor U42084 (N_42084,N_41634,N_40329);
nor U42085 (N_42085,N_40597,N_41028);
nand U42086 (N_42086,N_40930,N_41834);
or U42087 (N_42087,N_41898,N_41556);
nor U42088 (N_42088,N_40224,N_40051);
nor U42089 (N_42089,N_40967,N_40899);
nor U42090 (N_42090,N_40802,N_40208);
nand U42091 (N_42091,N_40830,N_41250);
nor U42092 (N_42092,N_40657,N_41370);
and U42093 (N_42093,N_41156,N_40637);
and U42094 (N_42094,N_40602,N_40617);
nand U42095 (N_42095,N_40308,N_41127);
or U42096 (N_42096,N_41438,N_41671);
and U42097 (N_42097,N_41244,N_40756);
xor U42098 (N_42098,N_40266,N_40731);
and U42099 (N_42099,N_41920,N_41318);
and U42100 (N_42100,N_41773,N_40501);
nand U42101 (N_42101,N_40698,N_41819);
and U42102 (N_42102,N_40927,N_40355);
nand U42103 (N_42103,N_41619,N_41521);
or U42104 (N_42104,N_41102,N_41426);
or U42105 (N_42105,N_40576,N_40406);
and U42106 (N_42106,N_41691,N_40073);
nand U42107 (N_42107,N_41889,N_40211);
nor U42108 (N_42108,N_40910,N_40144);
nand U42109 (N_42109,N_41650,N_40350);
and U42110 (N_42110,N_40837,N_40087);
nor U42111 (N_42111,N_41110,N_40419);
and U42112 (N_42112,N_41558,N_40024);
nor U42113 (N_42113,N_41162,N_41519);
or U42114 (N_42114,N_40499,N_40824);
or U42115 (N_42115,N_41714,N_40264);
and U42116 (N_42116,N_41282,N_40256);
nand U42117 (N_42117,N_41407,N_40046);
nor U42118 (N_42118,N_41228,N_41317);
nor U42119 (N_42119,N_41179,N_40487);
nor U42120 (N_42120,N_41717,N_40992);
and U42121 (N_42121,N_40294,N_41437);
or U42122 (N_42122,N_40077,N_41188);
nand U42123 (N_42123,N_40993,N_41160);
nor U42124 (N_42124,N_41658,N_41660);
and U42125 (N_42125,N_41479,N_41141);
xor U42126 (N_42126,N_41832,N_40623);
nor U42127 (N_42127,N_40287,N_40639);
or U42128 (N_42128,N_40734,N_41947);
and U42129 (N_42129,N_41398,N_41961);
nand U42130 (N_42130,N_40122,N_40564);
or U42131 (N_42131,N_41200,N_40067);
or U42132 (N_42132,N_41286,N_41950);
or U42133 (N_42133,N_41118,N_40761);
nor U42134 (N_42134,N_40649,N_41214);
nand U42135 (N_42135,N_41475,N_41376);
nand U42136 (N_42136,N_40903,N_40235);
xor U42137 (N_42137,N_41021,N_40199);
and U42138 (N_42138,N_41723,N_40606);
nor U42139 (N_42139,N_41683,N_41905);
nand U42140 (N_42140,N_40622,N_40444);
nor U42141 (N_42141,N_41578,N_41331);
or U42142 (N_42142,N_41613,N_41962);
or U42143 (N_42143,N_40360,N_40197);
or U42144 (N_42144,N_41570,N_41978);
xor U42145 (N_42145,N_41579,N_41125);
and U42146 (N_42146,N_41280,N_41821);
nand U42147 (N_42147,N_40716,N_40953);
nand U42148 (N_42148,N_40083,N_40042);
or U42149 (N_42149,N_41590,N_41232);
and U42150 (N_42150,N_40542,N_41554);
nand U42151 (N_42151,N_40794,N_41722);
xnor U42152 (N_42152,N_40749,N_41595);
nand U42153 (N_42153,N_41013,N_41409);
and U42154 (N_42154,N_40409,N_40026);
nand U42155 (N_42155,N_41150,N_41851);
and U42156 (N_42156,N_40828,N_40684);
nand U42157 (N_42157,N_40165,N_40679);
nor U42158 (N_42158,N_40584,N_40395);
xor U42159 (N_42159,N_40520,N_40354);
nor U42160 (N_42160,N_40902,N_40300);
nand U42161 (N_42161,N_41296,N_40838);
nor U42162 (N_42162,N_41857,N_40214);
nor U42163 (N_42163,N_41042,N_40777);
nor U42164 (N_42164,N_41858,N_41912);
nor U42165 (N_42165,N_41353,N_41176);
nand U42166 (N_42166,N_40531,N_41472);
nand U42167 (N_42167,N_41606,N_41977);
or U42168 (N_42168,N_40634,N_40254);
and U42169 (N_42169,N_41704,N_41796);
or U42170 (N_42170,N_40527,N_40218);
or U42171 (N_42171,N_40901,N_40833);
nor U42172 (N_42172,N_40714,N_40505);
or U42173 (N_42173,N_40252,N_41825);
nor U42174 (N_42174,N_40028,N_41984);
and U42175 (N_42175,N_41864,N_40996);
or U42176 (N_42176,N_40203,N_40507);
or U42177 (N_42177,N_41698,N_40269);
and U42178 (N_42178,N_40785,N_41066);
nor U42179 (N_42179,N_41276,N_41523);
and U42180 (N_42180,N_40962,N_41378);
nor U42181 (N_42181,N_41955,N_40441);
nand U42182 (N_42182,N_40226,N_41194);
nand U42183 (N_42183,N_41838,N_40394);
nor U42184 (N_42184,N_40886,N_41443);
nand U42185 (N_42185,N_41059,N_40808);
nor U42186 (N_42186,N_40255,N_41685);
nor U42187 (N_42187,N_40317,N_40480);
and U42188 (N_42188,N_40844,N_40291);
and U42189 (N_42189,N_40160,N_40286);
nand U42190 (N_42190,N_40082,N_40889);
nor U42191 (N_42191,N_40221,N_40868);
nand U42192 (N_42192,N_41369,N_40703);
and U42193 (N_42193,N_41534,N_40772);
nor U42194 (N_42194,N_40941,N_41540);
nor U42195 (N_42195,N_41289,N_41842);
nand U42196 (N_42196,N_40687,N_40006);
nand U42197 (N_42197,N_41420,N_41245);
and U42198 (N_42198,N_40654,N_41447);
and U42199 (N_42199,N_40645,N_41573);
and U42200 (N_42200,N_40948,N_41284);
nor U42201 (N_42201,N_41622,N_41140);
nand U42202 (N_42202,N_41966,N_40096);
or U42203 (N_42203,N_40016,N_40589);
nand U42204 (N_42204,N_40245,N_41406);
and U42205 (N_42205,N_41433,N_41004);
or U42206 (N_42206,N_40385,N_41908);
nor U42207 (N_42207,N_41526,N_41795);
or U42208 (N_42208,N_40474,N_41180);
or U42209 (N_42209,N_40448,N_40279);
or U42210 (N_42210,N_40601,N_40883);
nand U42211 (N_42211,N_41929,N_41873);
nor U42212 (N_42212,N_41949,N_41053);
nor U42213 (N_42213,N_40757,N_40608);
and U42214 (N_42214,N_41549,N_41602);
and U42215 (N_42215,N_41396,N_41751);
and U42216 (N_42216,N_40829,N_41060);
and U42217 (N_42217,N_40053,N_40359);
nor U42218 (N_42218,N_40957,N_40549);
nor U42219 (N_42219,N_40164,N_40989);
and U42220 (N_42220,N_41645,N_40153);
nand U42221 (N_42221,N_40007,N_41840);
and U42222 (N_42222,N_40348,N_41597);
and U42223 (N_42223,N_41390,N_40939);
or U42224 (N_42224,N_41439,N_40260);
and U42225 (N_42225,N_40753,N_41301);
nor U42226 (N_42226,N_41446,N_40888);
or U42227 (N_42227,N_40855,N_40560);
and U42228 (N_42228,N_41738,N_41235);
nor U42229 (N_42229,N_41215,N_40012);
nand U42230 (N_42230,N_40625,N_41278);
or U42231 (N_42231,N_41395,N_41109);
nand U42232 (N_42232,N_41823,N_41361);
xnor U42233 (N_42233,N_41580,N_41678);
and U42234 (N_42234,N_40518,N_40988);
and U42235 (N_42235,N_40201,N_40880);
nand U42236 (N_42236,N_41863,N_40069);
nor U42237 (N_42237,N_40823,N_40454);
or U42238 (N_42238,N_40356,N_41514);
or U42239 (N_42239,N_41191,N_41875);
or U42240 (N_42240,N_41237,N_40653);
or U42241 (N_42241,N_41006,N_40238);
nand U42242 (N_42242,N_41781,N_40156);
nor U42243 (N_42243,N_41868,N_40632);
nand U42244 (N_42244,N_41485,N_41919);
and U42245 (N_42245,N_41720,N_40726);
and U42246 (N_42246,N_41072,N_41183);
nor U42247 (N_42247,N_41213,N_40915);
or U42248 (N_42248,N_40878,N_41681);
xor U42249 (N_42249,N_41675,N_40352);
nand U42250 (N_42250,N_41826,N_41538);
nand U42251 (N_42251,N_41414,N_40545);
or U42252 (N_42252,N_41551,N_41352);
nor U42253 (N_42253,N_41989,N_41186);
xnor U42254 (N_42254,N_40532,N_40189);
and U42255 (N_42255,N_41829,N_40010);
nor U42256 (N_42256,N_40693,N_40090);
nand U42257 (N_42257,N_40037,N_41148);
or U42258 (N_42258,N_41217,N_41777);
nor U42259 (N_42259,N_41459,N_40876);
or U42260 (N_42260,N_41766,N_40556);
nor U42261 (N_42261,N_40852,N_40751);
xnor U42262 (N_42262,N_40299,N_41575);
or U42263 (N_42263,N_40947,N_41258);
or U42264 (N_42264,N_41725,N_40276);
or U42265 (N_42265,N_40316,N_40768);
nand U42266 (N_42266,N_40267,N_40674);
and U42267 (N_42267,N_41356,N_40477);
or U42268 (N_42268,N_40437,N_40140);
and U42269 (N_42269,N_41982,N_41498);
nor U42270 (N_42270,N_40169,N_41609);
nand U42271 (N_42271,N_41227,N_41708);
nand U42272 (N_42272,N_41524,N_41705);
or U42273 (N_42273,N_41394,N_40762);
nand U42274 (N_42274,N_41218,N_40055);
nand U42275 (N_42275,N_41513,N_40666);
and U42276 (N_42276,N_40708,N_41543);
and U42277 (N_42277,N_40859,N_41097);
nor U42278 (N_42278,N_40810,N_40449);
and U42279 (N_42279,N_41931,N_41801);
and U42280 (N_42280,N_40374,N_40574);
nand U42281 (N_42281,N_41389,N_40273);
nand U42282 (N_42282,N_40017,N_40161);
nor U42283 (N_42283,N_41116,N_41147);
and U42284 (N_42284,N_40200,N_40371);
nand U42285 (N_42285,N_41495,N_40389);
nor U42286 (N_42286,N_41144,N_41882);
nand U42287 (N_42287,N_41168,N_41605);
nand U42288 (N_42288,N_40604,N_41921);
and U42289 (N_42289,N_40863,N_40538);
nor U42290 (N_42290,N_40472,N_40407);
nor U42291 (N_42291,N_40033,N_40324);
nand U42292 (N_42292,N_40585,N_41380);
nor U42293 (N_42293,N_40318,N_40537);
and U42294 (N_42294,N_41327,N_41956);
and U42295 (N_42295,N_40198,N_41695);
or U42296 (N_42296,N_41862,N_41651);
nand U42297 (N_42297,N_41780,N_41533);
nor U42298 (N_42298,N_41582,N_41288);
or U42299 (N_42299,N_41221,N_40476);
nand U42300 (N_42300,N_41264,N_41743);
and U42301 (N_42301,N_40541,N_41778);
nand U42302 (N_42302,N_40289,N_41164);
nand U42303 (N_42303,N_41262,N_41088);
nor U42304 (N_42304,N_40175,N_40463);
xor U42305 (N_42305,N_40896,N_40467);
or U42306 (N_42306,N_41739,N_41366);
or U42307 (N_42307,N_41362,N_41745);
and U42308 (N_42308,N_40712,N_41324);
nor U42309 (N_42309,N_40661,N_41926);
and U42310 (N_42310,N_41528,N_41688);
and U42311 (N_42311,N_40964,N_40038);
nor U42312 (N_42312,N_41322,N_41259);
or U42313 (N_42313,N_40904,N_41436);
and U42314 (N_42314,N_40686,N_40831);
nand U42315 (N_42315,N_40121,N_40400);
or U42316 (N_42316,N_40108,N_40008);
nand U42317 (N_42317,N_40280,N_41625);
or U42318 (N_42318,N_41640,N_40072);
and U42319 (N_42319,N_41545,N_41051);
nor U42320 (N_42320,N_41510,N_40384);
and U42321 (N_42321,N_40041,N_40555);
and U42322 (N_42322,N_40523,N_40725);
nor U42323 (N_42323,N_40702,N_41499);
nor U42324 (N_42324,N_41944,N_40966);
nor U42325 (N_42325,N_41174,N_41642);
and U42326 (N_42326,N_41910,N_40516);
or U42327 (N_42327,N_41326,N_41488);
and U42328 (N_42328,N_41656,N_41486);
and U42329 (N_42329,N_41049,N_41783);
nor U42330 (N_42330,N_40853,N_41776);
nor U42331 (N_42331,N_40729,N_40220);
or U42332 (N_42332,N_41017,N_41363);
or U42333 (N_42333,N_41098,N_41270);
or U42334 (N_42334,N_41968,N_40298);
or U42335 (N_42335,N_41303,N_40701);
nand U42336 (N_42336,N_40767,N_40334);
nand U42337 (N_42337,N_41467,N_41044);
nand U42338 (N_42338,N_41065,N_40650);
or U42339 (N_42339,N_40142,N_41112);
and U42340 (N_42340,N_40750,N_40420);
and U42341 (N_42341,N_41031,N_41025);
nor U42342 (N_42342,N_41768,N_41490);
nand U42343 (N_42343,N_41294,N_40502);
or U42344 (N_42344,N_40265,N_41121);
nand U42345 (N_42345,N_40191,N_40397);
nor U42346 (N_42346,N_41124,N_40446);
nor U42347 (N_42347,N_41274,N_41061);
nand U42348 (N_42348,N_40559,N_40680);
nand U42349 (N_42349,N_40434,N_40994);
or U42350 (N_42350,N_40022,N_41037);
nor U42351 (N_42351,N_40075,N_40614);
nand U42352 (N_42352,N_40282,N_40227);
nor U42353 (N_42353,N_40094,N_41835);
or U42354 (N_42354,N_41405,N_40942);
nor U42355 (N_42355,N_41461,N_41105);
and U42356 (N_42356,N_41948,N_40548);
or U42357 (N_42357,N_41793,N_40825);
and U42358 (N_42358,N_40095,N_41581);
or U42359 (N_42359,N_41177,N_40633);
and U42360 (N_42360,N_41342,N_41569);
and U42361 (N_42361,N_41803,N_40135);
and U42362 (N_42362,N_41292,N_41349);
and U42363 (N_42363,N_40177,N_40155);
or U42364 (N_42364,N_40402,N_41383);
and U42365 (N_42365,N_40586,N_40871);
or U42366 (N_42366,N_41209,N_41740);
nand U42367 (N_42367,N_40764,N_41680);
nand U42368 (N_42368,N_40735,N_41410);
and U42369 (N_42369,N_40862,N_41063);
xnor U42370 (N_42370,N_41727,N_41149);
or U42371 (N_42371,N_40473,N_40596);
or U42372 (N_42372,N_41030,N_41987);
nand U42373 (N_42373,N_41752,N_41530);
nand U42374 (N_42374,N_41576,N_40922);
or U42375 (N_42375,N_40178,N_40568);
and U42376 (N_42376,N_40656,N_40166);
and U42377 (N_42377,N_40070,N_41337);
or U42378 (N_42378,N_41208,N_40304);
or U42379 (N_42379,N_41813,N_41735);
nand U42380 (N_42380,N_40881,N_40566);
nand U42381 (N_42381,N_41465,N_40869);
or U42382 (N_42382,N_40743,N_41869);
nand U42383 (N_42383,N_41789,N_40035);
and U42384 (N_42384,N_41421,N_40707);
and U42385 (N_42385,N_40030,N_40344);
nor U42386 (N_42386,N_41849,N_41381);
and U42387 (N_42387,N_40133,N_40987);
and U42388 (N_42388,N_41553,N_41113);
and U42389 (N_42389,N_40700,N_40933);
nand U42390 (N_42390,N_40076,N_41430);
or U42391 (N_42391,N_40945,N_41999);
nand U42392 (N_42392,N_41784,N_41320);
nand U42393 (N_42393,N_41083,N_41856);
and U42394 (N_42394,N_41566,N_40314);
and U42395 (N_42395,N_41364,N_40333);
or U42396 (N_42396,N_41670,N_40635);
or U42397 (N_42397,N_40188,N_40430);
xor U42398 (N_42398,N_41425,N_40872);
or U42399 (N_42399,N_41253,N_40944);
and U42400 (N_42400,N_40020,N_41589);
nand U42401 (N_42401,N_40399,N_41418);
nand U42402 (N_42402,N_40938,N_41598);
or U42403 (N_42403,N_41557,N_40919);
and U42404 (N_42404,N_40553,N_40847);
nand U42405 (N_42405,N_41608,N_40353);
and U42406 (N_42406,N_41638,N_41469);
nor U42407 (N_42407,N_40268,N_41079);
or U42408 (N_42408,N_40840,N_41633);
nand U42409 (N_42409,N_41070,N_40746);
or U42410 (N_42410,N_40219,N_40074);
and U42411 (N_42411,N_41623,N_40345);
or U42412 (N_42412,N_41611,N_40858);
nand U42413 (N_42413,N_41988,N_40682);
nor U42414 (N_42414,N_40139,N_40897);
and U42415 (N_42415,N_41263,N_41428);
nand U42416 (N_42416,N_40061,N_41441);
or U42417 (N_42417,N_41041,N_41480);
xnor U42418 (N_42418,N_41010,N_40277);
or U42419 (N_42419,N_41035,N_40949);
nand U42420 (N_42420,N_41732,N_41871);
and U42421 (N_42421,N_40683,N_40064);
nor U42422 (N_42422,N_41427,N_41552);
and U42423 (N_42423,N_40438,N_41792);
and U42424 (N_42424,N_41588,N_40429);
and U42425 (N_42425,N_41101,N_41812);
and U42426 (N_42426,N_41131,N_41607);
or U42427 (N_42427,N_41592,N_41841);
nor U42428 (N_42428,N_41515,N_40503);
or U42429 (N_42429,N_41536,N_40068);
and U42430 (N_42430,N_41612,N_41744);
or U42431 (N_42431,N_40421,N_41184);
or U42432 (N_42432,N_41711,N_41087);
or U42433 (N_42433,N_41811,N_41969);
nand U42434 (N_42434,N_40425,N_40445);
and U42435 (N_42435,N_41046,N_40427);
nand U42436 (N_42436,N_41542,N_40044);
or U42437 (N_42437,N_41747,N_41073);
or U42438 (N_42438,N_40950,N_40029);
nand U42439 (N_42439,N_41541,N_41285);
and U42440 (N_42440,N_41830,N_40417);
or U42441 (N_42441,N_41600,N_40851);
or U42442 (N_42442,N_40630,N_41998);
or U42443 (N_42443,N_40752,N_41039);
nor U42444 (N_42444,N_40811,N_40592);
or U42445 (N_42445,N_40848,N_41466);
or U42446 (N_42446,N_41064,N_40544);
nand U42447 (N_42447,N_40775,N_41637);
nor U42448 (N_42448,N_40442,N_40479);
xnor U42449 (N_42449,N_40117,N_41584);
or U42450 (N_42450,N_41885,N_41120);
nor U42451 (N_42451,N_41509,N_41325);
nor U42452 (N_42452,N_41076,N_40789);
nor U42453 (N_42453,N_41730,N_41128);
and U42454 (N_42454,N_40815,N_41531);
nor U42455 (N_42455,N_41248,N_41807);
nor U42456 (N_42456,N_41701,N_40112);
or U42457 (N_42457,N_41367,N_40040);
or U42458 (N_42458,N_40103,N_40065);
xnor U42459 (N_42459,N_40985,N_40159);
and U42460 (N_42460,N_41210,N_41462);
nand U42461 (N_42461,N_41769,N_40337);
nor U42462 (N_42462,N_40742,N_41497);
nor U42463 (N_42463,N_41005,N_40447);
and U42464 (N_42464,N_41810,N_41511);
nor U42465 (N_42465,N_40894,N_40968);
nand U42466 (N_42466,N_41755,N_40511);
or U42467 (N_42467,N_41532,N_40458);
and U42468 (N_42468,N_40484,N_40489);
nor U42469 (N_42469,N_40521,N_40873);
nand U42470 (N_42470,N_41458,N_40704);
nand U42471 (N_42471,N_40711,N_40998);
or U42472 (N_42472,N_40335,N_40882);
or U42473 (N_42473,N_40141,N_41193);
nor U42474 (N_42474,N_41134,N_41315);
nand U42475 (N_42475,N_41058,N_41516);
and U42476 (N_42476,N_41505,N_40670);
or U42477 (N_42477,N_41332,N_41484);
and U42478 (N_42478,N_40491,N_41697);
and U42479 (N_42479,N_40327,N_40628);
and U42480 (N_42480,N_41496,N_41254);
nand U42481 (N_42481,N_41809,N_41391);
nor U42482 (N_42482,N_40496,N_40195);
xnor U42483 (N_42483,N_40595,N_40357);
or U42484 (N_42484,N_40673,N_40913);
and U42485 (N_42485,N_41023,N_41473);
or U42486 (N_42486,N_41306,N_41694);
or U42487 (N_42487,N_40561,N_41764);
and U42488 (N_42488,N_40054,N_40331);
or U42489 (N_42489,N_41976,N_40583);
nor U42490 (N_42490,N_40125,N_41453);
nand U42491 (N_42491,N_40926,N_41311);
xnor U42492 (N_42492,N_40916,N_41733);
and U42493 (N_42493,N_40079,N_41900);
nor U42494 (N_42494,N_40222,N_40478);
nor U42495 (N_42495,N_41266,N_40795);
nand U42496 (N_42496,N_40820,N_41452);
or U42497 (N_42497,N_41724,N_40128);
and U42498 (N_42498,N_40049,N_40627);
nand U42499 (N_42499,N_40997,N_41603);
nor U42500 (N_42500,N_41937,N_40104);
xor U42501 (N_42501,N_40781,N_41828);
xnor U42502 (N_42502,N_40805,N_41631);
and U42503 (N_42503,N_41478,N_40835);
or U42504 (N_42504,N_40558,N_41161);
and U42505 (N_42505,N_40618,N_41935);
nand U42506 (N_42506,N_41360,N_41663);
nor U42507 (N_42507,N_40870,N_41876);
or U42508 (N_42508,N_41020,N_41537);
nand U42509 (N_42509,N_40975,N_40307);
or U42510 (N_42510,N_40194,N_41056);
nor U42511 (N_42511,N_40792,N_40793);
nand U42512 (N_42512,N_41676,N_40804);
nand U42513 (N_42513,N_41236,N_40546);
and U42514 (N_42514,N_41628,N_41255);
or U42515 (N_42515,N_40658,N_40167);
nor U42516 (N_42516,N_41489,N_41699);
and U42517 (N_42517,N_40923,N_41504);
nor U42518 (N_42518,N_40508,N_41024);
or U42519 (N_42519,N_40573,N_40059);
or U42520 (N_42520,N_41448,N_40084);
and U42521 (N_42521,N_40168,N_41130);
nand U42522 (N_42522,N_40149,N_40864);
nand U42523 (N_42523,N_40891,N_41451);
or U42524 (N_42524,N_41715,N_40342);
and U42525 (N_42525,N_41758,N_41983);
nand U42526 (N_42526,N_40367,N_41074);
and U42527 (N_42527,N_40130,N_40495);
or U42528 (N_42528,N_41242,N_40972);
and U42529 (N_42529,N_41995,N_41754);
xnor U42530 (N_42530,N_40170,N_40619);
nor U42531 (N_42531,N_40744,N_41736);
nand U42532 (N_42532,N_41195,N_41973);
nand U42533 (N_42533,N_41108,N_40431);
nand U42534 (N_42534,N_41172,N_41295);
nor U42535 (N_42535,N_41852,N_40797);
and U42536 (N_42536,N_41918,N_41827);
or U42537 (N_42537,N_40816,N_40771);
or U42538 (N_42538,N_41158,N_40925);
nand U42539 (N_42539,N_40557,N_40215);
nor U42540 (N_42540,N_41562,N_40292);
nand U42541 (N_42541,N_40667,N_40278);
nand U42542 (N_42542,N_41507,N_40097);
or U42543 (N_42543,N_40295,N_41340);
and U42544 (N_42544,N_41159,N_40526);
and U42545 (N_42545,N_40710,N_40483);
nand U42546 (N_42546,N_41702,N_40624);
nand U42547 (N_42547,N_40415,N_40718);
nor U42548 (N_42548,N_40209,N_40107);
nor U42549 (N_42549,N_40014,N_41089);
or U42550 (N_42550,N_41560,N_40313);
and U42551 (N_42551,N_41655,N_40572);
nor U42552 (N_42552,N_41474,N_40671);
nand U42553 (N_42553,N_41942,N_40469);
or U42554 (N_42554,N_40193,N_40723);
nor U42555 (N_42555,N_41879,N_40270);
nor U42556 (N_42556,N_41287,N_40403);
nor U42557 (N_42557,N_40646,N_40983);
nand U42558 (N_42558,N_41716,N_41224);
and U42559 (N_42559,N_41175,N_40488);
and U42560 (N_42560,N_40323,N_41431);
and U42561 (N_42561,N_40905,N_41312);
or U42562 (N_42562,N_40285,N_41710);
or U42563 (N_42563,N_41954,N_41219);
or U42564 (N_42564,N_40970,N_40206);
and U42565 (N_42565,N_41881,N_40439);
nor U42566 (N_42566,N_41482,N_40593);
and U42567 (N_42567,N_41707,N_40050);
and U42568 (N_42568,N_40379,N_41100);
or U42569 (N_42569,N_41341,N_41867);
nand U42570 (N_42570,N_41335,N_40290);
nor U42571 (N_42571,N_40765,N_41036);
or U42572 (N_42572,N_41742,N_41038);
nor U42573 (N_42573,N_41913,N_40677);
or U42574 (N_42574,N_41659,N_41045);
or U42575 (N_42575,N_40563,N_41114);
nor U42576 (N_42576,N_40364,N_40728);
and U42577 (N_42577,N_41762,N_41043);
and U42578 (N_42578,N_41052,N_41212);
nor U42579 (N_42579,N_41729,N_40283);
nor U42580 (N_42580,N_40060,N_41915);
or U42581 (N_42581,N_40813,N_41016);
nor U42582 (N_42582,N_41572,N_41146);
and U42583 (N_42583,N_41069,N_40115);
and U42584 (N_42584,N_40123,N_40387);
or U42585 (N_42585,N_41231,N_40696);
nand U42586 (N_42586,N_41385,N_41196);
nor U42587 (N_42587,N_40233,N_41365);
and U42588 (N_42588,N_41972,N_41855);
nand U42589 (N_42589,N_41774,N_40730);
nor U42590 (N_42590,N_40554,N_41782);
nand U42591 (N_42591,N_41154,N_40748);
nor U42592 (N_42592,N_40127,N_41805);
and U42593 (N_42593,N_40281,N_40867);
or U42594 (N_42594,N_41567,N_40253);
and U42595 (N_42595,N_40110,N_40971);
and U42596 (N_42596,N_41806,N_41649);
or U42597 (N_42597,N_40580,N_40570);
and U42598 (N_42598,N_40132,N_40216);
nor U42599 (N_42599,N_40783,N_41899);
and U42600 (N_42600,N_41138,N_40796);
nand U42601 (N_42601,N_40101,N_40309);
or U42602 (N_42602,N_41085,N_41343);
and U42603 (N_42603,N_41233,N_40665);
and U42604 (N_42604,N_41119,N_40343);
nand U42605 (N_42605,N_40741,N_40358);
or U42606 (N_42606,N_40984,N_41297);
nand U42607 (N_42607,N_40611,N_40152);
nor U42608 (N_42608,N_41644,N_41464);
or U42609 (N_42609,N_41178,N_40043);
xnor U42610 (N_42610,N_40080,N_41506);
nor U42611 (N_42611,N_40760,N_40321);
nand U42612 (N_42612,N_41170,N_41071);
and U42613 (N_42613,N_40958,N_40588);
and U42614 (N_42614,N_40917,N_41351);
and U42615 (N_42615,N_40914,N_41413);
nor U42616 (N_42616,N_40305,N_41861);
and U42617 (N_42617,N_41963,N_40443);
nor U42618 (N_42618,N_41082,N_41887);
nor U42619 (N_42619,N_40362,N_41316);
and U42620 (N_42620,N_40500,N_40845);
nor U42621 (N_42621,N_41571,N_41345);
nand U42622 (N_42622,N_40453,N_40414);
xor U42623 (N_42623,N_40540,N_41964);
or U42624 (N_42624,N_41002,N_40302);
nor U42625 (N_42625,N_41620,N_40577);
nand U42626 (N_42626,N_40591,N_40699);
nand U42627 (N_42627,N_40861,N_40773);
nor U42628 (N_42628,N_40212,N_40713);
and U42629 (N_42629,N_41143,N_40247);
or U42630 (N_42630,N_40363,N_40229);
nand U42631 (N_42631,N_40147,N_41990);
and U42632 (N_42632,N_40369,N_41939);
or U42633 (N_42633,N_41895,N_41477);
nand U42634 (N_42634,N_41388,N_40780);
nand U42635 (N_42635,N_40724,N_41000);
nor U42636 (N_42636,N_40325,N_41800);
nor U42637 (N_42637,N_40401,N_41372);
and U42638 (N_42638,N_41890,N_40695);
nand U42639 (N_42639,N_40924,N_41512);
and U42640 (N_42640,N_40404,N_41155);
and U42641 (N_42641,N_40432,N_41012);
or U42642 (N_42642,N_40995,N_40579);
nor U42643 (N_42643,N_41818,N_41096);
and U42644 (N_42644,N_40642,N_40733);
or U42645 (N_42645,N_40423,N_40912);
nor U42646 (N_42646,N_41741,N_41137);
nand U42647 (N_42647,N_40740,N_40411);
and U42648 (N_42648,N_41587,N_41308);
nor U42649 (N_42649,N_41350,N_40056);
nor U42650 (N_42650,N_40715,N_41014);
nor U42651 (N_42651,N_40536,N_40482);
nand U42652 (N_42652,N_40692,N_40582);
nand U42653 (N_42653,N_40361,N_41403);
and U42654 (N_42654,N_40539,N_41726);
nor U42655 (N_42655,N_40150,N_40599);
and U42656 (N_42656,N_40138,N_41077);
and U42657 (N_42657,N_41015,N_41081);
or U42658 (N_42658,N_40187,N_40236);
nand U42659 (N_42659,N_41054,N_41896);
or U42660 (N_42660,N_41877,N_40929);
and U42661 (N_42661,N_41518,N_40529);
nand U42662 (N_42662,N_40005,N_40424);
or U42663 (N_42663,N_40965,N_40755);
and U42664 (N_42664,N_40973,N_40099);
or U42665 (N_42665,N_40301,N_41249);
and U42666 (N_42666,N_40412,N_41432);
nand U42667 (N_42667,N_41222,N_41375);
and U42668 (N_42668,N_40143,N_41652);
nand U42669 (N_42669,N_41003,N_41456);
nor U42670 (N_42670,N_41055,N_41357);
nand U42671 (N_42671,N_41206,N_41445);
nand U42672 (N_42672,N_40946,N_40659);
and U42673 (N_42673,N_40481,N_40257);
nor U42674 (N_42674,N_40509,N_41936);
or U42675 (N_42675,N_40799,N_40745);
and U42676 (N_42676,N_41415,N_40102);
nand U42677 (N_42677,N_41185,N_40310);
nand U42678 (N_42678,N_40550,N_41152);
or U42679 (N_42679,N_40464,N_41641);
nand U42680 (N_42680,N_40525,N_41689);
nand U42681 (N_42681,N_40180,N_40205);
and U42682 (N_42682,N_41265,N_41904);
or U42683 (N_42683,N_40320,N_41481);
nand U42684 (N_42684,N_40937,N_40940);
nand U42685 (N_42685,N_41336,N_40990);
nor U42686 (N_42686,N_41922,N_40217);
xor U42687 (N_42687,N_41182,N_41892);
nand U42688 (N_42688,N_41673,N_41397);
nor U42689 (N_42689,N_41814,N_40907);
or U42690 (N_42690,N_40849,N_40720);
and U42691 (N_42691,N_40514,N_41086);
nand U42692 (N_42692,N_41009,N_41298);
nor U42693 (N_42693,N_41750,N_40565);
nand U42694 (N_42694,N_40935,N_40002);
and U42695 (N_42695,N_40651,N_40190);
and U42696 (N_42696,N_41423,N_41392);
or U42697 (N_42697,N_40631,N_40786);
nand U42698 (N_42698,N_40004,N_41953);
nor U42699 (N_42699,N_40727,N_40690);
or U42700 (N_42700,N_41123,N_41268);
and U42701 (N_42701,N_41787,N_41559);
or U42702 (N_42702,N_40754,N_41824);
nor U42703 (N_42703,N_40737,N_41914);
and U42704 (N_42704,N_41029,N_40451);
and U42705 (N_42705,N_41271,N_41493);
nand U42706 (N_42706,N_41040,N_40003);
and U42707 (N_42707,N_41047,N_41692);
or U42708 (N_42708,N_41535,N_41328);
and U42709 (N_42709,N_41772,N_41211);
nor U42710 (N_42710,N_41785,N_41330);
or U42711 (N_42711,N_40241,N_41958);
or U42712 (N_42712,N_40086,N_40638);
and U42713 (N_42713,N_40275,N_40250);
or U42714 (N_42714,N_41348,N_41546);
nand U42715 (N_42715,N_40875,N_41260);
or U42716 (N_42716,N_40315,N_41997);
nand U42717 (N_42717,N_41906,N_41226);
nor U42718 (N_42718,N_41804,N_40081);
or U42719 (N_42719,N_41501,N_41358);
and U42720 (N_42720,N_40390,N_40413);
or U42721 (N_42721,N_40262,N_40388);
nand U42722 (N_42722,N_41132,N_41181);
and U42723 (N_42723,N_41586,N_41075);
and U42724 (N_42724,N_41404,N_40052);
nand U42725 (N_42725,N_40936,N_41865);
nand U42726 (N_42726,N_40928,N_41563);
nand U42727 (N_42727,N_41974,N_40021);
or U42728 (N_42728,N_41402,N_41354);
nand U42729 (N_42729,N_40339,N_41677);
or U42730 (N_42730,N_41674,N_40662);
nand U42731 (N_42731,N_41664,N_41281);
and U42732 (N_42732,N_40846,N_41247);
and U42733 (N_42733,N_40109,N_41057);
nor U42734 (N_42734,N_40234,N_40498);
nand U42735 (N_42735,N_41886,N_41419);
or U42736 (N_42736,N_40185,N_41943);
nand U42737 (N_42737,N_41684,N_40600);
nand U42738 (N_42738,N_41522,N_40078);
nand U42739 (N_42739,N_40969,N_40636);
nand U42740 (N_42740,N_41980,N_41202);
and U42741 (N_42741,N_40534,N_41666);
nand U42742 (N_42742,N_41848,N_41737);
and U42743 (N_42743,N_40613,N_41959);
nand U42744 (N_42744,N_41709,N_41564);
nand U42745 (N_42745,N_40581,N_41690);
and U42746 (N_42746,N_41187,N_40732);
or U42747 (N_42747,N_41749,N_41199);
nand U42748 (N_42748,N_41334,N_40819);
nor U42749 (N_42749,N_40787,N_40812);
nand U42750 (N_42750,N_40426,N_41027);
or U42751 (N_42751,N_41721,N_40372);
nand U42752 (N_42752,N_40834,N_40089);
and U42753 (N_42753,N_40603,N_41679);
or U42754 (N_42754,N_41257,N_40782);
and U42755 (N_42755,N_41594,N_41201);
nand U42756 (N_42756,N_40898,N_40952);
nand U42757 (N_42757,N_41756,N_41463);
or U42758 (N_42758,N_41846,N_41269);
nor U42759 (N_42759,N_41574,N_40018);
or U42760 (N_42760,N_40513,N_41204);
nor U42761 (N_42761,N_41377,N_40163);
and U42762 (N_42762,N_40758,N_41878);
nor U42763 (N_42763,N_40675,N_40874);
and U42764 (N_42764,N_41517,N_41067);
and U42765 (N_42765,N_40836,N_41192);
nor U42766 (N_42766,N_41850,N_40246);
or U42767 (N_42767,N_41893,N_41991);
or U42768 (N_42768,N_41932,N_40763);
nand U42769 (N_42769,N_40248,N_41593);
and U42770 (N_42770,N_40906,N_41151);
nand U42771 (N_42771,N_41338,N_40615);
and U42772 (N_42772,N_41565,N_40934);
nor U42773 (N_42773,N_41610,N_41547);
nand U42774 (N_42774,N_41591,N_40457);
nor U42775 (N_42775,N_41731,N_41761);
nor U42776 (N_42776,N_41996,N_40322);
and U42777 (N_42777,N_41145,N_41843);
xor U42778 (N_42778,N_40232,N_41032);
and U42779 (N_42779,N_41500,N_40225);
or U42780 (N_42780,N_40460,N_41417);
nor U42781 (N_42781,N_40100,N_41836);
and U42782 (N_42782,N_40668,N_41621);
and U42783 (N_42783,N_40181,N_40598);
nor U42784 (N_42784,N_41313,N_41412);
or U42785 (N_42785,N_41169,N_41816);
or U42786 (N_42786,N_40173,N_41614);
nor U42787 (N_42787,N_40034,N_40986);
or U42788 (N_42788,N_40691,N_40174);
or U42789 (N_42789,N_40778,N_40485);
xnor U42790 (N_42790,N_41090,N_40817);
or U42791 (N_42791,N_40981,N_40114);
and U42792 (N_42792,N_41007,N_41355);
nor U42793 (N_42793,N_40519,N_40943);
nor U42794 (N_42794,N_41368,N_41310);
nand U42795 (N_42795,N_41632,N_41917);
and U42796 (N_42796,N_40366,N_40893);
xnor U42797 (N_42797,N_40184,N_41440);
nand U42798 (N_42798,N_41909,N_41577);
nor U42799 (N_42799,N_41095,N_41550);
nor U42800 (N_42800,N_41234,N_40376);
or U42801 (N_42801,N_40951,N_41760);
nor U42802 (N_42802,N_40066,N_41775);
and U42803 (N_42803,N_40288,N_40462);
or U42804 (N_42804,N_40784,N_41442);
nand U42805 (N_42805,N_40822,N_40641);
nand U42806 (N_42806,N_41117,N_40517);
nand U42807 (N_42807,N_40131,N_41639);
and U42808 (N_42808,N_41520,N_41457);
xnor U42809 (N_42809,N_40826,N_41084);
nand U42810 (N_42810,N_41106,N_40841);
nor U42811 (N_42811,N_41261,N_41902);
and U42812 (N_42812,N_40210,N_41967);
and U42813 (N_42813,N_40909,N_40621);
and U42814 (N_42814,N_40272,N_40106);
or U42815 (N_42815,N_40747,N_40148);
and U42816 (N_42816,N_41333,N_41718);
or U42817 (N_42817,N_41314,N_41616);
nand U42818 (N_42818,N_41669,N_41062);
and U42819 (N_42819,N_40857,N_40118);
nor U42820 (N_42820,N_40047,N_40230);
xor U42821 (N_42821,N_41429,N_40694);
or U42822 (N_42822,N_41945,N_41561);
and U42823 (N_42823,N_40791,N_41435);
and U42824 (N_42824,N_41993,N_40497);
or U42825 (N_42825,N_40814,N_40116);
or U42826 (N_42826,N_41985,N_41309);
or U42827 (N_42827,N_40980,N_40223);
and U42828 (N_42828,N_41883,N_41142);
or U42829 (N_42829,N_41275,N_40373);
or U42830 (N_42830,N_40146,N_40955);
or U42831 (N_42831,N_40091,N_41941);
nor U42832 (N_42832,N_41207,N_41411);
and U42833 (N_42833,N_40182,N_41596);
xor U42834 (N_42834,N_40383,N_41837);
nor U42835 (N_42835,N_41304,N_41107);
nand U42836 (N_42836,N_40678,N_40569);
nand U42837 (N_42837,N_41728,N_40134);
or U42838 (N_42838,N_40533,N_40689);
nor U42839 (N_42839,N_41880,N_40025);
nor U42840 (N_42840,N_40062,N_41759);
or U42841 (N_42841,N_41279,N_40092);
nand U42842 (N_42842,N_40722,N_40456);
or U42843 (N_42843,N_41854,N_41093);
xnor U42844 (N_42844,N_41382,N_40669);
nor U42845 (N_42845,N_40779,N_40976);
and U42846 (N_42846,N_40319,N_40126);
nand U42847 (N_42847,N_40932,N_41346);
or U42848 (N_42848,N_41129,N_40071);
nand U42849 (N_42849,N_40239,N_41099);
nor U42850 (N_42850,N_40524,N_40213);
or U42851 (N_42851,N_40956,N_40111);
and U42852 (N_42852,N_41648,N_41050);
nand U42853 (N_42853,N_40884,N_40058);
nand U42854 (N_42854,N_40408,N_40326);
xor U42855 (N_42855,N_41994,N_40045);
nor U42856 (N_42856,N_40151,N_40854);
and U42857 (N_42857,N_40879,N_40382);
nand U42858 (N_42858,N_41713,N_41548);
or U42859 (N_42859,N_40643,N_41373);
or U42860 (N_42860,N_41339,N_40418);
nor U42861 (N_42861,N_41167,N_40240);
and U42862 (N_42862,N_40465,N_40839);
or U42863 (N_42863,N_40528,N_41277);
and U42864 (N_42864,N_40386,N_41115);
nor U42865 (N_42865,N_41753,N_40179);
and U42866 (N_42866,N_41839,N_40717);
nand U42867 (N_42867,N_41307,N_41492);
nand U42868 (N_42868,N_41643,N_41894);
nand U42869 (N_42869,N_41815,N_40176);
and U42870 (N_42870,N_40249,N_40821);
and U42871 (N_42871,N_40818,N_40676);
and U42872 (N_42872,N_41636,N_41408);
and U42873 (N_42873,N_41703,N_40800);
nor U42874 (N_42874,N_40145,N_41668);
nor U42875 (N_42875,N_41952,N_40991);
or U42876 (N_42876,N_40032,N_40459);
nor U42877 (N_42877,N_40866,N_41847);
and U42878 (N_42878,N_41527,N_40931);
nor U42879 (N_42879,N_40380,N_41746);
nand U42880 (N_42880,N_40766,N_41903);
nand U42881 (N_42881,N_41471,N_40340);
or U42882 (N_42882,N_41163,N_40655);
and U42883 (N_42883,N_41779,N_41305);
nor U42884 (N_42884,N_41661,N_41319);
or U42885 (N_42885,N_41820,N_41011);
or U42886 (N_42886,N_41925,N_41757);
nand U42887 (N_42887,N_40297,N_41981);
nor U42888 (N_42888,N_41700,N_41986);
or U42889 (N_42889,N_41646,N_41133);
nor U42890 (N_42890,N_41933,N_41657);
nor U42891 (N_42891,N_40085,N_41629);
nor U42892 (N_42892,N_41916,N_41379);
and U42893 (N_42893,N_41359,N_41302);
and U42894 (N_42894,N_41765,N_41220);
or U42895 (N_42895,N_40258,N_40616);
nor U42896 (N_42896,N_40057,N_41874);
or U42897 (N_42897,N_41135,N_40790);
nor U42898 (N_42898,N_41483,N_41770);
nand U42899 (N_42899,N_40721,N_40137);
or U42900 (N_42900,N_41393,N_40705);
nor U42901 (N_42901,N_40961,N_40506);
nand U42902 (N_42902,N_41544,N_41946);
nand U42903 (N_42903,N_41139,N_40377);
and U42904 (N_42904,N_40918,N_40422);
nor U42905 (N_42905,N_41104,N_40900);
nand U42906 (N_42906,N_41216,N_40552);
or U42907 (N_42907,N_40311,N_41682);
nand U42908 (N_42908,N_40031,N_40842);
and U42909 (N_42909,N_40312,N_40435);
and U42910 (N_42910,N_40736,N_41290);
and U42911 (N_42911,N_40171,N_40978);
and U42912 (N_42912,N_40378,N_40640);
nor U42913 (N_42913,N_41712,N_41454);
and U42914 (N_42914,N_40492,N_41808);
or U42915 (N_42915,N_40346,N_40672);
xor U42916 (N_42916,N_41951,N_40979);
nand U42917 (N_42917,N_41252,N_40486);
nor U42918 (N_42918,N_41599,N_40237);
nor U42919 (N_42919,N_41938,N_40192);
or U42920 (N_42920,N_40157,N_40162);
nor U42921 (N_42921,N_40172,N_41831);
nand U42922 (N_42922,N_41153,N_40009);
nand U42923 (N_42923,N_40629,N_41626);
and U42924 (N_42924,N_41891,N_41870);
and U42925 (N_42925,N_40000,N_41401);
nor U42926 (N_42926,N_40607,N_41225);
nand U42927 (N_42927,N_40551,N_41604);
nand U42928 (N_42928,N_41930,N_40644);
and U42929 (N_42929,N_41907,N_40330);
nor U42930 (N_42930,N_41817,N_41238);
and U42931 (N_42931,N_41197,N_41601);
or U42932 (N_42932,N_41979,N_41654);
and U42933 (N_42933,N_40158,N_40274);
or U42934 (N_42934,N_41653,N_40349);
and U42935 (N_42935,N_41323,N_40510);
nor U42936 (N_42936,N_41901,N_40535);
nand U42937 (N_42937,N_40381,N_41911);
nand U42938 (N_42938,N_41444,N_41734);
and U42939 (N_42939,N_40512,N_40892);
nor U42940 (N_42940,N_41568,N_40370);
or U42941 (N_42941,N_40284,N_40470);
and U42942 (N_42942,N_40494,N_40428);
or U42943 (N_42943,N_40098,N_40468);
and U42944 (N_42944,N_40543,N_41665);
nor U42945 (N_42945,N_40063,N_40530);
nor U42946 (N_42946,N_41189,N_40578);
nor U42947 (N_42947,N_41272,N_40405);
nor U42948 (N_42948,N_41300,N_40036);
xnor U42949 (N_42949,N_40433,N_41001);
nand U42950 (N_42950,N_40590,N_40410);
or U42951 (N_42951,N_40196,N_40251);
or U42952 (N_42952,N_40626,N_41888);
or U42953 (N_42953,N_40850,N_41026);
nand U42954 (N_42954,N_40436,N_41136);
and U42955 (N_42955,N_41693,N_40798);
nand U42956 (N_42956,N_40093,N_41223);
nand U42957 (N_42957,N_40776,N_40877);
or U42958 (N_42958,N_41422,N_41198);
and U42959 (N_42959,N_41970,N_40493);
nand U42960 (N_42960,N_40023,N_40204);
xor U42961 (N_42961,N_41126,N_41291);
nand U42962 (N_42962,N_41487,N_41166);
nand U42963 (N_42963,N_41321,N_40303);
or U42964 (N_42964,N_40759,N_41384);
nor U42965 (N_42965,N_41241,N_40974);
nand U42966 (N_42966,N_41374,N_41347);
or U42967 (N_42967,N_41686,N_40011);
nand U42968 (N_42968,N_40827,N_41940);
nand U42969 (N_42969,N_41078,N_40612);
nand U42970 (N_42970,N_41923,N_40228);
and U42971 (N_42971,N_41662,N_41386);
nand U42972 (N_42972,N_40259,N_41329);
and U42973 (N_42973,N_40243,N_41555);
nor U42974 (N_42974,N_40039,N_40954);
nand U42975 (N_42975,N_41866,N_40959);
nor U42976 (N_42976,N_41627,N_41748);
nand U42977 (N_42977,N_41344,N_40885);
and U42978 (N_42978,N_40706,N_40375);
nor U42979 (N_42979,N_40231,N_41617);
and U42980 (N_42980,N_40960,N_41205);
and U42981 (N_42981,N_41034,N_40263);
nand U42982 (N_42982,N_40865,N_41696);
xnor U42983 (N_42983,N_41927,N_40660);
or U42984 (N_42984,N_41992,N_41468);
and U42985 (N_42985,N_41122,N_40338);
and U42986 (N_42986,N_41786,N_41503);
and U42987 (N_42987,N_40832,N_41833);
or U42988 (N_42988,N_41299,N_40306);
or U42989 (N_42989,N_41884,N_40999);
or U42990 (N_42990,N_41091,N_41799);
and U42991 (N_42991,N_41859,N_40774);
or U42992 (N_42992,N_41667,N_40562);
nor U42993 (N_42993,N_40719,N_41068);
or U42994 (N_42994,N_40105,N_41460);
nor U42995 (N_42995,N_41283,N_41171);
or U42996 (N_42996,N_41767,N_40019);
and U42997 (N_42997,N_40738,N_40963);
and U42998 (N_42998,N_41798,N_41387);
xor U42999 (N_42999,N_40547,N_41018);
nand U43000 (N_43000,N_41564,N_40179);
or U43001 (N_43001,N_40346,N_40929);
and U43002 (N_43002,N_41688,N_41258);
nand U43003 (N_43003,N_40033,N_41790);
or U43004 (N_43004,N_40897,N_41879);
nor U43005 (N_43005,N_41832,N_41550);
and U43006 (N_43006,N_40186,N_41510);
nor U43007 (N_43007,N_40231,N_41863);
and U43008 (N_43008,N_40856,N_40660);
nor U43009 (N_43009,N_40595,N_41112);
nand U43010 (N_43010,N_40052,N_40866);
nand U43011 (N_43011,N_41313,N_40377);
and U43012 (N_43012,N_41009,N_41197);
nand U43013 (N_43013,N_41813,N_40472);
nor U43014 (N_43014,N_41818,N_40264);
nand U43015 (N_43015,N_40608,N_41367);
or U43016 (N_43016,N_41305,N_40401);
and U43017 (N_43017,N_40439,N_40732);
nor U43018 (N_43018,N_40356,N_40038);
and U43019 (N_43019,N_41398,N_41675);
nand U43020 (N_43020,N_40931,N_41584);
and U43021 (N_43021,N_41832,N_40316);
nor U43022 (N_43022,N_41338,N_40107);
and U43023 (N_43023,N_41416,N_40944);
nand U43024 (N_43024,N_41943,N_40168);
nand U43025 (N_43025,N_41414,N_40217);
nor U43026 (N_43026,N_41327,N_40401);
or U43027 (N_43027,N_40095,N_41516);
and U43028 (N_43028,N_40437,N_40105);
xor U43029 (N_43029,N_41142,N_41014);
nand U43030 (N_43030,N_41831,N_41696);
nor U43031 (N_43031,N_41784,N_40523);
nor U43032 (N_43032,N_40161,N_41613);
nor U43033 (N_43033,N_40310,N_41319);
and U43034 (N_43034,N_40515,N_40645);
and U43035 (N_43035,N_40384,N_40517);
nand U43036 (N_43036,N_41320,N_40307);
and U43037 (N_43037,N_41996,N_41463);
nor U43038 (N_43038,N_41714,N_40031);
or U43039 (N_43039,N_41346,N_41832);
and U43040 (N_43040,N_41884,N_41345);
nand U43041 (N_43041,N_40292,N_40068);
nor U43042 (N_43042,N_40983,N_40065);
or U43043 (N_43043,N_40631,N_41791);
or U43044 (N_43044,N_41670,N_40352);
and U43045 (N_43045,N_40872,N_40887);
or U43046 (N_43046,N_40178,N_41893);
xor U43047 (N_43047,N_40405,N_41176);
or U43048 (N_43048,N_41956,N_40438);
nor U43049 (N_43049,N_40993,N_41768);
nor U43050 (N_43050,N_40856,N_40068);
xor U43051 (N_43051,N_41499,N_40550);
and U43052 (N_43052,N_40894,N_40298);
nand U43053 (N_43053,N_41498,N_40700);
nand U43054 (N_43054,N_41602,N_40390);
nand U43055 (N_43055,N_41633,N_41468);
or U43056 (N_43056,N_40735,N_40478);
or U43057 (N_43057,N_40493,N_41363);
or U43058 (N_43058,N_41715,N_40334);
or U43059 (N_43059,N_41559,N_41337);
nor U43060 (N_43060,N_40203,N_41308);
nor U43061 (N_43061,N_40786,N_41323);
nor U43062 (N_43062,N_41697,N_40367);
nand U43063 (N_43063,N_40445,N_40132);
or U43064 (N_43064,N_41889,N_40386);
nor U43065 (N_43065,N_41123,N_40537);
or U43066 (N_43066,N_41793,N_40678);
xnor U43067 (N_43067,N_41035,N_40184);
and U43068 (N_43068,N_40730,N_41276);
nor U43069 (N_43069,N_41805,N_40220);
xnor U43070 (N_43070,N_41944,N_40782);
and U43071 (N_43071,N_40654,N_41100);
nand U43072 (N_43072,N_40056,N_40271);
nor U43073 (N_43073,N_41494,N_40745);
nor U43074 (N_43074,N_41698,N_41807);
and U43075 (N_43075,N_40062,N_41737);
nor U43076 (N_43076,N_40927,N_41464);
and U43077 (N_43077,N_41171,N_41230);
nor U43078 (N_43078,N_40416,N_41578);
and U43079 (N_43079,N_40503,N_40550);
nand U43080 (N_43080,N_40835,N_41318);
or U43081 (N_43081,N_40879,N_41697);
nor U43082 (N_43082,N_40844,N_40300);
nor U43083 (N_43083,N_41855,N_40099);
nor U43084 (N_43084,N_41352,N_40717);
and U43085 (N_43085,N_40360,N_41628);
nand U43086 (N_43086,N_41469,N_41075);
nand U43087 (N_43087,N_40392,N_41744);
or U43088 (N_43088,N_41085,N_40580);
nor U43089 (N_43089,N_40364,N_40422);
nor U43090 (N_43090,N_41374,N_41128);
or U43091 (N_43091,N_40273,N_40167);
or U43092 (N_43092,N_40054,N_40951);
nor U43093 (N_43093,N_41968,N_41510);
or U43094 (N_43094,N_41951,N_40268);
and U43095 (N_43095,N_40646,N_41855);
nor U43096 (N_43096,N_40975,N_40225);
nand U43097 (N_43097,N_40870,N_41616);
nor U43098 (N_43098,N_41335,N_41385);
nand U43099 (N_43099,N_41371,N_41862);
and U43100 (N_43100,N_41470,N_40400);
and U43101 (N_43101,N_40450,N_41087);
and U43102 (N_43102,N_40765,N_40839);
xor U43103 (N_43103,N_40591,N_41460);
nor U43104 (N_43104,N_40670,N_40196);
and U43105 (N_43105,N_41500,N_41574);
nor U43106 (N_43106,N_41591,N_40524);
nand U43107 (N_43107,N_40236,N_40479);
nand U43108 (N_43108,N_41042,N_41607);
or U43109 (N_43109,N_41591,N_40316);
and U43110 (N_43110,N_41532,N_40927);
xor U43111 (N_43111,N_40899,N_41106);
nor U43112 (N_43112,N_41046,N_40193);
or U43113 (N_43113,N_41233,N_40423);
nand U43114 (N_43114,N_40708,N_41903);
or U43115 (N_43115,N_40035,N_40236);
or U43116 (N_43116,N_41734,N_41000);
nor U43117 (N_43117,N_41104,N_40736);
nor U43118 (N_43118,N_40929,N_41811);
nor U43119 (N_43119,N_41180,N_41235);
and U43120 (N_43120,N_40244,N_41807);
nand U43121 (N_43121,N_40163,N_40273);
or U43122 (N_43122,N_40622,N_41019);
nand U43123 (N_43123,N_40664,N_40681);
and U43124 (N_43124,N_40914,N_41802);
nand U43125 (N_43125,N_41468,N_40652);
or U43126 (N_43126,N_40412,N_40181);
nor U43127 (N_43127,N_40801,N_41494);
nor U43128 (N_43128,N_40411,N_41546);
nand U43129 (N_43129,N_40296,N_40415);
and U43130 (N_43130,N_41164,N_41496);
or U43131 (N_43131,N_40935,N_40592);
nor U43132 (N_43132,N_40244,N_40488);
or U43133 (N_43133,N_40520,N_40444);
and U43134 (N_43134,N_41811,N_40420);
and U43135 (N_43135,N_41884,N_40301);
nand U43136 (N_43136,N_41548,N_40595);
nand U43137 (N_43137,N_40803,N_41787);
nor U43138 (N_43138,N_41891,N_41094);
nor U43139 (N_43139,N_41279,N_41016);
nand U43140 (N_43140,N_41364,N_40998);
or U43141 (N_43141,N_41623,N_41166);
and U43142 (N_43142,N_41141,N_40388);
or U43143 (N_43143,N_40218,N_40576);
nand U43144 (N_43144,N_40604,N_41129);
xnor U43145 (N_43145,N_40433,N_41021);
or U43146 (N_43146,N_40870,N_41533);
nor U43147 (N_43147,N_40785,N_41937);
and U43148 (N_43148,N_40698,N_41414);
nor U43149 (N_43149,N_40840,N_41351);
and U43150 (N_43150,N_40904,N_41625);
nand U43151 (N_43151,N_41649,N_41194);
nor U43152 (N_43152,N_40254,N_40632);
or U43153 (N_43153,N_41757,N_40913);
and U43154 (N_43154,N_40766,N_40345);
nand U43155 (N_43155,N_40294,N_40961);
nand U43156 (N_43156,N_41485,N_40343);
nor U43157 (N_43157,N_40049,N_40892);
and U43158 (N_43158,N_40951,N_40813);
or U43159 (N_43159,N_40093,N_40816);
xnor U43160 (N_43160,N_41553,N_41416);
or U43161 (N_43161,N_41160,N_40386);
nand U43162 (N_43162,N_41777,N_41710);
nor U43163 (N_43163,N_41053,N_40084);
or U43164 (N_43164,N_41365,N_40574);
or U43165 (N_43165,N_41293,N_41610);
nand U43166 (N_43166,N_40829,N_41176);
nand U43167 (N_43167,N_40928,N_40190);
nor U43168 (N_43168,N_40762,N_41110);
nor U43169 (N_43169,N_41808,N_40311);
nor U43170 (N_43170,N_41063,N_41512);
nand U43171 (N_43171,N_40956,N_41165);
nor U43172 (N_43172,N_40246,N_41484);
nand U43173 (N_43173,N_40355,N_41390);
or U43174 (N_43174,N_41868,N_40110);
or U43175 (N_43175,N_40211,N_41618);
nand U43176 (N_43176,N_41320,N_41045);
and U43177 (N_43177,N_40933,N_40037);
nor U43178 (N_43178,N_40078,N_40259);
nor U43179 (N_43179,N_41827,N_41505);
or U43180 (N_43180,N_41833,N_40157);
nor U43181 (N_43181,N_41204,N_40407);
and U43182 (N_43182,N_41770,N_41868);
or U43183 (N_43183,N_41086,N_41114);
nor U43184 (N_43184,N_41172,N_40857);
and U43185 (N_43185,N_41162,N_40461);
or U43186 (N_43186,N_40247,N_40905);
or U43187 (N_43187,N_41698,N_41542);
or U43188 (N_43188,N_41197,N_40737);
and U43189 (N_43189,N_41213,N_41480);
nor U43190 (N_43190,N_40158,N_40199);
or U43191 (N_43191,N_41008,N_40304);
nand U43192 (N_43192,N_41653,N_41284);
and U43193 (N_43193,N_40933,N_40503);
and U43194 (N_43194,N_41352,N_41800);
nand U43195 (N_43195,N_41102,N_40374);
and U43196 (N_43196,N_40830,N_41388);
or U43197 (N_43197,N_40685,N_40878);
nand U43198 (N_43198,N_40556,N_41030);
or U43199 (N_43199,N_40810,N_40251);
nor U43200 (N_43200,N_40903,N_41266);
nand U43201 (N_43201,N_41111,N_41060);
or U43202 (N_43202,N_40291,N_40659);
nor U43203 (N_43203,N_40421,N_40870);
nand U43204 (N_43204,N_41305,N_40099);
nand U43205 (N_43205,N_41961,N_40327);
and U43206 (N_43206,N_40681,N_41510);
nand U43207 (N_43207,N_40964,N_40503);
or U43208 (N_43208,N_41097,N_40748);
xnor U43209 (N_43209,N_41060,N_40879);
nand U43210 (N_43210,N_41653,N_41805);
or U43211 (N_43211,N_41337,N_41845);
nor U43212 (N_43212,N_41056,N_41032);
nor U43213 (N_43213,N_40251,N_41156);
nand U43214 (N_43214,N_40010,N_41456);
nor U43215 (N_43215,N_40648,N_41143);
or U43216 (N_43216,N_41512,N_40560);
or U43217 (N_43217,N_41585,N_40180);
nor U43218 (N_43218,N_41348,N_40157);
or U43219 (N_43219,N_40196,N_40218);
or U43220 (N_43220,N_41483,N_40950);
nor U43221 (N_43221,N_41481,N_41579);
nand U43222 (N_43222,N_41418,N_41977);
and U43223 (N_43223,N_41397,N_41045);
nor U43224 (N_43224,N_40104,N_41513);
and U43225 (N_43225,N_41826,N_40192);
nor U43226 (N_43226,N_40720,N_40038);
nor U43227 (N_43227,N_40546,N_41683);
nand U43228 (N_43228,N_41916,N_40255);
nand U43229 (N_43229,N_40053,N_41547);
or U43230 (N_43230,N_41470,N_40710);
or U43231 (N_43231,N_40711,N_40090);
and U43232 (N_43232,N_41616,N_41809);
nor U43233 (N_43233,N_40084,N_40565);
nand U43234 (N_43234,N_40556,N_41451);
nor U43235 (N_43235,N_41941,N_41259);
nand U43236 (N_43236,N_41665,N_41968);
nand U43237 (N_43237,N_40270,N_40557);
nor U43238 (N_43238,N_41455,N_41553);
nand U43239 (N_43239,N_41233,N_41478);
nor U43240 (N_43240,N_40872,N_40684);
nand U43241 (N_43241,N_41455,N_41038);
nand U43242 (N_43242,N_41381,N_41180);
and U43243 (N_43243,N_40173,N_40001);
and U43244 (N_43244,N_40178,N_41751);
nor U43245 (N_43245,N_40214,N_40333);
and U43246 (N_43246,N_41050,N_40315);
or U43247 (N_43247,N_40757,N_41604);
nand U43248 (N_43248,N_40847,N_41468);
nand U43249 (N_43249,N_41583,N_40769);
or U43250 (N_43250,N_41137,N_40987);
nor U43251 (N_43251,N_40758,N_41557);
or U43252 (N_43252,N_41009,N_41732);
nor U43253 (N_43253,N_41680,N_41784);
nor U43254 (N_43254,N_40032,N_40045);
nand U43255 (N_43255,N_40315,N_41830);
nor U43256 (N_43256,N_40458,N_41247);
nand U43257 (N_43257,N_41330,N_40892);
and U43258 (N_43258,N_40021,N_41577);
or U43259 (N_43259,N_41158,N_41479);
nand U43260 (N_43260,N_40061,N_41496);
xnor U43261 (N_43261,N_41013,N_41531);
nor U43262 (N_43262,N_41492,N_41913);
or U43263 (N_43263,N_40857,N_41341);
nor U43264 (N_43264,N_41707,N_41666);
nand U43265 (N_43265,N_41139,N_40520);
or U43266 (N_43266,N_41378,N_40654);
nand U43267 (N_43267,N_40119,N_41304);
nand U43268 (N_43268,N_40705,N_40700);
and U43269 (N_43269,N_40609,N_41965);
nand U43270 (N_43270,N_41195,N_41349);
nand U43271 (N_43271,N_41363,N_40983);
and U43272 (N_43272,N_41636,N_41950);
and U43273 (N_43273,N_40557,N_40997);
and U43274 (N_43274,N_41083,N_40860);
or U43275 (N_43275,N_41704,N_40766);
or U43276 (N_43276,N_41409,N_41086);
xor U43277 (N_43277,N_41055,N_40078);
or U43278 (N_43278,N_40593,N_41956);
or U43279 (N_43279,N_40399,N_41809);
nor U43280 (N_43280,N_41633,N_41472);
xnor U43281 (N_43281,N_40324,N_40831);
or U43282 (N_43282,N_41384,N_40023);
xnor U43283 (N_43283,N_41209,N_41494);
nor U43284 (N_43284,N_41712,N_40338);
or U43285 (N_43285,N_41431,N_41273);
nand U43286 (N_43286,N_40903,N_41058);
nor U43287 (N_43287,N_41892,N_40269);
nand U43288 (N_43288,N_41076,N_40104);
nor U43289 (N_43289,N_40279,N_40871);
nor U43290 (N_43290,N_40067,N_41519);
nor U43291 (N_43291,N_40513,N_40183);
and U43292 (N_43292,N_40530,N_40551);
nor U43293 (N_43293,N_41171,N_41654);
nor U43294 (N_43294,N_40372,N_40329);
nor U43295 (N_43295,N_40616,N_40909);
nand U43296 (N_43296,N_40715,N_41361);
nor U43297 (N_43297,N_40287,N_41409);
nand U43298 (N_43298,N_41760,N_40274);
nor U43299 (N_43299,N_41265,N_40979);
or U43300 (N_43300,N_40831,N_41989);
nand U43301 (N_43301,N_40759,N_40334);
or U43302 (N_43302,N_40943,N_41142);
nor U43303 (N_43303,N_40530,N_41550);
nand U43304 (N_43304,N_41154,N_40152);
and U43305 (N_43305,N_41555,N_40480);
nor U43306 (N_43306,N_41786,N_40339);
nand U43307 (N_43307,N_41141,N_41775);
nand U43308 (N_43308,N_41569,N_40016);
or U43309 (N_43309,N_41541,N_41163);
nand U43310 (N_43310,N_40384,N_40534);
nand U43311 (N_43311,N_41436,N_41879);
nand U43312 (N_43312,N_41795,N_40961);
nor U43313 (N_43313,N_40370,N_41910);
and U43314 (N_43314,N_41141,N_41547);
nor U43315 (N_43315,N_41436,N_40145);
or U43316 (N_43316,N_41666,N_40592);
and U43317 (N_43317,N_41011,N_41051);
nand U43318 (N_43318,N_40485,N_40110);
or U43319 (N_43319,N_40159,N_41636);
nor U43320 (N_43320,N_41511,N_40721);
xnor U43321 (N_43321,N_40450,N_40923);
and U43322 (N_43322,N_40001,N_41293);
nor U43323 (N_43323,N_41723,N_40780);
and U43324 (N_43324,N_40691,N_41808);
nor U43325 (N_43325,N_41528,N_40766);
or U43326 (N_43326,N_40931,N_41651);
nand U43327 (N_43327,N_41569,N_40865);
nand U43328 (N_43328,N_40404,N_40569);
nand U43329 (N_43329,N_41703,N_41540);
and U43330 (N_43330,N_40300,N_41409);
nor U43331 (N_43331,N_41927,N_41281);
nand U43332 (N_43332,N_40558,N_40874);
nand U43333 (N_43333,N_40298,N_40305);
and U43334 (N_43334,N_41243,N_40855);
and U43335 (N_43335,N_40546,N_41841);
and U43336 (N_43336,N_41248,N_40866);
or U43337 (N_43337,N_40235,N_41207);
and U43338 (N_43338,N_40953,N_40908);
nand U43339 (N_43339,N_41689,N_40804);
xor U43340 (N_43340,N_41363,N_40712);
nand U43341 (N_43341,N_41913,N_41311);
and U43342 (N_43342,N_40932,N_41434);
and U43343 (N_43343,N_41597,N_41554);
and U43344 (N_43344,N_40592,N_40915);
nand U43345 (N_43345,N_40002,N_41594);
nor U43346 (N_43346,N_40457,N_41116);
and U43347 (N_43347,N_40351,N_40789);
and U43348 (N_43348,N_41664,N_41602);
nor U43349 (N_43349,N_40228,N_41930);
nor U43350 (N_43350,N_40716,N_41130);
or U43351 (N_43351,N_40583,N_41513);
nand U43352 (N_43352,N_40331,N_41664);
nor U43353 (N_43353,N_41016,N_40538);
nand U43354 (N_43354,N_41166,N_41879);
or U43355 (N_43355,N_40125,N_40798);
nor U43356 (N_43356,N_40641,N_41990);
nand U43357 (N_43357,N_41571,N_41722);
nor U43358 (N_43358,N_41338,N_40549);
and U43359 (N_43359,N_41938,N_40218);
or U43360 (N_43360,N_40789,N_41819);
nor U43361 (N_43361,N_40926,N_40107);
nor U43362 (N_43362,N_41006,N_41150);
nor U43363 (N_43363,N_40360,N_41160);
nor U43364 (N_43364,N_40058,N_41781);
nand U43365 (N_43365,N_41827,N_40214);
and U43366 (N_43366,N_40186,N_41138);
nor U43367 (N_43367,N_41334,N_41051);
or U43368 (N_43368,N_40568,N_41483);
and U43369 (N_43369,N_40065,N_40563);
nor U43370 (N_43370,N_41427,N_41324);
or U43371 (N_43371,N_40950,N_40836);
and U43372 (N_43372,N_41217,N_41090);
or U43373 (N_43373,N_41028,N_41147);
xnor U43374 (N_43374,N_41003,N_40383);
and U43375 (N_43375,N_40900,N_41170);
and U43376 (N_43376,N_40479,N_41728);
or U43377 (N_43377,N_41873,N_41343);
nor U43378 (N_43378,N_40449,N_40835);
nor U43379 (N_43379,N_41689,N_41722);
nor U43380 (N_43380,N_40887,N_41417);
and U43381 (N_43381,N_41713,N_41791);
nand U43382 (N_43382,N_40775,N_40730);
nor U43383 (N_43383,N_40222,N_40375);
or U43384 (N_43384,N_40305,N_40148);
and U43385 (N_43385,N_41308,N_40540);
nor U43386 (N_43386,N_41348,N_41446);
and U43387 (N_43387,N_41397,N_40366);
nand U43388 (N_43388,N_40473,N_41766);
nor U43389 (N_43389,N_40014,N_41713);
nand U43390 (N_43390,N_41946,N_40116);
and U43391 (N_43391,N_40383,N_40631);
and U43392 (N_43392,N_41622,N_41248);
nand U43393 (N_43393,N_41679,N_40843);
or U43394 (N_43394,N_40997,N_41934);
nor U43395 (N_43395,N_41321,N_41304);
and U43396 (N_43396,N_41073,N_40109);
and U43397 (N_43397,N_40995,N_40962);
nor U43398 (N_43398,N_40396,N_40678);
or U43399 (N_43399,N_40810,N_40887);
nor U43400 (N_43400,N_41911,N_40497);
nor U43401 (N_43401,N_41758,N_40445);
nor U43402 (N_43402,N_40178,N_41021);
and U43403 (N_43403,N_41668,N_41880);
nor U43404 (N_43404,N_40968,N_40417);
xor U43405 (N_43405,N_40546,N_41820);
nor U43406 (N_43406,N_41853,N_41413);
nor U43407 (N_43407,N_40531,N_40995);
and U43408 (N_43408,N_41280,N_41046);
or U43409 (N_43409,N_40412,N_40972);
and U43410 (N_43410,N_41506,N_41936);
and U43411 (N_43411,N_41087,N_41071);
and U43412 (N_43412,N_40075,N_41249);
or U43413 (N_43413,N_41715,N_41716);
nor U43414 (N_43414,N_41992,N_40752);
or U43415 (N_43415,N_41546,N_40242);
or U43416 (N_43416,N_40822,N_40241);
nand U43417 (N_43417,N_40402,N_41101);
nor U43418 (N_43418,N_40609,N_40308);
or U43419 (N_43419,N_40242,N_40002);
nand U43420 (N_43420,N_41241,N_41633);
nand U43421 (N_43421,N_40395,N_40840);
nand U43422 (N_43422,N_41038,N_40024);
or U43423 (N_43423,N_40452,N_41860);
or U43424 (N_43424,N_40151,N_41365);
nor U43425 (N_43425,N_41107,N_41600);
nor U43426 (N_43426,N_41460,N_41835);
nor U43427 (N_43427,N_41198,N_41070);
nor U43428 (N_43428,N_40782,N_40724);
or U43429 (N_43429,N_40219,N_41821);
and U43430 (N_43430,N_41518,N_40022);
and U43431 (N_43431,N_40550,N_41851);
and U43432 (N_43432,N_40772,N_40762);
nor U43433 (N_43433,N_41802,N_40694);
and U43434 (N_43434,N_41519,N_41895);
nor U43435 (N_43435,N_41856,N_41776);
or U43436 (N_43436,N_40247,N_40417);
and U43437 (N_43437,N_40988,N_41418);
nand U43438 (N_43438,N_40581,N_41182);
and U43439 (N_43439,N_40203,N_41603);
nand U43440 (N_43440,N_40245,N_41157);
nor U43441 (N_43441,N_41337,N_40138);
nand U43442 (N_43442,N_40873,N_41019);
and U43443 (N_43443,N_40379,N_40232);
nand U43444 (N_43444,N_41892,N_40314);
or U43445 (N_43445,N_41378,N_40162);
nor U43446 (N_43446,N_40537,N_41040);
nand U43447 (N_43447,N_40643,N_41851);
and U43448 (N_43448,N_40865,N_41505);
or U43449 (N_43449,N_40344,N_40158);
or U43450 (N_43450,N_41081,N_40416);
or U43451 (N_43451,N_40529,N_41243);
and U43452 (N_43452,N_41294,N_41059);
nor U43453 (N_43453,N_41166,N_41345);
and U43454 (N_43454,N_40663,N_41556);
nor U43455 (N_43455,N_40845,N_40188);
nor U43456 (N_43456,N_41901,N_41452);
nor U43457 (N_43457,N_41486,N_40020);
and U43458 (N_43458,N_40029,N_41926);
or U43459 (N_43459,N_40852,N_40981);
nor U43460 (N_43460,N_40341,N_41107);
nor U43461 (N_43461,N_40551,N_40754);
nor U43462 (N_43462,N_41142,N_40818);
nand U43463 (N_43463,N_40023,N_40071);
nand U43464 (N_43464,N_41832,N_41455);
and U43465 (N_43465,N_41948,N_40064);
and U43466 (N_43466,N_41578,N_41439);
or U43467 (N_43467,N_41367,N_41973);
nand U43468 (N_43468,N_41076,N_40518);
nor U43469 (N_43469,N_40547,N_41398);
or U43470 (N_43470,N_40111,N_41008);
or U43471 (N_43471,N_40105,N_41284);
nand U43472 (N_43472,N_41852,N_41777);
or U43473 (N_43473,N_41864,N_40920);
or U43474 (N_43474,N_41185,N_40206);
nor U43475 (N_43475,N_40914,N_41058);
nand U43476 (N_43476,N_40457,N_41434);
nand U43477 (N_43477,N_41571,N_40815);
nand U43478 (N_43478,N_41411,N_40534);
or U43479 (N_43479,N_40769,N_41626);
and U43480 (N_43480,N_41326,N_40077);
nand U43481 (N_43481,N_40915,N_41737);
nand U43482 (N_43482,N_40972,N_40657);
nor U43483 (N_43483,N_41839,N_40857);
or U43484 (N_43484,N_41819,N_41740);
nor U43485 (N_43485,N_40272,N_41321);
nand U43486 (N_43486,N_41808,N_41224);
nand U43487 (N_43487,N_41895,N_40239);
nand U43488 (N_43488,N_40444,N_40325);
nand U43489 (N_43489,N_41738,N_40921);
nor U43490 (N_43490,N_40290,N_41249);
or U43491 (N_43491,N_40722,N_40947);
nor U43492 (N_43492,N_41867,N_41319);
nor U43493 (N_43493,N_40390,N_41527);
xor U43494 (N_43494,N_40948,N_40418);
or U43495 (N_43495,N_41285,N_40549);
nor U43496 (N_43496,N_40554,N_40682);
or U43497 (N_43497,N_41664,N_41776);
nor U43498 (N_43498,N_40552,N_40936);
nand U43499 (N_43499,N_40521,N_41772);
nand U43500 (N_43500,N_40675,N_41225);
nor U43501 (N_43501,N_40812,N_41097);
nor U43502 (N_43502,N_41703,N_41319);
or U43503 (N_43503,N_41326,N_41188);
and U43504 (N_43504,N_41629,N_41620);
and U43505 (N_43505,N_40936,N_41523);
and U43506 (N_43506,N_40722,N_40499);
nand U43507 (N_43507,N_40746,N_41772);
or U43508 (N_43508,N_41543,N_41373);
or U43509 (N_43509,N_41473,N_41478);
and U43510 (N_43510,N_41627,N_40001);
or U43511 (N_43511,N_41423,N_40038);
nand U43512 (N_43512,N_40948,N_40762);
nor U43513 (N_43513,N_41018,N_41158);
nand U43514 (N_43514,N_41892,N_40120);
and U43515 (N_43515,N_40383,N_40916);
nor U43516 (N_43516,N_40613,N_40332);
and U43517 (N_43517,N_41212,N_41048);
and U43518 (N_43518,N_40045,N_40763);
and U43519 (N_43519,N_41226,N_41571);
or U43520 (N_43520,N_41734,N_41690);
nor U43521 (N_43521,N_41387,N_41562);
or U43522 (N_43522,N_41537,N_41306);
nand U43523 (N_43523,N_40472,N_40898);
nand U43524 (N_43524,N_40426,N_40391);
xnor U43525 (N_43525,N_41372,N_40384);
and U43526 (N_43526,N_41801,N_40022);
nor U43527 (N_43527,N_41178,N_40616);
nand U43528 (N_43528,N_41103,N_41534);
or U43529 (N_43529,N_40660,N_41183);
nor U43530 (N_43530,N_41146,N_41104);
nor U43531 (N_43531,N_41174,N_41383);
and U43532 (N_43532,N_41594,N_40405);
nand U43533 (N_43533,N_40870,N_40601);
or U43534 (N_43534,N_41802,N_41529);
nand U43535 (N_43535,N_40453,N_40673);
nand U43536 (N_43536,N_40067,N_40227);
nand U43537 (N_43537,N_41145,N_41783);
nand U43538 (N_43538,N_40597,N_40220);
and U43539 (N_43539,N_40440,N_40998);
or U43540 (N_43540,N_40772,N_41510);
nor U43541 (N_43541,N_40240,N_41930);
and U43542 (N_43542,N_40280,N_40254);
or U43543 (N_43543,N_41445,N_41805);
or U43544 (N_43544,N_41995,N_41760);
nand U43545 (N_43545,N_40888,N_40414);
or U43546 (N_43546,N_40805,N_40766);
nor U43547 (N_43547,N_40871,N_41429);
or U43548 (N_43548,N_40324,N_40602);
nor U43549 (N_43549,N_40220,N_41718);
nor U43550 (N_43550,N_40195,N_40166);
nor U43551 (N_43551,N_40386,N_41216);
and U43552 (N_43552,N_41932,N_40896);
and U43553 (N_43553,N_40218,N_41108);
nand U43554 (N_43554,N_41875,N_40100);
or U43555 (N_43555,N_41124,N_40792);
and U43556 (N_43556,N_41088,N_40560);
nor U43557 (N_43557,N_41916,N_40589);
and U43558 (N_43558,N_41831,N_40854);
or U43559 (N_43559,N_41545,N_40191);
nor U43560 (N_43560,N_41586,N_40905);
nor U43561 (N_43561,N_41354,N_40855);
nor U43562 (N_43562,N_41024,N_41565);
and U43563 (N_43563,N_41017,N_41804);
or U43564 (N_43564,N_40996,N_40532);
or U43565 (N_43565,N_40526,N_40298);
and U43566 (N_43566,N_40333,N_40372);
nor U43567 (N_43567,N_40870,N_41927);
nand U43568 (N_43568,N_40679,N_41603);
nand U43569 (N_43569,N_40818,N_40977);
or U43570 (N_43570,N_40149,N_40631);
nand U43571 (N_43571,N_40084,N_40633);
or U43572 (N_43572,N_41038,N_41143);
or U43573 (N_43573,N_41311,N_40702);
and U43574 (N_43574,N_40627,N_41685);
nand U43575 (N_43575,N_40354,N_41420);
and U43576 (N_43576,N_41344,N_40019);
or U43577 (N_43577,N_41951,N_40790);
xnor U43578 (N_43578,N_41407,N_40161);
and U43579 (N_43579,N_40382,N_41405);
and U43580 (N_43580,N_41304,N_40206);
xnor U43581 (N_43581,N_41849,N_41692);
nand U43582 (N_43582,N_41279,N_41129);
nor U43583 (N_43583,N_40867,N_41905);
nor U43584 (N_43584,N_41610,N_41254);
nor U43585 (N_43585,N_41546,N_40291);
nor U43586 (N_43586,N_41660,N_40764);
nand U43587 (N_43587,N_40960,N_41490);
and U43588 (N_43588,N_40050,N_41782);
nor U43589 (N_43589,N_41216,N_41379);
xnor U43590 (N_43590,N_41240,N_41213);
nor U43591 (N_43591,N_40711,N_40679);
nor U43592 (N_43592,N_41618,N_41234);
and U43593 (N_43593,N_40003,N_40946);
xor U43594 (N_43594,N_40967,N_41521);
nor U43595 (N_43595,N_40422,N_41990);
or U43596 (N_43596,N_41932,N_40670);
or U43597 (N_43597,N_41094,N_40747);
nand U43598 (N_43598,N_40628,N_40139);
or U43599 (N_43599,N_40647,N_40822);
nor U43600 (N_43600,N_41312,N_40364);
xor U43601 (N_43601,N_41464,N_40269);
or U43602 (N_43602,N_40899,N_41076);
nor U43603 (N_43603,N_41064,N_41710);
or U43604 (N_43604,N_40585,N_41207);
nand U43605 (N_43605,N_41536,N_40344);
nand U43606 (N_43606,N_41787,N_41647);
nand U43607 (N_43607,N_41171,N_41396);
or U43608 (N_43608,N_40518,N_41568);
and U43609 (N_43609,N_40302,N_40338);
and U43610 (N_43610,N_40603,N_40677);
and U43611 (N_43611,N_41758,N_40571);
and U43612 (N_43612,N_41502,N_40353);
nor U43613 (N_43613,N_41745,N_41010);
nand U43614 (N_43614,N_41972,N_41834);
and U43615 (N_43615,N_40767,N_40451);
and U43616 (N_43616,N_40873,N_40207);
or U43617 (N_43617,N_41331,N_40600);
and U43618 (N_43618,N_40951,N_40127);
and U43619 (N_43619,N_41986,N_41504);
xnor U43620 (N_43620,N_40117,N_40994);
nor U43621 (N_43621,N_41945,N_40239);
nand U43622 (N_43622,N_40981,N_40349);
nand U43623 (N_43623,N_41908,N_40953);
nor U43624 (N_43624,N_41256,N_41077);
or U43625 (N_43625,N_41025,N_41499);
and U43626 (N_43626,N_41963,N_41505);
nor U43627 (N_43627,N_40686,N_41019);
and U43628 (N_43628,N_41565,N_41179);
and U43629 (N_43629,N_40612,N_40047);
nor U43630 (N_43630,N_40696,N_41796);
and U43631 (N_43631,N_40594,N_41073);
and U43632 (N_43632,N_41014,N_41479);
nand U43633 (N_43633,N_40376,N_41826);
or U43634 (N_43634,N_40560,N_40924);
and U43635 (N_43635,N_40086,N_41399);
and U43636 (N_43636,N_41625,N_40926);
and U43637 (N_43637,N_40728,N_41905);
and U43638 (N_43638,N_41314,N_41191);
nand U43639 (N_43639,N_40983,N_41215);
nand U43640 (N_43640,N_41188,N_41316);
or U43641 (N_43641,N_40602,N_40467);
nand U43642 (N_43642,N_40125,N_40903);
xnor U43643 (N_43643,N_40268,N_41897);
or U43644 (N_43644,N_41072,N_40583);
or U43645 (N_43645,N_41091,N_40448);
nand U43646 (N_43646,N_41323,N_41314);
nand U43647 (N_43647,N_41809,N_41902);
and U43648 (N_43648,N_40845,N_40779);
or U43649 (N_43649,N_41370,N_41753);
nand U43650 (N_43650,N_41508,N_41213);
nand U43651 (N_43651,N_40319,N_41276);
nor U43652 (N_43652,N_40153,N_40767);
nand U43653 (N_43653,N_40326,N_40012);
nand U43654 (N_43654,N_41358,N_40707);
and U43655 (N_43655,N_40854,N_41330);
nand U43656 (N_43656,N_40635,N_40374);
nand U43657 (N_43657,N_40913,N_40346);
nor U43658 (N_43658,N_40292,N_40964);
xnor U43659 (N_43659,N_40741,N_41560);
and U43660 (N_43660,N_41986,N_41122);
or U43661 (N_43661,N_41854,N_41950);
or U43662 (N_43662,N_40156,N_40677);
or U43663 (N_43663,N_41761,N_40495);
nor U43664 (N_43664,N_40997,N_41305);
nor U43665 (N_43665,N_41665,N_40703);
nor U43666 (N_43666,N_40914,N_40316);
nand U43667 (N_43667,N_41524,N_40624);
or U43668 (N_43668,N_41711,N_41432);
or U43669 (N_43669,N_40050,N_40378);
or U43670 (N_43670,N_40943,N_41653);
nor U43671 (N_43671,N_40575,N_41794);
nor U43672 (N_43672,N_40408,N_40241);
or U43673 (N_43673,N_40164,N_40300);
nor U43674 (N_43674,N_40912,N_41209);
nor U43675 (N_43675,N_40175,N_41903);
nor U43676 (N_43676,N_40218,N_40059);
or U43677 (N_43677,N_41131,N_41324);
or U43678 (N_43678,N_40555,N_41070);
nand U43679 (N_43679,N_40108,N_40879);
or U43680 (N_43680,N_40439,N_41175);
nor U43681 (N_43681,N_41905,N_41008);
nand U43682 (N_43682,N_40028,N_41725);
nand U43683 (N_43683,N_40533,N_41383);
nand U43684 (N_43684,N_40144,N_41699);
or U43685 (N_43685,N_41750,N_40130);
and U43686 (N_43686,N_41746,N_41324);
and U43687 (N_43687,N_41689,N_40243);
xnor U43688 (N_43688,N_40843,N_41220);
or U43689 (N_43689,N_41233,N_41274);
and U43690 (N_43690,N_41708,N_41256);
nand U43691 (N_43691,N_41058,N_41071);
nor U43692 (N_43692,N_40404,N_41857);
and U43693 (N_43693,N_41002,N_41719);
nor U43694 (N_43694,N_40224,N_40626);
and U43695 (N_43695,N_40296,N_40576);
nand U43696 (N_43696,N_41680,N_41857);
nor U43697 (N_43697,N_41113,N_40029);
and U43698 (N_43698,N_40476,N_40052);
nand U43699 (N_43699,N_40762,N_41114);
nor U43700 (N_43700,N_40283,N_41921);
xor U43701 (N_43701,N_40532,N_41916);
nor U43702 (N_43702,N_41419,N_40932);
and U43703 (N_43703,N_41350,N_41236);
or U43704 (N_43704,N_40664,N_40354);
nand U43705 (N_43705,N_40094,N_41248);
nor U43706 (N_43706,N_40654,N_41340);
or U43707 (N_43707,N_40989,N_40000);
nor U43708 (N_43708,N_41772,N_41028);
or U43709 (N_43709,N_41223,N_40701);
or U43710 (N_43710,N_40521,N_40599);
nor U43711 (N_43711,N_40941,N_41964);
and U43712 (N_43712,N_41648,N_40503);
or U43713 (N_43713,N_40161,N_40593);
nor U43714 (N_43714,N_41240,N_40594);
and U43715 (N_43715,N_41859,N_40536);
nor U43716 (N_43716,N_40267,N_40404);
nor U43717 (N_43717,N_41475,N_40978);
nor U43718 (N_43718,N_40872,N_40605);
and U43719 (N_43719,N_41077,N_41751);
nand U43720 (N_43720,N_41430,N_40931);
nor U43721 (N_43721,N_41186,N_41024);
or U43722 (N_43722,N_40392,N_41785);
or U43723 (N_43723,N_41508,N_41583);
nand U43724 (N_43724,N_41149,N_41998);
and U43725 (N_43725,N_40498,N_41341);
and U43726 (N_43726,N_41915,N_41011);
nand U43727 (N_43727,N_41619,N_41886);
and U43728 (N_43728,N_40994,N_40350);
and U43729 (N_43729,N_40842,N_41597);
nor U43730 (N_43730,N_41236,N_41887);
nor U43731 (N_43731,N_41107,N_40598);
and U43732 (N_43732,N_40837,N_41963);
or U43733 (N_43733,N_41824,N_41915);
nor U43734 (N_43734,N_40019,N_41461);
or U43735 (N_43735,N_40273,N_41044);
or U43736 (N_43736,N_40643,N_40316);
or U43737 (N_43737,N_41654,N_41058);
nor U43738 (N_43738,N_40122,N_40706);
and U43739 (N_43739,N_40927,N_40839);
nand U43740 (N_43740,N_40628,N_41820);
and U43741 (N_43741,N_40705,N_41000);
or U43742 (N_43742,N_41130,N_41291);
and U43743 (N_43743,N_41061,N_40746);
nor U43744 (N_43744,N_40427,N_41401);
and U43745 (N_43745,N_41641,N_40961);
nor U43746 (N_43746,N_40006,N_41712);
and U43747 (N_43747,N_40887,N_40643);
nand U43748 (N_43748,N_41009,N_41174);
nand U43749 (N_43749,N_40340,N_41222);
or U43750 (N_43750,N_40659,N_41853);
nand U43751 (N_43751,N_41611,N_40500);
nand U43752 (N_43752,N_41767,N_41250);
nand U43753 (N_43753,N_40211,N_41112);
nand U43754 (N_43754,N_40835,N_40928);
nor U43755 (N_43755,N_41415,N_40935);
and U43756 (N_43756,N_40266,N_40288);
and U43757 (N_43757,N_40054,N_41952);
and U43758 (N_43758,N_41904,N_40258);
and U43759 (N_43759,N_40029,N_40195);
or U43760 (N_43760,N_40620,N_40594);
and U43761 (N_43761,N_41623,N_41348);
xor U43762 (N_43762,N_41613,N_40823);
and U43763 (N_43763,N_40092,N_41657);
or U43764 (N_43764,N_41497,N_41952);
nor U43765 (N_43765,N_41143,N_40908);
xor U43766 (N_43766,N_41199,N_41973);
nand U43767 (N_43767,N_41043,N_40100);
and U43768 (N_43768,N_41224,N_40526);
nand U43769 (N_43769,N_40611,N_40283);
or U43770 (N_43770,N_41185,N_41921);
nand U43771 (N_43771,N_41425,N_41747);
nand U43772 (N_43772,N_40206,N_41772);
or U43773 (N_43773,N_40887,N_41301);
or U43774 (N_43774,N_40269,N_41792);
xnor U43775 (N_43775,N_41894,N_41963);
nor U43776 (N_43776,N_40615,N_41202);
nand U43777 (N_43777,N_41386,N_40035);
or U43778 (N_43778,N_41597,N_41021);
and U43779 (N_43779,N_40936,N_40002);
or U43780 (N_43780,N_40172,N_40400);
nor U43781 (N_43781,N_41540,N_41644);
or U43782 (N_43782,N_40247,N_40887);
xor U43783 (N_43783,N_41909,N_40696);
or U43784 (N_43784,N_40329,N_41102);
and U43785 (N_43785,N_40209,N_40678);
nand U43786 (N_43786,N_40470,N_41875);
nand U43787 (N_43787,N_41247,N_40558);
nor U43788 (N_43788,N_40538,N_40035);
nor U43789 (N_43789,N_40214,N_40813);
nor U43790 (N_43790,N_40319,N_41805);
or U43791 (N_43791,N_40160,N_40021);
and U43792 (N_43792,N_40955,N_41702);
nor U43793 (N_43793,N_40783,N_40031);
or U43794 (N_43794,N_40796,N_40389);
or U43795 (N_43795,N_40561,N_40811);
or U43796 (N_43796,N_41620,N_41207);
nand U43797 (N_43797,N_40211,N_41638);
nand U43798 (N_43798,N_41300,N_40733);
and U43799 (N_43799,N_40289,N_40167);
nor U43800 (N_43800,N_41433,N_41218);
or U43801 (N_43801,N_40977,N_41580);
and U43802 (N_43802,N_41918,N_40161);
and U43803 (N_43803,N_40003,N_41419);
or U43804 (N_43804,N_40307,N_41059);
nand U43805 (N_43805,N_41974,N_41795);
nand U43806 (N_43806,N_41375,N_41645);
or U43807 (N_43807,N_41379,N_41583);
nand U43808 (N_43808,N_41996,N_41769);
or U43809 (N_43809,N_41353,N_40191);
and U43810 (N_43810,N_41080,N_41859);
nand U43811 (N_43811,N_40277,N_41493);
nand U43812 (N_43812,N_40246,N_41492);
or U43813 (N_43813,N_41704,N_41446);
nand U43814 (N_43814,N_40688,N_40504);
or U43815 (N_43815,N_41663,N_40937);
or U43816 (N_43816,N_40978,N_40577);
nand U43817 (N_43817,N_40379,N_40445);
nor U43818 (N_43818,N_40789,N_41142);
nor U43819 (N_43819,N_40932,N_40551);
nor U43820 (N_43820,N_41293,N_40478);
nand U43821 (N_43821,N_40588,N_41138);
nor U43822 (N_43822,N_40516,N_40266);
nand U43823 (N_43823,N_40232,N_41417);
nand U43824 (N_43824,N_40002,N_41890);
or U43825 (N_43825,N_40137,N_40175);
nand U43826 (N_43826,N_41553,N_40484);
nor U43827 (N_43827,N_41594,N_41617);
and U43828 (N_43828,N_40793,N_41243);
or U43829 (N_43829,N_41065,N_41006);
nand U43830 (N_43830,N_40325,N_41834);
nor U43831 (N_43831,N_41359,N_40572);
nor U43832 (N_43832,N_40876,N_41419);
or U43833 (N_43833,N_41838,N_41092);
nand U43834 (N_43834,N_40876,N_40252);
or U43835 (N_43835,N_40026,N_40597);
and U43836 (N_43836,N_41001,N_41008);
nor U43837 (N_43837,N_40524,N_41413);
and U43838 (N_43838,N_41649,N_40754);
nand U43839 (N_43839,N_40264,N_41833);
nor U43840 (N_43840,N_41268,N_41159);
and U43841 (N_43841,N_40988,N_41217);
nand U43842 (N_43842,N_41125,N_40553);
nand U43843 (N_43843,N_40435,N_40701);
or U43844 (N_43844,N_40202,N_40644);
nand U43845 (N_43845,N_41157,N_40830);
or U43846 (N_43846,N_40839,N_41978);
and U43847 (N_43847,N_41686,N_41945);
nor U43848 (N_43848,N_41955,N_41466);
nor U43849 (N_43849,N_40634,N_41253);
nand U43850 (N_43850,N_40739,N_40508);
and U43851 (N_43851,N_40840,N_41459);
or U43852 (N_43852,N_41507,N_40396);
nand U43853 (N_43853,N_41261,N_40290);
nor U43854 (N_43854,N_41378,N_40454);
and U43855 (N_43855,N_41913,N_40892);
nand U43856 (N_43856,N_40643,N_40451);
nand U43857 (N_43857,N_41936,N_40101);
nand U43858 (N_43858,N_41019,N_41526);
or U43859 (N_43859,N_40845,N_40325);
nand U43860 (N_43860,N_41097,N_40729);
nor U43861 (N_43861,N_41971,N_41367);
nor U43862 (N_43862,N_40200,N_40280);
nor U43863 (N_43863,N_41659,N_41755);
nand U43864 (N_43864,N_41988,N_41930);
and U43865 (N_43865,N_40772,N_40808);
nor U43866 (N_43866,N_40715,N_41171);
nor U43867 (N_43867,N_40606,N_41751);
or U43868 (N_43868,N_40795,N_41574);
and U43869 (N_43869,N_40117,N_40535);
nand U43870 (N_43870,N_41014,N_40265);
or U43871 (N_43871,N_41202,N_41172);
or U43872 (N_43872,N_40308,N_41455);
xor U43873 (N_43873,N_40372,N_40153);
and U43874 (N_43874,N_40369,N_41233);
nand U43875 (N_43875,N_41778,N_41136);
nor U43876 (N_43876,N_41731,N_41863);
nor U43877 (N_43877,N_41820,N_41503);
or U43878 (N_43878,N_40267,N_40375);
nor U43879 (N_43879,N_40035,N_41419);
nand U43880 (N_43880,N_40035,N_40758);
and U43881 (N_43881,N_41043,N_41595);
and U43882 (N_43882,N_41317,N_40181);
and U43883 (N_43883,N_40406,N_41961);
or U43884 (N_43884,N_40014,N_41755);
nand U43885 (N_43885,N_40027,N_41777);
nor U43886 (N_43886,N_41859,N_41089);
and U43887 (N_43887,N_41379,N_40474);
nor U43888 (N_43888,N_40370,N_41292);
or U43889 (N_43889,N_40165,N_40376);
nor U43890 (N_43890,N_41018,N_40563);
or U43891 (N_43891,N_40843,N_41435);
and U43892 (N_43892,N_41341,N_40713);
xor U43893 (N_43893,N_41716,N_40457);
nor U43894 (N_43894,N_40615,N_41805);
and U43895 (N_43895,N_40958,N_40324);
and U43896 (N_43896,N_41346,N_40197);
and U43897 (N_43897,N_41307,N_41680);
nor U43898 (N_43898,N_41417,N_40634);
nor U43899 (N_43899,N_41789,N_40645);
and U43900 (N_43900,N_41205,N_41442);
and U43901 (N_43901,N_40507,N_41098);
nor U43902 (N_43902,N_41197,N_41239);
nand U43903 (N_43903,N_40189,N_41813);
nand U43904 (N_43904,N_40457,N_40845);
and U43905 (N_43905,N_40686,N_40878);
nor U43906 (N_43906,N_40813,N_41236);
xnor U43907 (N_43907,N_41400,N_40593);
or U43908 (N_43908,N_40409,N_40103);
or U43909 (N_43909,N_40795,N_41233);
nand U43910 (N_43910,N_41366,N_40731);
and U43911 (N_43911,N_41153,N_41118);
nand U43912 (N_43912,N_41925,N_41921);
nor U43913 (N_43913,N_40404,N_40912);
nor U43914 (N_43914,N_40156,N_41975);
nand U43915 (N_43915,N_41895,N_40563);
and U43916 (N_43916,N_41390,N_40589);
nand U43917 (N_43917,N_40033,N_41676);
or U43918 (N_43918,N_40482,N_40432);
nor U43919 (N_43919,N_40411,N_41310);
or U43920 (N_43920,N_40075,N_41988);
or U43921 (N_43921,N_41489,N_40309);
or U43922 (N_43922,N_41651,N_40811);
nor U43923 (N_43923,N_41470,N_41059);
xor U43924 (N_43924,N_40101,N_40893);
nand U43925 (N_43925,N_41513,N_41305);
or U43926 (N_43926,N_41390,N_41506);
nand U43927 (N_43927,N_40069,N_40556);
or U43928 (N_43928,N_41377,N_40898);
nor U43929 (N_43929,N_41670,N_40794);
and U43930 (N_43930,N_40859,N_40432);
and U43931 (N_43931,N_40471,N_40153);
nand U43932 (N_43932,N_40802,N_41606);
or U43933 (N_43933,N_41341,N_40580);
nor U43934 (N_43934,N_41401,N_40672);
or U43935 (N_43935,N_40500,N_40331);
or U43936 (N_43936,N_40656,N_40604);
or U43937 (N_43937,N_40351,N_41630);
and U43938 (N_43938,N_40529,N_41288);
xor U43939 (N_43939,N_41954,N_40157);
and U43940 (N_43940,N_41099,N_40980);
or U43941 (N_43941,N_41038,N_40809);
or U43942 (N_43942,N_41953,N_40499);
or U43943 (N_43943,N_40679,N_40377);
nand U43944 (N_43944,N_41695,N_41232);
nor U43945 (N_43945,N_40338,N_41518);
nand U43946 (N_43946,N_41615,N_40897);
nor U43947 (N_43947,N_41951,N_40260);
and U43948 (N_43948,N_40561,N_40674);
or U43949 (N_43949,N_40456,N_40509);
nand U43950 (N_43950,N_41315,N_40443);
nor U43951 (N_43951,N_41992,N_40002);
nor U43952 (N_43952,N_40980,N_40656);
nand U43953 (N_43953,N_40211,N_40258);
and U43954 (N_43954,N_41759,N_40169);
nor U43955 (N_43955,N_41926,N_41925);
nor U43956 (N_43956,N_40570,N_41047);
or U43957 (N_43957,N_41237,N_40006);
nand U43958 (N_43958,N_41440,N_41213);
nor U43959 (N_43959,N_41699,N_40848);
nand U43960 (N_43960,N_40300,N_40858);
and U43961 (N_43961,N_41926,N_40602);
xnor U43962 (N_43962,N_41623,N_40311);
nor U43963 (N_43963,N_40878,N_40474);
or U43964 (N_43964,N_41028,N_40109);
and U43965 (N_43965,N_40244,N_41104);
and U43966 (N_43966,N_41449,N_40089);
nor U43967 (N_43967,N_40308,N_41481);
or U43968 (N_43968,N_40834,N_40892);
and U43969 (N_43969,N_40726,N_40646);
and U43970 (N_43970,N_41337,N_41104);
or U43971 (N_43971,N_40487,N_41059);
or U43972 (N_43972,N_40902,N_41977);
nor U43973 (N_43973,N_41228,N_40047);
nand U43974 (N_43974,N_41064,N_41565);
nand U43975 (N_43975,N_40789,N_41666);
nand U43976 (N_43976,N_41809,N_40338);
or U43977 (N_43977,N_41209,N_41178);
and U43978 (N_43978,N_40146,N_40749);
or U43979 (N_43979,N_41559,N_40961);
and U43980 (N_43980,N_40849,N_40128);
or U43981 (N_43981,N_40048,N_41381);
nor U43982 (N_43982,N_41839,N_40982);
and U43983 (N_43983,N_41455,N_40976);
nor U43984 (N_43984,N_41695,N_40881);
nand U43985 (N_43985,N_41013,N_41656);
nor U43986 (N_43986,N_40202,N_41648);
nand U43987 (N_43987,N_40910,N_41792);
nor U43988 (N_43988,N_41415,N_40429);
nand U43989 (N_43989,N_41964,N_41899);
or U43990 (N_43990,N_41088,N_41505);
and U43991 (N_43991,N_40752,N_41677);
or U43992 (N_43992,N_41397,N_41770);
and U43993 (N_43993,N_40130,N_41252);
nand U43994 (N_43994,N_41013,N_41200);
nor U43995 (N_43995,N_41286,N_40737);
nand U43996 (N_43996,N_40303,N_41883);
and U43997 (N_43997,N_40463,N_41928);
nand U43998 (N_43998,N_40942,N_41793);
nand U43999 (N_43999,N_41681,N_41206);
nor U44000 (N_44000,N_43917,N_42157);
nor U44001 (N_44001,N_43735,N_42913);
nand U44002 (N_44002,N_43931,N_43740);
or U44003 (N_44003,N_42156,N_42098);
nor U44004 (N_44004,N_42093,N_43833);
and U44005 (N_44005,N_43609,N_42878);
nor U44006 (N_44006,N_43975,N_43010);
and U44007 (N_44007,N_42396,N_42123);
or U44008 (N_44008,N_42781,N_42055);
xor U44009 (N_44009,N_42759,N_43845);
nand U44010 (N_44010,N_43046,N_43960);
nand U44011 (N_44011,N_42835,N_43172);
and U44012 (N_44012,N_43866,N_43313);
nor U44013 (N_44013,N_43196,N_43228);
nor U44014 (N_44014,N_42311,N_43851);
and U44015 (N_44015,N_43988,N_43547);
and U44016 (N_44016,N_43788,N_43443);
nand U44017 (N_44017,N_43958,N_42621);
and U44018 (N_44018,N_43572,N_43850);
nand U44019 (N_44019,N_43320,N_42625);
nand U44020 (N_44020,N_42280,N_42348);
nand U44021 (N_44021,N_43749,N_43865);
or U44022 (N_44022,N_43484,N_43289);
and U44023 (N_44023,N_43543,N_42673);
nor U44024 (N_44024,N_42198,N_42383);
nand U44025 (N_44025,N_43156,N_42530);
nor U44026 (N_44026,N_42392,N_43438);
nor U44027 (N_44027,N_42043,N_43981);
nand U44028 (N_44028,N_42889,N_42424);
or U44029 (N_44029,N_42062,N_42036);
or U44030 (N_44030,N_42379,N_42307);
nor U44031 (N_44031,N_43477,N_43369);
nand U44032 (N_44032,N_43149,N_42738);
or U44033 (N_44033,N_42146,N_42259);
xor U44034 (N_44034,N_43430,N_43863);
and U44035 (N_44035,N_43530,N_42532);
or U44036 (N_44036,N_43853,N_43508);
nand U44037 (N_44037,N_43295,N_42617);
and U44038 (N_44038,N_43654,N_42859);
nand U44039 (N_44039,N_43426,N_43246);
nor U44040 (N_44040,N_42124,N_42287);
or U44041 (N_44041,N_42543,N_43730);
or U44042 (N_44042,N_42829,N_42086);
nor U44043 (N_44043,N_42721,N_43445);
nand U44044 (N_44044,N_43005,N_42349);
or U44045 (N_44045,N_43110,N_42918);
nand U44046 (N_44046,N_42504,N_43413);
or U44047 (N_44047,N_42248,N_43009);
nor U44048 (N_44048,N_42095,N_42782);
or U44049 (N_44049,N_43684,N_43585);
nor U44050 (N_44050,N_42356,N_43551);
and U44051 (N_44051,N_42517,N_42097);
and U44052 (N_44052,N_42161,N_42616);
or U44053 (N_44053,N_43639,N_43029);
nor U44054 (N_44054,N_43444,N_42488);
and U44055 (N_44055,N_42393,N_43954);
nand U44056 (N_44056,N_42891,N_43271);
nand U44057 (N_44057,N_42813,N_42570);
or U44058 (N_44058,N_42810,N_43531);
nor U44059 (N_44059,N_42045,N_43347);
and U44060 (N_44060,N_43400,N_43679);
nand U44061 (N_44061,N_43063,N_42002);
or U44062 (N_44062,N_43283,N_43357);
nor U44063 (N_44063,N_42716,N_43948);
nand U44064 (N_44064,N_42176,N_42115);
and U44065 (N_44065,N_43300,N_42904);
nor U44066 (N_44066,N_42005,N_43433);
or U44067 (N_44067,N_43686,N_42523);
nand U44068 (N_44068,N_42887,N_43673);
nand U44069 (N_44069,N_42717,N_42141);
nand U44070 (N_44070,N_42578,N_43810);
and U44071 (N_44071,N_42037,N_43066);
and U44072 (N_44072,N_43586,N_42130);
xor U44073 (N_44073,N_43874,N_43200);
and U44074 (N_44074,N_42948,N_42221);
nor U44075 (N_44075,N_43742,N_42732);
or U44076 (N_44076,N_43145,N_43717);
nand U44077 (N_44077,N_43824,N_43549);
nor U44078 (N_44078,N_43902,N_42510);
nand U44079 (N_44079,N_42561,N_42257);
nor U44080 (N_44080,N_42049,N_42707);
nand U44081 (N_44081,N_42844,N_42126);
or U44082 (N_44082,N_43047,N_43823);
nand U44083 (N_44083,N_42206,N_43898);
or U44084 (N_44084,N_42085,N_42562);
and U44085 (N_44085,N_43457,N_42220);
and U44086 (N_44086,N_42678,N_42284);
and U44087 (N_44087,N_43532,N_43746);
and U44088 (N_44088,N_43521,N_43659);
nand U44089 (N_44089,N_42866,N_43640);
nand U44090 (N_44090,N_43809,N_43452);
nor U44091 (N_44091,N_42439,N_42529);
or U44092 (N_44092,N_43486,N_42806);
nand U44093 (N_44093,N_42010,N_43062);
and U44094 (N_44094,N_43577,N_42877);
nor U44095 (N_44095,N_42534,N_42652);
nor U44096 (N_44096,N_42648,N_43393);
or U44097 (N_44097,N_42177,N_42596);
and U44098 (N_44098,N_42870,N_42159);
and U44099 (N_44099,N_42201,N_42276);
or U44100 (N_44100,N_43178,N_43849);
xor U44101 (N_44101,N_42942,N_42091);
and U44102 (N_44102,N_43384,N_42317);
nand U44103 (N_44103,N_43260,N_42688);
nand U44104 (N_44104,N_43336,N_43995);
nand U44105 (N_44105,N_42399,N_43984);
and U44106 (N_44106,N_43937,N_42058);
and U44107 (N_44107,N_42905,N_42819);
nor U44108 (N_44108,N_42861,N_43195);
nor U44109 (N_44109,N_42594,N_43088);
nand U44110 (N_44110,N_42949,N_43424);
nor U44111 (N_44111,N_43672,N_42600);
nor U44112 (N_44112,N_42418,N_42729);
or U44113 (N_44113,N_42001,N_42660);
nand U44114 (N_44114,N_43461,N_42039);
nor U44115 (N_44115,N_43041,N_43277);
and U44116 (N_44116,N_43825,N_43170);
or U44117 (N_44117,N_42919,N_42193);
or U44118 (N_44118,N_43597,N_43500);
nand U44119 (N_44119,N_43364,N_42847);
nor U44120 (N_44120,N_42111,N_42962);
or U44121 (N_44121,N_42876,N_42929);
nor U44122 (N_44122,N_42644,N_42818);
nand U44123 (N_44123,N_43394,N_43253);
nor U44124 (N_44124,N_42726,N_43473);
and U44125 (N_44125,N_42295,N_42945);
nand U44126 (N_44126,N_42754,N_42983);
nand U44127 (N_44127,N_42746,N_43761);
nand U44128 (N_44128,N_42315,N_42546);
nand U44129 (N_44129,N_43692,N_42784);
or U44130 (N_44130,N_42793,N_43656);
nor U44131 (N_44131,N_43039,N_43732);
or U44132 (N_44132,N_43598,N_42492);
or U44133 (N_44133,N_43795,N_43959);
nor U44134 (N_44134,N_42432,N_43753);
nand U44135 (N_44135,N_43180,N_42106);
or U44136 (N_44136,N_43334,N_43385);
nand U44137 (N_44137,N_42387,N_43698);
nor U44138 (N_44138,N_43164,N_43647);
or U44139 (N_44139,N_42338,N_43829);
and U44140 (N_44140,N_42083,N_43186);
nor U44141 (N_44141,N_42635,N_42883);
or U44142 (N_44142,N_42382,N_43675);
or U44143 (N_44143,N_42417,N_43745);
or U44144 (N_44144,N_43620,N_42944);
nand U44145 (N_44145,N_42377,N_43250);
nand U44146 (N_44146,N_42266,N_43338);
nor U44147 (N_44147,N_42242,N_42080);
and U44148 (N_44148,N_43281,N_42737);
nor U44149 (N_44149,N_42419,N_43227);
or U44150 (N_44150,N_43933,N_43020);
or U44151 (N_44151,N_42473,N_42996);
and U44152 (N_44152,N_42760,N_42050);
or U44153 (N_44153,N_43564,N_42880);
nor U44154 (N_44154,N_42727,N_42826);
nand U44155 (N_44155,N_42502,N_43565);
nand U44156 (N_44156,N_42267,N_42512);
or U44157 (N_44157,N_43367,N_43723);
xnor U44158 (N_44158,N_42825,N_43789);
and U44159 (N_44159,N_43285,N_43867);
or U44160 (N_44160,N_43812,N_42371);
nor U44161 (N_44161,N_42458,N_42542);
nor U44162 (N_44162,N_42117,N_42636);
xnor U44163 (N_44163,N_43512,N_42327);
xor U44164 (N_44164,N_43026,N_42885);
and U44165 (N_44165,N_43807,N_43072);
and U44166 (N_44166,N_42511,N_42090);
nor U44167 (N_44167,N_42581,N_43923);
nor U44168 (N_44168,N_43463,N_43183);
nand U44169 (N_44169,N_42475,N_43095);
or U44170 (N_44170,N_43011,N_43217);
nor U44171 (N_44171,N_42306,N_43298);
nand U44172 (N_44172,N_43474,N_42369);
nand U44173 (N_44173,N_43569,N_43814);
nand U44174 (N_44174,N_43024,N_42351);
nand U44175 (N_44175,N_42397,N_43226);
nor U44176 (N_44176,N_42373,N_43575);
nor U44177 (N_44177,N_43361,N_42139);
and U44178 (N_44178,N_42375,N_42506);
nand U44179 (N_44179,N_42063,N_42898);
and U44180 (N_44180,N_42078,N_43398);
or U44181 (N_44181,N_42171,N_43117);
nand U44182 (N_44182,N_42467,N_43727);
nor U44183 (N_44183,N_42551,N_42838);
and U44184 (N_44184,N_42541,N_42074);
and U44185 (N_44185,N_43970,N_43202);
nor U44186 (N_44186,N_42548,N_42150);
or U44187 (N_44187,N_43816,N_42531);
or U44188 (N_44188,N_42990,N_42698);
nand U44189 (N_44189,N_42014,N_43151);
or U44190 (N_44190,N_43374,N_42857);
nor U44191 (N_44191,N_42102,N_43012);
and U44192 (N_44192,N_43506,N_42639);
or U44193 (N_44193,N_42910,N_42025);
nand U44194 (N_44194,N_42686,N_42586);
xnor U44195 (N_44195,N_42264,N_42282);
or U44196 (N_44196,N_42122,N_42185);
nand U44197 (N_44197,N_43124,N_42524);
and U44198 (N_44198,N_42019,N_42138);
or U44199 (N_44199,N_42997,N_43232);
or U44200 (N_44200,N_42004,N_43340);
or U44201 (N_44201,N_42359,N_43827);
and U44202 (N_44202,N_42195,N_42973);
and U44203 (N_44203,N_42426,N_42342);
or U44204 (N_44204,N_43466,N_42638);
nor U44205 (N_44205,N_42322,N_42238);
or U44206 (N_44206,N_43165,N_43160);
and U44207 (N_44207,N_43945,N_43328);
and U44208 (N_44208,N_43076,N_43587);
and U44209 (N_44209,N_42498,N_43633);
or U44210 (N_44210,N_42704,N_43768);
or U44211 (N_44211,N_42719,N_43096);
nor U44212 (N_44212,N_42258,N_43550);
and U44213 (N_44213,N_43614,N_43465);
and U44214 (N_44214,N_42977,N_43840);
or U44215 (N_44215,N_42935,N_43649);
nand U44216 (N_44216,N_43559,N_42766);
and U44217 (N_44217,N_42318,N_43125);
nand U44218 (N_44218,N_43420,N_42187);
nand U44219 (N_44219,N_43446,N_42775);
or U44220 (N_44220,N_42807,N_43650);
nand U44221 (N_44221,N_43513,N_43000);
nand U44222 (N_44222,N_42675,N_42491);
nand U44223 (N_44223,N_42030,N_42965);
or U44224 (N_44224,N_42101,N_42556);
nor U44225 (N_44225,N_42152,N_43225);
nor U44226 (N_44226,N_43891,N_42627);
or U44227 (N_44227,N_42909,N_43822);
nor U44228 (N_44228,N_42164,N_42940);
and U44229 (N_44229,N_42082,N_42076);
or U44230 (N_44230,N_43064,N_43671);
xor U44231 (N_44231,N_43333,N_43301);
nand U44232 (N_44232,N_43194,N_43478);
nand U44233 (N_44233,N_42302,N_43634);
or U44234 (N_44234,N_43952,N_43490);
nand U44235 (N_44235,N_43600,N_42901);
or U44236 (N_44236,N_42020,N_43126);
or U44237 (N_44237,N_43683,N_43159);
nand U44238 (N_44238,N_43601,N_43721);
or U44239 (N_44239,N_43001,N_43162);
nand U44240 (N_44240,N_43882,N_43023);
and U44241 (N_44241,N_42270,N_43188);
and U44242 (N_44242,N_43706,N_42113);
nand U44243 (N_44243,N_43419,N_42237);
or U44244 (N_44244,N_42231,N_43141);
and U44245 (N_44245,N_42699,N_43758);
nand U44246 (N_44246,N_43382,N_42182);
nor U44247 (N_44247,N_43499,N_42444);
and U44248 (N_44248,N_43909,N_43787);
and U44249 (N_44249,N_42742,N_43699);
nor U44250 (N_44250,N_42903,N_43806);
or U44251 (N_44251,N_43562,N_42034);
xor U44252 (N_44252,N_42319,N_42112);
nand U44253 (N_44253,N_43691,N_43034);
or U44254 (N_44254,N_43013,N_43501);
nand U44255 (N_44255,N_42725,N_43667);
or U44256 (N_44256,N_42469,N_42862);
nand U44257 (N_44257,N_42914,N_43366);
or U44258 (N_44258,N_42415,N_42733);
or U44259 (N_44259,N_42186,N_42692);
and U44260 (N_44260,N_42858,N_42681);
or U44261 (N_44261,N_42622,N_42026);
nand U44262 (N_44262,N_43555,N_43078);
nand U44263 (N_44263,N_43765,N_43440);
nand U44264 (N_44264,N_43546,N_42260);
nor U44265 (N_44265,N_43152,N_43083);
or U44266 (N_44266,N_42133,N_42199);
nand U44267 (N_44267,N_42212,N_42827);
nand U44268 (N_44268,N_43962,N_42344);
and U44269 (N_44269,N_43417,N_42951);
and U44270 (N_44270,N_43924,N_42028);
nor U44271 (N_44271,N_43397,N_42656);
or U44272 (N_44272,N_42526,N_43042);
or U44273 (N_44273,N_43515,N_43387);
nand U44274 (N_44274,N_43666,N_42430);
and U44275 (N_44275,N_42868,N_43748);
or U44276 (N_44276,N_42981,N_42824);
or U44277 (N_44277,N_42217,N_43762);
or U44278 (N_44278,N_43895,N_42851);
nor U44279 (N_44279,N_42277,N_43318);
or U44280 (N_44280,N_43939,N_42869);
nor U44281 (N_44281,N_43925,N_43834);
and U44282 (N_44282,N_43365,N_42966);
and U44283 (N_44283,N_42061,N_43747);
nor U44284 (N_44284,N_43056,N_43517);
and U44285 (N_44285,N_43264,N_43422);
nor U44286 (N_44286,N_42728,N_43617);
xnor U44287 (N_44287,N_43166,N_43224);
nand U44288 (N_44288,N_43099,N_43837);
or U44289 (N_44289,N_42852,N_42024);
and U44290 (N_44290,N_42335,N_43690);
nand U44291 (N_44291,N_42476,N_43004);
or U44292 (N_44292,N_42016,N_43557);
and U44293 (N_44293,N_42583,N_43657);
or U44294 (N_44294,N_43974,N_43838);
nor U44295 (N_44295,N_43714,N_42848);
xor U44296 (N_44296,N_43075,N_42105);
and U44297 (N_44297,N_43751,N_43638);
nor U44298 (N_44298,N_42730,N_42354);
nor U44299 (N_44299,N_42641,N_43903);
and U44300 (N_44300,N_42445,N_43233);
or U44301 (N_44301,N_43934,N_42381);
nand U44302 (N_44302,N_43835,N_43852);
and U44303 (N_44303,N_43901,N_43190);
nand U44304 (N_44304,N_42508,N_43629);
nand U44305 (N_44305,N_43969,N_43112);
nor U44306 (N_44306,N_43681,N_43791);
nand U44307 (N_44307,N_43003,N_42495);
nor U44308 (N_44308,N_43566,N_43870);
nor U44309 (N_44309,N_43910,N_42363);
and U44310 (N_44310,N_43329,N_43050);
nand U44311 (N_44311,N_43022,N_43571);
nand U44312 (N_44312,N_42679,N_43520);
or U44313 (N_44313,N_42285,N_42325);
or U44314 (N_44314,N_43883,N_42442);
or U44315 (N_44315,N_42613,N_43733);
or U44316 (N_44316,N_42575,N_43805);
nand U44317 (N_44317,N_43624,N_42573);
or U44318 (N_44318,N_43729,N_42433);
and U44319 (N_44319,N_43359,N_43935);
nand U44320 (N_44320,N_42537,N_42120);
and U44321 (N_44321,N_42740,N_43316);
xor U44322 (N_44322,N_42298,N_43932);
nand U44323 (N_44323,N_42682,N_43235);
nor U44324 (N_44324,N_42056,N_42449);
nor U44325 (N_44325,N_43709,N_43139);
nor U44326 (N_44326,N_43588,N_43203);
or U44327 (N_44327,N_43635,N_43381);
nor U44328 (N_44328,N_42214,N_42015);
and U44329 (N_44329,N_42247,N_42751);
nand U44330 (N_44330,N_42336,N_42821);
nor U44331 (N_44331,N_43947,N_42753);
and U44332 (N_44332,N_42017,N_43766);
nand U44333 (N_44333,N_42773,N_43375);
nand U44334 (N_44334,N_42855,N_42208);
and U44335 (N_44335,N_42374,N_42628);
xor U44336 (N_44336,N_43987,N_43157);
nand U44337 (N_44337,N_43198,N_42099);
or U44338 (N_44338,N_43102,N_43979);
nand U44339 (N_44339,N_43345,N_42047);
nand U44340 (N_44340,N_42203,N_42108);
nor U44341 (N_44341,N_42604,N_42837);
nand U44342 (N_44342,N_42646,N_43209);
nor U44343 (N_44343,N_43362,N_43350);
nand U44344 (N_44344,N_42448,N_42249);
or U44345 (N_44345,N_42364,N_42922);
nor U44346 (N_44346,N_43084,N_42576);
or U44347 (N_44347,N_42011,N_42454);
or U44348 (N_44348,N_43663,N_43137);
nor U44349 (N_44349,N_43689,N_43059);
nand U44350 (N_44350,N_42624,N_43997);
or U44351 (N_44351,N_42864,N_42988);
xor U44352 (N_44352,N_43857,N_42462);
or U44353 (N_44353,N_42170,N_43792);
and U44354 (N_44354,N_43563,N_42052);
nand U44355 (N_44355,N_42771,N_43608);
nand U44356 (N_44356,N_42455,N_42643);
and U44357 (N_44357,N_42118,N_43985);
nand U44358 (N_44358,N_43058,N_42494);
or U44359 (N_44359,N_43428,N_43841);
or U44360 (N_44360,N_42370,N_42987);
nand U44361 (N_44361,N_42230,N_42096);
or U44362 (N_44362,N_43282,N_43642);
or U44363 (N_44363,N_43242,N_42601);
nand U44364 (N_44364,N_43408,N_43539);
or U44365 (N_44365,N_42799,N_42674);
nand U44366 (N_44366,N_42143,N_43711);
nand U44367 (N_44367,N_42872,N_43383);
nor U44368 (N_44368,N_42933,N_42023);
nor U44369 (N_44369,N_43388,N_43319);
nor U44370 (N_44370,N_42599,N_43216);
nand U44371 (N_44371,N_43904,N_42691);
nand U44372 (N_44372,N_43580,N_42042);
nor U44373 (N_44373,N_43764,N_43469);
and U44374 (N_44374,N_42390,N_42867);
nor U44375 (N_44375,N_42846,N_42360);
nand U44376 (N_44376,N_42447,N_42464);
nor U44377 (N_44377,N_43286,N_42582);
or U44378 (N_44378,N_42057,N_42304);
or U44379 (N_44379,N_42155,N_42064);
nor U44380 (N_44380,N_43291,N_42985);
and U44381 (N_44381,N_42281,N_42459);
xnor U44382 (N_44382,N_43263,N_43222);
nand U44383 (N_44383,N_42489,N_42574);
nor U44384 (N_44384,N_43973,N_42653);
and U44385 (N_44385,N_43296,N_42693);
and U44386 (N_44386,N_42587,N_43950);
and U44387 (N_44387,N_42468,N_42589);
and U44388 (N_44388,N_42003,N_43254);
nand U44389 (N_44389,N_43492,N_43989);
nor U44390 (N_44390,N_42892,N_42553);
nand U44391 (N_44391,N_42979,N_43432);
nand U44392 (N_44392,N_42254,N_43770);
and U44393 (N_44393,N_42223,N_42006);
and U44394 (N_44394,N_42437,N_42993);
and U44395 (N_44395,N_43337,N_42896);
nor U44396 (N_44396,N_43237,N_43292);
nor U44397 (N_44397,N_42456,N_42768);
or U44398 (N_44398,N_43817,N_42046);
nand U44399 (N_44399,N_43467,N_43245);
xnor U44400 (N_44400,N_43140,N_42856);
or U44401 (N_44401,N_43037,N_43844);
or U44402 (N_44402,N_43406,N_42497);
nor U44403 (N_44403,N_43993,N_42712);
or U44404 (N_44404,N_42194,N_43472);
and U44405 (N_44405,N_42136,N_43953);
and U44406 (N_44406,N_43436,N_42368);
nand U44407 (N_44407,N_43583,N_42326);
nand U44408 (N_44408,N_42451,N_43705);
or U44409 (N_44409,N_42332,N_42525);
or U44410 (N_44410,N_43876,N_43485);
nor U44411 (N_44411,N_43670,N_43832);
nand U44412 (N_44412,N_42165,N_42547);
nor U44413 (N_44413,N_42772,N_43839);
xnor U44414 (N_44414,N_42107,N_42407);
nor U44415 (N_44415,N_43739,N_42347);
nor U44416 (N_44416,N_42372,N_42233);
nor U44417 (N_44417,N_42320,N_42022);
nand U44418 (N_44418,N_42995,N_42724);
nor U44419 (N_44419,N_43201,N_42478);
or U44420 (N_44420,N_42731,N_43694);
or U44421 (N_44421,N_43153,N_42228);
nand U44422 (N_44422,N_43644,N_42470);
and U44423 (N_44423,N_42816,N_43518);
nor U44424 (N_44424,N_43453,N_43405);
nand U44425 (N_44425,N_42752,N_42308);
and U44426 (N_44426,N_43674,N_43712);
nor U44427 (N_44427,N_42403,N_42252);
or U44428 (N_44428,N_43065,N_42466);
nand U44429 (N_44429,N_43621,N_43554);
nor U44430 (N_44430,N_43534,N_42767);
nand U44431 (N_44431,N_42190,N_42748);
or U44432 (N_44432,N_43980,N_42275);
and U44433 (N_44433,N_43977,N_43703);
nor U44434 (N_44434,N_43848,N_43100);
nor U44435 (N_44435,N_43085,N_42427);
and U44436 (N_44436,N_43109,N_43106);
nand U44437 (N_44437,N_43743,N_43113);
nand U44438 (N_44438,N_43135,N_42566);
nand U44439 (N_44439,N_43470,N_43726);
or U44440 (N_44440,N_43682,N_43793);
or U44441 (N_44441,N_43868,N_43875);
or U44442 (N_44442,N_43871,N_42196);
xor U44443 (N_44443,N_42761,N_42774);
and U44444 (N_44444,N_42804,N_42915);
and U44445 (N_44445,N_42272,N_43307);
nor U44446 (N_44446,N_43176,N_43459);
and U44447 (N_44447,N_43483,N_43312);
nor U44448 (N_44448,N_42565,N_43813);
and U44449 (N_44449,N_43391,N_43527);
and U44450 (N_44450,N_43578,N_43071);
nor U44451 (N_44451,N_43168,N_43881);
nor U44452 (N_44452,N_43314,N_42197);
or U44453 (N_44453,N_42480,N_42134);
or U44454 (N_44454,N_43158,N_43494);
nand U44455 (N_44455,N_43169,N_43779);
or U44456 (N_44456,N_42943,N_42103);
nor U44457 (N_44457,N_42135,N_42649);
nand U44458 (N_44458,N_43618,N_42978);
or U44459 (N_44459,N_43247,N_43258);
nor U44460 (N_44460,N_42038,N_42661);
or U44461 (N_44461,N_43368,N_42358);
or U44462 (N_44462,N_42817,N_42632);
and U44463 (N_44463,N_43294,N_43731);
or U44464 (N_44464,N_43595,N_43035);
nor U44465 (N_44465,N_43346,N_43567);
and U44466 (N_44466,N_43259,N_42923);
nand U44467 (N_44467,N_42597,N_42756);
or U44468 (N_44468,N_42406,N_43918);
nand U44469 (N_44469,N_43181,N_43048);
and U44470 (N_44470,N_42614,N_42414);
or U44471 (N_44471,N_43606,N_42833);
and U44472 (N_44472,N_42792,N_42013);
nor U44473 (N_44473,N_43218,N_43236);
and U44474 (N_44474,N_43045,N_42215);
and U44475 (N_44475,N_43107,N_43167);
and U44476 (N_44476,N_43028,N_42777);
nor U44477 (N_44477,N_42736,N_42592);
or U44478 (N_44478,N_43274,N_42202);
or U44479 (N_44479,N_43077,N_42314);
nor U44480 (N_44480,N_42316,N_43310);
and U44481 (N_44481,N_43700,N_43880);
or U44482 (N_44482,N_43630,N_43343);
nor U44483 (N_44483,N_42924,N_42972);
nor U44484 (N_44484,N_43842,N_42121);
or U44485 (N_44485,N_43653,N_42671);
and U44486 (N_44486,N_42808,N_43632);
nor U44487 (N_44487,N_43613,N_43308);
nor U44488 (N_44488,N_43309,N_43664);
and U44489 (N_44489,N_42702,N_42204);
or U44490 (N_44490,N_42416,N_42411);
nor U44491 (N_44491,N_42408,N_43786);
or U44492 (N_44492,N_43728,N_42953);
nor U44493 (N_44493,N_43067,N_43986);
or U44494 (N_44494,N_43576,N_42763);
nand U44495 (N_44495,N_43623,N_43171);
nor U44496 (N_44496,N_42181,N_42564);
nor U44497 (N_44497,N_43755,N_42685);
nand U44498 (N_44498,N_42645,N_43206);
nand U44499 (N_44499,N_43105,N_42404);
nand U44500 (N_44500,N_42324,N_43763);
nor U44501 (N_44501,N_42602,N_43146);
nand U44502 (N_44502,N_43799,N_42044);
nor U44503 (N_44503,N_42309,N_42800);
or U44504 (N_44504,N_43574,N_42168);
and U44505 (N_44505,N_43032,N_43138);
and U44506 (N_44506,N_43859,N_43774);
nor U44507 (N_44507,N_43121,N_42994);
or U44508 (N_44508,N_43404,N_43131);
and U44509 (N_44509,N_43482,N_43097);
nand U44510 (N_44510,N_42708,N_42588);
or U44511 (N_44511,N_42299,N_42687);
or U44512 (N_44512,N_42567,N_42474);
and U44513 (N_44513,N_42337,N_43493);
nor U44514 (N_44514,N_42192,N_42209);
xnor U44515 (N_44515,N_42422,N_42144);
nand U44516 (N_44516,N_42788,N_42269);
and U44517 (N_44517,N_43861,N_42747);
nand U44518 (N_44518,N_43458,N_42292);
nand U44519 (N_44519,N_42394,N_42585);
or U44520 (N_44520,N_43536,N_43266);
and U44521 (N_44521,N_42089,N_42384);
or U44522 (N_44522,N_42174,N_43489);
or U44523 (N_44523,N_42603,N_42321);
nand U44524 (N_44524,N_43017,N_43134);
and U44525 (N_44525,N_42059,N_42255);
and U44526 (N_44526,N_43702,N_43199);
xnor U44527 (N_44527,N_43229,N_43599);
nor U44528 (N_44528,N_43545,N_43115);
or U44529 (N_44529,N_43889,N_42009);
and U44530 (N_44530,N_43775,N_43284);
and U44531 (N_44531,N_42916,N_43790);
and U44532 (N_44532,N_42388,N_42631);
and U44533 (N_44533,N_42863,N_42907);
nor U44534 (N_44534,N_42580,N_43760);
or U44535 (N_44535,N_43377,N_43185);
nand U44536 (N_44536,N_43976,N_43631);
and U44537 (N_44537,N_42783,N_43556);
nor U44538 (N_44538,N_42770,N_42162);
or U44539 (N_44539,N_42874,N_42032);
and U44540 (N_44540,N_42323,N_42939);
and U44541 (N_44541,N_42402,N_43966);
nand U44542 (N_44542,N_43652,N_43290);
nor U44543 (N_44543,N_43685,N_43523);
and U44544 (N_44544,N_43495,N_42446);
and U44545 (N_44545,N_42440,N_43030);
or U44546 (N_44546,N_42584,N_43155);
nand U44547 (N_44547,N_43416,N_42412);
nand U44548 (N_44548,N_43234,N_43961);
or U44549 (N_44549,N_43884,N_43648);
nor U44550 (N_44550,N_42450,N_43992);
nand U44551 (N_44551,N_43193,N_43798);
nand U44552 (N_44552,N_43607,N_43352);
and U44553 (N_44553,N_42484,N_42895);
nor U44554 (N_44554,N_42471,N_42142);
nor U44555 (N_44555,N_43243,N_43676);
or U44556 (N_44556,N_42941,N_43794);
or U44557 (N_44557,N_43455,N_42590);
and U44558 (N_44558,N_43951,N_42303);
and U44559 (N_44559,N_43399,N_43864);
or U44560 (N_44560,N_43044,N_43912);
and U44561 (N_44561,N_43887,N_43800);
nor U44562 (N_44562,N_42927,N_43476);
and U44563 (N_44563,N_42608,N_42352);
nor U44564 (N_44564,N_42832,N_42743);
or U44565 (N_44565,N_42362,N_42180);
and U44566 (N_44566,N_42496,N_42033);
nor U44567 (N_44567,N_42791,N_42902);
nor U44568 (N_44568,N_43704,N_43287);
and U44569 (N_44569,N_43143,N_43847);
or U44570 (N_44570,N_43830,N_42936);
and U44571 (N_44571,N_42244,N_42288);
nor U44572 (N_44572,N_43205,N_42279);
nor U44573 (N_44573,N_42971,N_42148);
and U44574 (N_44574,N_43920,N_42071);
nand U44575 (N_44575,N_42184,N_42560);
nor U44576 (N_44576,N_42669,N_43269);
nor U44577 (N_44577,N_42956,N_43238);
nand U44578 (N_44578,N_42950,N_42605);
nor U44579 (N_44579,N_42389,N_43507);
and U44580 (N_44580,N_42479,N_42906);
xor U44581 (N_44581,N_42500,N_42522);
nand U44582 (N_44582,N_43349,N_43293);
nand U44583 (N_44583,N_43771,N_42501);
or U44584 (N_44584,N_42265,N_42420);
nor U44585 (N_44585,N_42718,N_43968);
nor U44586 (N_44586,N_43150,N_43561);
and U44587 (N_44587,N_42734,N_42251);
and U44588 (N_44588,N_43122,N_42723);
nand U44589 (N_44589,N_43687,N_42274);
nor U44590 (N_44590,N_43376,N_42172);
nand U44591 (N_44591,N_42018,N_42328);
and U44592 (N_44592,N_42234,N_43256);
or U44593 (N_44593,N_43544,N_43311);
or U44594 (N_44594,N_43991,N_42610);
nor U44595 (N_44595,N_43514,N_43900);
or U44596 (N_44596,N_43641,N_43724);
or U44597 (N_44597,N_43221,N_42831);
and U44598 (N_44598,N_43592,N_43080);
nor U44599 (N_44599,N_43244,N_42739);
nor U44600 (N_44600,N_42886,N_42129);
nand U44601 (N_44601,N_42409,N_42559);
nand U44602 (N_44602,N_43327,N_42917);
nand U44603 (N_44603,N_43701,N_42116);
nand U44604 (N_44604,N_42853,N_43815);
or U44605 (N_44605,N_43526,N_42930);
or U44606 (N_44606,N_43410,N_42183);
or U44607 (N_44607,N_42472,N_43906);
and U44608 (N_44608,N_43355,N_43360);
nand U44609 (N_44609,N_42296,N_43651);
or U44610 (N_44610,N_43371,N_43537);
nor U44611 (N_44611,N_42493,N_43390);
nand U44612 (N_44612,N_43038,N_42378);
nand U44613 (N_44613,N_43826,N_42518);
nand U44614 (N_44614,N_42765,N_42778);
or U44615 (N_44615,N_43480,N_42812);
xnor U44616 (N_44616,N_42769,N_43132);
and U44617 (N_44617,N_42934,N_43855);
nand U44618 (N_44618,N_42084,N_43491);
or U44619 (N_44619,N_43596,N_43801);
nand U44620 (N_44620,N_43270,N_43435);
nor U44621 (N_44621,N_43591,N_42957);
or U44622 (N_44622,N_42680,N_43332);
and U44623 (N_44623,N_42776,N_42568);
nor U44624 (N_44624,N_43054,N_43611);
and U44625 (N_44625,N_42178,N_43784);
nor U44626 (N_44626,N_43280,N_43091);
or U44627 (N_44627,N_43025,N_43315);
and U44628 (N_44628,N_43820,N_42571);
or U44629 (N_44629,N_43431,N_43052);
nor U44630 (N_44630,N_42087,N_43089);
nor U44631 (N_44631,N_43402,N_43177);
or U44632 (N_44632,N_43886,N_42920);
and U44633 (N_44633,N_43956,N_42505);
nand U44634 (N_44634,N_43916,N_43610);
nor U44635 (N_44635,N_42879,N_42485);
nand U44636 (N_44636,N_43718,N_43757);
nand U44637 (N_44637,N_43439,N_42779);
nand U44638 (N_44638,N_42947,N_43811);
nand U44639 (N_44639,N_43738,N_42147);
or U44640 (N_44640,N_43220,N_43379);
or U44641 (N_44641,N_43593,N_43819);
nor U44642 (N_44642,N_43570,N_42081);
or U44643 (N_44643,N_43488,N_42650);
nor U44644 (N_44644,N_43750,N_43836);
nand U44645 (N_44645,N_43214,N_42040);
or U44646 (N_44646,N_43358,N_43372);
or U44647 (N_44647,N_43767,N_43456);
and U44648 (N_44648,N_43878,N_43862);
and U44649 (N_44649,N_43516,N_43015);
or U44650 (N_44650,N_43060,N_42701);
nand U44651 (N_44651,N_42881,N_42744);
and U44652 (N_44652,N_42758,N_43447);
nor U44653 (N_44653,N_43451,N_43616);
nand U44654 (N_44654,N_43299,N_43584);
nor U44655 (N_44655,N_42514,N_43914);
or U44656 (N_44656,N_43860,N_43049);
xor U44657 (N_44657,N_42552,N_43785);
xor U44658 (N_44658,N_43248,N_42540);
xnor U44659 (N_44659,N_42151,N_42339);
or U44660 (N_44660,N_43856,N_43645);
or U44661 (N_44661,N_42606,N_43615);
or U44662 (N_44662,N_42888,N_42657);
xor U44663 (N_44663,N_43341,N_43304);
or U44664 (N_44664,N_42213,N_43073);
or U44665 (N_44665,N_42790,N_43708);
or U44666 (N_44666,N_43324,N_42519);
nor U44667 (N_44667,N_43619,N_42958);
nor U44668 (N_44668,N_42224,N_43154);
and U44669 (N_44669,N_43737,N_42569);
nand U44670 (N_44670,N_43602,N_42461);
nor U44671 (N_44671,N_42434,N_42283);
nor U44672 (N_44672,N_42175,N_42884);
nand U44673 (N_44673,N_42696,N_42520);
and U44674 (N_44674,N_43380,N_43581);
or U44675 (N_44675,N_42173,N_42579);
nor U44676 (N_44676,N_42486,N_42021);
nand U44677 (N_44677,N_42300,N_43251);
nor U44678 (N_44678,N_42598,N_43389);
and U44679 (N_44679,N_43873,N_43257);
and U44680 (N_44680,N_42069,N_43344);
nor U44681 (N_44681,N_42637,N_43722);
and U44682 (N_44682,N_42035,N_43018);
or U44683 (N_44683,N_43524,N_43752);
nand U44684 (N_44684,N_42897,N_43780);
nand U44685 (N_44685,N_42938,N_43978);
nor U44686 (N_44686,N_43462,N_42860);
or U44687 (N_44687,N_42713,N_42659);
and U44688 (N_44688,N_42253,N_42210);
and U44689 (N_44689,N_42114,N_43240);
nor U44690 (N_44690,N_42400,N_42550);
nor U44691 (N_44691,N_42854,N_43306);
and U44692 (N_44692,N_42822,N_43528);
nor U44693 (N_44693,N_42429,N_42391);
nand U44694 (N_44694,N_42528,N_42722);
or U44695 (N_44695,N_42357,N_42960);
nand U44696 (N_44696,N_43843,N_42545);
xnor U44697 (N_44697,N_43275,N_43877);
nand U44698 (N_44698,N_43637,N_42343);
nand U44699 (N_44699,N_42664,N_43086);
or U44700 (N_44700,N_42786,N_42554);
nor U44701 (N_44701,N_43831,N_43069);
nand U44702 (N_44702,N_43568,N_43129);
or U44703 (N_44703,N_42509,N_42235);
nand U44704 (N_44704,N_43090,N_43929);
nor U44705 (N_44705,N_43897,N_43016);
and U44706 (N_44706,N_42980,N_42787);
nor U44707 (N_44707,N_42755,N_42964);
and U44708 (N_44708,N_42615,N_42413);
nor U44709 (N_44709,N_43998,N_43305);
or U44710 (N_44710,N_42720,N_42507);
and U44711 (N_44711,N_42310,N_42205);
or U44712 (N_44712,N_43173,N_42460);
nand U44713 (N_44713,N_42054,N_42989);
xnor U44714 (N_44714,N_42395,N_42132);
nand U44715 (N_44715,N_42104,N_43707);
and U44716 (N_44716,N_42527,N_42672);
nor U44717 (N_44717,N_42834,N_42452);
or U44718 (N_44718,N_43223,N_43646);
and U44719 (N_44719,N_43212,N_42160);
nand U44720 (N_44720,N_42741,N_42263);
or U44721 (N_44721,N_42385,N_43342);
xor U44722 (N_44722,N_42246,N_42060);
nor U44723 (N_44723,N_43373,N_43429);
or U44724 (N_44724,N_43603,N_43885);
xnor U44725 (N_44725,N_43326,N_43074);
or U44726 (N_44726,N_42088,N_42557);
and U44727 (N_44727,N_43680,N_43662);
nand U44728 (N_44728,N_42154,N_42663);
nor U44729 (N_44729,N_43120,N_42273);
xor U44730 (N_44730,N_42595,N_43114);
or U44731 (N_44731,N_43108,N_43128);
nand U44732 (N_44732,N_43363,N_43696);
nand U44733 (N_44733,N_42976,N_43449);
and U44734 (N_44734,N_42365,N_43905);
or U44735 (N_44735,N_42757,N_43677);
nand U44736 (N_44736,N_43776,N_42477);
or U44737 (N_44737,N_42937,N_43144);
nand U44738 (N_44738,N_42268,N_43123);
nand U44739 (N_44739,N_42421,N_43027);
and U44740 (N_44740,N_42428,N_42431);
and U44741 (N_44741,N_43955,N_43055);
nand U44742 (N_44742,N_43418,N_42539);
nor U44743 (N_44743,N_42695,N_43111);
or U44744 (N_44744,N_43783,N_43803);
nand U44745 (N_44745,N_43197,N_43797);
and U44746 (N_44746,N_42079,N_42694);
and U44747 (N_44747,N_43441,N_42836);
nand U44748 (N_44748,N_43741,N_42710);
or U44749 (N_44749,N_42555,N_43401);
and U44750 (N_44750,N_43040,N_43031);
or U44751 (N_44751,N_42313,N_42331);
or U44752 (N_44752,N_43070,N_43262);
or U44753 (N_44753,N_42443,N_42441);
nand U44754 (N_44754,N_42536,N_43719);
nor U44755 (N_44755,N_43734,N_43092);
or U44756 (N_44756,N_42521,N_43660);
and U44757 (N_44757,N_43879,N_42236);
nor U44758 (N_44758,N_43622,N_43858);
nor U44759 (N_44759,N_42882,N_42207);
nor U44760 (N_44760,N_43872,N_43890);
nand U44761 (N_44761,N_43230,N_42286);
nor U44762 (N_44762,N_42908,N_43744);
nor U44763 (N_44763,N_43116,N_43468);
nor U44764 (N_44764,N_42801,N_43921);
xor U44765 (N_44765,N_42386,N_43940);
and U44766 (N_44766,N_43497,N_43655);
and U44767 (N_44767,N_42334,N_42841);
or U44768 (N_44768,N_42984,N_43033);
nand U44769 (N_44769,N_42503,N_42670);
nor U44770 (N_44770,N_42795,N_42435);
nor U44771 (N_44771,N_42952,N_43239);
nor U44772 (N_44772,N_42954,N_42640);
nand U44773 (N_44773,N_42191,N_42140);
and U44774 (N_44774,N_42366,N_42932);
and U44775 (N_44775,N_42077,N_42665);
xnor U44776 (N_44776,N_42839,N_42068);
xnor U44777 (N_44777,N_43437,N_43936);
nand U44778 (N_44778,N_43522,N_42802);
or U44779 (N_44779,N_42843,N_42762);
and U44780 (N_44780,N_42899,N_42425);
and U44781 (N_44781,N_42423,N_42667);
xnor U44782 (N_44782,N_42893,N_43321);
nand U44783 (N_44783,N_42007,N_43818);
and U44784 (N_44784,N_42609,N_43725);
nor U44785 (N_44785,N_43175,N_42262);
or U44786 (N_44786,N_43127,N_43104);
and U44787 (N_44787,N_43187,N_42179);
xnor U44788 (N_44788,N_42655,N_42072);
or U44789 (N_44789,N_43179,N_43302);
or U44790 (N_44790,N_42066,N_42218);
and U44791 (N_44791,N_43907,N_42703);
and U44792 (N_44792,N_42845,N_42239);
and U44793 (N_44793,N_43103,N_43915);
nand U44794 (N_44794,N_43192,N_42974);
nor U44795 (N_44795,N_43943,N_43423);
nand U44796 (N_44796,N_42607,N_43395);
or U44797 (N_44797,N_42127,N_43136);
xor U44798 (N_44798,N_42745,N_42232);
and U44799 (N_44799,N_42341,N_43896);
or U44800 (N_44800,N_43777,N_43990);
xor U44801 (N_44801,N_43094,N_43370);
nor U44802 (N_44802,N_42634,N_43249);
nand U44803 (N_44803,N_42031,N_42294);
or U44804 (N_44804,N_42900,N_43604);
nand U44805 (N_44805,N_42662,N_43828);
or U44806 (N_44806,N_42481,N_43053);
nand U44807 (N_44807,N_42153,N_43782);
nor U44808 (N_44808,N_42073,N_43854);
nand U44809 (N_44809,N_42245,N_43821);
or U44810 (N_44810,N_43781,N_43983);
nor U44811 (N_44811,N_43019,N_42626);
nand U44812 (N_44812,N_42463,N_43043);
nand U44813 (N_44813,N_42794,N_43911);
nor U44814 (N_44814,N_42535,N_43590);
and U44815 (N_44815,N_42305,N_42549);
nand U44816 (N_44816,N_42750,N_42538);
nor U44817 (N_44817,N_43392,N_43208);
and U44818 (N_44818,N_43511,N_42955);
nand U44819 (N_44819,N_42873,N_42658);
and U44820 (N_44820,N_42931,N_43093);
and U44821 (N_44821,N_42690,N_43335);
and U44822 (N_44822,N_43323,N_42968);
nor U44823 (N_44823,N_43533,N_43331);
nand U44824 (N_44824,N_43926,N_42842);
or U44825 (N_44825,N_42312,N_42975);
or U44826 (N_44826,N_43710,N_42572);
nand U44827 (N_44827,N_43573,N_43189);
and U44828 (N_44828,N_43265,N_43475);
and U44829 (N_44829,N_42340,N_43353);
or U44830 (N_44830,N_42533,N_43356);
nor U44831 (N_44831,N_43450,N_43594);
nor U44832 (N_44832,N_42515,N_43147);
nand U44833 (N_44833,N_42137,N_43322);
or U44834 (N_44834,N_43231,N_43403);
nor U44835 (N_44835,N_42828,N_42293);
and U44836 (N_44836,N_42158,N_42946);
or U44837 (N_44837,N_42128,N_42629);
and U44838 (N_44838,N_43464,N_42271);
nand U44839 (N_44839,N_42516,N_43715);
and U44840 (N_44840,N_42051,N_43802);
and U44841 (N_44841,N_42992,N_42840);
nor U44842 (N_44842,N_42000,N_42591);
or U44843 (N_44843,N_42167,N_43498);
or U44844 (N_44844,N_42329,N_43448);
nor U44845 (N_44845,N_42642,N_42809);
and U44846 (N_44846,N_42094,N_43720);
nand U44847 (N_44847,N_43427,N_42405);
nor U44848 (N_44848,N_42145,N_42706);
and U44849 (N_44849,N_42697,N_42291);
and U44850 (N_44850,N_42921,N_42243);
nor U44851 (N_44851,N_43688,N_42225);
and U44852 (N_44852,N_43605,N_43261);
or U44853 (N_44853,N_43421,N_43036);
xnor U44854 (N_44854,N_43061,N_43273);
or U44855 (N_44855,N_42297,N_43317);
and U44856 (N_44856,N_43627,N_42991);
nor U44857 (N_44857,N_43938,N_43272);
nand U44858 (N_44858,N_43542,N_43057);
and U44859 (N_44859,N_43087,N_43999);
nor U44860 (N_44860,N_43949,N_43553);
nor U44861 (N_44861,N_42048,N_42261);
and U44862 (N_44862,N_42705,N_42820);
nor U44863 (N_44863,N_42109,N_43207);
or U44864 (N_44864,N_42611,N_43268);
and U44865 (N_44865,N_42749,N_43669);
and U44866 (N_44866,N_43552,N_43716);
and U44867 (N_44867,N_42457,N_43213);
and U44868 (N_44868,N_43928,N_42709);
or U44869 (N_44869,N_43756,N_43101);
nor U44870 (N_44870,N_42998,N_43908);
or U44871 (N_44871,N_43893,N_42711);
or U44872 (N_44872,N_43519,N_42222);
nor U44873 (N_44873,N_43548,N_42008);
nor U44874 (N_44874,N_42677,N_43267);
or U44875 (N_44875,N_43481,N_43927);
nor U44876 (N_44876,N_42070,N_43007);
or U44877 (N_44877,N_43348,N_43479);
or U44878 (N_44878,N_43796,N_42067);
nor U44879 (N_44879,N_42131,N_42894);
nor U44880 (N_44880,N_43098,N_43582);
nand U44881 (N_44881,N_43414,N_42163);
nand U44882 (N_44882,N_42982,N_42544);
nand U44883 (N_44883,N_43942,N_43219);
and U44884 (N_44884,N_43930,N_42410);
nand U44885 (N_44885,N_43210,N_43759);
or U44886 (N_44886,N_43215,N_43396);
or U44887 (N_44887,N_42620,N_43002);
or U44888 (N_44888,N_43509,N_42499);
nand U44889 (N_44889,N_43964,N_42815);
or U44890 (N_44890,N_42689,N_43276);
nand U44891 (N_44891,N_42633,N_42959);
and U44892 (N_44892,N_42780,N_43161);
or U44893 (N_44893,N_42811,N_42092);
nor U44894 (N_44894,N_43804,N_43008);
or U44895 (N_44895,N_43118,N_42200);
nor U44896 (N_44896,N_42256,N_42345);
nor U44897 (N_44897,N_42398,N_43081);
nand U44898 (N_44898,N_42911,N_42041);
and U44899 (N_44899,N_43665,N_42890);
nand U44900 (N_44900,N_42482,N_43579);
or U44901 (N_44901,N_42355,N_42676);
nand U44902 (N_44902,N_43589,N_42166);
and U44903 (N_44903,N_43965,N_43994);
and U44904 (N_44904,N_42353,N_42465);
nand U44905 (N_44905,N_42612,N_42012);
and U44906 (N_44906,N_43386,N_43021);
or U44907 (N_44907,N_42219,N_43693);
nand U44908 (N_44908,N_43899,N_42619);
nand U44909 (N_44909,N_43668,N_43888);
and U44910 (N_44910,N_42967,N_43325);
or U44911 (N_44911,N_42169,N_43487);
nand U44912 (N_44912,N_42823,N_43411);
or U44913 (N_44913,N_42593,N_43425);
nor U44914 (N_44914,N_42875,N_42986);
nand U44915 (N_44915,N_42871,N_43407);
xnor U44916 (N_44916,N_42053,N_42330);
nand U44917 (N_44917,N_42805,N_43846);
and U44918 (N_44918,N_43628,N_42654);
nor U44919 (N_44919,N_43535,N_42803);
nand U44920 (N_44920,N_43625,N_43529);
and U44921 (N_44921,N_43378,N_43996);
nor U44922 (N_44922,N_42735,N_42290);
nand U44923 (N_44923,N_43354,N_43079);
nand U44924 (N_44924,N_43241,N_43303);
nor U44925 (N_44925,N_43944,N_42350);
and U44926 (N_44926,N_42216,N_43941);
nor U44927 (N_44927,N_43082,N_43252);
or U44928 (N_44928,N_43191,N_42229);
nand U44929 (N_44929,N_42125,N_43504);
and U44930 (N_44930,N_43148,N_43736);
nand U44931 (N_44931,N_42487,N_43163);
or U44932 (N_44932,N_43051,N_42333);
nand U44933 (N_44933,N_43460,N_43658);
nand U44934 (N_44934,N_42969,N_43713);
and U44935 (N_44935,N_43538,N_42027);
or U44936 (N_44936,N_42490,N_43636);
nand U44937 (N_44937,N_43130,N_43496);
and U44938 (N_44938,N_43434,N_43278);
nand U44939 (N_44939,N_42226,N_43279);
nor U44940 (N_44940,N_42865,N_42912);
or U44941 (N_44941,N_43142,N_43454);
or U44942 (N_44942,N_43503,N_42100);
nor U44943 (N_44943,N_42797,N_42715);
nand U44944 (N_44944,N_42630,N_43288);
nor U44945 (N_44945,N_43894,N_43772);
or U44946 (N_44946,N_43695,N_43502);
nand U44947 (N_44947,N_42618,N_42850);
nor U44948 (N_44948,N_42189,N_42563);
and U44949 (N_44949,N_42963,N_42814);
or U44950 (N_44950,N_42789,N_43971);
and U44951 (N_44951,N_43184,N_43558);
nor U44952 (N_44952,N_43626,N_43525);
or U44953 (N_44953,N_43769,N_42651);
and U44954 (N_44954,N_42438,N_43678);
or U44955 (N_44955,N_43351,N_43442);
nand U44956 (N_44956,N_43133,N_43661);
xor U44957 (N_44957,N_42684,N_43808);
nand U44958 (N_44958,N_42240,N_43560);
or U44959 (N_44959,N_43255,N_43922);
or U44960 (N_44960,N_43892,N_43773);
or U44961 (N_44961,N_42211,N_43068);
or U44962 (N_44962,N_42250,N_42110);
nor U44963 (N_44963,N_43982,N_42367);
nand U44964 (N_44964,N_42764,N_43204);
nand U44965 (N_44965,N_42577,N_42436);
nor U44966 (N_44966,N_43014,N_42289);
nand U44967 (N_44967,N_43643,N_42798);
or U44968 (N_44968,N_42647,N_42075);
nor U44969 (N_44969,N_43339,N_43963);
nor U44970 (N_44970,N_43869,N_43119);
and U44971 (N_44971,N_43297,N_43330);
or U44972 (N_44972,N_43697,N_43182);
or U44973 (N_44973,N_42065,N_42668);
and U44974 (N_44974,N_42926,N_42376);
nand U44975 (N_44975,N_42513,N_42483);
nand U44976 (N_44976,N_42666,N_42380);
and U44977 (N_44977,N_42830,N_42188);
or U44978 (N_44978,N_43612,N_42849);
nand U44979 (N_44979,N_43412,N_42925);
or U44980 (N_44980,N_43211,N_43972);
nand U44981 (N_44981,N_42401,N_42785);
nand U44982 (N_44982,N_43540,N_42301);
or U44983 (N_44983,N_42558,N_42700);
or U44984 (N_44984,N_42683,N_42796);
or U44985 (N_44985,N_42241,N_43754);
and U44986 (N_44986,N_42961,N_42453);
nand U44987 (N_44987,N_42119,N_42227);
nor U44988 (N_44988,N_42346,N_43946);
and U44989 (N_44989,N_42623,N_43778);
or U44990 (N_44990,N_42928,N_43006);
nand U44991 (N_44991,N_42278,N_43541);
and U44992 (N_44992,N_43967,N_43409);
nor U44993 (N_44993,N_43510,N_43471);
xor U44994 (N_44994,N_43174,N_43957);
nor U44995 (N_44995,N_42999,N_43919);
and U44996 (N_44996,N_42970,N_42361);
or U44997 (N_44997,N_43415,N_43913);
nand U44998 (N_44998,N_42029,N_42149);
and U44999 (N_44999,N_43505,N_42714);
or U45000 (N_45000,N_42278,N_43583);
and U45001 (N_45001,N_43669,N_43374);
or U45002 (N_45002,N_42727,N_42355);
or U45003 (N_45003,N_42897,N_42345);
or U45004 (N_45004,N_43442,N_43715);
xnor U45005 (N_45005,N_43427,N_42724);
or U45006 (N_45006,N_42028,N_43290);
nand U45007 (N_45007,N_43784,N_42664);
or U45008 (N_45008,N_42364,N_42885);
or U45009 (N_45009,N_42187,N_43633);
and U45010 (N_45010,N_43975,N_42274);
nand U45011 (N_45011,N_43466,N_43975);
nand U45012 (N_45012,N_43809,N_42003);
nor U45013 (N_45013,N_43743,N_42855);
and U45014 (N_45014,N_43852,N_42166);
nand U45015 (N_45015,N_43626,N_42606);
or U45016 (N_45016,N_43000,N_42428);
nor U45017 (N_45017,N_42493,N_43961);
and U45018 (N_45018,N_43893,N_42132);
or U45019 (N_45019,N_43111,N_42839);
or U45020 (N_45020,N_42456,N_42825);
nor U45021 (N_45021,N_43047,N_43669);
nand U45022 (N_45022,N_42518,N_42679);
nand U45023 (N_45023,N_42938,N_43483);
nand U45024 (N_45024,N_42059,N_43154);
or U45025 (N_45025,N_43914,N_43482);
nand U45026 (N_45026,N_43733,N_42149);
nor U45027 (N_45027,N_42922,N_42851);
and U45028 (N_45028,N_43191,N_43808);
or U45029 (N_45029,N_42545,N_43687);
and U45030 (N_45030,N_42428,N_42412);
nand U45031 (N_45031,N_42217,N_42074);
nand U45032 (N_45032,N_43286,N_43429);
or U45033 (N_45033,N_43414,N_42700);
and U45034 (N_45034,N_43317,N_42908);
nand U45035 (N_45035,N_42177,N_42906);
nand U45036 (N_45036,N_43875,N_42230);
xor U45037 (N_45037,N_43838,N_43706);
xor U45038 (N_45038,N_42450,N_43723);
nand U45039 (N_45039,N_42089,N_42933);
nand U45040 (N_45040,N_42080,N_42758);
nor U45041 (N_45041,N_42572,N_43081);
and U45042 (N_45042,N_42292,N_43955);
or U45043 (N_45043,N_43178,N_43024);
and U45044 (N_45044,N_42357,N_42412);
and U45045 (N_45045,N_42464,N_42846);
or U45046 (N_45046,N_43806,N_43841);
nor U45047 (N_45047,N_43450,N_42420);
nand U45048 (N_45048,N_43081,N_42186);
nor U45049 (N_45049,N_42963,N_43115);
nor U45050 (N_45050,N_42741,N_42268);
nor U45051 (N_45051,N_43347,N_43236);
and U45052 (N_45052,N_43617,N_42033);
nand U45053 (N_45053,N_42101,N_43499);
and U45054 (N_45054,N_42595,N_43119);
and U45055 (N_45055,N_42225,N_42032);
or U45056 (N_45056,N_42031,N_42957);
nand U45057 (N_45057,N_42546,N_43598);
nor U45058 (N_45058,N_42142,N_43439);
nand U45059 (N_45059,N_42361,N_43449);
and U45060 (N_45060,N_42432,N_43296);
nor U45061 (N_45061,N_42831,N_43379);
or U45062 (N_45062,N_42372,N_43844);
nor U45063 (N_45063,N_42186,N_43638);
or U45064 (N_45064,N_43626,N_42219);
or U45065 (N_45065,N_42089,N_43080);
nor U45066 (N_45066,N_43559,N_43677);
and U45067 (N_45067,N_42443,N_43715);
nor U45068 (N_45068,N_43333,N_42601);
nor U45069 (N_45069,N_42493,N_43511);
nand U45070 (N_45070,N_42759,N_43021);
and U45071 (N_45071,N_43074,N_43475);
or U45072 (N_45072,N_42927,N_42914);
nand U45073 (N_45073,N_43413,N_42889);
nor U45074 (N_45074,N_43607,N_42294);
nand U45075 (N_45075,N_42448,N_43581);
nor U45076 (N_45076,N_43866,N_43061);
nor U45077 (N_45077,N_43121,N_42131);
nand U45078 (N_45078,N_43463,N_43760);
and U45079 (N_45079,N_43721,N_43904);
and U45080 (N_45080,N_42306,N_42455);
and U45081 (N_45081,N_43446,N_42336);
nor U45082 (N_45082,N_43857,N_42055);
or U45083 (N_45083,N_43515,N_42654);
and U45084 (N_45084,N_42162,N_43009);
nand U45085 (N_45085,N_43482,N_43445);
and U45086 (N_45086,N_42040,N_43357);
nand U45087 (N_45087,N_42909,N_43126);
or U45088 (N_45088,N_43638,N_43078);
or U45089 (N_45089,N_42065,N_42057);
or U45090 (N_45090,N_42755,N_43570);
and U45091 (N_45091,N_43091,N_43651);
nand U45092 (N_45092,N_42409,N_42247);
nor U45093 (N_45093,N_42687,N_43499);
and U45094 (N_45094,N_42975,N_43304);
and U45095 (N_45095,N_42054,N_42314);
xor U45096 (N_45096,N_42294,N_42864);
nand U45097 (N_45097,N_43850,N_43581);
and U45098 (N_45098,N_43169,N_43222);
nand U45099 (N_45099,N_43396,N_42763);
or U45100 (N_45100,N_43029,N_43433);
nor U45101 (N_45101,N_42214,N_42407);
or U45102 (N_45102,N_42948,N_42440);
nor U45103 (N_45103,N_42365,N_43211);
and U45104 (N_45104,N_43060,N_42297);
nand U45105 (N_45105,N_42177,N_42351);
nor U45106 (N_45106,N_42722,N_43277);
nand U45107 (N_45107,N_42491,N_42790);
nor U45108 (N_45108,N_43394,N_42438);
and U45109 (N_45109,N_42579,N_43326);
or U45110 (N_45110,N_43097,N_42412);
or U45111 (N_45111,N_42947,N_42203);
nor U45112 (N_45112,N_43787,N_42997);
nor U45113 (N_45113,N_43161,N_42929);
nand U45114 (N_45114,N_43112,N_42589);
nand U45115 (N_45115,N_42655,N_42829);
or U45116 (N_45116,N_43682,N_43090);
nor U45117 (N_45117,N_43200,N_43990);
nor U45118 (N_45118,N_43537,N_42094);
nor U45119 (N_45119,N_43292,N_42375);
and U45120 (N_45120,N_43087,N_42401);
nor U45121 (N_45121,N_42180,N_42801);
nor U45122 (N_45122,N_43212,N_43358);
nor U45123 (N_45123,N_43234,N_42125);
nor U45124 (N_45124,N_42676,N_43975);
nor U45125 (N_45125,N_43850,N_42270);
or U45126 (N_45126,N_43443,N_42968);
nor U45127 (N_45127,N_42390,N_43531);
nand U45128 (N_45128,N_42278,N_42799);
xor U45129 (N_45129,N_43671,N_42853);
nand U45130 (N_45130,N_43471,N_43401);
nand U45131 (N_45131,N_43598,N_42898);
nand U45132 (N_45132,N_42634,N_42774);
or U45133 (N_45133,N_43616,N_43648);
and U45134 (N_45134,N_43536,N_42060);
nand U45135 (N_45135,N_43975,N_43104);
and U45136 (N_45136,N_42132,N_42980);
or U45137 (N_45137,N_42962,N_43465);
nand U45138 (N_45138,N_43070,N_43603);
nand U45139 (N_45139,N_43085,N_43956);
or U45140 (N_45140,N_43769,N_42855);
and U45141 (N_45141,N_42621,N_42035);
or U45142 (N_45142,N_43644,N_42091);
nand U45143 (N_45143,N_43662,N_43600);
nor U45144 (N_45144,N_42254,N_43984);
xnor U45145 (N_45145,N_43615,N_43777);
and U45146 (N_45146,N_42642,N_43199);
or U45147 (N_45147,N_42403,N_43130);
or U45148 (N_45148,N_43999,N_43196);
or U45149 (N_45149,N_43000,N_42269);
nand U45150 (N_45150,N_42995,N_43013);
nand U45151 (N_45151,N_43351,N_43130);
or U45152 (N_45152,N_42690,N_42410);
nand U45153 (N_45153,N_42947,N_42405);
or U45154 (N_45154,N_42019,N_43310);
nor U45155 (N_45155,N_42587,N_43667);
or U45156 (N_45156,N_42208,N_42654);
nand U45157 (N_45157,N_43866,N_43637);
nand U45158 (N_45158,N_43600,N_42524);
and U45159 (N_45159,N_42947,N_42242);
and U45160 (N_45160,N_42408,N_43813);
nor U45161 (N_45161,N_43831,N_42202);
and U45162 (N_45162,N_43339,N_42089);
nor U45163 (N_45163,N_42865,N_42746);
nor U45164 (N_45164,N_42402,N_43392);
nand U45165 (N_45165,N_42338,N_43663);
or U45166 (N_45166,N_43374,N_42498);
nand U45167 (N_45167,N_42607,N_42889);
nor U45168 (N_45168,N_42490,N_42765);
and U45169 (N_45169,N_42095,N_42275);
or U45170 (N_45170,N_43833,N_42381);
or U45171 (N_45171,N_42748,N_42060);
nor U45172 (N_45172,N_43088,N_42931);
and U45173 (N_45173,N_43805,N_43668);
nor U45174 (N_45174,N_42993,N_42306);
nor U45175 (N_45175,N_43333,N_42111);
or U45176 (N_45176,N_42343,N_43210);
and U45177 (N_45177,N_42915,N_43738);
nand U45178 (N_45178,N_43005,N_43799);
and U45179 (N_45179,N_43778,N_43950);
or U45180 (N_45180,N_42354,N_42296);
and U45181 (N_45181,N_43647,N_42874);
nor U45182 (N_45182,N_42327,N_43648);
and U45183 (N_45183,N_42453,N_43542);
nand U45184 (N_45184,N_43431,N_42616);
or U45185 (N_45185,N_42951,N_42228);
nand U45186 (N_45186,N_43324,N_42108);
nand U45187 (N_45187,N_42558,N_43719);
and U45188 (N_45188,N_43243,N_43813);
or U45189 (N_45189,N_43944,N_42133);
nor U45190 (N_45190,N_43876,N_43005);
nand U45191 (N_45191,N_43396,N_42123);
nand U45192 (N_45192,N_43605,N_42923);
nor U45193 (N_45193,N_43028,N_42742);
nand U45194 (N_45194,N_43676,N_42105);
nor U45195 (N_45195,N_43518,N_43841);
or U45196 (N_45196,N_43670,N_43419);
nand U45197 (N_45197,N_43121,N_42958);
and U45198 (N_45198,N_42740,N_42663);
or U45199 (N_45199,N_42795,N_43167);
nor U45200 (N_45200,N_43166,N_42038);
or U45201 (N_45201,N_43072,N_43933);
and U45202 (N_45202,N_43250,N_43429);
nor U45203 (N_45203,N_42009,N_42455);
or U45204 (N_45204,N_42807,N_43133);
or U45205 (N_45205,N_43905,N_43472);
or U45206 (N_45206,N_43626,N_43297);
nor U45207 (N_45207,N_42524,N_43359);
nand U45208 (N_45208,N_42150,N_42659);
or U45209 (N_45209,N_43992,N_43791);
or U45210 (N_45210,N_43224,N_42663);
or U45211 (N_45211,N_43331,N_43692);
or U45212 (N_45212,N_42209,N_43696);
nand U45213 (N_45213,N_43275,N_42703);
and U45214 (N_45214,N_42187,N_42910);
nand U45215 (N_45215,N_43497,N_43868);
nand U45216 (N_45216,N_43644,N_43135);
or U45217 (N_45217,N_42376,N_42303);
and U45218 (N_45218,N_43267,N_42045);
nand U45219 (N_45219,N_42585,N_42849);
or U45220 (N_45220,N_43951,N_42656);
nor U45221 (N_45221,N_43664,N_43488);
or U45222 (N_45222,N_43365,N_43534);
and U45223 (N_45223,N_43884,N_43919);
and U45224 (N_45224,N_42792,N_42308);
nand U45225 (N_45225,N_43361,N_43931);
and U45226 (N_45226,N_43367,N_43736);
and U45227 (N_45227,N_43994,N_42593);
nor U45228 (N_45228,N_43373,N_42528);
nor U45229 (N_45229,N_43293,N_42383);
or U45230 (N_45230,N_43240,N_43071);
nor U45231 (N_45231,N_42743,N_43687);
or U45232 (N_45232,N_42673,N_42115);
nand U45233 (N_45233,N_42848,N_43556);
nor U45234 (N_45234,N_42068,N_43323);
nand U45235 (N_45235,N_42099,N_42285);
nand U45236 (N_45236,N_42528,N_43651);
nand U45237 (N_45237,N_42849,N_42580);
nor U45238 (N_45238,N_43765,N_42875);
and U45239 (N_45239,N_42862,N_43919);
nand U45240 (N_45240,N_42251,N_43116);
and U45241 (N_45241,N_42831,N_42619);
nand U45242 (N_45242,N_42107,N_42058);
nand U45243 (N_45243,N_42231,N_42976);
nor U45244 (N_45244,N_43030,N_43522);
nor U45245 (N_45245,N_42091,N_43224);
or U45246 (N_45246,N_42959,N_43587);
and U45247 (N_45247,N_42135,N_43356);
nor U45248 (N_45248,N_43561,N_42015);
or U45249 (N_45249,N_42740,N_43248);
and U45250 (N_45250,N_42118,N_43849);
and U45251 (N_45251,N_43371,N_43237);
nand U45252 (N_45252,N_42057,N_43117);
nor U45253 (N_45253,N_43186,N_43039);
or U45254 (N_45254,N_42773,N_43270);
and U45255 (N_45255,N_42436,N_43821);
or U45256 (N_45256,N_43113,N_43969);
nor U45257 (N_45257,N_42996,N_43174);
nand U45258 (N_45258,N_42415,N_42374);
xor U45259 (N_45259,N_42163,N_43391);
nor U45260 (N_45260,N_43858,N_43036);
nor U45261 (N_45261,N_42555,N_43649);
nand U45262 (N_45262,N_43954,N_43211);
nor U45263 (N_45263,N_42131,N_42807);
nor U45264 (N_45264,N_43124,N_43688);
nand U45265 (N_45265,N_42906,N_42179);
nor U45266 (N_45266,N_43507,N_43993);
nand U45267 (N_45267,N_43643,N_43700);
xor U45268 (N_45268,N_43688,N_42411);
nor U45269 (N_45269,N_43319,N_42228);
or U45270 (N_45270,N_43853,N_42867);
nand U45271 (N_45271,N_43609,N_42139);
and U45272 (N_45272,N_42086,N_43812);
or U45273 (N_45273,N_42138,N_43750);
or U45274 (N_45274,N_42493,N_43127);
and U45275 (N_45275,N_42600,N_42716);
nor U45276 (N_45276,N_42781,N_43833);
nand U45277 (N_45277,N_42132,N_43768);
nand U45278 (N_45278,N_42053,N_43305);
nand U45279 (N_45279,N_43744,N_42207);
nand U45280 (N_45280,N_43096,N_43774);
or U45281 (N_45281,N_43592,N_42968);
nand U45282 (N_45282,N_43629,N_43123);
nor U45283 (N_45283,N_42667,N_43241);
and U45284 (N_45284,N_42891,N_43237);
nor U45285 (N_45285,N_42832,N_42655);
or U45286 (N_45286,N_43454,N_42811);
and U45287 (N_45287,N_43149,N_42705);
nand U45288 (N_45288,N_43963,N_43029);
and U45289 (N_45289,N_43120,N_42037);
nand U45290 (N_45290,N_42237,N_42801);
nand U45291 (N_45291,N_42240,N_42442);
nand U45292 (N_45292,N_43000,N_42824);
nand U45293 (N_45293,N_42387,N_43951);
and U45294 (N_45294,N_42515,N_43757);
nor U45295 (N_45295,N_42345,N_42024);
nor U45296 (N_45296,N_43529,N_42787);
nand U45297 (N_45297,N_42759,N_42272);
nand U45298 (N_45298,N_43805,N_43725);
and U45299 (N_45299,N_42555,N_42104);
or U45300 (N_45300,N_42328,N_43455);
or U45301 (N_45301,N_43517,N_42340);
and U45302 (N_45302,N_42161,N_42982);
nand U45303 (N_45303,N_43945,N_43000);
nor U45304 (N_45304,N_42512,N_42697);
xnor U45305 (N_45305,N_42993,N_42255);
and U45306 (N_45306,N_43947,N_42025);
and U45307 (N_45307,N_43351,N_43490);
and U45308 (N_45308,N_43516,N_43447);
nand U45309 (N_45309,N_43702,N_42000);
nor U45310 (N_45310,N_43164,N_42834);
xor U45311 (N_45311,N_43422,N_42273);
or U45312 (N_45312,N_43872,N_42747);
nor U45313 (N_45313,N_42464,N_42739);
nor U45314 (N_45314,N_43320,N_42644);
and U45315 (N_45315,N_42546,N_43860);
nand U45316 (N_45316,N_42571,N_43320);
nor U45317 (N_45317,N_42332,N_43798);
or U45318 (N_45318,N_42629,N_43395);
nor U45319 (N_45319,N_42626,N_43929);
or U45320 (N_45320,N_42642,N_43122);
nor U45321 (N_45321,N_42638,N_43603);
nor U45322 (N_45322,N_42760,N_43473);
or U45323 (N_45323,N_42707,N_42324);
and U45324 (N_45324,N_42708,N_43903);
and U45325 (N_45325,N_43186,N_43785);
nand U45326 (N_45326,N_43031,N_42455);
nor U45327 (N_45327,N_42170,N_43303);
nor U45328 (N_45328,N_43378,N_43331);
nand U45329 (N_45329,N_42600,N_43590);
nor U45330 (N_45330,N_43622,N_43760);
nand U45331 (N_45331,N_43847,N_43229);
xnor U45332 (N_45332,N_42931,N_43412);
and U45333 (N_45333,N_43490,N_42919);
nand U45334 (N_45334,N_42111,N_43706);
nor U45335 (N_45335,N_43415,N_42108);
nor U45336 (N_45336,N_43237,N_43822);
and U45337 (N_45337,N_42594,N_42051);
and U45338 (N_45338,N_43882,N_43810);
or U45339 (N_45339,N_43290,N_42210);
nor U45340 (N_45340,N_43511,N_43482);
nand U45341 (N_45341,N_43887,N_43549);
xor U45342 (N_45342,N_43676,N_43852);
nand U45343 (N_45343,N_42977,N_43742);
and U45344 (N_45344,N_43188,N_42041);
nand U45345 (N_45345,N_42443,N_42003);
and U45346 (N_45346,N_43240,N_43076);
nand U45347 (N_45347,N_43740,N_42203);
nand U45348 (N_45348,N_42004,N_42820);
or U45349 (N_45349,N_43140,N_42841);
or U45350 (N_45350,N_43964,N_42176);
or U45351 (N_45351,N_43489,N_43391);
nor U45352 (N_45352,N_42844,N_43872);
nand U45353 (N_45353,N_43757,N_43032);
nor U45354 (N_45354,N_42322,N_42567);
or U45355 (N_45355,N_42402,N_43195);
or U45356 (N_45356,N_43625,N_42713);
nor U45357 (N_45357,N_43457,N_42242);
or U45358 (N_45358,N_43708,N_43485);
and U45359 (N_45359,N_43351,N_43589);
or U45360 (N_45360,N_43653,N_42423);
nor U45361 (N_45361,N_43471,N_43362);
nand U45362 (N_45362,N_43861,N_43906);
nand U45363 (N_45363,N_42300,N_43350);
or U45364 (N_45364,N_42956,N_43016);
or U45365 (N_45365,N_43878,N_43900);
nand U45366 (N_45366,N_43023,N_42468);
and U45367 (N_45367,N_42950,N_43866);
and U45368 (N_45368,N_42630,N_42312);
nand U45369 (N_45369,N_42105,N_43476);
and U45370 (N_45370,N_43564,N_43444);
and U45371 (N_45371,N_43745,N_42159);
or U45372 (N_45372,N_43196,N_43333);
xnor U45373 (N_45373,N_42170,N_42019);
xnor U45374 (N_45374,N_42738,N_42179);
nor U45375 (N_45375,N_42998,N_42323);
nand U45376 (N_45376,N_42083,N_43206);
nand U45377 (N_45377,N_42244,N_43150);
nand U45378 (N_45378,N_42574,N_43532);
nand U45379 (N_45379,N_42144,N_42923);
and U45380 (N_45380,N_43370,N_42532);
and U45381 (N_45381,N_43721,N_43626);
and U45382 (N_45382,N_43661,N_43511);
nand U45383 (N_45383,N_42296,N_43639);
or U45384 (N_45384,N_42904,N_42843);
nor U45385 (N_45385,N_43858,N_42958);
and U45386 (N_45386,N_43885,N_43224);
or U45387 (N_45387,N_42926,N_43407);
and U45388 (N_45388,N_43537,N_42665);
and U45389 (N_45389,N_42967,N_43120);
and U45390 (N_45390,N_42809,N_43538);
and U45391 (N_45391,N_42873,N_43344);
nor U45392 (N_45392,N_43053,N_43327);
or U45393 (N_45393,N_43648,N_43290);
or U45394 (N_45394,N_43915,N_43560);
nor U45395 (N_45395,N_42533,N_42438);
nor U45396 (N_45396,N_43381,N_43785);
nand U45397 (N_45397,N_42278,N_42692);
or U45398 (N_45398,N_43970,N_42866);
or U45399 (N_45399,N_43195,N_43483);
and U45400 (N_45400,N_42873,N_42994);
nand U45401 (N_45401,N_42996,N_42026);
or U45402 (N_45402,N_42278,N_43410);
and U45403 (N_45403,N_43912,N_42190);
and U45404 (N_45404,N_43313,N_42544);
nand U45405 (N_45405,N_43279,N_43660);
nand U45406 (N_45406,N_42119,N_43565);
nor U45407 (N_45407,N_42827,N_42131);
nor U45408 (N_45408,N_42935,N_42039);
and U45409 (N_45409,N_42538,N_43080);
and U45410 (N_45410,N_43066,N_42984);
nor U45411 (N_45411,N_43895,N_43822);
and U45412 (N_45412,N_42909,N_43614);
nand U45413 (N_45413,N_42602,N_42287);
and U45414 (N_45414,N_42170,N_42519);
nor U45415 (N_45415,N_43384,N_43499);
and U45416 (N_45416,N_42550,N_42124);
and U45417 (N_45417,N_42766,N_43130);
or U45418 (N_45418,N_42549,N_43636);
and U45419 (N_45419,N_43014,N_42108);
nand U45420 (N_45420,N_42865,N_42982);
nand U45421 (N_45421,N_42443,N_43479);
and U45422 (N_45422,N_42238,N_43628);
or U45423 (N_45423,N_43079,N_42373);
or U45424 (N_45424,N_42548,N_42790);
and U45425 (N_45425,N_43728,N_42285);
xnor U45426 (N_45426,N_42914,N_43446);
nor U45427 (N_45427,N_43413,N_42334);
and U45428 (N_45428,N_42598,N_43151);
and U45429 (N_45429,N_43574,N_42550);
or U45430 (N_45430,N_42491,N_43664);
and U45431 (N_45431,N_42754,N_43290);
or U45432 (N_45432,N_43368,N_42360);
nand U45433 (N_45433,N_42340,N_43317);
nor U45434 (N_45434,N_42877,N_42764);
nor U45435 (N_45435,N_43801,N_43794);
nor U45436 (N_45436,N_42643,N_43024);
xnor U45437 (N_45437,N_42576,N_42670);
or U45438 (N_45438,N_42551,N_43772);
or U45439 (N_45439,N_42786,N_43226);
nand U45440 (N_45440,N_43525,N_43414);
nor U45441 (N_45441,N_42912,N_42221);
or U45442 (N_45442,N_43702,N_42122);
nand U45443 (N_45443,N_43948,N_43475);
nor U45444 (N_45444,N_43697,N_42944);
nor U45445 (N_45445,N_43545,N_42090);
xor U45446 (N_45446,N_43407,N_42794);
nand U45447 (N_45447,N_42897,N_43174);
or U45448 (N_45448,N_42742,N_42293);
nand U45449 (N_45449,N_43969,N_42438);
nor U45450 (N_45450,N_43495,N_43903);
or U45451 (N_45451,N_43190,N_42788);
nand U45452 (N_45452,N_42008,N_42245);
nor U45453 (N_45453,N_42937,N_43072);
or U45454 (N_45454,N_43698,N_42132);
and U45455 (N_45455,N_43442,N_42135);
or U45456 (N_45456,N_43049,N_43260);
nor U45457 (N_45457,N_43482,N_43043);
nor U45458 (N_45458,N_43807,N_43141);
nor U45459 (N_45459,N_42727,N_43012);
and U45460 (N_45460,N_42794,N_42680);
nand U45461 (N_45461,N_42119,N_43223);
and U45462 (N_45462,N_43336,N_42982);
nor U45463 (N_45463,N_42659,N_42416);
or U45464 (N_45464,N_42580,N_43644);
or U45465 (N_45465,N_42858,N_43072);
nor U45466 (N_45466,N_42188,N_42072);
or U45467 (N_45467,N_42353,N_42142);
and U45468 (N_45468,N_43090,N_43577);
nand U45469 (N_45469,N_43609,N_42667);
and U45470 (N_45470,N_43916,N_43403);
nand U45471 (N_45471,N_43448,N_42841);
or U45472 (N_45472,N_43879,N_43348);
nand U45473 (N_45473,N_42954,N_43274);
or U45474 (N_45474,N_43073,N_43495);
and U45475 (N_45475,N_42170,N_43840);
nand U45476 (N_45476,N_43109,N_43583);
and U45477 (N_45477,N_42167,N_43443);
and U45478 (N_45478,N_42476,N_43681);
and U45479 (N_45479,N_43151,N_43407);
and U45480 (N_45480,N_43864,N_42945);
and U45481 (N_45481,N_42011,N_43095);
xor U45482 (N_45482,N_43169,N_43949);
or U45483 (N_45483,N_43343,N_43574);
nand U45484 (N_45484,N_43745,N_42254);
and U45485 (N_45485,N_42435,N_42157);
nand U45486 (N_45486,N_43581,N_43262);
and U45487 (N_45487,N_42082,N_43159);
nor U45488 (N_45488,N_42705,N_42630);
nor U45489 (N_45489,N_43234,N_43009);
nand U45490 (N_45490,N_43894,N_43412);
nand U45491 (N_45491,N_43625,N_42383);
nand U45492 (N_45492,N_43983,N_42252);
and U45493 (N_45493,N_42357,N_43988);
nor U45494 (N_45494,N_42499,N_42489);
and U45495 (N_45495,N_43233,N_42708);
or U45496 (N_45496,N_42049,N_43101);
or U45497 (N_45497,N_43985,N_42706);
and U45498 (N_45498,N_43760,N_43986);
nor U45499 (N_45499,N_43468,N_42606);
xnor U45500 (N_45500,N_43278,N_43937);
and U45501 (N_45501,N_43187,N_42495);
xnor U45502 (N_45502,N_43672,N_43521);
and U45503 (N_45503,N_42501,N_43754);
or U45504 (N_45504,N_43506,N_42005);
or U45505 (N_45505,N_43520,N_42306);
and U45506 (N_45506,N_43285,N_42608);
and U45507 (N_45507,N_42142,N_42682);
and U45508 (N_45508,N_42534,N_42759);
nand U45509 (N_45509,N_42320,N_42691);
and U45510 (N_45510,N_43895,N_43273);
and U45511 (N_45511,N_43700,N_42830);
nand U45512 (N_45512,N_43982,N_42437);
nand U45513 (N_45513,N_42667,N_43321);
nand U45514 (N_45514,N_42395,N_43337);
or U45515 (N_45515,N_42060,N_43199);
or U45516 (N_45516,N_42363,N_42019);
nand U45517 (N_45517,N_42050,N_43103);
and U45518 (N_45518,N_42687,N_43292);
nand U45519 (N_45519,N_43095,N_43247);
nor U45520 (N_45520,N_42637,N_43840);
nor U45521 (N_45521,N_43607,N_42218);
and U45522 (N_45522,N_43785,N_42599);
nor U45523 (N_45523,N_42049,N_42365);
nor U45524 (N_45524,N_42607,N_42549);
and U45525 (N_45525,N_42424,N_43800);
nand U45526 (N_45526,N_43508,N_42002);
or U45527 (N_45527,N_43357,N_43371);
nor U45528 (N_45528,N_43455,N_43517);
nand U45529 (N_45529,N_42398,N_42002);
nand U45530 (N_45530,N_42618,N_43198);
nor U45531 (N_45531,N_43663,N_43192);
nor U45532 (N_45532,N_43274,N_43888);
nor U45533 (N_45533,N_42477,N_43875);
nand U45534 (N_45534,N_43935,N_42140);
or U45535 (N_45535,N_43667,N_43703);
nor U45536 (N_45536,N_42555,N_42739);
and U45537 (N_45537,N_43830,N_42050);
or U45538 (N_45538,N_42760,N_43144);
nor U45539 (N_45539,N_43750,N_42058);
and U45540 (N_45540,N_42325,N_43517);
xnor U45541 (N_45541,N_42756,N_43415);
nand U45542 (N_45542,N_42257,N_42512);
or U45543 (N_45543,N_43567,N_43291);
and U45544 (N_45544,N_42485,N_43340);
nand U45545 (N_45545,N_43416,N_42802);
and U45546 (N_45546,N_43454,N_42131);
nor U45547 (N_45547,N_42959,N_43694);
or U45548 (N_45548,N_42738,N_42835);
nor U45549 (N_45549,N_43645,N_43356);
or U45550 (N_45550,N_42832,N_43720);
nand U45551 (N_45551,N_43040,N_43239);
nand U45552 (N_45552,N_43799,N_43368);
nand U45553 (N_45553,N_43948,N_43615);
or U45554 (N_45554,N_43828,N_42221);
nand U45555 (N_45555,N_43990,N_43671);
or U45556 (N_45556,N_43347,N_42333);
and U45557 (N_45557,N_43939,N_43911);
or U45558 (N_45558,N_42454,N_43384);
and U45559 (N_45559,N_42185,N_43310);
or U45560 (N_45560,N_43889,N_42328);
nor U45561 (N_45561,N_42613,N_43954);
nand U45562 (N_45562,N_42489,N_43162);
nand U45563 (N_45563,N_42513,N_43013);
and U45564 (N_45564,N_42554,N_42593);
and U45565 (N_45565,N_42993,N_42300);
or U45566 (N_45566,N_43470,N_42470);
and U45567 (N_45567,N_42326,N_42912);
nand U45568 (N_45568,N_43673,N_42515);
nand U45569 (N_45569,N_43900,N_42138);
and U45570 (N_45570,N_43172,N_43309);
nor U45571 (N_45571,N_43341,N_42604);
or U45572 (N_45572,N_42253,N_42063);
and U45573 (N_45573,N_43126,N_42904);
nor U45574 (N_45574,N_42347,N_42271);
or U45575 (N_45575,N_43139,N_42808);
nand U45576 (N_45576,N_42103,N_42493);
nor U45577 (N_45577,N_42874,N_43963);
nor U45578 (N_45578,N_43253,N_42173);
nand U45579 (N_45579,N_42772,N_43828);
or U45580 (N_45580,N_42333,N_43909);
nand U45581 (N_45581,N_42807,N_42073);
nor U45582 (N_45582,N_43221,N_42115);
nor U45583 (N_45583,N_42796,N_42824);
or U45584 (N_45584,N_43266,N_43985);
and U45585 (N_45585,N_42940,N_42798);
nand U45586 (N_45586,N_42501,N_42961);
nor U45587 (N_45587,N_43675,N_42961);
xor U45588 (N_45588,N_42740,N_43952);
and U45589 (N_45589,N_42803,N_43539);
nor U45590 (N_45590,N_42801,N_43357);
nand U45591 (N_45591,N_43164,N_42894);
and U45592 (N_45592,N_42821,N_42261);
nor U45593 (N_45593,N_42065,N_43975);
or U45594 (N_45594,N_42187,N_42918);
or U45595 (N_45595,N_43399,N_43306);
or U45596 (N_45596,N_42171,N_43390);
or U45597 (N_45597,N_42734,N_42468);
nand U45598 (N_45598,N_42312,N_42055);
nor U45599 (N_45599,N_43780,N_42020);
or U45600 (N_45600,N_42538,N_42947);
or U45601 (N_45601,N_43783,N_42665);
nor U45602 (N_45602,N_43907,N_42613);
or U45603 (N_45603,N_42441,N_43913);
nand U45604 (N_45604,N_43047,N_42789);
and U45605 (N_45605,N_43495,N_43111);
nand U45606 (N_45606,N_43262,N_43835);
nand U45607 (N_45607,N_42225,N_42632);
nand U45608 (N_45608,N_42613,N_43378);
and U45609 (N_45609,N_43147,N_42041);
or U45610 (N_45610,N_42477,N_43919);
nand U45611 (N_45611,N_43808,N_42768);
nor U45612 (N_45612,N_42103,N_43546);
or U45613 (N_45613,N_42504,N_43013);
nand U45614 (N_45614,N_42358,N_43421);
nor U45615 (N_45615,N_42622,N_42038);
nand U45616 (N_45616,N_43730,N_42751);
nor U45617 (N_45617,N_43825,N_43077);
nor U45618 (N_45618,N_43252,N_43645);
nand U45619 (N_45619,N_42229,N_43126);
and U45620 (N_45620,N_43807,N_42312);
nor U45621 (N_45621,N_42361,N_42089);
and U45622 (N_45622,N_43524,N_43624);
or U45623 (N_45623,N_42150,N_43172);
nand U45624 (N_45624,N_42132,N_42536);
nor U45625 (N_45625,N_42472,N_43147);
or U45626 (N_45626,N_43984,N_42204);
nand U45627 (N_45627,N_42260,N_43647);
or U45628 (N_45628,N_42889,N_42213);
and U45629 (N_45629,N_42425,N_43376);
and U45630 (N_45630,N_43106,N_43615);
nor U45631 (N_45631,N_42661,N_43080);
and U45632 (N_45632,N_42317,N_42748);
nand U45633 (N_45633,N_42680,N_43417);
or U45634 (N_45634,N_42336,N_42913);
nor U45635 (N_45635,N_42183,N_43936);
nor U45636 (N_45636,N_42343,N_42269);
nor U45637 (N_45637,N_42688,N_42250);
nor U45638 (N_45638,N_43143,N_42113);
or U45639 (N_45639,N_42269,N_43122);
nor U45640 (N_45640,N_43588,N_42722);
nor U45641 (N_45641,N_43502,N_43973);
or U45642 (N_45642,N_42952,N_43918);
nand U45643 (N_45643,N_42368,N_43485);
nor U45644 (N_45644,N_42395,N_42978);
and U45645 (N_45645,N_42927,N_42774);
nand U45646 (N_45646,N_43518,N_42429);
nor U45647 (N_45647,N_43074,N_42442);
nor U45648 (N_45648,N_42224,N_42613);
nor U45649 (N_45649,N_42062,N_43791);
nand U45650 (N_45650,N_42616,N_43614);
nand U45651 (N_45651,N_42574,N_43347);
nand U45652 (N_45652,N_43912,N_43029);
and U45653 (N_45653,N_43581,N_43498);
nand U45654 (N_45654,N_42276,N_42564);
nand U45655 (N_45655,N_43386,N_42622);
or U45656 (N_45656,N_42325,N_42788);
or U45657 (N_45657,N_42690,N_42832);
nand U45658 (N_45658,N_42903,N_42633);
or U45659 (N_45659,N_43229,N_42061);
nor U45660 (N_45660,N_43962,N_43161);
xnor U45661 (N_45661,N_42397,N_42842);
and U45662 (N_45662,N_43064,N_43456);
nor U45663 (N_45663,N_43685,N_42177);
or U45664 (N_45664,N_42312,N_43792);
or U45665 (N_45665,N_43402,N_42152);
nand U45666 (N_45666,N_42362,N_42095);
or U45667 (N_45667,N_42295,N_43713);
and U45668 (N_45668,N_43994,N_43438);
nand U45669 (N_45669,N_43466,N_43842);
or U45670 (N_45670,N_42884,N_42198);
and U45671 (N_45671,N_43614,N_42389);
nand U45672 (N_45672,N_43463,N_43132);
nand U45673 (N_45673,N_42290,N_43277);
nor U45674 (N_45674,N_42399,N_43783);
and U45675 (N_45675,N_43022,N_43485);
nor U45676 (N_45676,N_42787,N_43834);
nor U45677 (N_45677,N_43216,N_43421);
nor U45678 (N_45678,N_42831,N_43639);
nand U45679 (N_45679,N_42910,N_42369);
or U45680 (N_45680,N_42300,N_43085);
or U45681 (N_45681,N_42955,N_43917);
xnor U45682 (N_45682,N_43712,N_43485);
nor U45683 (N_45683,N_43816,N_42170);
nand U45684 (N_45684,N_43992,N_42814);
nor U45685 (N_45685,N_42059,N_42758);
nand U45686 (N_45686,N_43393,N_43848);
or U45687 (N_45687,N_42624,N_43762);
nor U45688 (N_45688,N_42666,N_43424);
nor U45689 (N_45689,N_42402,N_43984);
nand U45690 (N_45690,N_43600,N_42407);
or U45691 (N_45691,N_42410,N_43202);
or U45692 (N_45692,N_43053,N_43988);
or U45693 (N_45693,N_42381,N_42246);
and U45694 (N_45694,N_42992,N_42549);
or U45695 (N_45695,N_43808,N_42774);
nand U45696 (N_45696,N_43401,N_42212);
or U45697 (N_45697,N_42857,N_43134);
or U45698 (N_45698,N_43440,N_42727);
or U45699 (N_45699,N_43130,N_43609);
nand U45700 (N_45700,N_43882,N_42277);
nor U45701 (N_45701,N_43910,N_42955);
nor U45702 (N_45702,N_42287,N_42659);
and U45703 (N_45703,N_43178,N_43279);
nor U45704 (N_45704,N_42763,N_43779);
and U45705 (N_45705,N_42746,N_43420);
and U45706 (N_45706,N_43157,N_43015);
nor U45707 (N_45707,N_42413,N_43129);
and U45708 (N_45708,N_43849,N_43617);
and U45709 (N_45709,N_42938,N_42618);
and U45710 (N_45710,N_42458,N_43648);
nor U45711 (N_45711,N_42272,N_42078);
nor U45712 (N_45712,N_43756,N_43974);
or U45713 (N_45713,N_42365,N_42000);
or U45714 (N_45714,N_42231,N_42964);
nand U45715 (N_45715,N_42152,N_42871);
and U45716 (N_45716,N_43536,N_43052);
or U45717 (N_45717,N_42473,N_42157);
nor U45718 (N_45718,N_43420,N_42289);
and U45719 (N_45719,N_42576,N_43297);
or U45720 (N_45720,N_42783,N_43248);
nor U45721 (N_45721,N_42291,N_43599);
or U45722 (N_45722,N_43890,N_42786);
nand U45723 (N_45723,N_42039,N_43057);
nand U45724 (N_45724,N_43902,N_43816);
or U45725 (N_45725,N_42609,N_43701);
nand U45726 (N_45726,N_43202,N_43265);
nand U45727 (N_45727,N_42919,N_42734);
nor U45728 (N_45728,N_43175,N_42758);
nor U45729 (N_45729,N_42906,N_42885);
nand U45730 (N_45730,N_42034,N_43813);
nor U45731 (N_45731,N_43190,N_43016);
or U45732 (N_45732,N_43514,N_43922);
xnor U45733 (N_45733,N_43980,N_42318);
nand U45734 (N_45734,N_43946,N_42196);
nand U45735 (N_45735,N_42293,N_42712);
and U45736 (N_45736,N_42856,N_43778);
nor U45737 (N_45737,N_43725,N_43419);
nand U45738 (N_45738,N_43294,N_42737);
nand U45739 (N_45739,N_42434,N_42349);
or U45740 (N_45740,N_42379,N_43896);
or U45741 (N_45741,N_42411,N_43325);
or U45742 (N_45742,N_43388,N_43451);
or U45743 (N_45743,N_43801,N_43183);
or U45744 (N_45744,N_43613,N_43157);
nor U45745 (N_45745,N_43181,N_42653);
and U45746 (N_45746,N_42844,N_43636);
xor U45747 (N_45747,N_42311,N_42977);
and U45748 (N_45748,N_43660,N_42861);
nor U45749 (N_45749,N_42228,N_43922);
or U45750 (N_45750,N_42793,N_43970);
or U45751 (N_45751,N_42078,N_43365);
or U45752 (N_45752,N_43832,N_43463);
or U45753 (N_45753,N_42234,N_43684);
and U45754 (N_45754,N_43315,N_42198);
or U45755 (N_45755,N_43962,N_43940);
nand U45756 (N_45756,N_43571,N_43802);
nand U45757 (N_45757,N_42640,N_42464);
nor U45758 (N_45758,N_43870,N_43584);
xor U45759 (N_45759,N_42421,N_43548);
and U45760 (N_45760,N_42856,N_42876);
nor U45761 (N_45761,N_43698,N_42165);
nand U45762 (N_45762,N_43699,N_42735);
or U45763 (N_45763,N_42606,N_43953);
and U45764 (N_45764,N_43254,N_43299);
or U45765 (N_45765,N_43616,N_43655);
or U45766 (N_45766,N_42378,N_43483);
nor U45767 (N_45767,N_42594,N_42630);
nand U45768 (N_45768,N_43639,N_42317);
nand U45769 (N_45769,N_43231,N_42089);
or U45770 (N_45770,N_43801,N_43753);
nor U45771 (N_45771,N_43441,N_43417);
and U45772 (N_45772,N_43120,N_42244);
nand U45773 (N_45773,N_43775,N_42890);
or U45774 (N_45774,N_43192,N_43493);
and U45775 (N_45775,N_43716,N_42480);
nor U45776 (N_45776,N_42311,N_42331);
and U45777 (N_45777,N_42790,N_42545);
nor U45778 (N_45778,N_43414,N_43179);
xnor U45779 (N_45779,N_43758,N_42925);
and U45780 (N_45780,N_43217,N_42883);
nand U45781 (N_45781,N_42528,N_43894);
or U45782 (N_45782,N_42601,N_42649);
and U45783 (N_45783,N_42481,N_42864);
nand U45784 (N_45784,N_43264,N_42597);
nor U45785 (N_45785,N_42472,N_42279);
nor U45786 (N_45786,N_43315,N_43863);
nand U45787 (N_45787,N_42204,N_42769);
nand U45788 (N_45788,N_43335,N_42711);
nand U45789 (N_45789,N_43933,N_42400);
and U45790 (N_45790,N_42538,N_43125);
nor U45791 (N_45791,N_42263,N_43754);
nor U45792 (N_45792,N_42155,N_43732);
nor U45793 (N_45793,N_42187,N_42293);
nand U45794 (N_45794,N_42618,N_43703);
nand U45795 (N_45795,N_42361,N_43476);
and U45796 (N_45796,N_43542,N_42786);
or U45797 (N_45797,N_43031,N_42027);
and U45798 (N_45798,N_43854,N_43273);
or U45799 (N_45799,N_43434,N_42913);
or U45800 (N_45800,N_43298,N_42692);
or U45801 (N_45801,N_42826,N_42548);
and U45802 (N_45802,N_43514,N_43559);
or U45803 (N_45803,N_42697,N_43102);
or U45804 (N_45804,N_43239,N_42930);
nand U45805 (N_45805,N_42057,N_43001);
nor U45806 (N_45806,N_42010,N_43708);
nor U45807 (N_45807,N_42359,N_43013);
nand U45808 (N_45808,N_42394,N_43422);
and U45809 (N_45809,N_43249,N_42613);
or U45810 (N_45810,N_43896,N_42077);
nand U45811 (N_45811,N_42905,N_43290);
nand U45812 (N_45812,N_42491,N_42672);
nand U45813 (N_45813,N_42815,N_42640);
nand U45814 (N_45814,N_42707,N_42403);
nand U45815 (N_45815,N_42591,N_43799);
nand U45816 (N_45816,N_42502,N_43775);
nand U45817 (N_45817,N_42046,N_42062);
nor U45818 (N_45818,N_42061,N_42260);
or U45819 (N_45819,N_42157,N_43264);
and U45820 (N_45820,N_42840,N_42598);
and U45821 (N_45821,N_43310,N_42098);
nor U45822 (N_45822,N_43486,N_43165);
nand U45823 (N_45823,N_42906,N_42066);
and U45824 (N_45824,N_42444,N_42450);
nor U45825 (N_45825,N_43173,N_42609);
nand U45826 (N_45826,N_42098,N_42919);
and U45827 (N_45827,N_42021,N_42785);
or U45828 (N_45828,N_43312,N_42878);
and U45829 (N_45829,N_42626,N_43093);
nand U45830 (N_45830,N_42455,N_43725);
or U45831 (N_45831,N_42865,N_43565);
or U45832 (N_45832,N_42454,N_42903);
or U45833 (N_45833,N_43703,N_43766);
and U45834 (N_45834,N_42306,N_42737);
nor U45835 (N_45835,N_42242,N_42691);
nand U45836 (N_45836,N_42042,N_43477);
and U45837 (N_45837,N_42489,N_43650);
nor U45838 (N_45838,N_42180,N_43618);
or U45839 (N_45839,N_43516,N_43097);
nor U45840 (N_45840,N_42754,N_43920);
nor U45841 (N_45841,N_42168,N_43423);
nand U45842 (N_45842,N_42989,N_43965);
nor U45843 (N_45843,N_43058,N_42407);
or U45844 (N_45844,N_42363,N_42114);
and U45845 (N_45845,N_42049,N_43861);
or U45846 (N_45846,N_42307,N_43801);
nand U45847 (N_45847,N_42528,N_43553);
nor U45848 (N_45848,N_42239,N_43446);
nor U45849 (N_45849,N_42718,N_42221);
or U45850 (N_45850,N_42410,N_43523);
nand U45851 (N_45851,N_43995,N_43193);
or U45852 (N_45852,N_43414,N_43228);
xor U45853 (N_45853,N_42762,N_42019);
or U45854 (N_45854,N_42236,N_42002);
and U45855 (N_45855,N_42609,N_43999);
nand U45856 (N_45856,N_43801,N_42504);
nor U45857 (N_45857,N_43577,N_42159);
nor U45858 (N_45858,N_42233,N_43067);
nor U45859 (N_45859,N_43855,N_43921);
or U45860 (N_45860,N_43008,N_42969);
nor U45861 (N_45861,N_42980,N_43449);
xor U45862 (N_45862,N_43465,N_42685);
nand U45863 (N_45863,N_43730,N_43253);
or U45864 (N_45864,N_42790,N_43055);
or U45865 (N_45865,N_43396,N_42427);
and U45866 (N_45866,N_42266,N_43097);
xnor U45867 (N_45867,N_43479,N_43158);
nor U45868 (N_45868,N_42609,N_43439);
and U45869 (N_45869,N_43478,N_42138);
nor U45870 (N_45870,N_42400,N_43446);
and U45871 (N_45871,N_43582,N_42953);
and U45872 (N_45872,N_42915,N_42986);
nand U45873 (N_45873,N_42429,N_42825);
and U45874 (N_45874,N_42311,N_43118);
or U45875 (N_45875,N_43818,N_43958);
and U45876 (N_45876,N_43234,N_42717);
or U45877 (N_45877,N_42895,N_43383);
and U45878 (N_45878,N_42896,N_42328);
nand U45879 (N_45879,N_43621,N_43614);
or U45880 (N_45880,N_42424,N_42486);
and U45881 (N_45881,N_43655,N_42491);
nand U45882 (N_45882,N_43615,N_42972);
nor U45883 (N_45883,N_43693,N_42581);
or U45884 (N_45884,N_43681,N_43065);
or U45885 (N_45885,N_43656,N_42308);
and U45886 (N_45886,N_43683,N_43501);
nand U45887 (N_45887,N_43518,N_43344);
or U45888 (N_45888,N_43579,N_43933);
nor U45889 (N_45889,N_42279,N_42461);
and U45890 (N_45890,N_43114,N_43315);
nand U45891 (N_45891,N_42757,N_43769);
and U45892 (N_45892,N_42056,N_43601);
nor U45893 (N_45893,N_42926,N_42295);
or U45894 (N_45894,N_43050,N_43453);
nor U45895 (N_45895,N_43314,N_42911);
or U45896 (N_45896,N_43319,N_42591);
xnor U45897 (N_45897,N_42170,N_42853);
nor U45898 (N_45898,N_43892,N_42046);
nand U45899 (N_45899,N_43956,N_43782);
nand U45900 (N_45900,N_42072,N_42955);
or U45901 (N_45901,N_42805,N_42674);
and U45902 (N_45902,N_42025,N_43358);
nor U45903 (N_45903,N_42418,N_42103);
nor U45904 (N_45904,N_42673,N_43221);
nor U45905 (N_45905,N_42095,N_43229);
or U45906 (N_45906,N_43989,N_43447);
or U45907 (N_45907,N_42427,N_43897);
nand U45908 (N_45908,N_42544,N_43672);
or U45909 (N_45909,N_43739,N_42224);
nand U45910 (N_45910,N_43948,N_42391);
and U45911 (N_45911,N_42140,N_42001);
or U45912 (N_45912,N_42012,N_43439);
or U45913 (N_45913,N_42441,N_43323);
or U45914 (N_45914,N_43568,N_43713);
and U45915 (N_45915,N_43404,N_42018);
nor U45916 (N_45916,N_42061,N_43669);
and U45917 (N_45917,N_43886,N_42278);
nand U45918 (N_45918,N_42993,N_42801);
nor U45919 (N_45919,N_42901,N_43582);
and U45920 (N_45920,N_43536,N_43728);
and U45921 (N_45921,N_43024,N_43585);
or U45922 (N_45922,N_43399,N_42295);
and U45923 (N_45923,N_43493,N_43931);
nand U45924 (N_45924,N_43596,N_42023);
nand U45925 (N_45925,N_43942,N_42790);
and U45926 (N_45926,N_42535,N_42238);
and U45927 (N_45927,N_42283,N_43579);
or U45928 (N_45928,N_43714,N_42208);
xor U45929 (N_45929,N_43857,N_42883);
and U45930 (N_45930,N_42788,N_42455);
or U45931 (N_45931,N_43235,N_43113);
or U45932 (N_45932,N_43331,N_43577);
nand U45933 (N_45933,N_42750,N_43559);
nand U45934 (N_45934,N_43850,N_43381);
nor U45935 (N_45935,N_42766,N_43736);
and U45936 (N_45936,N_42280,N_43086);
and U45937 (N_45937,N_43231,N_43195);
and U45938 (N_45938,N_42348,N_43477);
nor U45939 (N_45939,N_42721,N_42467);
nand U45940 (N_45940,N_42012,N_42907);
nor U45941 (N_45941,N_43562,N_43871);
and U45942 (N_45942,N_43902,N_43054);
nand U45943 (N_45943,N_43709,N_42700);
nor U45944 (N_45944,N_42428,N_43308);
nand U45945 (N_45945,N_43323,N_43898);
nor U45946 (N_45946,N_42703,N_42898);
or U45947 (N_45947,N_42480,N_43668);
xor U45948 (N_45948,N_42395,N_43298);
and U45949 (N_45949,N_42897,N_42797);
and U45950 (N_45950,N_43451,N_43385);
nor U45951 (N_45951,N_42254,N_42624);
nand U45952 (N_45952,N_42708,N_42643);
nor U45953 (N_45953,N_42642,N_43017);
nand U45954 (N_45954,N_43550,N_43883);
xor U45955 (N_45955,N_43608,N_42558);
or U45956 (N_45956,N_43952,N_42920);
and U45957 (N_45957,N_42059,N_43314);
nor U45958 (N_45958,N_43480,N_42110);
or U45959 (N_45959,N_43165,N_42875);
nor U45960 (N_45960,N_42550,N_43773);
nor U45961 (N_45961,N_42506,N_43649);
nor U45962 (N_45962,N_43641,N_43998);
or U45963 (N_45963,N_42001,N_43357);
nor U45964 (N_45964,N_43124,N_43270);
and U45965 (N_45965,N_42985,N_42564);
and U45966 (N_45966,N_42958,N_43863);
and U45967 (N_45967,N_42316,N_42889);
and U45968 (N_45968,N_42021,N_43834);
nand U45969 (N_45969,N_42396,N_42550);
and U45970 (N_45970,N_43066,N_43491);
and U45971 (N_45971,N_43496,N_43419);
nor U45972 (N_45972,N_43480,N_42425);
and U45973 (N_45973,N_43091,N_42342);
or U45974 (N_45974,N_43755,N_43564);
nand U45975 (N_45975,N_42736,N_43470);
nand U45976 (N_45976,N_42848,N_43428);
nand U45977 (N_45977,N_42387,N_43415);
nand U45978 (N_45978,N_43466,N_42863);
and U45979 (N_45979,N_42338,N_43764);
nand U45980 (N_45980,N_42237,N_42537);
or U45981 (N_45981,N_42871,N_42080);
or U45982 (N_45982,N_43130,N_42271);
or U45983 (N_45983,N_42624,N_43200);
or U45984 (N_45984,N_43175,N_42650);
nand U45985 (N_45985,N_42511,N_42348);
and U45986 (N_45986,N_43856,N_42874);
nand U45987 (N_45987,N_43899,N_42744);
and U45988 (N_45988,N_43899,N_42372);
nor U45989 (N_45989,N_42177,N_42866);
and U45990 (N_45990,N_42396,N_42574);
and U45991 (N_45991,N_42301,N_42602);
and U45992 (N_45992,N_42338,N_43381);
and U45993 (N_45993,N_42917,N_42818);
nand U45994 (N_45994,N_43615,N_43966);
and U45995 (N_45995,N_42416,N_42934);
or U45996 (N_45996,N_43703,N_42027);
nand U45997 (N_45997,N_43963,N_42388);
nor U45998 (N_45998,N_42991,N_42362);
or U45999 (N_45999,N_42852,N_42272);
xnor U46000 (N_46000,N_44652,N_44038);
nor U46001 (N_46001,N_44947,N_44369);
nor U46002 (N_46002,N_44164,N_45119);
nor U46003 (N_46003,N_45989,N_45364);
nand U46004 (N_46004,N_45736,N_44791);
or U46005 (N_46005,N_44967,N_45444);
nor U46006 (N_46006,N_44013,N_45828);
nand U46007 (N_46007,N_45913,N_45904);
or U46008 (N_46008,N_44601,N_44669);
or U46009 (N_46009,N_44372,N_45422);
or U46010 (N_46010,N_45966,N_44896);
or U46011 (N_46011,N_44066,N_45584);
or U46012 (N_46012,N_44322,N_44981);
or U46013 (N_46013,N_45852,N_44099);
or U46014 (N_46014,N_45661,N_45432);
and U46015 (N_46015,N_44235,N_44408);
nand U46016 (N_46016,N_45211,N_45405);
or U46017 (N_46017,N_45954,N_45361);
nand U46018 (N_46018,N_45461,N_45009);
or U46019 (N_46019,N_44763,N_45513);
and U46020 (N_46020,N_44506,N_45698);
nand U46021 (N_46021,N_44116,N_45688);
or U46022 (N_46022,N_44646,N_44142);
nand U46023 (N_46023,N_45214,N_45097);
and U46024 (N_46024,N_44217,N_44173);
and U46025 (N_46025,N_45535,N_44167);
or U46026 (N_46026,N_45762,N_44618);
nand U46027 (N_46027,N_45402,N_45225);
nor U46028 (N_46028,N_44027,N_45370);
and U46029 (N_46029,N_45007,N_44931);
nor U46030 (N_46030,N_44089,N_45223);
nor U46031 (N_46031,N_44163,N_44531);
or U46032 (N_46032,N_44168,N_44835);
nand U46033 (N_46033,N_44297,N_44499);
nor U46034 (N_46034,N_45678,N_45433);
and U46035 (N_46035,N_44501,N_45070);
and U46036 (N_46036,N_45343,N_44907);
nand U46037 (N_46037,N_44630,N_44537);
and U46038 (N_46038,N_44274,N_44416);
and U46039 (N_46039,N_44747,N_45887);
nand U46040 (N_46040,N_45118,N_45052);
nor U46041 (N_46041,N_45006,N_44381);
nor U46042 (N_46042,N_44852,N_45266);
and U46043 (N_46043,N_44882,N_44880);
nand U46044 (N_46044,N_44782,N_44776);
nor U46045 (N_46045,N_45699,N_44358);
and U46046 (N_46046,N_44014,N_45991);
or U46047 (N_46047,N_44304,N_44445);
nor U46048 (N_46048,N_44562,N_45808);
nand U46049 (N_46049,N_45591,N_45403);
nor U46050 (N_46050,N_45157,N_44341);
or U46051 (N_46051,N_44334,N_44664);
xnor U46052 (N_46052,N_44197,N_45191);
nor U46053 (N_46053,N_45986,N_44615);
nor U46054 (N_46054,N_44223,N_45572);
nor U46055 (N_46055,N_44527,N_44814);
nor U46056 (N_46056,N_44658,N_45624);
and U46057 (N_46057,N_44177,N_45997);
nand U46058 (N_46058,N_45041,N_45293);
or U46059 (N_46059,N_44820,N_44570);
nand U46060 (N_46060,N_45834,N_45942);
and U46061 (N_46061,N_45278,N_44002);
or U46062 (N_46062,N_45121,N_44312);
nand U46063 (N_46063,N_45716,N_44489);
and U46064 (N_46064,N_45603,N_44236);
and U46065 (N_46065,N_44113,N_44962);
nor U46066 (N_46066,N_45031,N_45084);
nor U46067 (N_46067,N_45515,N_45162);
and U46068 (N_46068,N_44935,N_44143);
nor U46069 (N_46069,N_44017,N_45764);
nor U46070 (N_46070,N_45639,N_45151);
or U46071 (N_46071,N_44022,N_45171);
or U46072 (N_46072,N_45044,N_45181);
nand U46073 (N_46073,N_44873,N_44564);
nand U46074 (N_46074,N_44775,N_44659);
nand U46075 (N_46075,N_45632,N_45496);
nor U46076 (N_46076,N_44594,N_44928);
and U46077 (N_46077,N_44172,N_45096);
nor U46078 (N_46078,N_45105,N_45917);
and U46079 (N_46079,N_45089,N_44878);
or U46080 (N_46080,N_44244,N_45288);
or U46081 (N_46081,N_45216,N_45256);
or U46082 (N_46082,N_44753,N_44488);
or U46083 (N_46083,N_45028,N_45780);
nor U46084 (N_46084,N_44353,N_45335);
and U46085 (N_46085,N_44221,N_44779);
nor U46086 (N_46086,N_44303,N_44342);
and U46087 (N_46087,N_44437,N_45429);
nand U46088 (N_46088,N_44308,N_44587);
nor U46089 (N_46089,N_44714,N_45271);
nor U46090 (N_46090,N_44667,N_45165);
nand U46091 (N_46091,N_44176,N_44491);
or U46092 (N_46092,N_45564,N_45691);
nor U46093 (N_46093,N_44700,N_44202);
nor U46094 (N_46094,N_44592,N_44617);
nand U46095 (N_46095,N_45619,N_44529);
and U46096 (N_46096,N_45366,N_45082);
nand U46097 (N_46097,N_45609,N_45988);
nand U46098 (N_46098,N_45883,N_44711);
and U46099 (N_46099,N_45640,N_45571);
nor U46100 (N_46100,N_45880,N_45693);
and U46101 (N_46101,N_45514,N_44670);
nand U46102 (N_46102,N_44407,N_45312);
nor U46103 (N_46103,N_44251,N_44533);
nor U46104 (N_46104,N_45772,N_45455);
nor U46105 (N_46105,N_44141,N_44378);
or U46106 (N_46106,N_45004,N_45566);
and U46107 (N_46107,N_44530,N_45824);
nand U46108 (N_46108,N_44455,N_45526);
and U46109 (N_46109,N_44641,N_45134);
nand U46110 (N_46110,N_45098,N_44734);
nand U46111 (N_46111,N_44541,N_44335);
or U46112 (N_46112,N_45302,N_44858);
nand U46113 (N_46113,N_44628,N_45941);
nand U46114 (N_46114,N_45295,N_45919);
or U46115 (N_46115,N_45759,N_44538);
or U46116 (N_46116,N_45166,N_45099);
nor U46117 (N_46117,N_45039,N_45869);
xnor U46118 (N_46118,N_44319,N_45814);
or U46119 (N_46119,N_45818,N_44532);
nor U46120 (N_46120,N_44808,N_45209);
nor U46121 (N_46121,N_44123,N_44605);
nand U46122 (N_46122,N_44316,N_45113);
nor U46123 (N_46123,N_44079,N_44082);
and U46124 (N_46124,N_45717,N_44115);
and U46125 (N_46125,N_45695,N_44879);
or U46126 (N_46126,N_44192,N_44213);
or U46127 (N_46127,N_45835,N_45350);
nand U46128 (N_46128,N_44588,N_44366);
nor U46129 (N_46129,N_44229,N_44560);
nor U46130 (N_46130,N_45077,N_44602);
nor U46131 (N_46131,N_45649,N_45809);
nand U46132 (N_46132,N_45358,N_45864);
nand U46133 (N_46133,N_45086,N_45376);
or U46134 (N_46134,N_44902,N_45465);
nand U46135 (N_46135,N_44903,N_44277);
nand U46136 (N_46136,N_44867,N_44625);
and U46137 (N_46137,N_44603,N_44806);
nor U46138 (N_46138,N_44078,N_44462);
nand U46139 (N_46139,N_45657,N_45848);
nor U46140 (N_46140,N_45215,N_45999);
and U46141 (N_46141,N_44200,N_45888);
xnor U46142 (N_46142,N_44466,N_45352);
and U46143 (N_46143,N_44050,N_45222);
and U46144 (N_46144,N_45645,N_45635);
nand U46145 (N_46145,N_44243,N_44608);
nor U46146 (N_46146,N_44152,N_44004);
and U46147 (N_46147,N_44886,N_45479);
nor U46148 (N_46148,N_44222,N_44227);
and U46149 (N_46149,N_45643,N_44616);
nor U46150 (N_46150,N_44490,N_44075);
or U46151 (N_46151,N_45971,N_44346);
or U46152 (N_46152,N_45017,N_44619);
nor U46153 (N_46153,N_44999,N_45247);
nor U46154 (N_46154,N_44895,N_44479);
and U46155 (N_46155,N_44969,N_44385);
nand U46156 (N_46156,N_45368,N_45608);
nor U46157 (N_46157,N_45633,N_45996);
or U46158 (N_46158,N_45722,N_45036);
and U46159 (N_46159,N_45858,N_44812);
and U46160 (N_46160,N_45525,N_45146);
and U46161 (N_46161,N_44629,N_44337);
nor U46162 (N_46162,N_44140,N_45159);
nand U46163 (N_46163,N_45831,N_45062);
nor U46164 (N_46164,N_45682,N_45318);
and U46165 (N_46165,N_45967,N_44803);
and U46166 (N_46166,N_45095,N_45252);
nand U46167 (N_46167,N_45807,N_45180);
and U46168 (N_46168,N_44766,N_44710);
and U46169 (N_46169,N_45841,N_45022);
nand U46170 (N_46170,N_45451,N_45748);
and U46171 (N_46171,N_44675,N_44138);
or U46172 (N_46172,N_45079,N_44118);
and U46173 (N_46173,N_45424,N_45602);
and U46174 (N_46174,N_44047,N_45475);
and U46175 (N_46175,N_44283,N_44190);
nand U46176 (N_46176,N_44522,N_45385);
nor U46177 (N_46177,N_44510,N_45174);
or U46178 (N_46178,N_44175,N_44476);
and U46179 (N_46179,N_44136,N_44211);
or U46180 (N_46180,N_45035,N_44745);
or U46181 (N_46181,N_44234,N_45787);
nor U46182 (N_46182,N_44732,N_45188);
nor U46183 (N_46183,N_45784,N_44707);
or U46184 (N_46184,N_45458,N_45738);
nand U46185 (N_46185,N_45254,N_45933);
nor U46186 (N_46186,N_44733,N_44104);
nand U46187 (N_46187,N_45927,N_45790);
nor U46188 (N_46188,N_44318,N_44454);
nand U46189 (N_46189,N_44627,N_44819);
nand U46190 (N_46190,N_45877,N_44845);
nand U46191 (N_46191,N_44752,N_44925);
or U46192 (N_46192,N_44984,N_44870);
or U46193 (N_46193,N_45969,N_44003);
nor U46194 (N_46194,N_44582,N_45510);
and U46195 (N_46195,N_45241,N_44551);
or U46196 (N_46196,N_45328,N_44827);
nand U46197 (N_46197,N_44585,N_44633);
nand U46198 (N_46198,N_45172,N_45173);
or U46199 (N_46199,N_44860,N_45542);
nand U46200 (N_46200,N_45143,N_45426);
nor U46201 (N_46201,N_44053,N_45186);
nor U46202 (N_46202,N_45272,N_45763);
or U46203 (N_46203,N_45056,N_44150);
nand U46204 (N_46204,N_44894,N_45321);
or U46205 (N_46205,N_44039,N_44284);
or U46206 (N_46206,N_44117,N_44685);
nor U46207 (N_46207,N_45304,N_44362);
nand U46208 (N_46208,N_44974,N_45550);
nand U46209 (N_46209,N_44958,N_45224);
nand U46210 (N_46210,N_45061,N_45894);
nand U46211 (N_46211,N_45504,N_45217);
or U46212 (N_46212,N_45154,N_44414);
and U46213 (N_46213,N_44964,N_44101);
nand U46214 (N_46214,N_44210,N_45248);
or U46215 (N_46215,N_45265,N_44415);
and U46216 (N_46216,N_45005,N_44206);
and U46217 (N_46217,N_45543,N_44948);
and U46218 (N_46218,N_45646,N_45131);
nor U46219 (N_46219,N_45559,N_44924);
or U46220 (N_46220,N_45538,N_45723);
or U46221 (N_46221,N_45604,N_44821);
nand U46222 (N_46222,N_45568,N_44232);
nor U46223 (N_46223,N_44653,N_44281);
or U46224 (N_46224,N_44575,N_45187);
nand U46225 (N_46225,N_44420,N_44373);
and U46226 (N_46226,N_44996,N_44552);
nand U46227 (N_46227,N_44556,N_45669);
nand U46228 (N_46228,N_44398,N_45839);
and U46229 (N_46229,N_45177,N_45727);
or U46230 (N_46230,N_45593,N_44477);
nand U46231 (N_46231,N_44517,N_45903);
nand U46232 (N_46232,N_44239,N_45440);
or U46233 (N_46233,N_44945,N_45298);
nor U46234 (N_46234,N_45779,N_44323);
nand U46235 (N_46235,N_44688,N_44044);
or U46236 (N_46236,N_45218,N_44286);
xnor U46237 (N_46237,N_45970,N_45488);
nor U46238 (N_46238,N_45129,N_45355);
and U46239 (N_46239,N_45711,N_44120);
nor U46240 (N_46240,N_45910,N_45726);
nand U46241 (N_46241,N_44306,N_45946);
nand U46242 (N_46242,N_44650,N_45371);
xnor U46243 (N_46243,N_44822,N_44875);
or U46244 (N_46244,N_44324,N_44704);
or U46245 (N_46245,N_45331,N_45554);
nand U46246 (N_46246,N_45582,N_45753);
nor U46247 (N_46247,N_44139,N_44995);
nand U46248 (N_46248,N_45250,N_44713);
and U46249 (N_46249,N_45008,N_45502);
nand U46250 (N_46250,N_45949,N_44986);
or U46251 (N_46251,N_45430,N_45276);
nor U46252 (N_46252,N_45932,N_44660);
nand U46253 (N_46253,N_44702,N_44638);
and U46254 (N_46254,N_45863,N_44718);
nor U46255 (N_46255,N_44509,N_45414);
and U46256 (N_46256,N_44205,N_44781);
and U46257 (N_46257,N_44149,N_44165);
xnor U46258 (N_46258,N_44057,N_44125);
nand U46259 (N_46259,N_45108,N_44926);
or U46260 (N_46260,N_45704,N_44487);
and U46261 (N_46261,N_44418,N_45378);
nand U46262 (N_46262,N_44481,N_44310);
or U46263 (N_46263,N_44406,N_45742);
nand U46264 (N_46264,N_45629,N_44072);
nor U46265 (N_46265,N_45577,N_45512);
and U46266 (N_46266,N_44112,N_44010);
and U46267 (N_46267,N_44502,N_45494);
nor U46268 (N_46268,N_45655,N_44598);
nor U46269 (N_46269,N_45275,N_45937);
or U46270 (N_46270,N_45911,N_44228);
and U46271 (N_46271,N_44727,N_45387);
or U46272 (N_46272,N_44106,N_44130);
nor U46273 (N_46273,N_44215,N_45322);
nand U46274 (N_46274,N_44467,N_45524);
and U46275 (N_46275,N_45239,N_44196);
or U46276 (N_46276,N_44409,N_44187);
or U46277 (N_46277,N_45957,N_45590);
and U46278 (N_46278,N_44393,N_45269);
nor U46279 (N_46279,N_45194,N_45397);
nor U46280 (N_46280,N_45040,N_44811);
or U46281 (N_46281,N_44518,N_45075);
nand U46282 (N_46282,N_44387,N_44723);
nand U46283 (N_46283,N_44938,N_45487);
nand U46284 (N_46284,N_45558,N_44275);
and U46285 (N_46285,N_44427,N_45963);
nor U46286 (N_46286,N_45102,N_45263);
and U46287 (N_46287,N_45701,N_45588);
xor U46288 (N_46288,N_44203,N_45220);
nor U46289 (N_46289,N_45054,N_45516);
nand U46290 (N_46290,N_45408,N_44842);
nand U46291 (N_46291,N_45483,N_45485);
or U46292 (N_46292,N_45340,N_45020);
or U46293 (N_46293,N_45138,N_45418);
or U46294 (N_46294,N_44258,N_44073);
or U46295 (N_46295,N_44376,N_44290);
nor U46296 (N_46296,N_45536,N_45630);
nand U46297 (N_46297,N_45939,N_45905);
or U46298 (N_46298,N_45560,N_45240);
nand U46299 (N_46299,N_44578,N_45205);
or U46300 (N_46300,N_45115,N_45838);
nand U46301 (N_46301,N_45872,N_45749);
nor U46302 (N_46302,N_45735,N_44500);
nand U46303 (N_46303,N_44549,N_45308);
and U46304 (N_46304,N_44000,N_45406);
nand U46305 (N_46305,N_44024,N_44891);
and U46306 (N_46306,N_44662,N_44829);
xor U46307 (N_46307,N_44268,N_44769);
and U46308 (N_46308,N_44857,N_44679);
or U46309 (N_46309,N_44330,N_44982);
nand U46310 (N_46310,N_44975,N_45766);
and U46311 (N_46311,N_45442,N_45206);
or U46312 (N_46312,N_44729,N_45087);
or U46313 (N_46313,N_44621,N_45407);
and U46314 (N_46314,N_45132,N_45016);
or U46315 (N_46315,N_45931,N_44607);
nand U46316 (N_46316,N_45955,N_45972);
nor U46317 (N_46317,N_44861,N_45384);
nor U46318 (N_46318,N_45725,N_44349);
and U46319 (N_46319,N_45627,N_44712);
nand U46320 (N_46320,N_44987,N_44313);
nand U46321 (N_46321,N_44444,N_45270);
nand U46322 (N_46322,N_45803,N_44034);
and U46323 (N_46323,N_44634,N_45672);
nor U46324 (N_46324,N_44442,N_44350);
nor U46325 (N_46325,N_44831,N_45628);
nor U46326 (N_46326,N_45198,N_44465);
nand U46327 (N_46327,N_45565,N_44171);
nand U46328 (N_46328,N_44657,N_44114);
nand U46329 (N_46329,N_44338,N_44859);
or U46330 (N_46330,N_44897,N_45567);
nand U46331 (N_46331,N_45968,N_44802);
nor U46332 (N_46332,N_44789,N_44755);
nor U46333 (N_46333,N_45169,N_45768);
or U46334 (N_46334,N_45109,N_44065);
nor U46335 (N_46335,N_45100,N_45306);
nand U46336 (N_46336,N_45330,N_44411);
or U46337 (N_46337,N_44833,N_44102);
nor U46338 (N_46338,N_44071,N_44508);
nand U46339 (N_46339,N_44750,N_44944);
nand U46340 (N_46340,N_45032,N_44788);
nand U46341 (N_46341,N_45093,N_45317);
and U46342 (N_46342,N_44435,N_44054);
and U46343 (N_46343,N_45936,N_44119);
and U46344 (N_46344,N_45078,N_44085);
nand U46345 (N_46345,N_44771,N_45066);
xor U46346 (N_46346,N_44854,N_45003);
nor U46347 (N_46347,N_45719,N_44642);
xnor U46348 (N_46348,N_45531,N_45046);
nand U46349 (N_46349,N_44161,N_45897);
nand U46350 (N_46350,N_44193,N_45273);
nor U46351 (N_46351,N_45718,N_45973);
or U46352 (N_46352,N_45987,N_45163);
and U46353 (N_46353,N_45491,N_44365);
nand U46354 (N_46354,N_44890,N_45012);
or U46355 (N_46355,N_44395,N_45601);
nor U46356 (N_46356,N_45319,N_45666);
nand U46357 (N_46357,N_44813,N_45898);
or U46358 (N_46358,N_44514,N_45419);
and U46359 (N_46359,N_45656,N_45092);
nor U46360 (N_46360,N_45325,N_45423);
nor U46361 (N_46361,N_45659,N_45517);
nand U46362 (N_46362,N_44815,N_45329);
nand U46363 (N_46363,N_44741,N_45401);
or U46364 (N_46364,N_44512,N_44298);
and U46365 (N_46365,N_44474,N_44291);
or U46366 (N_46366,N_45421,N_45622);
nand U46367 (N_46367,N_45472,N_45579);
and U46368 (N_46368,N_45416,N_45859);
nand U46369 (N_46369,N_44368,N_45747);
nor U46370 (N_46370,N_45776,N_45679);
nand U46371 (N_46371,N_45861,N_44262);
nor U46372 (N_46372,N_45037,N_45802);
and U46373 (N_46373,N_45156,N_44447);
and U46374 (N_46374,N_45179,N_45739);
nor U46375 (N_46375,N_45333,N_45111);
and U46376 (N_46376,N_44953,N_44147);
nor U46377 (N_46377,N_44916,N_45342);
nand U46378 (N_46378,N_45553,N_44862);
nand U46379 (N_46379,N_44098,N_45389);
nand U46380 (N_46380,N_44849,N_44473);
and U46381 (N_46381,N_45391,N_44965);
and U46382 (N_46382,N_44023,N_45409);
nor U46383 (N_46383,N_44033,N_44901);
and U46384 (N_46384,N_45696,N_45706);
nor U46385 (N_46385,N_45832,N_44932);
or U46386 (N_46386,N_44949,N_45221);
or U46387 (N_46387,N_45529,N_44148);
nand U46388 (N_46388,N_44220,N_45786);
and U46389 (N_46389,N_45375,N_44355);
and U46390 (N_46390,N_44526,N_45482);
nand U46391 (N_46391,N_44425,N_44495);
and U46392 (N_46392,N_45644,N_44269);
nor U46393 (N_46393,N_44485,N_44145);
or U46394 (N_46394,N_45615,N_45168);
nand U46395 (N_46395,N_44701,N_44238);
or U46396 (N_46396,N_45354,N_45120);
nand U46397 (N_46397,N_45404,N_45703);
nor U46398 (N_46398,N_44826,N_44333);
or U46399 (N_46399,N_44056,N_44364);
nand U46400 (N_46400,N_45074,N_44893);
and U46401 (N_46401,N_45654,N_45956);
nor U46402 (N_46402,N_45801,N_44680);
or U46403 (N_46403,N_44441,N_45382);
nor U46404 (N_46404,N_44793,N_44542);
or U46405 (N_46405,N_44955,N_45984);
nand U46406 (N_46406,N_45279,N_45462);
or U46407 (N_46407,N_45773,N_45960);
nand U46408 (N_46408,N_45800,N_45519);
nor U46409 (N_46409,N_45277,N_45653);
nand U46410 (N_46410,N_45122,N_45923);
or U46411 (N_46411,N_45740,N_45744);
and U46412 (N_46412,N_45309,N_45359);
or U46413 (N_46413,N_44272,N_45357);
nand U46414 (N_46414,N_44255,N_45621);
nand U46415 (N_46415,N_44809,N_45561);
nor U46416 (N_46416,N_45842,N_45977);
nor U46417 (N_46417,N_44389,N_44131);
xor U46418 (N_46418,N_45058,N_45799);
nor U46419 (N_46419,N_44716,N_44440);
and U46420 (N_46420,N_44048,N_45822);
or U46421 (N_46421,N_44486,N_45201);
and U46422 (N_46422,N_45332,N_44884);
and U46423 (N_46423,N_44801,N_45815);
and U46424 (N_46424,N_44637,N_45616);
nor U46425 (N_46425,N_45446,N_44064);
or U46426 (N_46426,N_44020,N_45125);
nand U46427 (N_46427,N_44794,N_45344);
or U46428 (N_46428,N_45520,N_45648);
or U46429 (N_46429,N_44108,N_45449);
and U46430 (N_46430,N_45091,N_45733);
nand U46431 (N_46431,N_44746,N_44946);
nor U46432 (N_46432,N_44352,N_45051);
or U46433 (N_46433,N_45985,N_44699);
nand U46434 (N_46434,N_44840,N_44636);
or U46435 (N_46435,N_44844,N_45314);
nand U46436 (N_46436,N_45316,N_44452);
or U46437 (N_46437,N_45895,N_44503);
nor U46438 (N_46438,N_45300,N_44068);
nor U46439 (N_46439,N_45369,N_44158);
nor U46440 (N_46440,N_45025,N_45879);
nand U46441 (N_46441,N_45072,N_44754);
and U46442 (N_46442,N_45994,N_44770);
nor U46443 (N_46443,N_44631,N_45110);
and U46444 (N_46444,N_44865,N_45501);
nor U46445 (N_46445,N_45310,N_44838);
and U46446 (N_46446,N_45785,N_44348);
nor U46447 (N_46447,N_44386,N_44889);
or U46448 (N_46448,N_44124,N_44548);
or U46449 (N_46449,N_45892,N_44070);
nor U46450 (N_46450,N_44841,N_45126);
and U46451 (N_46451,N_45694,N_45088);
nand U46452 (N_46452,N_44345,N_44326);
and U46453 (N_46453,N_45144,N_44683);
nor U46454 (N_46454,N_45618,N_45677);
nand U46455 (N_46455,N_45024,N_45460);
and U46456 (N_46456,N_44980,N_44983);
nand U46457 (N_46457,N_44749,N_45757);
nor U46458 (N_46458,N_44218,N_45683);
and U46459 (N_46459,N_45207,N_44816);
or U46460 (N_46460,N_44302,N_45027);
and U46461 (N_46461,N_44818,N_45843);
or U46462 (N_46462,N_45614,N_44371);
and U46463 (N_46463,N_44122,N_44720);
nand U46464 (N_46464,N_44590,N_45238);
xor U46465 (N_46465,N_45876,N_45208);
or U46466 (N_46466,N_44908,N_44497);
nor U46467 (N_46467,N_45761,N_45523);
nand U46468 (N_46468,N_45063,N_45901);
and U46469 (N_46469,N_44804,N_44824);
nor U46470 (N_46470,N_44706,N_44600);
and U46471 (N_46471,N_45292,N_44558);
or U46472 (N_46472,N_44087,N_44736);
and U46473 (N_46473,N_44709,N_45562);
nand U46474 (N_46474,N_44654,N_45782);
nor U46475 (N_46475,N_44647,N_45244);
nor U46476 (N_46476,N_44520,N_45468);
nand U46477 (N_46477,N_44913,N_44460);
or U46478 (N_46478,N_44757,N_45865);
or U46479 (N_46479,N_45104,N_44383);
nand U46480 (N_46480,N_44606,N_45914);
nor U46481 (N_46481,N_45522,N_44049);
and U46482 (N_46482,N_44651,N_44271);
nor U46483 (N_46483,N_45018,N_44344);
nor U46484 (N_46484,N_45658,N_45705);
and U46485 (N_46485,N_44513,N_44241);
xor U46486 (N_46486,N_45415,N_44478);
nor U46487 (N_46487,N_45990,N_45383);
or U46488 (N_46488,N_45164,N_45867);
nor U46489 (N_46489,N_44001,N_45073);
and U46490 (N_46490,N_44956,N_45160);
or U46491 (N_46491,N_44469,N_45396);
or U46492 (N_46492,N_45544,N_45721);
and U46493 (N_46493,N_45549,N_45612);
or U46494 (N_46494,N_44760,N_44877);
nor U46495 (N_46495,N_44876,N_45975);
or U46496 (N_46496,N_44359,N_44580);
nor U46497 (N_46497,N_44671,N_44567);
nor U46498 (N_46498,N_45282,N_44155);
and U46499 (N_46499,N_44674,N_44129);
nor U46500 (N_46500,N_44851,N_45489);
or U46501 (N_46501,N_44074,N_45611);
and U46502 (N_46502,N_44963,N_44092);
or U46503 (N_46503,N_45230,N_45586);
nor U46504 (N_46504,N_44100,N_44758);
or U46505 (N_46505,N_44263,N_45000);
or U46506 (N_46506,N_45926,N_45650);
or U46507 (N_46507,N_44909,N_45175);
nand U46508 (N_46508,N_44966,N_44086);
or U46509 (N_46509,N_45798,N_44379);
nand U46510 (N_46510,N_45665,N_45459);
and U46511 (N_46511,N_44036,N_44097);
nand U46512 (N_46512,N_45038,N_44620);
and U46513 (N_46513,N_45540,N_45943);
and U46514 (N_46514,N_45065,N_44007);
or U46515 (N_46515,N_44843,N_45953);
or U46516 (N_46516,N_44058,N_45114);
nand U46517 (N_46517,N_44866,N_44640);
and U46518 (N_46518,N_45107,N_44936);
and U46519 (N_46519,N_45057,N_44311);
and U46520 (N_46520,N_44314,N_45837);
or U46521 (N_46521,N_44287,N_45878);
and U46522 (N_46522,N_44692,N_44374);
or U46523 (N_46523,N_45507,N_45234);
nor U46524 (N_46524,N_45147,N_45259);
or U46525 (N_46525,N_44018,N_44059);
nor U46526 (N_46526,N_44848,N_45049);
nor U46527 (N_46527,N_44265,N_45925);
nand U46528 (N_46528,N_44863,N_44786);
and U46529 (N_46529,N_45261,N_45813);
and U46530 (N_46530,N_44246,N_45530);
nor U46531 (N_46531,N_45518,N_44550);
or U46532 (N_46532,N_44971,N_44402);
nand U46533 (N_46533,N_44367,N_45229);
or U46534 (N_46534,N_45885,N_44855);
nand U46535 (N_46535,N_45896,N_44162);
nor U46536 (N_46536,N_45064,N_44032);
and U46537 (N_46537,N_44553,N_44422);
and U46538 (N_46538,N_45992,N_45043);
and U46539 (N_46539,N_44599,N_45023);
and U46540 (N_46540,N_44401,N_45133);
and U46541 (N_46541,N_44546,N_44426);
nor U46542 (N_46542,N_44705,N_44528);
nor U46543 (N_46543,N_45995,N_44030);
or U46544 (N_46544,N_45202,N_44708);
and U46545 (N_46545,N_45532,N_45606);
or U46546 (N_46546,N_44471,N_45882);
nor U46547 (N_46547,N_45924,N_45145);
nand U46548 (N_46548,N_45982,N_45210);
and U46549 (N_46549,N_45908,N_45840);
nor U46550 (N_46550,N_44761,N_45707);
or U46551 (N_46551,N_45581,N_45469);
nand U46552 (N_46552,N_44377,N_44396);
nand U46553 (N_46553,N_44250,N_44604);
nor U46554 (N_46554,N_45527,N_44233);
nand U46555 (N_46555,N_44110,N_45339);
xor U46556 (N_46556,N_44428,N_44224);
nor U46557 (N_46557,N_44219,N_44237);
xnor U46558 (N_46558,N_45103,N_45728);
and U46559 (N_46559,N_45770,N_44189);
or U46560 (N_46560,N_44690,N_45713);
or U46561 (N_46561,N_44774,N_45431);
and U46562 (N_46562,N_45286,N_45441);
nor U46563 (N_46563,N_44293,N_44561);
and U46564 (N_46564,N_45236,N_45870);
nand U46565 (N_46565,N_45687,N_44439);
and U46566 (N_46566,N_44613,N_45817);
nor U46567 (N_46567,N_44691,N_44008);
xnor U46568 (N_46568,N_44195,N_44201);
nand U46569 (N_46569,N_44507,N_44740);
nor U46570 (N_46570,N_44060,N_44951);
nor U46571 (N_46571,N_45373,N_45720);
and U46572 (N_46572,N_45909,N_45280);
or U46573 (N_46573,N_45347,N_45081);
nand U46574 (N_46574,N_44245,N_45466);
nand U46575 (N_46575,N_44037,N_44083);
nor U46576 (N_46576,N_44912,N_44340);
nor U46577 (N_46577,N_45345,N_44317);
or U46578 (N_46578,N_45958,N_45219);
or U46579 (N_46579,N_44109,N_44810);
or U46580 (N_46580,N_45866,N_44950);
or U46581 (N_46581,N_45506,N_44446);
nor U46582 (N_46582,N_44157,N_45737);
nor U46583 (N_46583,N_44035,N_45856);
or U46584 (N_46584,N_45486,N_45456);
nor U46585 (N_46585,N_45819,N_45594);
nand U46586 (N_46586,N_44207,N_45664);
nor U46587 (N_46587,N_44392,N_44388);
nor U46588 (N_46588,N_45673,N_44649);
or U46589 (N_46589,N_44534,N_45771);
or U46590 (N_46590,N_45670,N_44574);
nor U46591 (N_46591,N_45702,N_44762);
and U46592 (N_46592,N_45874,N_44961);
nand U46593 (N_46593,N_44126,N_45313);
and U46594 (N_46594,N_45573,N_44307);
nor U46595 (N_46595,N_45233,N_44156);
nand U46596 (N_46596,N_44724,N_45849);
or U46597 (N_46597,N_45847,N_44656);
or U46598 (N_46598,N_44458,N_45284);
and U46599 (N_46599,N_44009,N_44081);
or U46600 (N_46600,N_45379,N_45124);
nor U46601 (N_46601,N_44360,N_45569);
nand U46602 (N_46602,N_44026,N_45400);
and U46603 (N_46603,N_45681,N_45534);
nor U46604 (N_46604,N_44985,N_45021);
nand U46605 (N_46605,N_45480,N_44170);
and U46606 (N_46606,N_44041,N_45556);
nor U46607 (N_46607,N_44673,N_44273);
nor U46608 (N_46608,N_45474,N_45150);
and U46609 (N_46609,N_44914,N_44850);
nor U46610 (N_46610,N_45756,N_45412);
nor U46611 (N_46611,N_44260,N_44834);
nand U46612 (N_46612,N_45029,N_44703);
nand U46613 (N_46613,N_45551,N_44686);
nand U46614 (N_46614,N_44028,N_45855);
and U46615 (N_46615,N_44301,N_44327);
or U46616 (N_46616,N_44133,N_45945);
nand U46617 (N_46617,N_44461,N_45290);
or U46618 (N_46618,N_44796,N_44519);
nor U46619 (N_46619,N_45047,N_44648);
nand U46620 (N_46620,N_44419,N_45578);
or U46621 (N_46621,N_45090,N_44231);
or U46622 (N_46622,N_44391,N_44256);
nor U46623 (N_46623,N_45101,N_44412);
nand U46624 (N_46624,N_44992,N_45258);
nor U46625 (N_46625,N_44449,N_45792);
nor U46626 (N_46626,N_44780,N_45734);
nand U46627 (N_46627,N_44095,N_44611);
nor U46628 (N_46628,N_45136,N_45710);
and U46629 (N_46629,N_45583,N_45434);
and U46630 (N_46630,N_44132,N_44792);
and U46631 (N_46631,N_44093,N_44463);
and U46632 (N_46632,N_44997,N_45597);
and U46633 (N_46633,N_45048,N_44166);
nand U46634 (N_46634,N_45094,N_45242);
nand U46635 (N_46635,N_44410,N_44790);
and U46636 (N_46636,N_45580,N_45360);
and U46637 (N_46637,N_45916,N_44871);
and U46638 (N_46638,N_44021,N_45311);
or U46639 (N_46639,N_45651,N_44817);
or U46640 (N_46640,N_45123,N_44525);
nand U46641 (N_46641,N_44665,N_45724);
nand U46642 (N_46642,N_45563,N_45854);
nand U46643 (N_46643,N_45684,N_44954);
and U46644 (N_46644,N_45794,N_45576);
nand U46645 (N_46645,N_44635,N_45922);
nand U46646 (N_46646,N_44457,N_44472);
or U46647 (N_46647,N_44137,N_45348);
or U46648 (N_46648,N_44934,N_45503);
nand U46649 (N_46649,N_45393,N_45498);
nor U46650 (N_46650,N_45758,N_45978);
nor U46651 (N_46651,N_44748,N_44225);
or U46652 (N_46652,N_45299,N_45297);
or U46653 (N_46653,N_44178,N_44655);
or U46654 (N_46654,N_44846,N_44839);
nor U46655 (N_46655,N_44390,N_44915);
or U46656 (N_46656,N_45729,N_44063);
nor U46657 (N_46657,N_45961,N_45539);
or U46658 (N_46658,N_44153,N_44693);
nand U46659 (N_46659,N_45437,N_45826);
nand U46660 (N_46660,N_45853,N_45552);
or U46661 (N_46661,N_45690,N_44596);
nand U46662 (N_46662,N_44885,N_44942);
nor U46663 (N_46663,N_44429,N_45775);
and U46664 (N_46664,N_45668,N_44404);
or U46665 (N_46665,N_44728,N_44354);
nor U46666 (N_46666,N_44025,N_44188);
nand U46667 (N_46667,N_45425,N_45274);
nor U46668 (N_46668,N_45700,N_44433);
or U46669 (N_46669,N_44676,N_45034);
nor U46670 (N_46670,N_45463,N_44403);
nand U46671 (N_46671,N_45410,N_44384);
and U46672 (N_46672,N_44257,N_45918);
nand U46673 (N_46673,N_45964,N_44464);
nand U46674 (N_46674,N_44917,N_44544);
or U46675 (N_46675,N_44719,N_45743);
nor U46676 (N_46676,N_45190,N_45010);
or U46677 (N_46677,N_45625,N_45363);
nor U46678 (N_46678,N_45769,N_44547);
or U46679 (N_46679,N_45069,N_45712);
or U46680 (N_46680,N_45184,N_45014);
and U46681 (N_46681,N_44626,N_44248);
nand U46682 (N_46682,N_44181,N_45326);
or U46683 (N_46683,N_44571,N_45754);
nand U46684 (N_46684,N_45938,N_45899);
nor U46685 (N_46685,N_44576,N_44830);
nor U46686 (N_46686,N_45365,N_45767);
nand U46687 (N_46687,N_45731,N_45196);
and U46688 (N_46688,N_45158,N_45857);
nand U46689 (N_46689,N_45490,N_45155);
and U46690 (N_46690,N_44357,N_45447);
and U46691 (N_46691,N_45253,N_44127);
or U46692 (N_46692,N_45499,N_44677);
nand U46693 (N_46693,N_45367,N_44423);
nand U46694 (N_46694,N_45192,N_45438);
nor U46695 (N_46695,N_45294,N_44807);
or U46696 (N_46696,N_45116,N_45574);
and U46697 (N_46697,N_44663,N_45652);
nor U46698 (N_46698,N_45890,N_45613);
nand U46699 (N_46699,N_45183,N_45993);
nor U46700 (N_46700,N_44040,N_45255);
or U46701 (N_46701,N_45541,N_44184);
and U46702 (N_46702,N_44067,N_44212);
and U46703 (N_46703,N_45127,N_44643);
nand U46704 (N_46704,N_44055,N_45338);
nand U46705 (N_46705,N_44998,N_44523);
or U46706 (N_46706,N_44151,N_45481);
and U46707 (N_46707,N_45751,N_44887);
nor U46708 (N_46708,N_45671,N_45471);
and U46709 (N_46709,N_45212,N_45450);
nand U46710 (N_46710,N_44421,N_44778);
and U46711 (N_46711,N_45830,N_44765);
and U46712 (N_46712,N_44622,N_45495);
nor U46713 (N_46713,N_44689,N_45493);
and U46714 (N_46714,N_45200,N_44159);
nor U46715 (N_46715,N_44883,N_44972);
and U46716 (N_46716,N_45500,N_44242);
nor U46717 (N_46717,N_44744,N_45634);
nand U46718 (N_46718,N_45796,N_44483);
nand U46719 (N_46719,N_44105,N_45860);
and U46720 (N_46720,N_45019,N_45497);
or U46721 (N_46721,N_45820,N_44498);
nand U46722 (N_46722,N_45714,N_45059);
nor U46723 (N_46723,N_44666,N_44591);
or U46724 (N_46724,N_45732,N_45912);
nand U46725 (N_46725,N_44535,N_44413);
and U46726 (N_46726,N_44743,N_45781);
or U46727 (N_46727,N_45372,N_45600);
and U46728 (N_46728,N_45998,N_45708);
nand U46729 (N_46729,N_45301,N_44432);
nand U46730 (N_46730,N_44230,N_45777);
and U46731 (N_46731,N_44185,N_44289);
nand U46732 (N_46732,N_44198,N_44279);
nor U46733 (N_46733,N_44276,N_45083);
xnor U46734 (N_46734,N_44989,N_45002);
nor U46735 (N_46735,N_44328,N_44751);
and U46736 (N_46736,N_44730,N_45142);
nand U46737 (N_46737,N_45816,N_44612);
nor U46738 (N_46738,N_44695,N_44991);
or U46739 (N_46739,N_45026,N_44566);
and U46740 (N_46740,N_44595,N_44759);
or U46741 (N_46741,N_44722,N_45589);
or U46742 (N_46742,N_45592,N_44768);
and U46743 (N_46743,N_44448,N_44836);
nor U46744 (N_46744,N_45327,N_45829);
and U46745 (N_46745,N_45380,N_45915);
and U46746 (N_46746,N_44336,N_44016);
nor U46747 (N_46747,N_45033,N_44569);
nor U46748 (N_46748,N_45203,N_45962);
and U46749 (N_46749,N_45011,N_45875);
or U46750 (N_46750,N_44456,N_45934);
nor U46751 (N_46751,N_44103,N_44929);
nor U46752 (N_46752,N_45137,N_45388);
nor U46753 (N_46753,N_45509,N_44043);
nor U46754 (N_46754,N_44480,N_44756);
or U46755 (N_46755,N_44589,N_45030);
or U46756 (N_46756,N_45053,N_44920);
and U46757 (N_46757,N_45685,N_44940);
and U46758 (N_46758,N_45185,N_45246);
or U46759 (N_46759,N_45307,N_45902);
nor U46760 (N_46760,N_45153,N_45140);
nand U46761 (N_46761,N_44267,N_45920);
xnor U46762 (N_46762,N_45470,N_45417);
or U46763 (N_46763,N_44278,N_45871);
nand U46764 (N_46764,N_44405,N_45760);
and U46765 (N_46765,N_44394,N_45076);
nand U46766 (N_46766,N_44668,N_44672);
and U46767 (N_46767,N_44180,N_44259);
and U46768 (N_46768,N_45980,N_45804);
or U46769 (N_46769,N_44990,N_45595);
and U46770 (N_46770,N_45420,N_45055);
or U46771 (N_46771,N_44042,N_45390);
and U46772 (N_46772,N_45929,N_44459);
or U46773 (N_46773,N_44555,N_44343);
nor U46774 (N_46774,N_44717,N_44494);
nand U46775 (N_46775,N_45001,N_44453);
and U46776 (N_46776,N_44905,N_45930);
nor U46777 (N_46777,N_44795,N_45399);
nand U46778 (N_46778,N_44933,N_45952);
nor U46779 (N_46779,N_45686,N_45610);
nor U46780 (N_46780,N_44545,N_44111);
nor U46781 (N_46781,N_45647,N_44417);
nor U46782 (N_46782,N_44511,N_45845);
and U46783 (N_46783,N_44742,N_44644);
nor U46784 (N_46784,N_45130,N_44973);
nand U46785 (N_46785,N_44084,N_45362);
and U46786 (N_46786,N_44696,N_44825);
nor U46787 (N_46787,N_44593,N_45394);
nand U46788 (N_46788,N_45436,N_44247);
and U46789 (N_46789,N_44943,N_44639);
nor U46790 (N_46790,N_44451,N_44261);
and U46791 (N_46791,N_44563,N_45427);
and U46792 (N_46792,N_44096,N_45891);
and U46793 (N_46793,N_44179,N_45453);
nor U46794 (N_46794,N_45492,N_45598);
nand U46795 (N_46795,N_44557,N_45846);
xnor U46796 (N_46796,N_44309,N_45015);
or U46797 (N_46797,N_45085,N_44976);
or U46798 (N_46798,N_44496,N_44698);
or U46799 (N_46799,N_45452,N_44731);
and U46800 (N_46800,N_44475,N_45951);
nand U46801 (N_46801,N_45979,N_45128);
nor U46802 (N_46802,N_44682,N_44543);
xor U46803 (N_46803,N_44584,N_45249);
or U46804 (N_46804,N_45674,N_44524);
or U46805 (N_46805,N_45795,N_44772);
nor U46806 (N_46806,N_44315,N_45473);
xor U46807 (N_46807,N_44226,N_45599);
nor U46808 (N_46808,N_44090,N_45921);
xor U46809 (N_46809,N_44076,N_45139);
nand U46810 (N_46810,N_45283,N_44694);
nor U46811 (N_46811,N_45228,N_44012);
or U46812 (N_46812,N_45730,N_44295);
nand U46813 (N_46813,N_45285,N_44554);
nor U46814 (N_46814,N_44375,N_44434);
nor U46815 (N_46815,N_45398,N_44154);
and U46816 (N_46816,N_45467,N_44253);
and U46817 (N_46817,N_44282,N_45570);
nor U46818 (N_46818,N_45227,N_45605);
nor U46819 (N_46819,N_44978,N_45235);
or U46820 (N_46820,N_45268,N_45377);
and U46821 (N_46821,N_44805,N_44568);
nor U46822 (N_46822,N_44993,N_45413);
nor U46823 (N_46823,N_44370,N_45448);
nor U46824 (N_46824,N_44320,N_44536);
or U46825 (N_46825,N_44382,N_44431);
nand U46826 (N_46826,N_45454,N_45680);
or U46827 (N_46827,N_45245,N_45346);
and U46828 (N_46828,N_44684,N_45850);
nand U46829 (N_46829,N_44169,N_45636);
or U46830 (N_46830,N_45981,N_45893);
nor U46831 (N_46831,N_44174,N_45262);
nor U46832 (N_46832,N_44339,N_44450);
xnor U46833 (N_46833,N_45149,N_44988);
or U46834 (N_46834,N_45323,N_44128);
nor U46835 (N_46835,N_44923,N_44565);
and U46836 (N_46836,N_45213,N_45797);
or U46837 (N_46837,N_45199,N_44031);
nand U46838 (N_46838,N_44351,N_45161);
nand U46839 (N_46839,N_45195,N_44191);
nor U46840 (N_46840,N_44011,N_44052);
nor U46841 (N_46841,N_45783,N_44182);
nand U46842 (N_46842,N_44252,N_44930);
or U46843 (N_46843,N_44186,N_45555);
nor U46844 (N_46844,N_44869,N_45476);
nand U46845 (N_46845,N_44094,N_45287);
nor U46846 (N_46846,N_45545,N_45965);
nand U46847 (N_46847,N_44868,N_44881);
and U46848 (N_46848,N_45944,N_45141);
nand U46849 (N_46849,N_45193,N_44121);
nand U46850 (N_46850,N_44828,N_44784);
xnor U46851 (N_46851,N_44146,N_45013);
nand U46852 (N_46852,N_45585,N_44853);
nor U46853 (N_46853,N_44468,N_44735);
nor U46854 (N_46854,N_45715,N_44739);
nand U46855 (N_46855,N_44624,N_45521);
or U46856 (N_46856,N_44356,N_44296);
nand U46857 (N_46857,N_45948,N_44077);
nand U46858 (N_46858,N_44919,N_45789);
nor U46859 (N_46859,N_44539,N_44632);
nand U46860 (N_46860,N_44847,N_44069);
nor U46861 (N_46861,N_45868,N_44921);
or U46862 (N_46862,N_45257,N_45623);
nand U46863 (N_46863,N_45778,N_45428);
and U46864 (N_46864,N_45435,N_45642);
nand U46865 (N_46865,N_45303,N_44493);
nor U46866 (N_46866,N_44515,N_44721);
and U46867 (N_46867,N_45464,N_44204);
nand U46868 (N_46868,N_45443,N_44134);
and U46869 (N_46869,N_44783,N_45662);
and U46870 (N_46870,N_44363,N_45907);
nand U46871 (N_46871,N_45477,N_44968);
or U46872 (N_46872,N_44209,N_45697);
nor U46873 (N_46873,N_45264,N_45548);
nand U46874 (N_46874,N_44091,N_45660);
or U46875 (N_46875,N_44798,N_45755);
nand U46876 (N_46876,N_45152,N_44505);
nand U46877 (N_46877,N_45900,N_44299);
and U46878 (N_46878,N_45825,N_44199);
or U46879 (N_46879,N_45148,N_45935);
or U46880 (N_46880,N_45774,N_45827);
and U46881 (N_46881,N_44160,N_44773);
nand U46882 (N_46882,N_44872,N_45356);
or U46883 (N_46883,N_44725,N_44577);
nor U46884 (N_46884,N_44957,N_44959);
nand U46885 (N_46885,N_45296,N_45267);
nor U46886 (N_46886,N_45631,N_44911);
nor U46887 (N_46887,N_44300,N_45176);
and U46888 (N_46888,N_44697,N_44332);
or U46889 (N_46889,N_45231,N_45508);
nand U46890 (N_46890,N_44424,N_45976);
or U46891 (N_46891,N_44994,N_45547);
or U46892 (N_46892,N_45511,N_45291);
or U46893 (N_46893,N_45663,N_45884);
and U46894 (N_46894,N_44888,N_45626);
nor U46895 (N_46895,N_44280,N_45505);
nor U46896 (N_46896,N_45042,N_44006);
nand U46897 (N_46897,N_44610,N_44979);
or U46898 (N_46898,N_44484,N_44046);
or U46899 (N_46899,N_44952,N_45806);
or U46900 (N_46900,N_44321,N_45689);
and U46901 (N_46901,N_45045,N_45315);
nor U46902 (N_46902,N_45226,N_44438);
nand U46903 (N_46903,N_45533,N_45823);
nand U46904 (N_46904,N_44623,N_45862);
or U46905 (N_46905,N_45940,N_45745);
and U46906 (N_46906,N_45112,N_45752);
or U46907 (N_46907,N_44687,N_45793);
nand U46908 (N_46908,N_45675,N_44144);
and U46909 (N_46909,N_44436,N_45341);
and U46910 (N_46910,N_45289,N_45439);
and U46911 (N_46911,N_44586,N_45305);
nor U46912 (N_46912,N_45060,N_44572);
nor U46913 (N_46913,N_45237,N_45068);
or U46914 (N_46914,N_45765,N_45620);
or U46915 (N_46915,N_45546,N_45320);
or U46916 (N_46916,N_45607,N_44107);
nand U46917 (N_46917,N_45478,N_44941);
nor U46918 (N_46918,N_44521,N_45182);
and U46919 (N_46919,N_44785,N_44579);
nor U46920 (N_46920,N_44019,N_44504);
nand U46921 (N_46921,N_45178,N_45484);
xor U46922 (N_46922,N_45537,N_44937);
nor U46923 (N_46923,N_45873,N_44874);
or U46924 (N_46924,N_45197,N_44080);
xor U46925 (N_46925,N_45950,N_45189);
and U46926 (N_46926,N_44285,N_44264);
nand U46927 (N_46927,N_44194,N_44906);
or U46928 (N_46928,N_44678,N_44767);
and U46929 (N_46929,N_45336,N_45886);
nand U46930 (N_46930,N_45750,N_44764);
nor U46931 (N_46931,N_45821,N_45667);
nand U46932 (N_46932,N_44292,N_45374);
and U46933 (N_46933,N_44681,N_44399);
or U46934 (N_46934,N_44015,N_44208);
nor U46935 (N_46935,N_44347,N_44266);
and U46936 (N_46936,N_44061,N_44977);
nor U46937 (N_46937,N_44540,N_44240);
nor U46938 (N_46938,N_44005,N_44799);
nand U46939 (N_46939,N_45974,N_44892);
nor U46940 (N_46940,N_45889,N_45080);
or U46941 (N_46941,N_44135,N_45324);
and U46942 (N_46942,N_45392,N_44305);
nor U46943 (N_46943,N_44270,N_45528);
nand U46944 (N_46944,N_44910,N_45457);
and U46945 (N_46945,N_44645,N_45709);
and U46946 (N_46946,N_45353,N_45638);
or U46947 (N_46947,N_45334,N_44939);
nand U46948 (N_46948,N_44088,N_44400);
or U46949 (N_46949,N_44900,N_45251);
nand U46950 (N_46950,N_45959,N_44581);
or U46951 (N_46951,N_45349,N_45617);
nand U46952 (N_46952,N_44661,N_45676);
nand U46953 (N_46953,N_45260,N_45811);
and U46954 (N_46954,N_44797,N_44960);
xnor U46955 (N_46955,N_44516,N_45445);
nand U46956 (N_46956,N_45810,N_44904);
xor U46957 (N_46957,N_44294,N_45337);
or U46958 (N_46958,N_44492,N_44470);
nor U46959 (N_46959,N_44609,N_45411);
and U46960 (N_46960,N_44927,N_45351);
nor U46961 (N_46961,N_44837,N_45170);
nor U46962 (N_46962,N_44331,N_44214);
and U46963 (N_46963,N_44583,N_45692);
nor U46964 (N_46964,N_44597,N_44482);
nor U46965 (N_46965,N_45596,N_44922);
or U46966 (N_46966,N_44361,N_44737);
and U46967 (N_46967,N_45812,N_44329);
xor U46968 (N_46968,N_45906,N_45587);
nor U46969 (N_46969,N_45071,N_44856);
nand U46970 (N_46970,N_45805,N_44430);
nand U46971 (N_46971,N_44045,N_44062);
nor U46972 (N_46972,N_45395,N_45741);
and U46973 (N_46973,N_44573,N_44800);
or U46974 (N_46974,N_45791,N_45836);
xor U46975 (N_46975,N_44918,N_45575);
nor U46976 (N_46976,N_44443,N_45117);
nand U46977 (N_46977,N_44325,N_44288);
and U46978 (N_46978,N_45381,N_45135);
or U46979 (N_46979,N_45928,N_45833);
or U46980 (N_46980,N_44614,N_44380);
nand U46981 (N_46981,N_45983,N_45050);
and U46982 (N_46982,N_44254,N_45881);
nor U46983 (N_46983,N_45641,N_44397);
and U46984 (N_46984,N_44715,N_45386);
nor U46985 (N_46985,N_44183,N_45844);
nor U46986 (N_46986,N_44738,N_44823);
nand U46987 (N_46987,N_45204,N_44777);
or U46988 (N_46988,N_44726,N_45232);
nand U46989 (N_46989,N_44029,N_45637);
and U46990 (N_46990,N_44832,N_44898);
and U46991 (N_46991,N_44559,N_45746);
nor U46992 (N_46992,N_44787,N_44216);
and U46993 (N_46993,N_45106,N_44970);
nand U46994 (N_46994,N_45947,N_44899);
and U46995 (N_46995,N_45243,N_45167);
nand U46996 (N_46996,N_45067,N_45557);
nand U46997 (N_46997,N_44864,N_45281);
nand U46998 (N_46998,N_45788,N_44249);
or U46999 (N_46999,N_45851,N_44051);
nand U47000 (N_47000,N_45488,N_44897);
nand U47001 (N_47001,N_45146,N_44565);
or U47002 (N_47002,N_44239,N_45900);
nand U47003 (N_47003,N_45875,N_44115);
or U47004 (N_47004,N_45323,N_44204);
nand U47005 (N_47005,N_45875,N_44529);
and U47006 (N_47006,N_45633,N_44116);
or U47007 (N_47007,N_44062,N_44058);
nor U47008 (N_47008,N_44600,N_45287);
nor U47009 (N_47009,N_45891,N_45419);
xor U47010 (N_47010,N_45165,N_45609);
nand U47011 (N_47011,N_45606,N_44330);
and U47012 (N_47012,N_45809,N_44631);
nand U47013 (N_47013,N_44661,N_45842);
and U47014 (N_47014,N_45968,N_44671);
or U47015 (N_47015,N_44059,N_44272);
nand U47016 (N_47016,N_45742,N_44532);
nand U47017 (N_47017,N_45334,N_44457);
and U47018 (N_47018,N_45408,N_44091);
and U47019 (N_47019,N_44735,N_45681);
and U47020 (N_47020,N_45360,N_44449);
or U47021 (N_47021,N_44771,N_45909);
or U47022 (N_47022,N_44748,N_44863);
nand U47023 (N_47023,N_45914,N_45572);
nor U47024 (N_47024,N_45167,N_45467);
or U47025 (N_47025,N_45732,N_44363);
or U47026 (N_47026,N_44323,N_45725);
nor U47027 (N_47027,N_45897,N_44772);
nor U47028 (N_47028,N_44249,N_44367);
nand U47029 (N_47029,N_44630,N_44645);
nor U47030 (N_47030,N_44397,N_44851);
or U47031 (N_47031,N_45005,N_44241);
or U47032 (N_47032,N_45551,N_44950);
or U47033 (N_47033,N_44129,N_45038);
nor U47034 (N_47034,N_44470,N_45706);
and U47035 (N_47035,N_44693,N_44614);
nand U47036 (N_47036,N_44201,N_44991);
nor U47037 (N_47037,N_45668,N_45580);
or U47038 (N_47038,N_45854,N_44171);
nor U47039 (N_47039,N_44114,N_44154);
nor U47040 (N_47040,N_45881,N_45337);
nand U47041 (N_47041,N_44701,N_44667);
nor U47042 (N_47042,N_45479,N_44970);
or U47043 (N_47043,N_45116,N_45792);
nor U47044 (N_47044,N_45317,N_45940);
nand U47045 (N_47045,N_45170,N_44026);
nand U47046 (N_47046,N_45968,N_44795);
or U47047 (N_47047,N_44158,N_45750);
nand U47048 (N_47048,N_44178,N_44552);
or U47049 (N_47049,N_45662,N_45705);
nand U47050 (N_47050,N_45867,N_45787);
nor U47051 (N_47051,N_44058,N_44279);
or U47052 (N_47052,N_44908,N_44661);
and U47053 (N_47053,N_45695,N_45266);
nand U47054 (N_47054,N_44048,N_44774);
nand U47055 (N_47055,N_44772,N_44854);
or U47056 (N_47056,N_45992,N_44360);
nand U47057 (N_47057,N_44362,N_44102);
or U47058 (N_47058,N_44435,N_45226);
nor U47059 (N_47059,N_44535,N_44756);
nor U47060 (N_47060,N_44749,N_45030);
and U47061 (N_47061,N_45278,N_44605);
and U47062 (N_47062,N_45365,N_44121);
and U47063 (N_47063,N_45515,N_44348);
nand U47064 (N_47064,N_45148,N_44881);
nor U47065 (N_47065,N_44898,N_45190);
nor U47066 (N_47066,N_44390,N_44906);
nand U47067 (N_47067,N_44830,N_45573);
or U47068 (N_47068,N_44484,N_45162);
nand U47069 (N_47069,N_45125,N_44086);
nor U47070 (N_47070,N_44112,N_44516);
and U47071 (N_47071,N_45043,N_44437);
nor U47072 (N_47072,N_44534,N_45308);
and U47073 (N_47073,N_44907,N_44811);
nor U47074 (N_47074,N_44739,N_45208);
nor U47075 (N_47075,N_45104,N_45636);
and U47076 (N_47076,N_44670,N_44863);
nor U47077 (N_47077,N_45291,N_44622);
nor U47078 (N_47078,N_45568,N_44882);
and U47079 (N_47079,N_44468,N_45999);
xor U47080 (N_47080,N_45090,N_45116);
or U47081 (N_47081,N_44563,N_44325);
or U47082 (N_47082,N_45517,N_45361);
or U47083 (N_47083,N_45331,N_45667);
and U47084 (N_47084,N_44611,N_45431);
xor U47085 (N_47085,N_45327,N_45217);
or U47086 (N_47086,N_45832,N_45916);
nor U47087 (N_47087,N_44074,N_45006);
and U47088 (N_47088,N_44310,N_44862);
nand U47089 (N_47089,N_45101,N_45736);
and U47090 (N_47090,N_45227,N_44326);
and U47091 (N_47091,N_44237,N_45103);
and U47092 (N_47092,N_44369,N_44736);
nand U47093 (N_47093,N_44036,N_45864);
and U47094 (N_47094,N_44159,N_44764);
nor U47095 (N_47095,N_45390,N_45850);
or U47096 (N_47096,N_45087,N_45293);
nor U47097 (N_47097,N_45973,N_44781);
and U47098 (N_47098,N_45423,N_45938);
nand U47099 (N_47099,N_45198,N_44299);
nor U47100 (N_47100,N_44714,N_44353);
and U47101 (N_47101,N_44931,N_44333);
nand U47102 (N_47102,N_45931,N_44125);
nand U47103 (N_47103,N_45892,N_44995);
or U47104 (N_47104,N_44646,N_45674);
nand U47105 (N_47105,N_44176,N_45364);
and U47106 (N_47106,N_45512,N_44359);
or U47107 (N_47107,N_45402,N_45195);
nand U47108 (N_47108,N_44173,N_45616);
or U47109 (N_47109,N_44506,N_44143);
or U47110 (N_47110,N_44489,N_44641);
or U47111 (N_47111,N_44151,N_44803);
and U47112 (N_47112,N_45855,N_44974);
or U47113 (N_47113,N_45404,N_45018);
nor U47114 (N_47114,N_44314,N_45430);
nor U47115 (N_47115,N_44466,N_45475);
or U47116 (N_47116,N_45326,N_44577);
nand U47117 (N_47117,N_44759,N_45899);
or U47118 (N_47118,N_44840,N_45285);
nand U47119 (N_47119,N_45667,N_44274);
and U47120 (N_47120,N_44008,N_45206);
nand U47121 (N_47121,N_44440,N_44931);
nand U47122 (N_47122,N_45341,N_44859);
or U47123 (N_47123,N_44421,N_44231);
and U47124 (N_47124,N_45993,N_44901);
nor U47125 (N_47125,N_44635,N_45928);
nor U47126 (N_47126,N_44731,N_44310);
or U47127 (N_47127,N_44297,N_44891);
and U47128 (N_47128,N_44020,N_45442);
and U47129 (N_47129,N_44776,N_44411);
and U47130 (N_47130,N_44946,N_45178);
nor U47131 (N_47131,N_45443,N_45526);
nand U47132 (N_47132,N_45312,N_45480);
xor U47133 (N_47133,N_44676,N_45601);
nand U47134 (N_47134,N_44316,N_45993);
nand U47135 (N_47135,N_45396,N_44756);
and U47136 (N_47136,N_44458,N_44866);
or U47137 (N_47137,N_44525,N_44181);
and U47138 (N_47138,N_44297,N_45202);
or U47139 (N_47139,N_45177,N_45948);
nor U47140 (N_47140,N_45680,N_44172);
and U47141 (N_47141,N_44730,N_44750);
and U47142 (N_47142,N_45475,N_45693);
nor U47143 (N_47143,N_44537,N_45452);
and U47144 (N_47144,N_44418,N_45597);
or U47145 (N_47145,N_44707,N_44959);
or U47146 (N_47146,N_44640,N_45934);
or U47147 (N_47147,N_44850,N_45729);
or U47148 (N_47148,N_45727,N_44650);
and U47149 (N_47149,N_45816,N_45355);
nor U47150 (N_47150,N_45775,N_45394);
or U47151 (N_47151,N_45730,N_44364);
nor U47152 (N_47152,N_45762,N_44810);
and U47153 (N_47153,N_45556,N_45135);
nand U47154 (N_47154,N_44029,N_44466);
and U47155 (N_47155,N_44776,N_44308);
nor U47156 (N_47156,N_45632,N_45298);
and U47157 (N_47157,N_45269,N_44552);
or U47158 (N_47158,N_45536,N_44998);
nor U47159 (N_47159,N_45062,N_45936);
nand U47160 (N_47160,N_45227,N_44278);
nand U47161 (N_47161,N_44925,N_44727);
nor U47162 (N_47162,N_45829,N_44018);
xor U47163 (N_47163,N_44258,N_44877);
nor U47164 (N_47164,N_45521,N_45341);
and U47165 (N_47165,N_45984,N_44028);
and U47166 (N_47166,N_44174,N_44562);
nor U47167 (N_47167,N_44844,N_45256);
or U47168 (N_47168,N_44372,N_44889);
nand U47169 (N_47169,N_44217,N_44094);
nor U47170 (N_47170,N_44944,N_44532);
nand U47171 (N_47171,N_44389,N_44939);
nand U47172 (N_47172,N_44739,N_45276);
nand U47173 (N_47173,N_44439,N_45993);
nor U47174 (N_47174,N_44720,N_44916);
and U47175 (N_47175,N_45929,N_44618);
nand U47176 (N_47176,N_45318,N_44837);
and U47177 (N_47177,N_45410,N_45953);
or U47178 (N_47178,N_44710,N_45617);
and U47179 (N_47179,N_44469,N_45572);
or U47180 (N_47180,N_45070,N_44857);
and U47181 (N_47181,N_45816,N_45096);
or U47182 (N_47182,N_45478,N_44101);
nand U47183 (N_47183,N_44065,N_45043);
or U47184 (N_47184,N_44245,N_45525);
nor U47185 (N_47185,N_44985,N_45822);
nor U47186 (N_47186,N_44271,N_45439);
or U47187 (N_47187,N_45660,N_44650);
or U47188 (N_47188,N_44961,N_44387);
or U47189 (N_47189,N_44558,N_44768);
or U47190 (N_47190,N_45005,N_44311);
and U47191 (N_47191,N_44434,N_45939);
nand U47192 (N_47192,N_45515,N_45916);
nor U47193 (N_47193,N_44596,N_45062);
nand U47194 (N_47194,N_45186,N_45696);
and U47195 (N_47195,N_44814,N_45260);
and U47196 (N_47196,N_44715,N_44845);
and U47197 (N_47197,N_45524,N_44810);
or U47198 (N_47198,N_45251,N_45439);
and U47199 (N_47199,N_44041,N_45769);
nor U47200 (N_47200,N_45167,N_44009);
xnor U47201 (N_47201,N_45956,N_44371);
nor U47202 (N_47202,N_44304,N_45327);
nor U47203 (N_47203,N_45818,N_44543);
and U47204 (N_47204,N_45257,N_44953);
nand U47205 (N_47205,N_45691,N_45938);
or U47206 (N_47206,N_45503,N_45913);
nor U47207 (N_47207,N_45914,N_45713);
nor U47208 (N_47208,N_45755,N_44409);
nand U47209 (N_47209,N_45402,N_45956);
or U47210 (N_47210,N_45095,N_45737);
nand U47211 (N_47211,N_45560,N_44917);
nand U47212 (N_47212,N_44443,N_44354);
nand U47213 (N_47213,N_44170,N_45234);
nand U47214 (N_47214,N_45548,N_45671);
or U47215 (N_47215,N_44694,N_44571);
or U47216 (N_47216,N_44265,N_45919);
nor U47217 (N_47217,N_44309,N_44615);
and U47218 (N_47218,N_45921,N_44047);
nand U47219 (N_47219,N_44891,N_44529);
nor U47220 (N_47220,N_45798,N_44674);
or U47221 (N_47221,N_44021,N_44110);
xor U47222 (N_47222,N_45961,N_45033);
nand U47223 (N_47223,N_45071,N_44308);
nor U47224 (N_47224,N_44740,N_44625);
xor U47225 (N_47225,N_45566,N_44638);
and U47226 (N_47226,N_44469,N_45363);
nor U47227 (N_47227,N_45951,N_44855);
nand U47228 (N_47228,N_44948,N_45712);
or U47229 (N_47229,N_45252,N_45278);
nand U47230 (N_47230,N_44540,N_44672);
and U47231 (N_47231,N_45462,N_45039);
or U47232 (N_47232,N_45144,N_44976);
xor U47233 (N_47233,N_44586,N_45242);
nor U47234 (N_47234,N_44321,N_45790);
or U47235 (N_47235,N_44635,N_45112);
or U47236 (N_47236,N_45892,N_44072);
and U47237 (N_47237,N_44384,N_44772);
nor U47238 (N_47238,N_44679,N_44620);
or U47239 (N_47239,N_44717,N_44782);
nor U47240 (N_47240,N_44090,N_45491);
nand U47241 (N_47241,N_44547,N_45300);
nand U47242 (N_47242,N_44805,N_44888);
nand U47243 (N_47243,N_44256,N_44801);
nand U47244 (N_47244,N_44635,N_45142);
or U47245 (N_47245,N_45895,N_45071);
and U47246 (N_47246,N_45836,N_44826);
nand U47247 (N_47247,N_45480,N_45292);
nor U47248 (N_47248,N_44107,N_44695);
nand U47249 (N_47249,N_45627,N_45305);
xnor U47250 (N_47250,N_44633,N_44582);
or U47251 (N_47251,N_45929,N_44311);
xnor U47252 (N_47252,N_45716,N_45515);
and U47253 (N_47253,N_44527,N_45407);
nand U47254 (N_47254,N_44609,N_45726);
nand U47255 (N_47255,N_44271,N_45944);
and U47256 (N_47256,N_45581,N_45973);
or U47257 (N_47257,N_45924,N_45993);
nand U47258 (N_47258,N_45023,N_44211);
nand U47259 (N_47259,N_45568,N_45262);
or U47260 (N_47260,N_44842,N_45576);
nor U47261 (N_47261,N_45452,N_45958);
nor U47262 (N_47262,N_44530,N_44411);
nand U47263 (N_47263,N_45800,N_45132);
or U47264 (N_47264,N_44702,N_44603);
or U47265 (N_47265,N_44302,N_45988);
nand U47266 (N_47266,N_44211,N_45253);
and U47267 (N_47267,N_45357,N_45828);
nor U47268 (N_47268,N_44821,N_44104);
or U47269 (N_47269,N_44574,N_45776);
nand U47270 (N_47270,N_44894,N_45788);
and U47271 (N_47271,N_44016,N_45756);
and U47272 (N_47272,N_45484,N_44724);
nor U47273 (N_47273,N_44384,N_44099);
nor U47274 (N_47274,N_45666,N_45917);
nor U47275 (N_47275,N_44372,N_45338);
nor U47276 (N_47276,N_45209,N_45010);
and U47277 (N_47277,N_44133,N_45674);
or U47278 (N_47278,N_44065,N_44357);
nor U47279 (N_47279,N_45957,N_44274);
and U47280 (N_47280,N_44941,N_44011);
and U47281 (N_47281,N_45617,N_44194);
or U47282 (N_47282,N_45115,N_45399);
and U47283 (N_47283,N_45997,N_45973);
or U47284 (N_47284,N_45032,N_45112);
or U47285 (N_47285,N_45885,N_45009);
and U47286 (N_47286,N_44004,N_44029);
nand U47287 (N_47287,N_45717,N_44308);
and U47288 (N_47288,N_45975,N_45679);
nor U47289 (N_47289,N_44015,N_44746);
nand U47290 (N_47290,N_44593,N_44191);
nor U47291 (N_47291,N_45362,N_44215);
and U47292 (N_47292,N_44079,N_44850);
nor U47293 (N_47293,N_44462,N_45276);
xor U47294 (N_47294,N_44953,N_45151);
or U47295 (N_47295,N_45500,N_44249);
or U47296 (N_47296,N_44221,N_44659);
and U47297 (N_47297,N_45811,N_44696);
or U47298 (N_47298,N_45600,N_45758);
nand U47299 (N_47299,N_44925,N_45527);
nor U47300 (N_47300,N_44699,N_45737);
nor U47301 (N_47301,N_45373,N_44075);
or U47302 (N_47302,N_45726,N_44547);
xor U47303 (N_47303,N_44131,N_44775);
nand U47304 (N_47304,N_44212,N_45365);
nand U47305 (N_47305,N_45094,N_44489);
nor U47306 (N_47306,N_44894,N_44184);
nand U47307 (N_47307,N_45409,N_45834);
or U47308 (N_47308,N_45769,N_45777);
nand U47309 (N_47309,N_45596,N_45190);
nor U47310 (N_47310,N_44059,N_45471);
or U47311 (N_47311,N_44019,N_44074);
or U47312 (N_47312,N_44052,N_45034);
and U47313 (N_47313,N_44506,N_44552);
or U47314 (N_47314,N_45877,N_45271);
or U47315 (N_47315,N_44414,N_45782);
nand U47316 (N_47316,N_45623,N_44326);
and U47317 (N_47317,N_44573,N_45574);
nand U47318 (N_47318,N_44734,N_45679);
nand U47319 (N_47319,N_44001,N_44587);
nor U47320 (N_47320,N_45783,N_44889);
and U47321 (N_47321,N_45526,N_44934);
and U47322 (N_47322,N_44701,N_44025);
nand U47323 (N_47323,N_44107,N_44013);
nor U47324 (N_47324,N_45116,N_45397);
nand U47325 (N_47325,N_45277,N_45122);
nand U47326 (N_47326,N_45924,N_45875);
or U47327 (N_47327,N_44121,N_45272);
nor U47328 (N_47328,N_45791,N_45302);
nor U47329 (N_47329,N_44611,N_44509);
nor U47330 (N_47330,N_45255,N_44208);
nor U47331 (N_47331,N_45730,N_45880);
nor U47332 (N_47332,N_45042,N_45318);
nor U47333 (N_47333,N_44469,N_45181);
nand U47334 (N_47334,N_45181,N_44217);
and U47335 (N_47335,N_45821,N_45844);
or U47336 (N_47336,N_45900,N_45448);
and U47337 (N_47337,N_45532,N_44725);
xnor U47338 (N_47338,N_45424,N_44755);
nor U47339 (N_47339,N_45311,N_45770);
nand U47340 (N_47340,N_44946,N_44209);
and U47341 (N_47341,N_44702,N_44692);
nor U47342 (N_47342,N_45564,N_44620);
xor U47343 (N_47343,N_45253,N_44924);
nand U47344 (N_47344,N_44159,N_45617);
nor U47345 (N_47345,N_45828,N_44856);
or U47346 (N_47346,N_45460,N_45056);
and U47347 (N_47347,N_44052,N_45555);
nor U47348 (N_47348,N_45372,N_44467);
and U47349 (N_47349,N_44323,N_44213);
or U47350 (N_47350,N_44523,N_44317);
nand U47351 (N_47351,N_44867,N_45762);
and U47352 (N_47352,N_45840,N_44683);
or U47353 (N_47353,N_45044,N_44514);
and U47354 (N_47354,N_45107,N_44869);
nor U47355 (N_47355,N_45372,N_44485);
or U47356 (N_47356,N_44137,N_45644);
and U47357 (N_47357,N_44875,N_44361);
or U47358 (N_47358,N_44837,N_45643);
or U47359 (N_47359,N_45581,N_45752);
nor U47360 (N_47360,N_44341,N_45530);
or U47361 (N_47361,N_45043,N_45141);
nor U47362 (N_47362,N_44918,N_45613);
nor U47363 (N_47363,N_45805,N_45405);
nor U47364 (N_47364,N_44890,N_44830);
nand U47365 (N_47365,N_45406,N_45625);
or U47366 (N_47366,N_44940,N_44684);
and U47367 (N_47367,N_44523,N_44366);
nand U47368 (N_47368,N_45415,N_44858);
nor U47369 (N_47369,N_45302,N_45184);
or U47370 (N_47370,N_45935,N_44285);
nor U47371 (N_47371,N_44575,N_44634);
nand U47372 (N_47372,N_44292,N_44466);
and U47373 (N_47373,N_44644,N_45132);
or U47374 (N_47374,N_44789,N_44229);
nor U47375 (N_47375,N_45105,N_45770);
nor U47376 (N_47376,N_44030,N_45442);
and U47377 (N_47377,N_45864,N_44796);
nand U47378 (N_47378,N_44594,N_45540);
nor U47379 (N_47379,N_45095,N_45434);
and U47380 (N_47380,N_45081,N_44994);
nor U47381 (N_47381,N_45115,N_44873);
or U47382 (N_47382,N_45827,N_44926);
and U47383 (N_47383,N_44157,N_44813);
nand U47384 (N_47384,N_44811,N_45147);
and U47385 (N_47385,N_45551,N_44051);
or U47386 (N_47386,N_45181,N_45539);
or U47387 (N_47387,N_45949,N_44175);
or U47388 (N_47388,N_44921,N_45473);
nand U47389 (N_47389,N_45511,N_45981);
nor U47390 (N_47390,N_44751,N_44519);
or U47391 (N_47391,N_45063,N_44610);
nand U47392 (N_47392,N_45937,N_44451);
or U47393 (N_47393,N_45911,N_44802);
nor U47394 (N_47394,N_45778,N_45124);
nor U47395 (N_47395,N_45648,N_44903);
or U47396 (N_47396,N_45491,N_45357);
nand U47397 (N_47397,N_45031,N_44159);
nand U47398 (N_47398,N_45237,N_45086);
and U47399 (N_47399,N_44424,N_45370);
nand U47400 (N_47400,N_45701,N_45603);
or U47401 (N_47401,N_45712,N_44086);
nor U47402 (N_47402,N_44789,N_45637);
xor U47403 (N_47403,N_44670,N_45866);
or U47404 (N_47404,N_45056,N_44579);
xnor U47405 (N_47405,N_44527,N_44183);
and U47406 (N_47406,N_45737,N_45798);
or U47407 (N_47407,N_44719,N_45753);
or U47408 (N_47408,N_44819,N_44440);
nand U47409 (N_47409,N_45198,N_45541);
nand U47410 (N_47410,N_44694,N_45908);
and U47411 (N_47411,N_45119,N_45368);
nand U47412 (N_47412,N_44237,N_45432);
nor U47413 (N_47413,N_45468,N_45224);
and U47414 (N_47414,N_44293,N_44780);
nor U47415 (N_47415,N_44842,N_45708);
or U47416 (N_47416,N_45648,N_44699);
and U47417 (N_47417,N_44237,N_44447);
or U47418 (N_47418,N_44799,N_45331);
nand U47419 (N_47419,N_44658,N_44832);
nand U47420 (N_47420,N_45528,N_45462);
and U47421 (N_47421,N_45469,N_45479);
and U47422 (N_47422,N_45387,N_44214);
nor U47423 (N_47423,N_44089,N_44823);
and U47424 (N_47424,N_44212,N_44853);
or U47425 (N_47425,N_45730,N_44823);
and U47426 (N_47426,N_45054,N_45903);
or U47427 (N_47427,N_45922,N_44115);
nand U47428 (N_47428,N_44914,N_44067);
nand U47429 (N_47429,N_45425,N_44429);
and U47430 (N_47430,N_45715,N_44211);
nor U47431 (N_47431,N_44165,N_44833);
and U47432 (N_47432,N_45072,N_44593);
or U47433 (N_47433,N_45518,N_45560);
and U47434 (N_47434,N_44803,N_45874);
nand U47435 (N_47435,N_45592,N_45838);
nor U47436 (N_47436,N_44668,N_45441);
and U47437 (N_47437,N_45500,N_45438);
nand U47438 (N_47438,N_44332,N_45314);
nand U47439 (N_47439,N_45219,N_45234);
or U47440 (N_47440,N_44284,N_45703);
or U47441 (N_47441,N_44003,N_44533);
nand U47442 (N_47442,N_45992,N_45970);
or U47443 (N_47443,N_44816,N_45316);
nor U47444 (N_47444,N_45351,N_44805);
and U47445 (N_47445,N_44349,N_45092);
nor U47446 (N_47446,N_45848,N_44137);
xnor U47447 (N_47447,N_44568,N_45158);
nand U47448 (N_47448,N_45757,N_45987);
or U47449 (N_47449,N_45593,N_45741);
nand U47450 (N_47450,N_44690,N_44962);
nand U47451 (N_47451,N_44795,N_44129);
nor U47452 (N_47452,N_45537,N_45706);
nand U47453 (N_47453,N_44843,N_45902);
nor U47454 (N_47454,N_44943,N_44237);
xor U47455 (N_47455,N_45152,N_44916);
and U47456 (N_47456,N_45809,N_45706);
nor U47457 (N_47457,N_44290,N_45775);
or U47458 (N_47458,N_45107,N_44436);
nor U47459 (N_47459,N_45161,N_45747);
or U47460 (N_47460,N_45787,N_45923);
and U47461 (N_47461,N_45218,N_44058);
nand U47462 (N_47462,N_45240,N_44294);
or U47463 (N_47463,N_44623,N_44970);
nand U47464 (N_47464,N_44006,N_45985);
and U47465 (N_47465,N_44542,N_44883);
nand U47466 (N_47466,N_44968,N_44662);
or U47467 (N_47467,N_44507,N_44403);
and U47468 (N_47468,N_44052,N_44785);
nand U47469 (N_47469,N_45023,N_45089);
and U47470 (N_47470,N_45518,N_45452);
and U47471 (N_47471,N_44550,N_44512);
nor U47472 (N_47472,N_44487,N_45346);
or U47473 (N_47473,N_44662,N_45221);
or U47474 (N_47474,N_45375,N_44963);
and U47475 (N_47475,N_45031,N_44334);
nor U47476 (N_47476,N_44780,N_44115);
or U47477 (N_47477,N_44624,N_44535);
nand U47478 (N_47478,N_45857,N_44535);
xor U47479 (N_47479,N_44480,N_45106);
or U47480 (N_47480,N_44167,N_45137);
and U47481 (N_47481,N_45329,N_45648);
nand U47482 (N_47482,N_44735,N_44355);
and U47483 (N_47483,N_45206,N_45920);
nor U47484 (N_47484,N_44547,N_44852);
nand U47485 (N_47485,N_45499,N_44834);
nand U47486 (N_47486,N_44231,N_45478);
nand U47487 (N_47487,N_44599,N_44066);
and U47488 (N_47488,N_44331,N_44701);
and U47489 (N_47489,N_45733,N_44841);
nand U47490 (N_47490,N_44638,N_44684);
and U47491 (N_47491,N_44733,N_44430);
nand U47492 (N_47492,N_44158,N_45612);
or U47493 (N_47493,N_44619,N_44078);
nand U47494 (N_47494,N_44043,N_44972);
nor U47495 (N_47495,N_44042,N_44510);
or U47496 (N_47496,N_44113,N_45747);
and U47497 (N_47497,N_44793,N_44279);
or U47498 (N_47498,N_44424,N_45550);
nor U47499 (N_47499,N_45306,N_45836);
nand U47500 (N_47500,N_44117,N_45788);
nand U47501 (N_47501,N_45815,N_44586);
nand U47502 (N_47502,N_45652,N_44931);
nand U47503 (N_47503,N_44248,N_44681);
nor U47504 (N_47504,N_44616,N_44920);
and U47505 (N_47505,N_44874,N_44745);
or U47506 (N_47506,N_45568,N_44943);
nand U47507 (N_47507,N_44161,N_45040);
nor U47508 (N_47508,N_45791,N_45382);
or U47509 (N_47509,N_44935,N_44899);
nand U47510 (N_47510,N_45440,N_44422);
nand U47511 (N_47511,N_45630,N_45774);
and U47512 (N_47512,N_44251,N_44332);
or U47513 (N_47513,N_44459,N_45114);
and U47514 (N_47514,N_45789,N_45487);
nor U47515 (N_47515,N_45782,N_44990);
and U47516 (N_47516,N_44652,N_44375);
and U47517 (N_47517,N_44782,N_45840);
nand U47518 (N_47518,N_45092,N_45697);
or U47519 (N_47519,N_45479,N_45539);
and U47520 (N_47520,N_45803,N_45162);
nand U47521 (N_47521,N_44249,N_44866);
nor U47522 (N_47522,N_44101,N_45858);
and U47523 (N_47523,N_44540,N_44621);
or U47524 (N_47524,N_45171,N_44649);
nor U47525 (N_47525,N_44364,N_44820);
or U47526 (N_47526,N_44715,N_44337);
or U47527 (N_47527,N_45783,N_44320);
nand U47528 (N_47528,N_45463,N_45236);
and U47529 (N_47529,N_45660,N_45940);
and U47530 (N_47530,N_44876,N_44361);
nor U47531 (N_47531,N_44701,N_45270);
and U47532 (N_47532,N_44142,N_44245);
and U47533 (N_47533,N_45043,N_44150);
or U47534 (N_47534,N_45386,N_44184);
nor U47535 (N_47535,N_45818,N_44463);
and U47536 (N_47536,N_44159,N_44770);
nand U47537 (N_47537,N_44798,N_45118);
or U47538 (N_47538,N_45527,N_45864);
nor U47539 (N_47539,N_45622,N_44588);
nand U47540 (N_47540,N_45556,N_44851);
nor U47541 (N_47541,N_45788,N_45384);
nand U47542 (N_47542,N_45870,N_44263);
nor U47543 (N_47543,N_45826,N_45763);
or U47544 (N_47544,N_44441,N_44520);
nand U47545 (N_47545,N_44579,N_44081);
or U47546 (N_47546,N_44915,N_44886);
or U47547 (N_47547,N_44511,N_45814);
or U47548 (N_47548,N_45849,N_44718);
nor U47549 (N_47549,N_45331,N_45379);
or U47550 (N_47550,N_45469,N_45950);
and U47551 (N_47551,N_44399,N_45998);
or U47552 (N_47552,N_44283,N_44622);
nand U47553 (N_47553,N_45932,N_44998);
nand U47554 (N_47554,N_44872,N_44104);
or U47555 (N_47555,N_44179,N_44418);
and U47556 (N_47556,N_45472,N_44895);
and U47557 (N_47557,N_44377,N_45251);
or U47558 (N_47558,N_44945,N_45385);
and U47559 (N_47559,N_45520,N_44346);
and U47560 (N_47560,N_44412,N_45860);
or U47561 (N_47561,N_45352,N_44576);
and U47562 (N_47562,N_44525,N_45473);
and U47563 (N_47563,N_45522,N_45853);
nand U47564 (N_47564,N_44580,N_45221);
nor U47565 (N_47565,N_44404,N_44409);
or U47566 (N_47566,N_44100,N_45247);
nor U47567 (N_47567,N_45451,N_45629);
nor U47568 (N_47568,N_45167,N_44222);
nand U47569 (N_47569,N_45251,N_45045);
nand U47570 (N_47570,N_45133,N_44284);
and U47571 (N_47571,N_44182,N_45422);
and U47572 (N_47572,N_45291,N_44590);
nor U47573 (N_47573,N_45824,N_45272);
and U47574 (N_47574,N_44622,N_44426);
nor U47575 (N_47575,N_44556,N_44210);
and U47576 (N_47576,N_44873,N_44868);
or U47577 (N_47577,N_45736,N_45430);
nor U47578 (N_47578,N_44337,N_44917);
nand U47579 (N_47579,N_44097,N_45237);
or U47580 (N_47580,N_44798,N_44511);
nand U47581 (N_47581,N_45975,N_44304);
nand U47582 (N_47582,N_44217,N_45723);
nor U47583 (N_47583,N_45720,N_44442);
and U47584 (N_47584,N_44026,N_44342);
nand U47585 (N_47585,N_45084,N_45814);
and U47586 (N_47586,N_44313,N_45275);
nor U47587 (N_47587,N_45360,N_44575);
or U47588 (N_47588,N_45917,N_44870);
nand U47589 (N_47589,N_44735,N_44589);
or U47590 (N_47590,N_45115,N_44635);
and U47591 (N_47591,N_44911,N_44169);
and U47592 (N_47592,N_44851,N_45865);
nor U47593 (N_47593,N_44709,N_44668);
xnor U47594 (N_47594,N_45917,N_44141);
nand U47595 (N_47595,N_44089,N_45395);
or U47596 (N_47596,N_44630,N_44370);
nand U47597 (N_47597,N_45091,N_45349);
or U47598 (N_47598,N_45535,N_44963);
nor U47599 (N_47599,N_44648,N_44222);
nand U47600 (N_47600,N_45734,N_44353);
and U47601 (N_47601,N_44954,N_45969);
or U47602 (N_47602,N_45545,N_44881);
nand U47603 (N_47603,N_45768,N_45432);
nand U47604 (N_47604,N_45613,N_45624);
nand U47605 (N_47605,N_44931,N_45044);
nor U47606 (N_47606,N_44393,N_45119);
nor U47607 (N_47607,N_45918,N_45861);
or U47608 (N_47608,N_45885,N_45262);
or U47609 (N_47609,N_44841,N_44671);
and U47610 (N_47610,N_45910,N_44834);
nor U47611 (N_47611,N_44028,N_44205);
nand U47612 (N_47612,N_45872,N_45464);
or U47613 (N_47613,N_44381,N_44355);
nor U47614 (N_47614,N_45945,N_44694);
nand U47615 (N_47615,N_45320,N_44865);
or U47616 (N_47616,N_44400,N_44052);
nand U47617 (N_47617,N_44518,N_44767);
and U47618 (N_47618,N_45679,N_44126);
nor U47619 (N_47619,N_45876,N_44090);
and U47620 (N_47620,N_44225,N_45520);
or U47621 (N_47621,N_45031,N_45141);
or U47622 (N_47622,N_45481,N_45492);
and U47623 (N_47623,N_45804,N_45484);
nor U47624 (N_47624,N_45769,N_45207);
and U47625 (N_47625,N_45752,N_45519);
nor U47626 (N_47626,N_44965,N_44445);
and U47627 (N_47627,N_44175,N_45416);
nor U47628 (N_47628,N_44006,N_44357);
and U47629 (N_47629,N_44917,N_45835);
nand U47630 (N_47630,N_44551,N_44211);
nand U47631 (N_47631,N_44836,N_44535);
nand U47632 (N_47632,N_44649,N_45531);
or U47633 (N_47633,N_44972,N_44545);
nand U47634 (N_47634,N_44890,N_44328);
nor U47635 (N_47635,N_44547,N_45099);
or U47636 (N_47636,N_45564,N_45184);
or U47637 (N_47637,N_44693,N_45234);
nor U47638 (N_47638,N_45729,N_44570);
or U47639 (N_47639,N_45078,N_45497);
or U47640 (N_47640,N_44710,N_45152);
nand U47641 (N_47641,N_44717,N_45418);
nand U47642 (N_47642,N_44460,N_44497);
and U47643 (N_47643,N_44212,N_44060);
and U47644 (N_47644,N_44295,N_44546);
and U47645 (N_47645,N_45562,N_44093);
and U47646 (N_47646,N_44101,N_45704);
or U47647 (N_47647,N_44951,N_44764);
or U47648 (N_47648,N_44932,N_45797);
nand U47649 (N_47649,N_44688,N_44852);
nand U47650 (N_47650,N_45291,N_44446);
xor U47651 (N_47651,N_45873,N_44138);
nor U47652 (N_47652,N_44088,N_45080);
and U47653 (N_47653,N_45362,N_44512);
and U47654 (N_47654,N_45359,N_44190);
nand U47655 (N_47655,N_44181,N_44784);
nor U47656 (N_47656,N_44815,N_45851);
nor U47657 (N_47657,N_44733,N_44532);
or U47658 (N_47658,N_44041,N_45367);
nor U47659 (N_47659,N_44587,N_45192);
and U47660 (N_47660,N_44272,N_45058);
nor U47661 (N_47661,N_44892,N_44492);
nand U47662 (N_47662,N_44939,N_45729);
and U47663 (N_47663,N_45966,N_45800);
or U47664 (N_47664,N_44532,N_44058);
nand U47665 (N_47665,N_44876,N_44823);
or U47666 (N_47666,N_44457,N_44553);
nand U47667 (N_47667,N_45858,N_44387);
nand U47668 (N_47668,N_45738,N_45958);
or U47669 (N_47669,N_44814,N_44844);
and U47670 (N_47670,N_45356,N_44729);
nor U47671 (N_47671,N_45926,N_44767);
and U47672 (N_47672,N_45100,N_44388);
or U47673 (N_47673,N_44562,N_45620);
nand U47674 (N_47674,N_44028,N_45225);
or U47675 (N_47675,N_45034,N_44978);
and U47676 (N_47676,N_44776,N_44937);
or U47677 (N_47677,N_44112,N_44794);
or U47678 (N_47678,N_44551,N_44746);
or U47679 (N_47679,N_45436,N_45601);
xnor U47680 (N_47680,N_45822,N_45978);
nand U47681 (N_47681,N_45947,N_44901);
and U47682 (N_47682,N_45654,N_44745);
or U47683 (N_47683,N_44808,N_45339);
nor U47684 (N_47684,N_45690,N_45773);
and U47685 (N_47685,N_44009,N_44128);
xor U47686 (N_47686,N_44694,N_45268);
and U47687 (N_47687,N_44378,N_45138);
nor U47688 (N_47688,N_44144,N_44852);
nand U47689 (N_47689,N_45303,N_44072);
nand U47690 (N_47690,N_44547,N_45337);
nor U47691 (N_47691,N_45607,N_44781);
nand U47692 (N_47692,N_44129,N_44914);
or U47693 (N_47693,N_45567,N_45018);
or U47694 (N_47694,N_45710,N_44507);
nand U47695 (N_47695,N_45272,N_45363);
nand U47696 (N_47696,N_44306,N_44976);
nand U47697 (N_47697,N_44140,N_44172);
nor U47698 (N_47698,N_44767,N_45755);
or U47699 (N_47699,N_44476,N_44038);
or U47700 (N_47700,N_44671,N_45922);
or U47701 (N_47701,N_45179,N_44354);
nand U47702 (N_47702,N_44394,N_44976);
and U47703 (N_47703,N_45695,N_45965);
nor U47704 (N_47704,N_44606,N_45123);
nor U47705 (N_47705,N_44205,N_45338);
xor U47706 (N_47706,N_45208,N_44711);
nand U47707 (N_47707,N_44600,N_45481);
nand U47708 (N_47708,N_44358,N_44696);
and U47709 (N_47709,N_44803,N_44365);
and U47710 (N_47710,N_45579,N_45986);
and U47711 (N_47711,N_44560,N_45766);
and U47712 (N_47712,N_45658,N_45332);
nand U47713 (N_47713,N_44645,N_45525);
or U47714 (N_47714,N_44443,N_45546);
or U47715 (N_47715,N_44273,N_44512);
nand U47716 (N_47716,N_44875,N_45068);
nor U47717 (N_47717,N_45407,N_44196);
and U47718 (N_47718,N_45750,N_45814);
nand U47719 (N_47719,N_45091,N_44361);
nand U47720 (N_47720,N_44423,N_45873);
and U47721 (N_47721,N_44422,N_44292);
nand U47722 (N_47722,N_45274,N_45428);
nand U47723 (N_47723,N_45678,N_44121);
nand U47724 (N_47724,N_45026,N_45253);
nor U47725 (N_47725,N_45560,N_44117);
and U47726 (N_47726,N_44220,N_44951);
nor U47727 (N_47727,N_45798,N_45446);
or U47728 (N_47728,N_44355,N_44202);
nor U47729 (N_47729,N_44304,N_45516);
or U47730 (N_47730,N_44411,N_45464);
and U47731 (N_47731,N_45117,N_44126);
nand U47732 (N_47732,N_45842,N_45645);
nand U47733 (N_47733,N_45208,N_45300);
or U47734 (N_47734,N_45722,N_44386);
and U47735 (N_47735,N_45310,N_45188);
xor U47736 (N_47736,N_45005,N_45950);
nand U47737 (N_47737,N_44825,N_45401);
and U47738 (N_47738,N_45512,N_44238);
nand U47739 (N_47739,N_45668,N_44694);
nand U47740 (N_47740,N_44570,N_44253);
or U47741 (N_47741,N_45103,N_44106);
nor U47742 (N_47742,N_44544,N_44843);
and U47743 (N_47743,N_45771,N_45373);
nand U47744 (N_47744,N_44467,N_45236);
nand U47745 (N_47745,N_44593,N_45179);
or U47746 (N_47746,N_45429,N_44576);
nor U47747 (N_47747,N_45976,N_45253);
or U47748 (N_47748,N_45665,N_45441);
xnor U47749 (N_47749,N_45460,N_44853);
nor U47750 (N_47750,N_45291,N_44128);
nor U47751 (N_47751,N_44474,N_44548);
nand U47752 (N_47752,N_45155,N_44455);
and U47753 (N_47753,N_45941,N_44005);
or U47754 (N_47754,N_45205,N_45290);
nand U47755 (N_47755,N_45309,N_44943);
and U47756 (N_47756,N_45881,N_44584);
and U47757 (N_47757,N_44394,N_45064);
or U47758 (N_47758,N_45131,N_44487);
and U47759 (N_47759,N_44012,N_44667);
nor U47760 (N_47760,N_44422,N_45706);
nand U47761 (N_47761,N_45439,N_45147);
or U47762 (N_47762,N_44327,N_44056);
and U47763 (N_47763,N_44450,N_45198);
nor U47764 (N_47764,N_44695,N_44953);
nor U47765 (N_47765,N_44637,N_44511);
or U47766 (N_47766,N_44508,N_44871);
nand U47767 (N_47767,N_45459,N_44442);
nor U47768 (N_47768,N_45754,N_44741);
nand U47769 (N_47769,N_45615,N_44961);
xor U47770 (N_47770,N_45185,N_44174);
or U47771 (N_47771,N_44984,N_45148);
or U47772 (N_47772,N_45798,N_44821);
or U47773 (N_47773,N_44233,N_44843);
xor U47774 (N_47774,N_45087,N_44027);
nor U47775 (N_47775,N_44191,N_44707);
and U47776 (N_47776,N_44482,N_44929);
or U47777 (N_47777,N_45502,N_45374);
or U47778 (N_47778,N_45156,N_44853);
or U47779 (N_47779,N_45557,N_45436);
and U47780 (N_47780,N_45428,N_45465);
nand U47781 (N_47781,N_44016,N_45001);
nor U47782 (N_47782,N_45565,N_44690);
nand U47783 (N_47783,N_44514,N_45849);
nand U47784 (N_47784,N_44513,N_44540);
nor U47785 (N_47785,N_45008,N_45207);
and U47786 (N_47786,N_44352,N_44807);
nor U47787 (N_47787,N_44188,N_44381);
and U47788 (N_47788,N_44186,N_44103);
or U47789 (N_47789,N_45557,N_45994);
and U47790 (N_47790,N_45840,N_45251);
and U47791 (N_47791,N_44726,N_45327);
nor U47792 (N_47792,N_45600,N_44289);
nand U47793 (N_47793,N_44342,N_45894);
and U47794 (N_47794,N_45354,N_44581);
and U47795 (N_47795,N_45961,N_44227);
or U47796 (N_47796,N_44555,N_44585);
nand U47797 (N_47797,N_45410,N_44124);
or U47798 (N_47798,N_45933,N_45265);
or U47799 (N_47799,N_44231,N_45850);
nand U47800 (N_47800,N_44025,N_45907);
nor U47801 (N_47801,N_45750,N_44983);
or U47802 (N_47802,N_44528,N_45802);
xnor U47803 (N_47803,N_45896,N_44377);
nand U47804 (N_47804,N_44022,N_44304);
and U47805 (N_47805,N_45200,N_44818);
and U47806 (N_47806,N_45616,N_44541);
nand U47807 (N_47807,N_45700,N_44854);
or U47808 (N_47808,N_44363,N_45305);
or U47809 (N_47809,N_45195,N_45264);
nand U47810 (N_47810,N_44168,N_44968);
or U47811 (N_47811,N_45620,N_45096);
and U47812 (N_47812,N_44591,N_45824);
or U47813 (N_47813,N_45596,N_44994);
nor U47814 (N_47814,N_45333,N_45134);
xor U47815 (N_47815,N_45226,N_45770);
nor U47816 (N_47816,N_44011,N_45893);
nand U47817 (N_47817,N_44508,N_45712);
nand U47818 (N_47818,N_45718,N_44541);
or U47819 (N_47819,N_45574,N_45932);
or U47820 (N_47820,N_44403,N_45066);
or U47821 (N_47821,N_45325,N_44225);
nand U47822 (N_47822,N_44684,N_45316);
or U47823 (N_47823,N_45522,N_44029);
or U47824 (N_47824,N_45699,N_45872);
or U47825 (N_47825,N_45748,N_44065);
or U47826 (N_47826,N_44942,N_44981);
nand U47827 (N_47827,N_45836,N_45078);
nor U47828 (N_47828,N_44595,N_45504);
or U47829 (N_47829,N_44809,N_44906);
nand U47830 (N_47830,N_45931,N_45064);
and U47831 (N_47831,N_45796,N_44275);
nor U47832 (N_47832,N_45195,N_44157);
nand U47833 (N_47833,N_44268,N_44114);
and U47834 (N_47834,N_44344,N_44194);
or U47835 (N_47835,N_45418,N_45694);
nor U47836 (N_47836,N_44702,N_44898);
nor U47837 (N_47837,N_45832,N_45484);
nand U47838 (N_47838,N_45037,N_44989);
and U47839 (N_47839,N_44036,N_44253);
nand U47840 (N_47840,N_44092,N_44621);
and U47841 (N_47841,N_44892,N_44568);
and U47842 (N_47842,N_44484,N_44275);
nand U47843 (N_47843,N_45684,N_45148);
and U47844 (N_47844,N_44973,N_45456);
nor U47845 (N_47845,N_44550,N_44408);
or U47846 (N_47846,N_45077,N_45695);
and U47847 (N_47847,N_44916,N_45870);
and U47848 (N_47848,N_44860,N_44622);
nor U47849 (N_47849,N_44151,N_44231);
nand U47850 (N_47850,N_44187,N_45554);
and U47851 (N_47851,N_44110,N_45665);
or U47852 (N_47852,N_45113,N_44397);
and U47853 (N_47853,N_45584,N_44989);
or U47854 (N_47854,N_45017,N_44616);
and U47855 (N_47855,N_45732,N_45627);
nor U47856 (N_47856,N_44073,N_44199);
or U47857 (N_47857,N_45246,N_45948);
and U47858 (N_47858,N_44855,N_44244);
nor U47859 (N_47859,N_44913,N_44132);
or U47860 (N_47860,N_44366,N_44565);
and U47861 (N_47861,N_45405,N_45000);
and U47862 (N_47862,N_45935,N_45385);
nor U47863 (N_47863,N_44427,N_44641);
nand U47864 (N_47864,N_44930,N_45105);
nor U47865 (N_47865,N_45744,N_44577);
nor U47866 (N_47866,N_45414,N_45110);
and U47867 (N_47867,N_45701,N_44942);
xor U47868 (N_47868,N_45674,N_45911);
or U47869 (N_47869,N_45425,N_45157);
or U47870 (N_47870,N_45171,N_45462);
nand U47871 (N_47871,N_45304,N_45808);
or U47872 (N_47872,N_44692,N_44829);
nand U47873 (N_47873,N_44914,N_45904);
and U47874 (N_47874,N_45438,N_45592);
or U47875 (N_47875,N_45156,N_45907);
nor U47876 (N_47876,N_44361,N_45800);
nand U47877 (N_47877,N_45591,N_44088);
and U47878 (N_47878,N_45211,N_44362);
nor U47879 (N_47879,N_44474,N_45623);
or U47880 (N_47880,N_44465,N_45157);
nand U47881 (N_47881,N_45916,N_45398);
and U47882 (N_47882,N_44422,N_45274);
nand U47883 (N_47883,N_45728,N_44742);
nand U47884 (N_47884,N_44548,N_45954);
nor U47885 (N_47885,N_45512,N_44074);
nand U47886 (N_47886,N_44122,N_45051);
nor U47887 (N_47887,N_44491,N_44031);
or U47888 (N_47888,N_44925,N_45691);
nand U47889 (N_47889,N_44946,N_44822);
nand U47890 (N_47890,N_45292,N_44585);
or U47891 (N_47891,N_45246,N_45266);
nand U47892 (N_47892,N_45373,N_45733);
or U47893 (N_47893,N_44269,N_45867);
and U47894 (N_47894,N_45647,N_44761);
nand U47895 (N_47895,N_44599,N_44482);
xnor U47896 (N_47896,N_45515,N_44987);
or U47897 (N_47897,N_44003,N_45177);
or U47898 (N_47898,N_44481,N_44182);
nand U47899 (N_47899,N_44099,N_44289);
nand U47900 (N_47900,N_44749,N_45992);
nand U47901 (N_47901,N_44626,N_44749);
and U47902 (N_47902,N_44171,N_44323);
nand U47903 (N_47903,N_44807,N_45129);
or U47904 (N_47904,N_44011,N_45114);
and U47905 (N_47905,N_44695,N_44178);
nand U47906 (N_47906,N_45864,N_44605);
nor U47907 (N_47907,N_44725,N_45395);
nand U47908 (N_47908,N_44987,N_44586);
or U47909 (N_47909,N_44953,N_45086);
and U47910 (N_47910,N_44484,N_45703);
nor U47911 (N_47911,N_45173,N_45358);
or U47912 (N_47912,N_44747,N_45538);
and U47913 (N_47913,N_45560,N_45545);
or U47914 (N_47914,N_45333,N_44145);
nand U47915 (N_47915,N_45534,N_45185);
and U47916 (N_47916,N_44333,N_44747);
xnor U47917 (N_47917,N_45296,N_44385);
nand U47918 (N_47918,N_44744,N_45053);
or U47919 (N_47919,N_45203,N_45220);
nand U47920 (N_47920,N_44010,N_44672);
nand U47921 (N_47921,N_44768,N_45937);
nand U47922 (N_47922,N_44851,N_44151);
xor U47923 (N_47923,N_44128,N_44025);
and U47924 (N_47924,N_44731,N_44033);
nand U47925 (N_47925,N_44656,N_44717);
or U47926 (N_47926,N_44961,N_45241);
nor U47927 (N_47927,N_45557,N_45307);
nor U47928 (N_47928,N_45795,N_44406);
nand U47929 (N_47929,N_44110,N_44540);
and U47930 (N_47930,N_44478,N_45182);
nand U47931 (N_47931,N_44722,N_44373);
and U47932 (N_47932,N_45206,N_45675);
nor U47933 (N_47933,N_45825,N_44177);
or U47934 (N_47934,N_45906,N_45555);
or U47935 (N_47935,N_44046,N_45739);
nor U47936 (N_47936,N_44349,N_45626);
and U47937 (N_47937,N_44259,N_45973);
or U47938 (N_47938,N_44392,N_44258);
nand U47939 (N_47939,N_45044,N_45160);
and U47940 (N_47940,N_44287,N_45818);
nor U47941 (N_47941,N_44931,N_45646);
and U47942 (N_47942,N_45915,N_44498);
nor U47943 (N_47943,N_45744,N_45824);
and U47944 (N_47944,N_44945,N_45427);
or U47945 (N_47945,N_44345,N_45491);
and U47946 (N_47946,N_44056,N_44064);
nand U47947 (N_47947,N_45200,N_45672);
nor U47948 (N_47948,N_45637,N_44930);
or U47949 (N_47949,N_44744,N_45704);
or U47950 (N_47950,N_45668,N_45994);
nor U47951 (N_47951,N_44739,N_45683);
nor U47952 (N_47952,N_44195,N_45117);
and U47953 (N_47953,N_45054,N_45039);
or U47954 (N_47954,N_44202,N_44338);
and U47955 (N_47955,N_45406,N_45479);
and U47956 (N_47956,N_45422,N_44658);
nor U47957 (N_47957,N_44932,N_44822);
or U47958 (N_47958,N_45239,N_44578);
and U47959 (N_47959,N_45585,N_45750);
nand U47960 (N_47960,N_45188,N_44125);
xnor U47961 (N_47961,N_45618,N_44361);
or U47962 (N_47962,N_45087,N_44634);
xor U47963 (N_47963,N_44450,N_44488);
and U47964 (N_47964,N_44005,N_45052);
nor U47965 (N_47965,N_45013,N_45011);
nand U47966 (N_47966,N_44248,N_45591);
nor U47967 (N_47967,N_45154,N_44996);
and U47968 (N_47968,N_44767,N_44744);
xnor U47969 (N_47969,N_45137,N_45131);
or U47970 (N_47970,N_45762,N_44866);
nand U47971 (N_47971,N_45820,N_45631);
and U47972 (N_47972,N_45506,N_45039);
nand U47973 (N_47973,N_45788,N_44216);
and U47974 (N_47974,N_44966,N_45483);
and U47975 (N_47975,N_44682,N_45316);
or U47976 (N_47976,N_44960,N_44765);
nand U47977 (N_47977,N_44200,N_44700);
nor U47978 (N_47978,N_44671,N_44995);
or U47979 (N_47979,N_44802,N_45566);
nand U47980 (N_47980,N_45740,N_45553);
and U47981 (N_47981,N_45951,N_44794);
and U47982 (N_47982,N_44419,N_44015);
or U47983 (N_47983,N_44053,N_44835);
and U47984 (N_47984,N_44407,N_45945);
and U47985 (N_47985,N_45347,N_44561);
and U47986 (N_47986,N_44110,N_44481);
xnor U47987 (N_47987,N_45382,N_44487);
nand U47988 (N_47988,N_44606,N_44148);
or U47989 (N_47989,N_45316,N_44358);
xor U47990 (N_47990,N_45779,N_44663);
nor U47991 (N_47991,N_44239,N_44203);
nor U47992 (N_47992,N_44156,N_45281);
nand U47993 (N_47993,N_45292,N_45839);
nor U47994 (N_47994,N_45077,N_45578);
nand U47995 (N_47995,N_45478,N_44393);
nand U47996 (N_47996,N_44149,N_44021);
and U47997 (N_47997,N_45615,N_45749);
and U47998 (N_47998,N_44806,N_44354);
nor U47999 (N_47999,N_44060,N_44458);
nor U48000 (N_48000,N_46902,N_46328);
and U48001 (N_48001,N_47762,N_47476);
or U48002 (N_48002,N_47807,N_47205);
nor U48003 (N_48003,N_47688,N_46154);
nor U48004 (N_48004,N_47801,N_47847);
or U48005 (N_48005,N_47073,N_47568);
and U48006 (N_48006,N_47882,N_46913);
nor U48007 (N_48007,N_47005,N_46065);
nor U48008 (N_48008,N_47958,N_47109);
and U48009 (N_48009,N_46653,N_47028);
nand U48010 (N_48010,N_47698,N_47630);
xnor U48011 (N_48011,N_47475,N_46311);
or U48012 (N_48012,N_46051,N_46658);
and U48013 (N_48013,N_46216,N_47692);
nand U48014 (N_48014,N_47327,N_46246);
and U48015 (N_48015,N_46650,N_46222);
nand U48016 (N_48016,N_46025,N_46043);
or U48017 (N_48017,N_46735,N_47591);
nor U48018 (N_48018,N_46001,N_47237);
nor U48019 (N_48019,N_46260,N_47751);
nand U48020 (N_48020,N_46022,N_46402);
nand U48021 (N_48021,N_47395,N_46869);
nor U48022 (N_48022,N_47238,N_47673);
nor U48023 (N_48023,N_47022,N_47548);
nand U48024 (N_48024,N_47935,N_46122);
or U48025 (N_48025,N_47521,N_47045);
or U48026 (N_48026,N_46310,N_46605);
and U48027 (N_48027,N_47485,N_47153);
or U48028 (N_48028,N_47438,N_47160);
xor U48029 (N_48029,N_46860,N_47681);
nor U48030 (N_48030,N_46232,N_47718);
nor U48031 (N_48031,N_46331,N_46689);
nor U48032 (N_48032,N_47985,N_46964);
nand U48033 (N_48033,N_46489,N_47457);
nand U48034 (N_48034,N_46821,N_46018);
nand U48035 (N_48035,N_46743,N_47785);
nand U48036 (N_48036,N_47744,N_47366);
and U48037 (N_48037,N_47081,N_46600);
nand U48038 (N_48038,N_47381,N_47023);
and U48039 (N_48039,N_47804,N_47497);
nand U48040 (N_48040,N_46110,N_46569);
nor U48041 (N_48041,N_46713,N_47855);
nor U48042 (N_48042,N_46295,N_47709);
and U48043 (N_48043,N_47931,N_47062);
or U48044 (N_48044,N_46158,N_46731);
and U48045 (N_48045,N_46140,N_46736);
or U48046 (N_48046,N_46875,N_47333);
nor U48047 (N_48047,N_47654,N_47553);
nand U48048 (N_48048,N_47006,N_47064);
or U48049 (N_48049,N_47021,N_47639);
and U48050 (N_48050,N_47295,N_47836);
nand U48051 (N_48051,N_46505,N_47072);
nor U48052 (N_48052,N_47307,N_46917);
or U48053 (N_48053,N_46789,N_47802);
or U48054 (N_48054,N_47504,N_47375);
or U48055 (N_48055,N_46725,N_46879);
or U48056 (N_48056,N_47010,N_46360);
nand U48057 (N_48057,N_46189,N_47458);
and U48058 (N_48058,N_47133,N_47125);
and U48059 (N_48059,N_46738,N_47279);
nor U48060 (N_48060,N_47254,N_47661);
nand U48061 (N_48061,N_47247,N_46292);
nand U48062 (N_48062,N_46485,N_46803);
nor U48063 (N_48063,N_47649,N_46013);
nand U48064 (N_48064,N_46159,N_47215);
and U48065 (N_48065,N_47530,N_46830);
nor U48066 (N_48066,N_46698,N_47165);
and U48067 (N_48067,N_47077,N_47092);
nand U48068 (N_48068,N_46834,N_46703);
nand U48069 (N_48069,N_46574,N_46589);
nand U48070 (N_48070,N_47490,N_46268);
or U48071 (N_48071,N_47594,N_47309);
and U48072 (N_48072,N_46291,N_46612);
nand U48073 (N_48073,N_46135,N_47896);
nor U48074 (N_48074,N_47047,N_47027);
or U48075 (N_48075,N_47441,N_47505);
nand U48076 (N_48076,N_46802,N_46628);
or U48077 (N_48077,N_46123,N_46363);
and U48078 (N_48078,N_47872,N_46290);
and U48079 (N_48079,N_46339,N_47905);
nor U48080 (N_48080,N_47976,N_46987);
or U48081 (N_48081,N_47465,N_47204);
and U48082 (N_48082,N_46053,N_47748);
and U48083 (N_48083,N_46206,N_46027);
or U48084 (N_48084,N_46835,N_46308);
or U48085 (N_48085,N_46488,N_46412);
nand U48086 (N_48086,N_46444,N_47735);
nand U48087 (N_48087,N_46817,N_46033);
nor U48088 (N_48088,N_46225,N_46724);
nor U48089 (N_48089,N_47991,N_46376);
nor U48090 (N_48090,N_47199,N_46465);
nand U48091 (N_48091,N_47920,N_47910);
nand U48092 (N_48092,N_47763,N_46639);
or U48093 (N_48093,N_47912,N_46867);
nor U48094 (N_48094,N_46252,N_47518);
nor U48095 (N_48095,N_46336,N_46066);
or U48096 (N_48096,N_47294,N_47603);
nor U48097 (N_48097,N_46071,N_47184);
nor U48098 (N_48098,N_47755,N_46192);
or U48099 (N_48099,N_46769,N_46666);
nor U48100 (N_48100,N_46818,N_47058);
nor U48101 (N_48101,N_46358,N_47429);
and U48102 (N_48102,N_47103,N_46634);
or U48103 (N_48103,N_47054,N_47357);
and U48104 (N_48104,N_47312,N_47601);
nor U48105 (N_48105,N_47837,N_46576);
nand U48106 (N_48106,N_47456,N_47406);
nand U48107 (N_48107,N_47454,N_47819);
nand U48108 (N_48108,N_46956,N_46498);
xnor U48109 (N_48109,N_46200,N_47641);
nor U48110 (N_48110,N_46971,N_46037);
nand U48111 (N_48111,N_47059,N_46688);
nand U48112 (N_48112,N_47445,N_47296);
and U48113 (N_48113,N_46909,N_46915);
nor U48114 (N_48114,N_47493,N_47282);
nor U48115 (N_48115,N_46923,N_46142);
xor U48116 (N_48116,N_46756,N_47759);
and U48117 (N_48117,N_46409,N_46259);
xor U48118 (N_48118,N_46824,N_47304);
nand U48119 (N_48119,N_47724,N_47245);
nor U48120 (N_48120,N_47579,N_46531);
or U48121 (N_48121,N_46809,N_47849);
and U48122 (N_48122,N_46642,N_47037);
and U48123 (N_48123,N_47672,N_47795);
and U48124 (N_48124,N_46244,N_46313);
and U48125 (N_48125,N_47960,N_47275);
or U48126 (N_48126,N_46541,N_47933);
nor U48127 (N_48127,N_46795,N_46712);
and U48128 (N_48128,N_46808,N_46329);
nand U48129 (N_48129,N_46030,N_47030);
nor U48130 (N_48130,N_46947,N_47330);
and U48131 (N_48131,N_46935,N_47217);
and U48132 (N_48132,N_47788,N_47886);
nand U48133 (N_48133,N_47089,N_47830);
or U48134 (N_48134,N_46606,N_46315);
nor U48135 (N_48135,N_46721,N_47586);
nand U48136 (N_48136,N_46381,N_47640);
nand U48137 (N_48137,N_46385,N_46750);
nand U48138 (N_48138,N_47564,N_47244);
nor U48139 (N_48139,N_46578,N_47897);
nand U48140 (N_48140,N_47015,N_47565);
nor U48141 (N_48141,N_46718,N_46579);
nand U48142 (N_48142,N_47981,N_47123);
or U48143 (N_48143,N_46182,N_46684);
and U48144 (N_48144,N_47183,N_46325);
xnor U48145 (N_48145,N_47007,N_46111);
nand U48146 (N_48146,N_46139,N_47039);
and U48147 (N_48147,N_46029,N_47214);
or U48148 (N_48148,N_46581,N_46038);
nand U48149 (N_48149,N_47340,N_47368);
nor U48150 (N_48150,N_47303,N_47838);
nand U48151 (N_48151,N_47699,N_46473);
nor U48152 (N_48152,N_46016,N_47335);
nor U48153 (N_48153,N_46660,N_46491);
nand U48154 (N_48154,N_46480,N_46865);
nor U48155 (N_48155,N_47447,N_46458);
and U48156 (N_48156,N_47192,N_46878);
or U48157 (N_48157,N_47900,N_47711);
or U48158 (N_48158,N_47746,N_46112);
nor U48159 (N_48159,N_47822,N_47116);
nor U48160 (N_48160,N_46633,N_47008);
nor U48161 (N_48161,N_47404,N_47501);
nand U48162 (N_48162,N_47210,N_47651);
and U48163 (N_48163,N_47632,N_47048);
or U48164 (N_48164,N_47474,N_46237);
nor U48165 (N_48165,N_47218,N_47970);
nor U48166 (N_48166,N_47211,N_47070);
nand U48167 (N_48167,N_46499,N_47251);
nand U48168 (N_48168,N_46883,N_47557);
nor U48169 (N_48169,N_46610,N_47894);
and U48170 (N_48170,N_46784,N_46350);
and U48171 (N_48171,N_46994,N_47220);
nor U48172 (N_48172,N_47388,N_46209);
and U48173 (N_48173,N_46431,N_47331);
or U48174 (N_48174,N_46050,N_47703);
and U48175 (N_48175,N_46486,N_47469);
or U48176 (N_48176,N_46299,N_46945);
nor U48177 (N_48177,N_47992,N_46717);
nand U48178 (N_48178,N_47575,N_47895);
nand U48179 (N_48179,N_46848,N_47043);
and U48180 (N_48180,N_47818,N_46266);
xor U48181 (N_48181,N_46919,N_46305);
nor U48182 (N_48182,N_47531,N_46287);
or U48183 (N_48183,N_46876,N_46249);
nor U48184 (N_48184,N_46966,N_47209);
or U48185 (N_48185,N_47656,N_47563);
or U48186 (N_48186,N_46101,N_46264);
nor U48187 (N_48187,N_46072,N_47877);
and U48188 (N_48188,N_46341,N_47980);
nand U48189 (N_48189,N_47362,N_46495);
nor U48190 (N_48190,N_46035,N_46972);
nand U48191 (N_48191,N_47500,N_47840);
nor U48192 (N_48192,N_46760,N_46423);
xnor U48193 (N_48193,N_47325,N_47108);
nor U48194 (N_48194,N_46852,N_47754);
and U48195 (N_48195,N_47843,N_46397);
or U48196 (N_48196,N_47203,N_46279);
and U48197 (N_48197,N_46286,N_46554);
and U48198 (N_48198,N_46088,N_47181);
nor U48199 (N_48199,N_47223,N_47236);
or U48200 (N_48200,N_46661,N_46114);
and U48201 (N_48201,N_47696,N_47433);
or U48202 (N_48202,N_46082,N_46034);
nor U48203 (N_48203,N_47577,N_46424);
and U48204 (N_48204,N_46276,N_47364);
nand U48205 (N_48205,N_47034,N_47927);
or U48206 (N_48206,N_46324,N_46833);
or U48207 (N_48207,N_46031,N_47947);
nor U48208 (N_48208,N_47923,N_46611);
or U48209 (N_48209,N_46400,N_47104);
nand U48210 (N_48210,N_47812,N_46483);
or U48211 (N_48211,N_46185,N_47256);
nor U48212 (N_48212,N_47879,N_46248);
and U48213 (N_48213,N_46457,N_46213);
or U48214 (N_48214,N_46882,N_46877);
or U48215 (N_48215,N_46952,N_46479);
nand U48216 (N_48216,N_46615,N_47988);
nor U48217 (N_48217,N_46847,N_46707);
xor U48218 (N_48218,N_46508,N_47370);
and U48219 (N_48219,N_47396,N_47851);
and U48220 (N_48220,N_47519,N_47913);
nor U48221 (N_48221,N_47908,N_46282);
or U48222 (N_48222,N_46391,N_46930);
nand U48223 (N_48223,N_47522,N_47378);
and U48224 (N_48224,N_47257,N_46356);
nor U48225 (N_48225,N_46680,N_46675);
nor U48226 (N_48226,N_47679,N_47202);
or U48227 (N_48227,N_46357,N_46487);
and U48228 (N_48228,N_46543,N_46410);
or U48229 (N_48229,N_46638,N_47997);
or U48230 (N_48230,N_47989,N_46077);
nor U48231 (N_48231,N_47858,N_46109);
and U48232 (N_48232,N_46822,N_47621);
or U48233 (N_48233,N_46474,N_46155);
nor U48234 (N_48234,N_47578,N_46899);
and U48235 (N_48235,N_46797,N_46662);
or U48236 (N_48236,N_47271,N_46303);
nor U48237 (N_48237,N_47983,N_47292);
nand U48238 (N_48238,N_46300,N_46434);
or U48239 (N_48239,N_46378,N_46438);
nand U48240 (N_48240,N_47401,N_47052);
xnor U48241 (N_48241,N_47188,N_46630);
or U48242 (N_48242,N_46861,N_46620);
nor U48243 (N_48243,N_46614,N_47410);
nor U48244 (N_48244,N_46418,N_46812);
nand U48245 (N_48245,N_47582,N_47112);
nor U48246 (N_48246,N_46384,N_47000);
nor U48247 (N_48247,N_46470,N_47277);
and U48248 (N_48248,N_47107,N_47029);
and U48249 (N_48249,N_47780,N_46218);
and U48250 (N_48250,N_46926,N_46096);
nor U48251 (N_48251,N_46404,N_46641);
or U48252 (N_48252,N_47228,N_46392);
or U48253 (N_48253,N_47173,N_46573);
and U48254 (N_48254,N_47241,N_47635);
or U48255 (N_48255,N_46318,N_46080);
and U48256 (N_48256,N_46863,N_47714);
or U48257 (N_48257,N_47570,N_46986);
or U48258 (N_48258,N_47336,N_47903);
nand U48259 (N_48259,N_47729,N_47371);
xnor U48260 (N_48260,N_47170,N_47393);
nand U48261 (N_48261,N_46501,N_46224);
nand U48262 (N_48262,N_47018,N_46790);
nor U48263 (N_48263,N_47154,N_47098);
nor U48264 (N_48264,N_47056,N_46250);
nand U48265 (N_48265,N_46567,N_46532);
or U48266 (N_48266,N_47157,N_47922);
xnor U48267 (N_48267,N_46740,N_47683);
nor U48268 (N_48268,N_46466,N_46635);
or U48269 (N_48269,N_46759,N_47142);
or U48270 (N_48270,N_46369,N_47722);
or U48271 (N_48271,N_47191,N_46399);
nand U48272 (N_48272,N_46715,N_46280);
nor U48273 (N_48273,N_46173,N_47937);
nor U48274 (N_48274,N_47562,N_46492);
nand U48275 (N_48275,N_47253,N_47479);
and U48276 (N_48276,N_47085,N_46621);
nand U48277 (N_48277,N_46429,N_47152);
nand U48278 (N_48278,N_47890,N_47462);
nand U48279 (N_48279,N_47156,N_46362);
and U48280 (N_48280,N_47794,N_47229);
nand U48281 (N_48281,N_47260,N_46649);
or U48282 (N_48282,N_47353,N_47911);
or U48283 (N_48283,N_47317,N_47706);
or U48284 (N_48284,N_47584,N_46060);
nand U48285 (N_48285,N_47118,N_46234);
or U48286 (N_48286,N_47715,N_47305);
and U48287 (N_48287,N_46220,N_46912);
and U48288 (N_48288,N_46996,N_47593);
and U48289 (N_48289,N_46102,N_46940);
or U48290 (N_48290,N_46699,N_47730);
nand U48291 (N_48291,N_47080,N_46332);
or U48292 (N_48292,N_46856,N_47796);
xor U48293 (N_48293,N_46496,N_47604);
nor U48294 (N_48294,N_46352,N_47131);
xnor U48295 (N_48295,N_47213,N_46028);
nand U48296 (N_48296,N_46380,N_47808);
nor U48297 (N_48297,N_47197,N_46723);
nand U48298 (N_48298,N_46623,N_47536);
or U48299 (N_48299,N_46230,N_47289);
and U48300 (N_48300,N_46163,N_47613);
or U48301 (N_48301,N_46608,N_46656);
nor U48302 (N_48302,N_46153,N_47032);
and U48303 (N_48303,N_47881,N_47685);
nand U48304 (N_48304,N_47399,N_46842);
and U48305 (N_48305,N_46477,N_46011);
nand U48306 (N_48306,N_47695,N_47999);
or U48307 (N_48307,N_47413,N_46849);
nand U48308 (N_48308,N_47982,N_46798);
or U48309 (N_48309,N_46165,N_47422);
and U48310 (N_48310,N_47246,N_47164);
nand U48311 (N_48311,N_46585,N_46598);
nor U48312 (N_48312,N_47605,N_47798);
and U48313 (N_48313,N_46730,N_47956);
nor U48314 (N_48314,N_46193,N_47207);
nor U48315 (N_48315,N_47473,N_47084);
and U48316 (N_48316,N_47971,N_47743);
or U48317 (N_48317,N_46309,N_47916);
nor U48318 (N_48318,N_47278,N_46125);
and U48319 (N_48319,N_46613,N_47471);
or U48320 (N_48320,N_47731,N_47221);
nor U48321 (N_48321,N_47431,N_46506);
or U48322 (N_48322,N_46106,N_47560);
and U48323 (N_48323,N_46233,N_47887);
nor U48324 (N_48324,N_47629,N_47200);
nand U48325 (N_48325,N_46348,N_47764);
or U48326 (N_48326,N_46898,N_46068);
nor U48327 (N_48327,N_47051,N_47537);
and U48328 (N_48328,N_47095,N_46704);
nor U48329 (N_48329,N_46124,N_46786);
or U48330 (N_48330,N_47171,N_47513);
and U48331 (N_48331,N_47324,N_46745);
nor U48332 (N_48332,N_47806,N_47952);
or U48333 (N_48333,N_46198,N_46979);
or U48334 (N_48334,N_46859,N_47182);
or U48335 (N_48335,N_46678,N_46463);
nand U48336 (N_48336,N_46105,N_46469);
nor U48337 (N_48337,N_46811,N_46910);
nand U48338 (N_48338,N_46223,N_47805);
and U48339 (N_48339,N_46632,N_47283);
nand U48340 (N_48340,N_46599,N_46646);
or U48341 (N_48341,N_46526,N_46188);
nand U48342 (N_48342,N_46548,N_46827);
nand U48343 (N_48343,N_47797,N_46655);
nand U48344 (N_48344,N_46373,N_47360);
nor U48345 (N_48345,N_47693,N_46507);
and U48346 (N_48346,N_46014,N_47839);
or U48347 (N_48347,N_47541,N_46162);
and U48348 (N_48348,N_47242,N_46596);
nor U48349 (N_48349,N_47509,N_47040);
or U48350 (N_48350,N_46896,N_46388);
nand U48351 (N_48351,N_46026,N_47155);
or U48352 (N_48352,N_47625,N_46166);
nor U48353 (N_48353,N_46382,N_47932);
or U48354 (N_48354,N_47719,N_47506);
nand U48355 (N_48355,N_47416,N_47784);
nand U48356 (N_48356,N_47883,N_46770);
nor U48357 (N_48357,N_46481,N_47139);
nand U48358 (N_48358,N_47770,N_47717);
xnor U48359 (N_48359,N_46781,N_47359);
nand U48360 (N_48360,N_47619,N_47176);
nand U48361 (N_48361,N_47372,N_47571);
nand U48362 (N_48362,N_46838,N_46958);
nand U48363 (N_48363,N_47878,N_46107);
or U48364 (N_48364,N_46367,N_47319);
or U48365 (N_48365,N_47655,N_47876);
xor U48366 (N_48366,N_46100,N_46074);
and U48367 (N_48367,N_47723,N_47595);
or U48368 (N_48368,N_46519,N_47898);
or U48369 (N_48369,N_46512,N_47114);
or U48370 (N_48370,N_47122,N_46513);
nor U48371 (N_48371,N_46251,N_46685);
nand U48372 (N_48372,N_47162,N_46379);
and U48373 (N_48373,N_46335,N_47195);
or U48374 (N_48374,N_46361,N_46099);
and U48375 (N_48375,N_47691,N_46330);
nor U48376 (N_48376,N_47082,N_47859);
and U48377 (N_48377,N_47090,N_46042);
nor U48378 (N_48378,N_47113,N_46523);
and U48379 (N_48379,N_46572,N_46010);
nand U48380 (N_48380,N_46005,N_47231);
and U48381 (N_48381,N_47533,N_47592);
nor U48382 (N_48382,N_47934,N_47823);
nor U48383 (N_48383,N_46478,N_47670);
nor U48384 (N_48384,N_46073,N_46070);
or U48385 (N_48385,N_47857,N_46081);
nor U48386 (N_48386,N_47815,N_46801);
and U48387 (N_48387,N_46127,N_47280);
nor U48388 (N_48388,N_47833,N_47208);
nor U48389 (N_48389,N_47606,N_46370);
and U48390 (N_48390,N_47373,N_46938);
nand U48391 (N_48391,N_47352,N_46459);
nor U48392 (N_48392,N_46436,N_46046);
nor U48393 (N_48393,N_47093,N_47669);
nor U48394 (N_48394,N_46408,N_46075);
and U48395 (N_48395,N_46277,N_46298);
and U48396 (N_48396,N_46733,N_46187);
nor U48397 (N_48397,N_46098,N_47824);
xor U48398 (N_48398,N_46890,N_47284);
nand U48399 (N_48399,N_46441,N_46217);
nand U48400 (N_48400,N_46191,N_46920);
nand U48401 (N_48401,N_47385,N_47166);
or U48402 (N_48402,N_47042,N_47068);
xnor U48403 (N_48403,N_46575,N_47001);
and U48404 (N_48404,N_47761,N_46806);
nor U48405 (N_48405,N_47534,N_46793);
nor U48406 (N_48406,N_46853,N_47350);
and U48407 (N_48407,N_46398,N_46746);
nand U48408 (N_48408,N_47790,N_47094);
xnor U48409 (N_48409,N_46905,N_46967);
nor U48410 (N_48410,N_46588,N_47167);
nor U48411 (N_48411,N_47392,N_47875);
or U48412 (N_48412,N_46067,N_46955);
and U48413 (N_48413,N_46236,N_46709);
or U48414 (N_48414,N_46749,N_47608);
nor U48415 (N_48415,N_47682,N_46959);
xor U48416 (N_48416,N_47346,N_47400);
nor U48417 (N_48417,N_47756,N_46447);
nor U48418 (N_48418,N_47674,N_47974);
nor U48419 (N_48419,N_47665,N_46052);
or U48420 (N_48420,N_47909,N_46442);
nand U48421 (N_48421,N_47694,N_47994);
nand U48422 (N_48422,N_46977,N_47511);
and U48423 (N_48423,N_47844,N_47659);
nand U48424 (N_48424,N_47558,N_47384);
xor U48425 (N_48425,N_47128,N_47856);
and U48426 (N_48426,N_46593,N_47444);
nor U48427 (N_48427,N_47782,N_46147);
nor U48428 (N_48428,N_46754,N_46416);
or U48429 (N_48429,N_46887,N_47628);
nor U48430 (N_48430,N_46643,N_46134);
nor U48431 (N_48431,N_47115,N_47127);
and U48432 (N_48432,N_47574,N_46427);
or U48433 (N_48433,N_47701,N_46629);
and U48434 (N_48434,N_46500,N_47687);
nand U48435 (N_48435,N_47274,N_47273);
nor U48436 (N_48436,N_47580,N_46338);
nand U48437 (N_48437,N_47720,N_46296);
nor U48438 (N_48438,N_46603,N_47138);
or U48439 (N_48439,N_47233,N_47261);
nand U48440 (N_48440,N_46862,N_47874);
or U48441 (N_48441,N_46561,N_46006);
and U48442 (N_48442,N_46411,N_46445);
nand U48443 (N_48443,N_47071,N_46651);
nand U48444 (N_48444,N_47546,N_47463);
or U48445 (N_48445,N_46254,N_46241);
and U48446 (N_48446,N_47676,N_46895);
nand U48447 (N_48447,N_47573,N_46464);
nand U48448 (N_48448,N_46211,N_47159);
or U48449 (N_48449,N_47966,N_47929);
and U48450 (N_48450,N_47145,N_46104);
and U48451 (N_48451,N_46916,N_47299);
nor U48452 (N_48452,N_47590,N_46804);
nor U48453 (N_48453,N_46776,N_46889);
nor U48454 (N_48454,N_47567,N_46871);
nand U48455 (N_48455,N_46918,N_47135);
nor U48456 (N_48456,N_47602,N_46873);
nand U48457 (N_48457,N_47320,N_47959);
and U48458 (N_48458,N_46936,N_47019);
or U48459 (N_48459,N_46462,N_46425);
nor U48460 (N_48460,N_47187,N_47821);
or U48461 (N_48461,N_46999,N_46533);
nand U48462 (N_48462,N_47101,N_47623);
or U48463 (N_48463,N_46265,N_46880);
nand U48464 (N_48464,N_47633,N_46064);
and U48465 (N_48465,N_46476,N_47297);
nor U48466 (N_48466,N_46008,N_47742);
nand U48467 (N_48467,N_46047,N_47678);
or U48468 (N_48468,N_47076,N_46845);
or U48469 (N_48469,N_46403,N_47528);
and U48470 (N_48470,N_47965,N_46056);
nand U48471 (N_48471,N_46547,N_46720);
and U48472 (N_48472,N_46768,N_47967);
nand U48473 (N_48473,N_46262,N_47436);
or U48474 (N_48474,N_46948,N_46183);
and U48475 (N_48475,N_46195,N_47620);
nand U48476 (N_48476,N_46239,N_46944);
nor U48477 (N_48477,N_47451,N_46706);
nor U48478 (N_48478,N_46969,N_47820);
nor U48479 (N_48479,N_47727,N_46383);
nand U48480 (N_48480,N_47117,N_46931);
or U48481 (N_48481,N_46454,N_47355);
nor U48482 (N_48482,N_46059,N_46467);
nor U48483 (N_48483,N_46118,N_47739);
nand U48484 (N_48484,N_47491,N_47705);
nor U48485 (N_48485,N_46235,N_46090);
or U48486 (N_48486,N_46764,N_47921);
or U48487 (N_48487,N_46925,N_46792);
nor U48488 (N_48488,N_47252,N_46040);
and U48489 (N_48489,N_46440,N_47940);
or U48490 (N_48490,N_47163,N_46767);
xnor U48491 (N_48491,N_46985,N_46844);
nor U48492 (N_48492,N_46870,N_47276);
or U48493 (N_48493,N_46647,N_46509);
or U48494 (N_48494,N_47334,N_46659);
nor U48495 (N_48495,N_46617,N_47492);
nand U48496 (N_48496,N_47732,N_47189);
nor U48497 (N_48497,N_47035,N_46366);
nand U48498 (N_48498,N_46592,N_47004);
and U48499 (N_48499,N_46734,N_46019);
nor U48500 (N_48500,N_46083,N_46009);
and U48501 (N_48501,N_47369,N_46371);
nor U48502 (N_48502,N_47969,N_47596);
nand U48503 (N_48503,N_47402,N_46184);
nand U48504 (N_48504,N_46669,N_47025);
nor U48505 (N_48505,N_46616,N_47597);
nand U48506 (N_48506,N_47539,N_46521);
or U48507 (N_48507,N_46992,N_46003);
nor U48508 (N_48508,N_46552,N_47488);
and U48509 (N_48509,N_47979,N_46805);
or U48510 (N_48510,N_47222,N_47452);
and U48511 (N_48511,N_47549,N_47942);
or U48512 (N_48512,N_46327,N_46933);
and U48513 (N_48513,N_47817,N_46131);
xor U48514 (N_48514,N_46432,N_46973);
nor U48515 (N_48515,N_46525,N_47901);
nand U48516 (N_48516,N_46884,N_46891);
and U48517 (N_48517,N_46901,N_46168);
or U48518 (N_48518,N_47753,N_47963);
and U48519 (N_48519,N_47459,N_47232);
or U48520 (N_48520,N_47885,N_47811);
nand U48521 (N_48521,N_47889,N_46452);
or U48522 (N_48522,N_46304,N_47800);
nor U48523 (N_48523,N_46607,N_47168);
nand U48524 (N_48524,N_46800,N_46085);
nand U48525 (N_48525,N_46156,N_46747);
nor U48526 (N_48526,N_47016,N_46670);
nand U48527 (N_48527,N_46020,N_47984);
nand U48528 (N_48528,N_47408,N_46517);
and U48529 (N_48529,N_46594,N_46888);
or U48530 (N_48530,N_46690,N_46839);
and U48531 (N_48531,N_46086,N_47150);
or U48532 (N_48532,N_46823,N_47250);
nand U48533 (N_48533,N_46212,N_46582);
nor U48534 (N_48534,N_46446,N_47177);
or U48535 (N_48535,N_47814,N_47419);
nor U48536 (N_48536,N_47442,N_47489);
xor U48537 (N_48537,N_47225,N_47264);
and U48538 (N_48538,N_46231,N_47239);
nand U48539 (N_48539,N_47599,N_46631);
or U48540 (N_48540,N_47009,N_47124);
and U48541 (N_48541,N_46129,N_47069);
and U48542 (N_48542,N_46850,N_46544);
or U48543 (N_48543,N_47990,N_47866);
nor U48544 (N_48544,N_47206,N_47230);
nor U48545 (N_48545,N_47663,N_47067);
nor U48546 (N_48546,N_46160,N_47356);
nor U48547 (N_48547,N_47930,N_46538);
and U48548 (N_48548,N_47995,N_46322);
and U48549 (N_48549,N_47382,N_46774);
nand U48550 (N_48550,N_47151,N_46044);
or U48551 (N_48551,N_46170,N_47892);
nand U48552 (N_48552,N_46435,N_46854);
nor U48553 (N_48553,N_46078,N_46333);
nor U48554 (N_48554,N_46121,N_46753);
nor U48555 (N_48555,N_46228,N_47810);
and U48556 (N_48556,N_46283,N_47517);
nand U48557 (N_48557,N_46682,N_47158);
nand U48558 (N_48558,N_47111,N_46255);
or U48559 (N_48559,N_46788,N_46157);
xor U48560 (N_48560,N_46138,N_46624);
and U48561 (N_48561,N_47216,N_47193);
xor U48562 (N_48562,N_46063,N_46494);
nand U48563 (N_48563,N_46974,N_46267);
or U48564 (N_48564,N_47914,N_46942);
or U48565 (N_48565,N_47951,N_46820);
xnor U48566 (N_48566,N_47179,N_47552);
xor U48567 (N_48567,N_46989,N_46991);
or U48568 (N_48568,N_47496,N_47779);
nand U48569 (N_48569,N_46269,N_47020);
and U48570 (N_48570,N_47666,N_47919);
or U48571 (N_48571,N_46537,N_47467);
or U48572 (N_48572,N_47637,N_47550);
or U48573 (N_48573,N_46729,N_47520);
nor U48574 (N_48574,N_46816,N_46726);
or U48575 (N_48575,N_47854,N_47443);
and U48576 (N_48576,N_47924,N_46253);
nor U48577 (N_48577,N_47842,N_46765);
and U48578 (N_48578,N_47765,N_46149);
or U48579 (N_48579,N_47394,N_47100);
and U48580 (N_48580,N_46701,N_47063);
and U48581 (N_48581,N_46443,N_46354);
or U48582 (N_48582,N_47470,N_47716);
nand U48583 (N_48583,N_47769,N_46167);
nand U48584 (N_48584,N_47540,N_46914);
nand U48585 (N_48585,N_47572,N_46637);
and U48586 (N_48586,N_46002,N_47852);
nor U48587 (N_48587,N_47760,N_47634);
or U48588 (N_48588,N_46258,N_47972);
nor U48589 (N_48589,N_46039,N_46143);
nor U48590 (N_48590,N_46148,N_46089);
nor U48591 (N_48591,N_46227,N_46428);
nor U48592 (N_48592,N_46036,N_46897);
nand U48593 (N_48593,N_47624,N_47495);
nor U48594 (N_48594,N_46095,N_46807);
and U48595 (N_48595,N_47226,N_47906);
nand U48596 (N_48596,N_47288,N_47038);
xnor U48597 (N_48597,N_47918,N_47148);
nor U48598 (N_48598,N_46627,N_47411);
or U48599 (N_48599,N_47468,N_46420);
and U48600 (N_48600,N_46389,N_46570);
nor U48601 (N_48601,N_46674,N_46221);
nand U48602 (N_48602,N_47658,N_46278);
nand U48603 (N_48603,N_46203,N_47290);
xnor U48604 (N_48604,N_47660,N_47792);
and U48605 (N_48605,N_47417,N_46535);
or U48606 (N_48606,N_47945,N_47308);
nand U48607 (N_48607,N_46214,N_47643);
xor U48608 (N_48608,N_47186,N_46557);
or U48609 (N_48609,N_47427,N_47532);
or U48610 (N_48610,N_47828,N_46007);
and U48611 (N_48611,N_47448,N_47012);
nand U48612 (N_48612,N_46421,N_47585);
or U48613 (N_48613,N_46472,N_47644);
or U48614 (N_48614,N_47680,N_46705);
or U48615 (N_48615,N_46796,N_46885);
xnor U48616 (N_48616,N_46215,N_46340);
nand U48617 (N_48617,N_46568,N_46828);
nor U48618 (N_48618,N_47065,N_46636);
and U48619 (N_48619,N_47850,N_46530);
and U48620 (N_48620,N_46980,N_47099);
or U48621 (N_48621,N_46055,N_46900);
nor U48622 (N_48622,N_46344,N_47786);
and U48623 (N_48623,N_47535,N_47365);
nor U48624 (N_48624,N_46094,N_46562);
or U48625 (N_48625,N_46069,N_46560);
nor U48626 (N_48626,N_46903,N_47343);
nand U48627 (N_48627,N_46619,N_46238);
nand U48628 (N_48628,N_46857,N_46904);
nor U48629 (N_48629,N_47936,N_47555);
nand U48630 (N_48630,N_46586,N_47622);
xnor U48631 (N_48631,N_46766,N_46676);
nor U48632 (N_48632,N_47367,N_47827);
and U48633 (N_48633,N_47328,N_47219);
and U48634 (N_48634,N_46702,N_47407);
and U48635 (N_48635,N_46312,N_47662);
nor U48636 (N_48636,N_47129,N_47904);
xnor U48637 (N_48637,N_46347,N_46386);
xor U48638 (N_48638,N_47120,N_47559);
and U48639 (N_48639,N_46461,N_46108);
or U48640 (N_48640,N_46504,N_46681);
nor U48641 (N_48641,N_46732,N_46728);
nor U48642 (N_48642,N_47863,N_46294);
or U48643 (N_48643,N_47609,N_46468);
or U48644 (N_48644,N_46136,N_47255);
or U48645 (N_48645,N_46957,N_46171);
xor U48646 (N_48646,N_46196,N_47583);
nor U48647 (N_48647,N_47767,N_46455);
and U48648 (N_48648,N_46306,N_46739);
nor U48649 (N_48649,N_46115,N_46093);
nor U48650 (N_48650,N_47414,N_46565);
nor U48651 (N_48651,N_47589,N_46048);
nor U48652 (N_48652,N_46694,N_46307);
nand U48653 (N_48653,N_47793,N_46484);
and U48654 (N_48654,N_46210,N_47269);
nor U48655 (N_48655,N_47861,N_46451);
and U48656 (N_48656,N_47341,N_47588);
nor U48657 (N_48657,N_47140,N_47348);
and U48658 (N_48658,N_46261,N_47561);
nand U48659 (N_48659,N_46772,N_46527);
nor U48660 (N_48660,N_47899,N_47146);
or U48661 (N_48661,N_47379,N_47566);
nor U48662 (N_48662,N_46953,N_47461);
nand U48663 (N_48663,N_46175,N_46406);
nor U48664 (N_48664,N_47086,N_47943);
nor U48665 (N_48665,N_47758,N_47865);
and U48666 (N_48666,N_46906,N_46528);
or U48667 (N_48667,N_46202,N_47031);
or U48668 (N_48668,N_46868,N_47234);
and U48669 (N_48669,N_46204,N_46057);
and U48670 (N_48670,N_47576,N_47646);
or U48671 (N_48671,N_46297,N_47736);
or U48672 (N_48672,N_46021,N_47105);
nand U48673 (N_48673,N_47938,N_47789);
nor U48674 (N_48674,N_47968,N_47598);
nor U48675 (N_48675,N_46667,N_46744);
and U48676 (N_48676,N_46493,N_47917);
or U48677 (N_48677,N_47829,N_47771);
xor U48678 (N_48678,N_47944,N_46284);
or U48679 (N_48679,N_46394,N_46686);
xor U48680 (N_48680,N_47612,N_47291);
and U48681 (N_48681,N_47144,N_46965);
nor U48682 (N_48682,N_47618,N_47668);
nor U48683 (N_48683,N_46128,N_47003);
nor U48684 (N_48684,N_47270,N_46079);
and U48685 (N_48685,N_46954,N_47106);
or U48686 (N_48686,N_47344,N_47415);
nor U48687 (N_48687,N_46146,N_46321);
nor U48688 (N_48688,N_46644,N_46076);
nor U48689 (N_48689,N_46393,N_47119);
or U48690 (N_48690,N_47873,N_46751);
nor U48691 (N_48691,N_47301,N_47862);
or U48692 (N_48692,N_46141,N_46625);
or U48693 (N_48693,N_46984,N_47224);
nor U48694 (N_48694,N_47321,N_46529);
nand U48695 (N_48695,N_46540,N_46061);
nor U48696 (N_48696,N_46864,N_46990);
and U48697 (N_48697,N_47645,N_46256);
nor U48698 (N_48698,N_47950,N_46293);
or U48699 (N_48699,N_47766,N_46652);
nor U48700 (N_48700,N_46949,N_46679);
nor U48701 (N_48701,N_46482,N_47337);
nor U48702 (N_48702,N_46794,N_46226);
nor U48703 (N_48703,N_47631,N_46032);
or U48704 (N_48704,N_46534,N_46993);
nand U48705 (N_48705,N_47689,N_47026);
or U48706 (N_48706,N_46243,N_47704);
nor U48707 (N_48707,N_47272,N_46762);
nand U48708 (N_48708,N_46539,N_47725);
and U48709 (N_48709,N_46414,N_46609);
or U48710 (N_48710,N_47781,N_47424);
nand U48711 (N_48711,N_47258,N_46584);
nand U48712 (N_48712,N_47939,N_46375);
nor U48713 (N_48713,N_46437,N_46549);
or U48714 (N_48714,N_47664,N_47174);
nor U48715 (N_48715,N_46317,N_46757);
or U48716 (N_48716,N_46355,N_47777);
nand U48717 (N_48717,N_46810,N_46190);
and U48718 (N_48718,N_47768,N_46490);
or U48719 (N_48719,N_47775,N_46132);
and U48720 (N_48720,N_46671,N_46866);
nor U48721 (N_48721,N_46169,N_46922);
nor U48722 (N_48722,N_46407,N_46813);
or U48723 (N_48723,N_47380,N_47529);
or U48724 (N_48724,N_46692,N_47266);
nor U48725 (N_48725,N_46091,N_47332);
or U48726 (N_48726,N_47543,N_47428);
or U48727 (N_48727,N_46597,N_46433);
nand U48728 (N_48728,N_47617,N_46126);
nand U48729 (N_48729,N_46872,N_46120);
nand U48730 (N_48730,N_46374,N_47198);
and U48731 (N_48731,N_46555,N_47494);
or U48732 (N_48732,N_47316,N_46219);
nand U48733 (N_48733,N_47600,N_46395);
or U48734 (N_48734,N_46604,N_47480);
xor U48735 (N_48735,N_46365,N_46426);
and U48736 (N_48736,N_46113,N_47915);
nand U48737 (N_48737,N_46932,N_46708);
and U48738 (N_48738,N_47926,N_47338);
nand U48739 (N_48739,N_47430,N_46242);
or U48740 (N_48740,N_47708,N_46186);
nor U48741 (N_48741,N_47390,N_47484);
and U48742 (N_48742,N_46886,N_46405);
and U48743 (N_48743,N_46775,N_47752);
nor U48744 (N_48744,N_46566,N_46983);
nand U48745 (N_48745,N_46894,N_46640);
nand U48746 (N_48746,N_47686,N_46456);
or U48747 (N_48747,N_47074,N_46881);
and U48748 (N_48748,N_47684,N_46323);
nand U48749 (N_48749,N_47243,N_47201);
or U48750 (N_48750,N_46997,N_46319);
nand U48751 (N_48751,N_46130,N_46771);
nand U48752 (N_48752,N_47481,N_47498);
nor U48753 (N_48753,N_47650,N_46908);
nand U48754 (N_48754,N_47626,N_47259);
nor U48755 (N_48755,N_47737,N_47841);
and U48756 (N_48756,N_47835,N_46152);
or U48757 (N_48757,N_46737,N_47750);
nor U48758 (N_48758,N_47831,N_47977);
and U48759 (N_48759,N_47172,N_46117);
nand U48760 (N_48760,N_47050,N_47542);
xnor U48761 (N_48761,N_47499,N_47143);
nand U48762 (N_48762,N_47432,N_47310);
and U48763 (N_48763,N_46780,N_47361);
or U48764 (N_48764,N_47697,N_46672);
nor U48765 (N_48765,N_47235,N_47514);
nand U48766 (N_48766,N_47791,N_46963);
nand U48767 (N_48767,N_47194,N_47383);
or U48768 (N_48768,N_47329,N_47961);
and U48769 (N_48769,N_47712,N_47057);
and U48770 (N_48770,N_47061,N_46791);
or U48771 (N_48771,N_47880,N_47391);
nand U48772 (N_48772,N_46591,N_46346);
nor U48773 (N_48773,N_46359,N_47893);
and U48774 (N_48774,N_47949,N_46161);
or U48775 (N_48775,N_47293,N_46982);
nand U48776 (N_48776,N_47314,N_46450);
and U48777 (N_48777,N_46275,N_47738);
nand U48778 (N_48778,N_46556,N_46855);
nor U48779 (N_48779,N_46563,N_47487);
and U48780 (N_48780,N_47196,N_47017);
and U48781 (N_48781,N_47941,N_46921);
nor U48782 (N_48782,N_46174,N_47581);
and U48783 (N_48783,N_46257,N_47946);
and U48784 (N_48784,N_47902,N_46103);
nor U48785 (N_48785,N_47648,N_46626);
nand U48786 (N_48786,N_47813,N_46205);
nor U48787 (N_48787,N_46511,N_47508);
nor U48788 (N_48788,N_47587,N_47955);
or U48789 (N_48789,N_46197,N_46841);
or U48790 (N_48790,N_46314,N_47169);
or U48791 (N_48791,N_46840,N_47339);
and U48792 (N_48792,N_46004,N_47349);
or U48793 (N_48793,N_47014,N_46041);
nor U48794 (N_48794,N_47925,N_46422);
and U48795 (N_48795,N_47547,N_47477);
and U48796 (N_48796,N_46665,N_47426);
and U48797 (N_48797,N_47075,N_47707);
nand U48798 (N_48798,N_46510,N_46577);
and U48799 (N_48799,N_47342,N_46893);
and U48800 (N_48800,N_46194,N_47351);
nand U48801 (N_48801,N_46201,N_47525);
and U48802 (N_48802,N_46316,N_47046);
nor U48803 (N_48803,N_46181,N_46564);
xor U48804 (N_48804,N_46892,N_46092);
nor U48805 (N_48805,N_47868,N_46911);
and U48806 (N_48806,N_47962,N_46545);
and U48807 (N_48807,N_46172,N_47435);
nor U48808 (N_48808,N_46058,N_47130);
nor U48809 (N_48809,N_46716,N_47249);
nand U48810 (N_48810,N_46645,N_47615);
nor U48811 (N_48811,N_46727,N_46837);
xnor U48812 (N_48812,N_47281,N_47078);
nand U48813 (N_48813,N_47011,N_46831);
nand U48814 (N_48814,N_47110,N_46430);
nor U48815 (N_48815,N_47287,N_46049);
or U48816 (N_48816,N_47507,N_46587);
nand U48817 (N_48817,N_47510,N_47345);
or U48818 (N_48818,N_47180,N_46351);
or U48819 (N_48819,N_47036,N_47776);
nand U48820 (N_48820,N_46396,N_46263);
nor U48821 (N_48821,N_46777,N_47055);
and U48822 (N_48822,N_46097,N_46023);
and U48823 (N_48823,N_47554,N_46515);
nand U48824 (N_48824,N_46654,N_46024);
and U48825 (N_48825,N_47726,N_46988);
nand U48826 (N_48826,N_47302,N_47741);
nor U48827 (N_48827,N_47973,N_47825);
nor U48828 (N_48828,N_46778,N_46981);
nand U48829 (N_48829,N_46697,N_47860);
and U48830 (N_48830,N_47734,N_47757);
nand U48831 (N_48831,N_46087,N_47066);
nand U48832 (N_48832,N_46542,N_46691);
nor U48833 (N_48833,N_46270,N_46700);
and U48834 (N_48834,N_47434,N_47638);
nand U48835 (N_48835,N_46722,N_47987);
nor U48836 (N_48836,N_46449,N_47846);
and U48837 (N_48837,N_46602,N_47538);
nor U48838 (N_48838,N_47888,N_47544);
nand U48839 (N_48839,N_47954,N_47907);
or U48840 (N_48840,N_46518,N_47998);
and U48841 (N_48841,N_46524,N_47137);
nand U48842 (N_48842,N_47423,N_46551);
xor U48843 (N_48843,N_47460,N_47149);
nand U48844 (N_48844,N_46349,N_46116);
and U48845 (N_48845,N_46151,N_46301);
nor U48846 (N_48846,N_47002,N_46826);
and U48847 (N_48847,N_47675,N_46326);
nand U48848 (N_48848,N_46343,N_47749);
nand U48849 (N_48849,N_46062,N_46015);
nand U48850 (N_48850,N_46978,N_47773);
or U48851 (N_48851,N_47053,N_47049);
or U48852 (N_48852,N_47627,N_47728);
nand U48853 (N_48853,N_47087,N_47551);
nor U48854 (N_48854,N_47453,N_46829);
nand U48855 (N_48855,N_46714,N_47263);
and U48856 (N_48856,N_46377,N_46761);
nand U48857 (N_48857,N_47141,N_46998);
or U48858 (N_48858,N_46550,N_46337);
or U48859 (N_48859,N_46668,N_47354);
xor U48860 (N_48860,N_46285,N_47867);
nor U48861 (N_48861,N_46497,N_46951);
nand U48862 (N_48862,N_46390,N_46364);
nand U48863 (N_48863,N_46858,N_46000);
or U48864 (N_48864,N_47472,N_46353);
nand U48865 (N_48865,N_46907,N_46677);
or U48866 (N_48866,N_47318,N_46229);
and U48867 (N_48867,N_46516,N_47248);
nor U48868 (N_48868,N_46460,N_47450);
and U48869 (N_48869,N_47652,N_47964);
nand U48870 (N_48870,N_46832,N_47799);
and U48871 (N_48871,N_47024,N_46755);
nor U48872 (N_48872,N_47700,N_46779);
and U48873 (N_48873,N_46176,N_47088);
nor U48874 (N_48874,N_47268,N_47482);
or U48875 (N_48875,N_47097,N_46514);
and U48876 (N_48876,N_47834,N_46943);
nor U48877 (N_48877,N_47446,N_46622);
nand U48878 (N_48878,N_47322,N_47315);
and U48879 (N_48879,N_47178,N_47091);
and U48880 (N_48880,N_47774,N_47569);
nor U48881 (N_48881,N_47376,N_46180);
and U48882 (N_48882,N_46144,N_46928);
or U48883 (N_48883,N_47267,N_46687);
nand U48884 (N_48884,N_46595,N_47870);
nand U48885 (N_48885,N_47832,N_47545);
and U48886 (N_48886,N_46413,N_47403);
or U48887 (N_48887,N_47033,N_47611);
nand U48888 (N_48888,N_47398,N_46874);
nand U48889 (N_48889,N_46929,N_47524);
nand U48890 (N_48890,N_46663,N_46084);
nand U48891 (N_48891,N_46150,N_46054);
nand U48892 (N_48892,N_46288,N_46851);
xnor U48893 (N_48893,N_46281,N_46289);
and U48894 (N_48894,N_47747,N_47190);
nand U48895 (N_48895,N_47869,N_47079);
and U48896 (N_48896,N_47358,N_47993);
and U48897 (N_48897,N_47871,N_46825);
nand U48898 (N_48898,N_47884,N_46648);
and U48899 (N_48899,N_47412,N_47386);
nand U48900 (N_48900,N_47483,N_47953);
or U48901 (N_48901,N_47323,N_47677);
and U48902 (N_48902,N_47647,N_47147);
or U48903 (N_48903,N_47772,N_46520);
nand U48904 (N_48904,N_47262,N_47363);
and U48905 (N_48905,N_47418,N_47409);
xnor U48906 (N_48906,N_47311,N_47134);
and U48907 (N_48907,N_47975,N_46178);
nor U48908 (N_48908,N_46815,N_46164);
nor U48909 (N_48909,N_47733,N_46664);
and U48910 (N_48910,N_47816,N_46133);
and U48911 (N_48911,N_46693,N_46719);
nor U48912 (N_48912,N_47845,N_47286);
and U48913 (N_48913,N_47783,N_46012);
nand U48914 (N_48914,N_47778,N_46657);
nand U48915 (N_48915,N_47041,N_47803);
or U48916 (N_48916,N_46199,N_47326);
or U48917 (N_48917,N_46417,N_46846);
nor U48918 (N_48918,N_47616,N_47642);
nor U48919 (N_48919,N_46503,N_46439);
and U48920 (N_48920,N_46927,N_47809);
nand U48921 (N_48921,N_47185,N_46448);
nand U48922 (N_48922,N_46245,N_46580);
and U48923 (N_48923,N_46946,N_46843);
or U48924 (N_48924,N_46934,N_46618);
or U48925 (N_48925,N_47240,N_46017);
or U48926 (N_48926,N_47300,N_46968);
or U48927 (N_48927,N_47212,N_46975);
nand U48928 (N_48928,N_47083,N_46783);
and U48929 (N_48929,N_47132,N_47667);
or U48930 (N_48930,N_47420,N_46475);
nor U48931 (N_48931,N_47126,N_47864);
or U48932 (N_48932,N_46961,N_46695);
nand U48933 (N_48933,N_46415,N_47721);
nand U48934 (N_48934,N_47313,N_46799);
nand U48935 (N_48935,N_46583,N_47437);
nor U48936 (N_48936,N_47745,N_47486);
nor U48937 (N_48937,N_47503,N_46601);
nand U48938 (N_48938,N_47636,N_46673);
and U48939 (N_48939,N_46536,N_46045);
nand U48940 (N_48940,N_46342,N_47657);
nand U48941 (N_48941,N_47347,N_47978);
xnor U48942 (N_48942,N_46995,N_46502);
and U48943 (N_48943,N_47466,N_47848);
and U48944 (N_48944,N_46334,N_47610);
and U48945 (N_48945,N_47527,N_46240);
and U48946 (N_48946,N_46207,N_46208);
or U48947 (N_48947,N_47397,N_46302);
nor U48948 (N_48948,N_46247,N_47787);
and U48949 (N_48949,N_47044,N_46558);
nand U48950 (N_48950,N_46683,N_46782);
or U48951 (N_48951,N_47523,N_46119);
or U48952 (N_48952,N_46937,N_46387);
or U48953 (N_48953,N_46748,N_47690);
or U48954 (N_48954,N_46471,N_46941);
nor U48955 (N_48955,N_46271,N_46741);
and U48956 (N_48956,N_47374,N_47096);
and U48957 (N_48957,N_47928,N_46546);
and U48958 (N_48958,N_46179,N_47405);
xor U48959 (N_48959,N_46752,N_47440);
or U48960 (N_48960,N_47556,N_47265);
nor U48961 (N_48961,N_46814,N_47710);
nand U48962 (N_48962,N_47060,N_47671);
and U48963 (N_48963,N_46787,N_46553);
xnor U48964 (N_48964,N_47455,N_47306);
or U48965 (N_48965,N_46401,N_47387);
or U48966 (N_48966,N_47161,N_46137);
or U48967 (N_48967,N_46419,N_47285);
nand U48968 (N_48968,N_46368,N_46763);
nor U48969 (N_48969,N_46590,N_47515);
and U48970 (N_48970,N_47377,N_47986);
xor U48971 (N_48971,N_47948,N_46272);
and U48972 (N_48972,N_47298,N_46962);
nand U48973 (N_48973,N_46939,N_46145);
or U48974 (N_48974,N_47614,N_47121);
or U48975 (N_48975,N_47389,N_46273);
and U48976 (N_48976,N_47449,N_46559);
or U48977 (N_48977,N_47853,N_46372);
nor U48978 (N_48978,N_47175,N_47502);
and U48979 (N_48979,N_46819,N_46274);
nor U48980 (N_48980,N_46785,N_46453);
nor U48981 (N_48981,N_46976,N_47013);
nor U48982 (N_48982,N_47996,N_47653);
and U48983 (N_48983,N_46571,N_46970);
nand U48984 (N_48984,N_46924,N_47439);
nor U48985 (N_48985,N_47740,N_46960);
or U48986 (N_48986,N_46742,N_47512);
nand U48987 (N_48987,N_46758,N_47826);
or U48988 (N_48988,N_46711,N_46773);
nor U48989 (N_48989,N_46696,N_47136);
nor U48990 (N_48990,N_47713,N_47102);
or U48991 (N_48991,N_47702,N_46836);
or U48992 (N_48992,N_46710,N_47421);
nor U48993 (N_48993,N_46320,N_47425);
nor U48994 (N_48994,N_47526,N_47891);
and U48995 (N_48995,N_47478,N_47464);
or U48996 (N_48996,N_46950,N_47227);
nor U48997 (N_48997,N_47516,N_47957);
nor U48998 (N_48998,N_46522,N_46177);
or U48999 (N_48999,N_47607,N_46345);
or U49000 (N_49000,N_47798,N_46660);
nor U49001 (N_49001,N_46881,N_47205);
or U49002 (N_49002,N_47099,N_47709);
nand U49003 (N_49003,N_46910,N_47581);
or U49004 (N_49004,N_47212,N_47238);
or U49005 (N_49005,N_46813,N_47267);
nand U49006 (N_49006,N_46661,N_46569);
nor U49007 (N_49007,N_46731,N_47333);
nand U49008 (N_49008,N_47055,N_47329);
or U49009 (N_49009,N_47510,N_46468);
nand U49010 (N_49010,N_46715,N_46040);
or U49011 (N_49011,N_47888,N_47253);
and U49012 (N_49012,N_47127,N_47045);
nor U49013 (N_49013,N_46762,N_47516);
nor U49014 (N_49014,N_47063,N_46328);
nor U49015 (N_49015,N_47060,N_47558);
or U49016 (N_49016,N_47305,N_47085);
xor U49017 (N_49017,N_46377,N_46568);
nand U49018 (N_49018,N_46777,N_47605);
nand U49019 (N_49019,N_47663,N_46845);
and U49020 (N_49020,N_46509,N_46015);
or U49021 (N_49021,N_46261,N_46381);
nand U49022 (N_49022,N_46641,N_47357);
and U49023 (N_49023,N_46809,N_47456);
xnor U49024 (N_49024,N_47012,N_47643);
and U49025 (N_49025,N_47244,N_47591);
xor U49026 (N_49026,N_47675,N_46466);
and U49027 (N_49027,N_46927,N_47440);
and U49028 (N_49028,N_47387,N_46297);
nand U49029 (N_49029,N_47393,N_47347);
nand U49030 (N_49030,N_46503,N_47051);
nor U49031 (N_49031,N_47803,N_46689);
nor U49032 (N_49032,N_47435,N_46599);
or U49033 (N_49033,N_46368,N_46204);
and U49034 (N_49034,N_46081,N_47663);
nand U49035 (N_49035,N_47730,N_46045);
nand U49036 (N_49036,N_47608,N_47724);
nand U49037 (N_49037,N_46834,N_46336);
and U49038 (N_49038,N_47650,N_47022);
nor U49039 (N_49039,N_47508,N_46156);
or U49040 (N_49040,N_46101,N_46387);
and U49041 (N_49041,N_46949,N_47088);
and U49042 (N_49042,N_47074,N_47856);
nor U49043 (N_49043,N_46871,N_46847);
nor U49044 (N_49044,N_46861,N_46416);
nor U49045 (N_49045,N_47311,N_46016);
and U49046 (N_49046,N_46933,N_47853);
nor U49047 (N_49047,N_47466,N_46939);
or U49048 (N_49048,N_47851,N_47037);
nand U49049 (N_49049,N_47309,N_46159);
nor U49050 (N_49050,N_46447,N_47532);
or U49051 (N_49051,N_47219,N_46512);
and U49052 (N_49052,N_46511,N_47201);
nor U49053 (N_49053,N_46723,N_47088);
or U49054 (N_49054,N_47189,N_46322);
nand U49055 (N_49055,N_47872,N_47085);
xor U49056 (N_49056,N_47829,N_46369);
nand U49057 (N_49057,N_46433,N_47877);
nor U49058 (N_49058,N_46509,N_47776);
nor U49059 (N_49059,N_46718,N_47272);
and U49060 (N_49060,N_47727,N_47830);
nand U49061 (N_49061,N_46451,N_46461);
nor U49062 (N_49062,N_46324,N_46188);
nand U49063 (N_49063,N_46796,N_47813);
or U49064 (N_49064,N_46596,N_47716);
nor U49065 (N_49065,N_47887,N_47197);
nor U49066 (N_49066,N_47123,N_46023);
or U49067 (N_49067,N_47214,N_47330);
or U49068 (N_49068,N_47030,N_46855);
and U49069 (N_49069,N_46067,N_46469);
nand U49070 (N_49070,N_46096,N_47767);
nand U49071 (N_49071,N_46569,N_47208);
and U49072 (N_49072,N_46343,N_47711);
or U49073 (N_49073,N_46850,N_47568);
and U49074 (N_49074,N_46270,N_46735);
nor U49075 (N_49075,N_46721,N_46148);
xnor U49076 (N_49076,N_47033,N_46797);
or U49077 (N_49077,N_47326,N_46738);
and U49078 (N_49078,N_47158,N_47150);
or U49079 (N_49079,N_46553,N_47757);
nor U49080 (N_49080,N_46392,N_46377);
and U49081 (N_49081,N_46920,N_47033);
or U49082 (N_49082,N_47588,N_46971);
nand U49083 (N_49083,N_46038,N_46363);
or U49084 (N_49084,N_47415,N_46750);
nand U49085 (N_49085,N_46065,N_46551);
nand U49086 (N_49086,N_46782,N_47350);
nand U49087 (N_49087,N_47932,N_47339);
or U49088 (N_49088,N_46030,N_46361);
or U49089 (N_49089,N_47367,N_46514);
or U49090 (N_49090,N_47868,N_46256);
or U49091 (N_49091,N_47788,N_46744);
or U49092 (N_49092,N_46293,N_46912);
nand U49093 (N_49093,N_46966,N_46915);
nand U49094 (N_49094,N_46731,N_46370);
nand U49095 (N_49095,N_47962,N_46422);
or U49096 (N_49096,N_47291,N_46902);
nor U49097 (N_49097,N_47206,N_47295);
and U49098 (N_49098,N_46480,N_47823);
nand U49099 (N_49099,N_46673,N_47850);
or U49100 (N_49100,N_46915,N_47915);
nor U49101 (N_49101,N_47264,N_47143);
and U49102 (N_49102,N_46524,N_47072);
and U49103 (N_49103,N_47497,N_46358);
xor U49104 (N_49104,N_46180,N_46787);
and U49105 (N_49105,N_47733,N_46541);
nor U49106 (N_49106,N_46612,N_47687);
and U49107 (N_49107,N_47551,N_47963);
xnor U49108 (N_49108,N_46270,N_47786);
or U49109 (N_49109,N_47618,N_47470);
nor U49110 (N_49110,N_47891,N_47836);
nand U49111 (N_49111,N_46429,N_47117);
nor U49112 (N_49112,N_47232,N_46708);
nor U49113 (N_49113,N_47681,N_46196);
or U49114 (N_49114,N_47802,N_47563);
nor U49115 (N_49115,N_47193,N_46963);
nor U49116 (N_49116,N_47700,N_46527);
nand U49117 (N_49117,N_46468,N_47118);
nor U49118 (N_49118,N_47586,N_47607);
and U49119 (N_49119,N_46056,N_47048);
nor U49120 (N_49120,N_46395,N_47889);
and U49121 (N_49121,N_46055,N_46905);
and U49122 (N_49122,N_47939,N_46710);
nand U49123 (N_49123,N_46738,N_47024);
or U49124 (N_49124,N_46879,N_47481);
nor U49125 (N_49125,N_46869,N_47965);
and U49126 (N_49126,N_46238,N_47351);
and U49127 (N_49127,N_46792,N_47224);
or U49128 (N_49128,N_46144,N_47659);
nand U49129 (N_49129,N_47997,N_46716);
xor U49130 (N_49130,N_47275,N_47093);
or U49131 (N_49131,N_47844,N_46055);
and U49132 (N_49132,N_47542,N_46249);
or U49133 (N_49133,N_47624,N_46575);
nor U49134 (N_49134,N_46139,N_47161);
or U49135 (N_49135,N_47417,N_47783);
and U49136 (N_49136,N_47441,N_46454);
nor U49137 (N_49137,N_46904,N_46180);
and U49138 (N_49138,N_47629,N_46700);
and U49139 (N_49139,N_46433,N_47991);
nand U49140 (N_49140,N_46362,N_47645);
and U49141 (N_49141,N_46961,N_46665);
nor U49142 (N_49142,N_47052,N_47142);
nor U49143 (N_49143,N_46079,N_47959);
and U49144 (N_49144,N_46164,N_47935);
and U49145 (N_49145,N_47007,N_47328);
nor U49146 (N_49146,N_46447,N_47062);
and U49147 (N_49147,N_47019,N_47339);
nand U49148 (N_49148,N_46149,N_46565);
and U49149 (N_49149,N_47071,N_47405);
nor U49150 (N_49150,N_47698,N_46037);
and U49151 (N_49151,N_46243,N_46595);
and U49152 (N_49152,N_46401,N_47762);
nand U49153 (N_49153,N_47543,N_47265);
and U49154 (N_49154,N_47278,N_47546);
nand U49155 (N_49155,N_46687,N_46279);
nor U49156 (N_49156,N_46187,N_47467);
nand U49157 (N_49157,N_47719,N_47467);
and U49158 (N_49158,N_47584,N_46243);
nand U49159 (N_49159,N_46787,N_47468);
nand U49160 (N_49160,N_47088,N_46603);
or U49161 (N_49161,N_46297,N_46919);
nor U49162 (N_49162,N_46932,N_47886);
nand U49163 (N_49163,N_47854,N_47710);
nand U49164 (N_49164,N_47141,N_47566);
nor U49165 (N_49165,N_47069,N_46867);
and U49166 (N_49166,N_47892,N_47173);
nor U49167 (N_49167,N_47386,N_46818);
and U49168 (N_49168,N_47364,N_47506);
nand U49169 (N_49169,N_46495,N_46888);
nand U49170 (N_49170,N_46102,N_47665);
nand U49171 (N_49171,N_46207,N_47723);
nor U49172 (N_49172,N_46063,N_46449);
nor U49173 (N_49173,N_46156,N_46072);
and U49174 (N_49174,N_46190,N_47260);
or U49175 (N_49175,N_47340,N_47503);
nor U49176 (N_49176,N_46916,N_46094);
and U49177 (N_49177,N_46453,N_47163);
nor U49178 (N_49178,N_46361,N_46155);
nand U49179 (N_49179,N_46866,N_46847);
and U49180 (N_49180,N_47325,N_47669);
and U49181 (N_49181,N_47236,N_46524);
and U49182 (N_49182,N_47978,N_46341);
nor U49183 (N_49183,N_46123,N_47435);
and U49184 (N_49184,N_46035,N_46898);
nor U49185 (N_49185,N_47760,N_47547);
xor U49186 (N_49186,N_47644,N_47094);
nand U49187 (N_49187,N_46875,N_47050);
nand U49188 (N_49188,N_46696,N_46749);
nor U49189 (N_49189,N_46154,N_46423);
nor U49190 (N_49190,N_46828,N_46169);
nor U49191 (N_49191,N_47158,N_47465);
and U49192 (N_49192,N_46097,N_47356);
nor U49193 (N_49193,N_46868,N_46940);
nor U49194 (N_49194,N_46397,N_46958);
nor U49195 (N_49195,N_47268,N_47610);
and U49196 (N_49196,N_47463,N_46877);
nand U49197 (N_49197,N_46225,N_46895);
nand U49198 (N_49198,N_46666,N_47136);
nand U49199 (N_49199,N_47954,N_47697);
xor U49200 (N_49200,N_47677,N_46703);
nand U49201 (N_49201,N_46767,N_46908);
nor U49202 (N_49202,N_47998,N_46960);
and U49203 (N_49203,N_47711,N_46286);
and U49204 (N_49204,N_47683,N_47070);
nand U49205 (N_49205,N_47632,N_47101);
and U49206 (N_49206,N_47108,N_46760);
nand U49207 (N_49207,N_47118,N_46703);
nor U49208 (N_49208,N_46854,N_46384);
nor U49209 (N_49209,N_46617,N_46508);
nand U49210 (N_49210,N_47038,N_47868);
nand U49211 (N_49211,N_46458,N_47651);
nand U49212 (N_49212,N_46367,N_47980);
or U49213 (N_49213,N_47062,N_47833);
nand U49214 (N_49214,N_47077,N_46404);
nor U49215 (N_49215,N_46477,N_47125);
and U49216 (N_49216,N_46524,N_47032);
nand U49217 (N_49217,N_46609,N_46203);
or U49218 (N_49218,N_46517,N_47665);
nor U49219 (N_49219,N_46928,N_46295);
nor U49220 (N_49220,N_47783,N_47821);
nand U49221 (N_49221,N_46268,N_46671);
and U49222 (N_49222,N_46935,N_46864);
or U49223 (N_49223,N_46203,N_47570);
and U49224 (N_49224,N_47137,N_47836);
nand U49225 (N_49225,N_47794,N_46940);
and U49226 (N_49226,N_47134,N_46884);
and U49227 (N_49227,N_47733,N_47086);
or U49228 (N_49228,N_46582,N_47256);
and U49229 (N_49229,N_46914,N_46699);
or U49230 (N_49230,N_47267,N_47711);
nand U49231 (N_49231,N_47449,N_47927);
nand U49232 (N_49232,N_46680,N_46455);
and U49233 (N_49233,N_46236,N_46902);
and U49234 (N_49234,N_47538,N_46636);
nor U49235 (N_49235,N_46362,N_46189);
xnor U49236 (N_49236,N_46254,N_47351);
and U49237 (N_49237,N_46018,N_47212);
or U49238 (N_49238,N_47404,N_46966);
and U49239 (N_49239,N_47463,N_46543);
and U49240 (N_49240,N_46462,N_46414);
or U49241 (N_49241,N_46407,N_47761);
or U49242 (N_49242,N_46002,N_46679);
or U49243 (N_49243,N_46105,N_47123);
nand U49244 (N_49244,N_46241,N_47307);
nor U49245 (N_49245,N_47374,N_47387);
nor U49246 (N_49246,N_46447,N_47531);
and U49247 (N_49247,N_47758,N_46653);
or U49248 (N_49248,N_46802,N_46788);
nand U49249 (N_49249,N_47280,N_47010);
or U49250 (N_49250,N_46726,N_47318);
nand U49251 (N_49251,N_47198,N_47840);
and U49252 (N_49252,N_46895,N_47482);
and U49253 (N_49253,N_47698,N_47219);
nand U49254 (N_49254,N_46342,N_47155);
or U49255 (N_49255,N_47328,N_46084);
nor U49256 (N_49256,N_46692,N_46108);
nor U49257 (N_49257,N_47089,N_46744);
nand U49258 (N_49258,N_46655,N_47641);
nor U49259 (N_49259,N_46360,N_46681);
and U49260 (N_49260,N_47005,N_46811);
nor U49261 (N_49261,N_47088,N_46440);
and U49262 (N_49262,N_47148,N_46396);
or U49263 (N_49263,N_46993,N_46292);
nor U49264 (N_49264,N_47628,N_46120);
and U49265 (N_49265,N_46552,N_46138);
nand U49266 (N_49266,N_46548,N_46278);
or U49267 (N_49267,N_47797,N_47004);
and U49268 (N_49268,N_46660,N_47151);
and U49269 (N_49269,N_47170,N_46352);
nor U49270 (N_49270,N_46048,N_47058);
or U49271 (N_49271,N_46855,N_47897);
nand U49272 (N_49272,N_46984,N_47830);
xnor U49273 (N_49273,N_46321,N_46074);
or U49274 (N_49274,N_47451,N_46372);
nor U49275 (N_49275,N_46285,N_46319);
or U49276 (N_49276,N_46216,N_46609);
and U49277 (N_49277,N_46641,N_46903);
nor U49278 (N_49278,N_47111,N_46158);
and U49279 (N_49279,N_46603,N_47445);
nand U49280 (N_49280,N_46767,N_46885);
and U49281 (N_49281,N_46300,N_47846);
nand U49282 (N_49282,N_47582,N_46101);
nand U49283 (N_49283,N_47461,N_46377);
nand U49284 (N_49284,N_47425,N_46344);
nand U49285 (N_49285,N_47581,N_46829);
nor U49286 (N_49286,N_46049,N_47302);
and U49287 (N_49287,N_46495,N_47346);
and U49288 (N_49288,N_47498,N_46552);
and U49289 (N_49289,N_47991,N_47234);
nand U49290 (N_49290,N_47223,N_46966);
or U49291 (N_49291,N_47204,N_47028);
nor U49292 (N_49292,N_47864,N_46688);
nand U49293 (N_49293,N_46660,N_47901);
nand U49294 (N_49294,N_46393,N_46598);
nand U49295 (N_49295,N_47702,N_46298);
or U49296 (N_49296,N_46724,N_46706);
nor U49297 (N_49297,N_46652,N_46004);
nor U49298 (N_49298,N_46897,N_47056);
and U49299 (N_49299,N_46608,N_46256);
or U49300 (N_49300,N_46454,N_46104);
and U49301 (N_49301,N_47924,N_46356);
or U49302 (N_49302,N_46825,N_47764);
and U49303 (N_49303,N_46422,N_47181);
nor U49304 (N_49304,N_46839,N_46629);
and U49305 (N_49305,N_47571,N_46497);
nor U49306 (N_49306,N_47195,N_47070);
or U49307 (N_49307,N_47605,N_46319);
xor U49308 (N_49308,N_47630,N_47499);
and U49309 (N_49309,N_47588,N_47750);
or U49310 (N_49310,N_46221,N_46470);
xnor U49311 (N_49311,N_46304,N_46956);
nand U49312 (N_49312,N_46828,N_46031);
nor U49313 (N_49313,N_46428,N_47680);
nand U49314 (N_49314,N_46045,N_46921);
nor U49315 (N_49315,N_47192,N_47114);
nor U49316 (N_49316,N_47144,N_47242);
and U49317 (N_49317,N_46012,N_46703);
or U49318 (N_49318,N_47615,N_46146);
or U49319 (N_49319,N_46449,N_46686);
or U49320 (N_49320,N_46920,N_47780);
nand U49321 (N_49321,N_47834,N_46603);
nor U49322 (N_49322,N_47608,N_47544);
nand U49323 (N_49323,N_46932,N_47290);
nor U49324 (N_49324,N_47666,N_47136);
or U49325 (N_49325,N_46794,N_47952);
or U49326 (N_49326,N_47258,N_46931);
and U49327 (N_49327,N_47672,N_46126);
or U49328 (N_49328,N_46352,N_47374);
nand U49329 (N_49329,N_47539,N_46511);
or U49330 (N_49330,N_47286,N_47477);
nand U49331 (N_49331,N_46544,N_47598);
or U49332 (N_49332,N_47303,N_47885);
nor U49333 (N_49333,N_47720,N_46203);
or U49334 (N_49334,N_47741,N_46372);
and U49335 (N_49335,N_47261,N_46383);
xnor U49336 (N_49336,N_47789,N_47818);
nand U49337 (N_49337,N_46865,N_47519);
or U49338 (N_49338,N_47704,N_46829);
or U49339 (N_49339,N_47776,N_46590);
xor U49340 (N_49340,N_47266,N_47329);
or U49341 (N_49341,N_46937,N_46179);
xor U49342 (N_49342,N_47991,N_47811);
and U49343 (N_49343,N_46610,N_46067);
xnor U49344 (N_49344,N_46349,N_46643);
nor U49345 (N_49345,N_47658,N_47910);
nor U49346 (N_49346,N_46830,N_47963);
and U49347 (N_49347,N_47943,N_46753);
nand U49348 (N_49348,N_47592,N_46022);
or U49349 (N_49349,N_46787,N_47912);
nand U49350 (N_49350,N_46177,N_47071);
and U49351 (N_49351,N_47990,N_46712);
nand U49352 (N_49352,N_46004,N_47475);
and U49353 (N_49353,N_46954,N_46891);
nor U49354 (N_49354,N_47798,N_47637);
nor U49355 (N_49355,N_46368,N_47424);
or U49356 (N_49356,N_47202,N_47018);
nor U49357 (N_49357,N_47873,N_47916);
or U49358 (N_49358,N_46737,N_47582);
and U49359 (N_49359,N_47184,N_47969);
nand U49360 (N_49360,N_46415,N_46082);
and U49361 (N_49361,N_47404,N_46819);
nor U49362 (N_49362,N_46891,N_46787);
nand U49363 (N_49363,N_47137,N_47896);
and U49364 (N_49364,N_46758,N_46790);
nand U49365 (N_49365,N_47694,N_47893);
nand U49366 (N_49366,N_46099,N_46057);
and U49367 (N_49367,N_46568,N_46794);
and U49368 (N_49368,N_47349,N_46658);
nand U49369 (N_49369,N_47120,N_47272);
nand U49370 (N_49370,N_46300,N_46793);
nor U49371 (N_49371,N_47579,N_47183);
nand U49372 (N_49372,N_46659,N_46479);
nand U49373 (N_49373,N_47580,N_47739);
nor U49374 (N_49374,N_46853,N_46807);
nand U49375 (N_49375,N_46043,N_47205);
nor U49376 (N_49376,N_46676,N_47576);
or U49377 (N_49377,N_47087,N_47426);
nor U49378 (N_49378,N_47191,N_46115);
and U49379 (N_49379,N_47616,N_46206);
nor U49380 (N_49380,N_47017,N_46164);
and U49381 (N_49381,N_46318,N_46243);
nand U49382 (N_49382,N_47658,N_47896);
or U49383 (N_49383,N_46562,N_47958);
nand U49384 (N_49384,N_46490,N_46165);
nor U49385 (N_49385,N_46618,N_46440);
nor U49386 (N_49386,N_46781,N_46844);
and U49387 (N_49387,N_46768,N_47247);
nor U49388 (N_49388,N_47779,N_46444);
nor U49389 (N_49389,N_46544,N_47670);
nor U49390 (N_49390,N_47135,N_46634);
and U49391 (N_49391,N_47649,N_47614);
nor U49392 (N_49392,N_47200,N_47770);
nor U49393 (N_49393,N_46417,N_47743);
nor U49394 (N_49394,N_46438,N_47362);
or U49395 (N_49395,N_47348,N_47067);
xnor U49396 (N_49396,N_46829,N_47637);
or U49397 (N_49397,N_47496,N_46085);
nor U49398 (N_49398,N_46413,N_46880);
nor U49399 (N_49399,N_46126,N_46489);
or U49400 (N_49400,N_47971,N_47256);
and U49401 (N_49401,N_46875,N_47638);
or U49402 (N_49402,N_46430,N_47966);
and U49403 (N_49403,N_47879,N_46523);
nand U49404 (N_49404,N_46649,N_46024);
nor U49405 (N_49405,N_47611,N_46038);
xnor U49406 (N_49406,N_47517,N_47713);
and U49407 (N_49407,N_46483,N_46479);
or U49408 (N_49408,N_46279,N_46885);
or U49409 (N_49409,N_46268,N_47283);
or U49410 (N_49410,N_47335,N_47560);
xnor U49411 (N_49411,N_47671,N_46307);
nand U49412 (N_49412,N_46847,N_46528);
nand U49413 (N_49413,N_46296,N_46094);
and U49414 (N_49414,N_47839,N_47821);
nor U49415 (N_49415,N_46605,N_47265);
nor U49416 (N_49416,N_47346,N_47808);
nor U49417 (N_49417,N_46760,N_47976);
and U49418 (N_49418,N_47460,N_46371);
nor U49419 (N_49419,N_46373,N_46875);
and U49420 (N_49420,N_47986,N_47267);
nand U49421 (N_49421,N_46817,N_47864);
and U49422 (N_49422,N_47026,N_47201);
or U49423 (N_49423,N_47543,N_46274);
nor U49424 (N_49424,N_46703,N_46736);
nand U49425 (N_49425,N_46760,N_46166);
nand U49426 (N_49426,N_46194,N_46506);
and U49427 (N_49427,N_46784,N_46653);
and U49428 (N_49428,N_47434,N_46685);
nor U49429 (N_49429,N_46231,N_46095);
nor U49430 (N_49430,N_46016,N_47951);
nor U49431 (N_49431,N_46789,N_46117);
nand U49432 (N_49432,N_46693,N_47470);
nand U49433 (N_49433,N_47751,N_47840);
or U49434 (N_49434,N_47777,N_47625);
or U49435 (N_49435,N_46729,N_46071);
and U49436 (N_49436,N_46740,N_47177);
or U49437 (N_49437,N_47551,N_46858);
nand U49438 (N_49438,N_46105,N_46205);
and U49439 (N_49439,N_46407,N_47528);
or U49440 (N_49440,N_46931,N_47591);
or U49441 (N_49441,N_46351,N_46430);
xor U49442 (N_49442,N_46468,N_46912);
nand U49443 (N_49443,N_47406,N_47274);
nor U49444 (N_49444,N_47436,N_46683);
nand U49445 (N_49445,N_46396,N_47278);
or U49446 (N_49446,N_47211,N_47678);
and U49447 (N_49447,N_46645,N_46317);
and U49448 (N_49448,N_47475,N_47444);
xnor U49449 (N_49449,N_46122,N_47451);
and U49450 (N_49450,N_46505,N_46193);
or U49451 (N_49451,N_46565,N_46423);
or U49452 (N_49452,N_47870,N_47658);
or U49453 (N_49453,N_47666,N_46255);
nor U49454 (N_49454,N_47261,N_47058);
nor U49455 (N_49455,N_47152,N_46114);
nand U49456 (N_49456,N_47505,N_46230);
nor U49457 (N_49457,N_47549,N_46441);
and U49458 (N_49458,N_47134,N_46047);
or U49459 (N_49459,N_47062,N_46594);
xnor U49460 (N_49460,N_46893,N_47310);
or U49461 (N_49461,N_47990,N_47875);
nor U49462 (N_49462,N_47737,N_46997);
nand U49463 (N_49463,N_46056,N_46396);
or U49464 (N_49464,N_47559,N_46171);
xor U49465 (N_49465,N_47994,N_46903);
or U49466 (N_49466,N_46436,N_46096);
nand U49467 (N_49467,N_46397,N_46589);
nor U49468 (N_49468,N_47755,N_46533);
nor U49469 (N_49469,N_46256,N_46845);
and U49470 (N_49470,N_47818,N_46437);
or U49471 (N_49471,N_46026,N_46549);
and U49472 (N_49472,N_47251,N_46096);
or U49473 (N_49473,N_47789,N_46885);
nor U49474 (N_49474,N_47672,N_47933);
and U49475 (N_49475,N_47912,N_47671);
and U49476 (N_49476,N_46272,N_47704);
nor U49477 (N_49477,N_46603,N_47506);
nor U49478 (N_49478,N_46638,N_46359);
nor U49479 (N_49479,N_47483,N_46971);
nor U49480 (N_49480,N_46990,N_47183);
nor U49481 (N_49481,N_47501,N_46761);
and U49482 (N_49482,N_47257,N_46679);
and U49483 (N_49483,N_46748,N_46349);
nand U49484 (N_49484,N_47461,N_47477);
and U49485 (N_49485,N_47831,N_46558);
nand U49486 (N_49486,N_46273,N_47803);
and U49487 (N_49487,N_47134,N_47211);
and U49488 (N_49488,N_46498,N_47192);
nor U49489 (N_49489,N_46140,N_46572);
or U49490 (N_49490,N_47599,N_47166);
nor U49491 (N_49491,N_46906,N_47773);
nand U49492 (N_49492,N_47741,N_47895);
nand U49493 (N_49493,N_46377,N_47806);
and U49494 (N_49494,N_47706,N_47013);
nand U49495 (N_49495,N_46808,N_47688);
and U49496 (N_49496,N_47751,N_46151);
nand U49497 (N_49497,N_47601,N_47826);
nor U49498 (N_49498,N_46981,N_47726);
nand U49499 (N_49499,N_46011,N_46116);
nor U49500 (N_49500,N_47390,N_47167);
and U49501 (N_49501,N_46565,N_46380);
nor U49502 (N_49502,N_46315,N_47535);
or U49503 (N_49503,N_46486,N_46498);
and U49504 (N_49504,N_46897,N_46431);
nand U49505 (N_49505,N_47053,N_46808);
and U49506 (N_49506,N_46250,N_46746);
or U49507 (N_49507,N_47474,N_47937);
or U49508 (N_49508,N_46149,N_47220);
nand U49509 (N_49509,N_47623,N_47664);
and U49510 (N_49510,N_46960,N_47690);
nand U49511 (N_49511,N_46044,N_47003);
nor U49512 (N_49512,N_47260,N_47062);
nand U49513 (N_49513,N_47999,N_47249);
or U49514 (N_49514,N_47693,N_46093);
and U49515 (N_49515,N_46879,N_47424);
and U49516 (N_49516,N_47189,N_47275);
or U49517 (N_49517,N_47540,N_46160);
nand U49518 (N_49518,N_47595,N_47715);
and U49519 (N_49519,N_47237,N_47528);
or U49520 (N_49520,N_46548,N_46952);
or U49521 (N_49521,N_46580,N_47204);
or U49522 (N_49522,N_46674,N_46735);
nand U49523 (N_49523,N_46103,N_46892);
and U49524 (N_49524,N_47576,N_47604);
nand U49525 (N_49525,N_47833,N_47849);
or U49526 (N_49526,N_46114,N_46159);
and U49527 (N_49527,N_47592,N_47101);
and U49528 (N_49528,N_46436,N_47123);
and U49529 (N_49529,N_46704,N_47477);
nand U49530 (N_49530,N_47267,N_47675);
nand U49531 (N_49531,N_46018,N_46637);
or U49532 (N_49532,N_47784,N_46281);
and U49533 (N_49533,N_46958,N_46532);
nor U49534 (N_49534,N_46872,N_47888);
and U49535 (N_49535,N_47440,N_46709);
or U49536 (N_49536,N_47610,N_47515);
or U49537 (N_49537,N_46790,N_47040);
xnor U49538 (N_49538,N_47263,N_46071);
nand U49539 (N_49539,N_46219,N_46584);
and U49540 (N_49540,N_47448,N_46801);
and U49541 (N_49541,N_46954,N_46636);
nor U49542 (N_49542,N_47763,N_47334);
or U49543 (N_49543,N_47167,N_47591);
or U49544 (N_49544,N_46092,N_47427);
xnor U49545 (N_49545,N_46724,N_47269);
and U49546 (N_49546,N_46224,N_46455);
and U49547 (N_49547,N_47741,N_47667);
nand U49548 (N_49548,N_46900,N_46079);
or U49549 (N_49549,N_46302,N_46890);
and U49550 (N_49550,N_46426,N_46332);
nand U49551 (N_49551,N_47350,N_47257);
nor U49552 (N_49552,N_46776,N_46305);
nand U49553 (N_49553,N_46413,N_46942);
or U49554 (N_49554,N_47363,N_46220);
or U49555 (N_49555,N_46031,N_46415);
nor U49556 (N_49556,N_46278,N_46894);
and U49557 (N_49557,N_47686,N_47918);
nand U49558 (N_49558,N_47495,N_47263);
nand U49559 (N_49559,N_47994,N_46684);
nand U49560 (N_49560,N_47897,N_47497);
and U49561 (N_49561,N_46141,N_46258);
nand U49562 (N_49562,N_46029,N_47835);
or U49563 (N_49563,N_47488,N_46019);
nand U49564 (N_49564,N_47356,N_46077);
nand U49565 (N_49565,N_46796,N_47698);
nor U49566 (N_49566,N_46066,N_47023);
nor U49567 (N_49567,N_47369,N_46486);
or U49568 (N_49568,N_47221,N_46300);
nand U49569 (N_49569,N_46725,N_46983);
or U49570 (N_49570,N_47006,N_47618);
or U49571 (N_49571,N_47503,N_47123);
nand U49572 (N_49572,N_46698,N_46693);
nor U49573 (N_49573,N_47211,N_46801);
and U49574 (N_49574,N_47540,N_47803);
and U49575 (N_49575,N_47100,N_47620);
or U49576 (N_49576,N_47349,N_47218);
nand U49577 (N_49577,N_47709,N_46721);
nand U49578 (N_49578,N_46254,N_46582);
nor U49579 (N_49579,N_47385,N_47321);
and U49580 (N_49580,N_47200,N_46846);
nor U49581 (N_49581,N_47442,N_46897);
and U49582 (N_49582,N_47753,N_47785);
nand U49583 (N_49583,N_46591,N_47304);
nand U49584 (N_49584,N_46088,N_47138);
or U49585 (N_49585,N_46735,N_47903);
and U49586 (N_49586,N_47262,N_46677);
and U49587 (N_49587,N_46227,N_47412);
xnor U49588 (N_49588,N_47693,N_46025);
nand U49589 (N_49589,N_47054,N_46983);
nand U49590 (N_49590,N_47740,N_46732);
or U49591 (N_49591,N_47745,N_46120);
nand U49592 (N_49592,N_47225,N_46511);
nand U49593 (N_49593,N_47796,N_47284);
nand U49594 (N_49594,N_47503,N_46754);
or U49595 (N_49595,N_46717,N_46359);
and U49596 (N_49596,N_47374,N_46645);
or U49597 (N_49597,N_47640,N_46817);
or U49598 (N_49598,N_47903,N_47555);
nand U49599 (N_49599,N_46109,N_47707);
nor U49600 (N_49600,N_46406,N_46595);
and U49601 (N_49601,N_46293,N_47102);
nor U49602 (N_49602,N_47021,N_47341);
nand U49603 (N_49603,N_46429,N_46256);
nor U49604 (N_49604,N_47669,N_47190);
nor U49605 (N_49605,N_47516,N_47780);
or U49606 (N_49606,N_47019,N_46169);
or U49607 (N_49607,N_46294,N_47804);
nand U49608 (N_49608,N_46844,N_47766);
nand U49609 (N_49609,N_47826,N_47204);
or U49610 (N_49610,N_47858,N_46830);
or U49611 (N_49611,N_47708,N_46913);
nand U49612 (N_49612,N_46363,N_46377);
nor U49613 (N_49613,N_47556,N_46528);
nor U49614 (N_49614,N_46546,N_46719);
or U49615 (N_49615,N_47523,N_46328);
or U49616 (N_49616,N_47394,N_46485);
nand U49617 (N_49617,N_46221,N_46492);
and U49618 (N_49618,N_46584,N_47888);
nor U49619 (N_49619,N_47198,N_47233);
nand U49620 (N_49620,N_47115,N_47043);
and U49621 (N_49621,N_47591,N_47297);
and U49622 (N_49622,N_47328,N_47024);
nand U49623 (N_49623,N_47483,N_46675);
or U49624 (N_49624,N_47216,N_46232);
nor U49625 (N_49625,N_46951,N_46644);
and U49626 (N_49626,N_46748,N_46246);
nand U49627 (N_49627,N_47968,N_47798);
nor U49628 (N_49628,N_46216,N_46890);
nand U49629 (N_49629,N_47062,N_47678);
and U49630 (N_49630,N_46311,N_47530);
or U49631 (N_49631,N_46814,N_47760);
or U49632 (N_49632,N_46030,N_46513);
and U49633 (N_49633,N_46638,N_46192);
and U49634 (N_49634,N_46122,N_46805);
or U49635 (N_49635,N_46437,N_46712);
or U49636 (N_49636,N_47821,N_47280);
and U49637 (N_49637,N_47232,N_47463);
and U49638 (N_49638,N_46845,N_46989);
nand U49639 (N_49639,N_47108,N_47106);
nand U49640 (N_49640,N_47792,N_47921);
or U49641 (N_49641,N_46293,N_47272);
or U49642 (N_49642,N_46499,N_46955);
nand U49643 (N_49643,N_47741,N_46143);
nand U49644 (N_49644,N_47726,N_46334);
or U49645 (N_49645,N_47308,N_47591);
nor U49646 (N_49646,N_46940,N_47618);
or U49647 (N_49647,N_46762,N_47006);
nor U49648 (N_49648,N_47884,N_47718);
nand U49649 (N_49649,N_47101,N_46545);
nor U49650 (N_49650,N_47439,N_46973);
and U49651 (N_49651,N_47561,N_47258);
nor U49652 (N_49652,N_46071,N_46935);
or U49653 (N_49653,N_46828,N_46344);
nand U49654 (N_49654,N_47080,N_46197);
or U49655 (N_49655,N_47717,N_46281);
nor U49656 (N_49656,N_46639,N_46492);
or U49657 (N_49657,N_47848,N_46480);
nand U49658 (N_49658,N_47648,N_47664);
nor U49659 (N_49659,N_47414,N_47405);
or U49660 (N_49660,N_46016,N_47850);
nor U49661 (N_49661,N_47995,N_47828);
and U49662 (N_49662,N_46077,N_47371);
and U49663 (N_49663,N_47531,N_47803);
nor U49664 (N_49664,N_46306,N_46190);
and U49665 (N_49665,N_47087,N_47771);
and U49666 (N_49666,N_46916,N_46667);
or U49667 (N_49667,N_46546,N_47313);
nand U49668 (N_49668,N_46681,N_46172);
nand U49669 (N_49669,N_47620,N_47897);
or U49670 (N_49670,N_46553,N_46045);
nor U49671 (N_49671,N_47711,N_47410);
or U49672 (N_49672,N_46217,N_47025);
and U49673 (N_49673,N_46656,N_46965);
or U49674 (N_49674,N_46530,N_46559);
and U49675 (N_49675,N_46120,N_47013);
nor U49676 (N_49676,N_46085,N_47539);
and U49677 (N_49677,N_47068,N_46248);
nor U49678 (N_49678,N_47566,N_46594);
nand U49679 (N_49679,N_46942,N_47759);
nor U49680 (N_49680,N_46854,N_46569);
or U49681 (N_49681,N_47270,N_46952);
nor U49682 (N_49682,N_47758,N_47407);
nor U49683 (N_49683,N_47930,N_47781);
nand U49684 (N_49684,N_47719,N_47689);
nor U49685 (N_49685,N_47463,N_47787);
and U49686 (N_49686,N_47722,N_47307);
nor U49687 (N_49687,N_47872,N_46496);
xnor U49688 (N_49688,N_47855,N_47040);
and U49689 (N_49689,N_47232,N_47440);
and U49690 (N_49690,N_47904,N_47985);
nand U49691 (N_49691,N_47622,N_47799);
nand U49692 (N_49692,N_47701,N_46752);
nand U49693 (N_49693,N_47288,N_46090);
nor U49694 (N_49694,N_46155,N_47044);
or U49695 (N_49695,N_47149,N_47561);
nand U49696 (N_49696,N_47237,N_46255);
and U49697 (N_49697,N_46463,N_46769);
nor U49698 (N_49698,N_46584,N_47592);
nand U49699 (N_49699,N_47661,N_46500);
nand U49700 (N_49700,N_46878,N_46956);
and U49701 (N_49701,N_46376,N_46614);
or U49702 (N_49702,N_46842,N_46537);
and U49703 (N_49703,N_46232,N_46238);
nor U49704 (N_49704,N_46630,N_47406);
and U49705 (N_49705,N_46347,N_47252);
nand U49706 (N_49706,N_47828,N_46908);
nand U49707 (N_49707,N_46883,N_46652);
nand U49708 (N_49708,N_46216,N_47014);
and U49709 (N_49709,N_47200,N_46894);
nor U49710 (N_49710,N_46814,N_47799);
and U49711 (N_49711,N_46975,N_46141);
or U49712 (N_49712,N_46824,N_47810);
xnor U49713 (N_49713,N_47877,N_46511);
nand U49714 (N_49714,N_47524,N_47164);
or U49715 (N_49715,N_47156,N_47019);
or U49716 (N_49716,N_46058,N_47080);
nand U49717 (N_49717,N_46096,N_46100);
nand U49718 (N_49718,N_47635,N_47640);
and U49719 (N_49719,N_47377,N_47915);
or U49720 (N_49720,N_47280,N_46031);
and U49721 (N_49721,N_47045,N_47961);
and U49722 (N_49722,N_47923,N_47560);
nor U49723 (N_49723,N_47563,N_47400);
nor U49724 (N_49724,N_46839,N_47325);
nand U49725 (N_49725,N_47990,N_47867);
or U49726 (N_49726,N_47421,N_46624);
and U49727 (N_49727,N_47846,N_46458);
nand U49728 (N_49728,N_47653,N_47431);
nand U49729 (N_49729,N_47721,N_47058);
and U49730 (N_49730,N_46980,N_47301);
or U49731 (N_49731,N_47313,N_46881);
nand U49732 (N_49732,N_46759,N_47795);
and U49733 (N_49733,N_46827,N_47106);
and U49734 (N_49734,N_46478,N_46929);
and U49735 (N_49735,N_47073,N_47926);
or U49736 (N_49736,N_46735,N_47016);
and U49737 (N_49737,N_47248,N_47659);
or U49738 (N_49738,N_47624,N_46342);
or U49739 (N_49739,N_47995,N_46824);
nand U49740 (N_49740,N_46734,N_46419);
or U49741 (N_49741,N_47302,N_46838);
and U49742 (N_49742,N_46418,N_47463);
nand U49743 (N_49743,N_46744,N_46486);
and U49744 (N_49744,N_46323,N_46766);
nand U49745 (N_49745,N_46124,N_46309);
nor U49746 (N_49746,N_46971,N_46591);
or U49747 (N_49747,N_47546,N_46197);
and U49748 (N_49748,N_46562,N_47088);
nor U49749 (N_49749,N_47249,N_46268);
or U49750 (N_49750,N_47918,N_47891);
nand U49751 (N_49751,N_47854,N_47642);
nor U49752 (N_49752,N_46584,N_46785);
and U49753 (N_49753,N_47900,N_47345);
nand U49754 (N_49754,N_46058,N_47453);
nand U49755 (N_49755,N_46756,N_46584);
or U49756 (N_49756,N_46981,N_47133);
nand U49757 (N_49757,N_46628,N_47612);
or U49758 (N_49758,N_46571,N_46265);
nor U49759 (N_49759,N_46327,N_47210);
nand U49760 (N_49760,N_46055,N_46929);
nand U49761 (N_49761,N_46899,N_46157);
nand U49762 (N_49762,N_47065,N_46997);
and U49763 (N_49763,N_46169,N_46893);
nand U49764 (N_49764,N_47977,N_47919);
nand U49765 (N_49765,N_46299,N_47828);
nor U49766 (N_49766,N_47793,N_47025);
nor U49767 (N_49767,N_47264,N_47663);
nand U49768 (N_49768,N_46379,N_46569);
nand U49769 (N_49769,N_47599,N_47996);
nor U49770 (N_49770,N_46046,N_47485);
nand U49771 (N_49771,N_46099,N_47129);
nor U49772 (N_49772,N_46828,N_46640);
and U49773 (N_49773,N_46818,N_46397);
and U49774 (N_49774,N_46080,N_46979);
and U49775 (N_49775,N_46449,N_46920);
and U49776 (N_49776,N_46444,N_46431);
nand U49777 (N_49777,N_47858,N_47047);
nand U49778 (N_49778,N_47209,N_46731);
nand U49779 (N_49779,N_47964,N_47109);
and U49780 (N_49780,N_47946,N_47037);
nor U49781 (N_49781,N_47325,N_46708);
nand U49782 (N_49782,N_46373,N_47983);
or U49783 (N_49783,N_47070,N_46482);
or U49784 (N_49784,N_47985,N_47774);
xnor U49785 (N_49785,N_46993,N_47722);
or U49786 (N_49786,N_46177,N_46722);
or U49787 (N_49787,N_47667,N_46051);
nand U49788 (N_49788,N_46167,N_46471);
or U49789 (N_49789,N_47090,N_47099);
nor U49790 (N_49790,N_46554,N_46072);
and U49791 (N_49791,N_47553,N_46290);
and U49792 (N_49792,N_47612,N_47914);
nand U49793 (N_49793,N_47769,N_46076);
nand U49794 (N_49794,N_47367,N_46279);
nand U49795 (N_49795,N_47150,N_47223);
nor U49796 (N_49796,N_46660,N_47998);
and U49797 (N_49797,N_47212,N_47630);
nand U49798 (N_49798,N_46954,N_47574);
or U49799 (N_49799,N_46393,N_46057);
and U49800 (N_49800,N_47246,N_46927);
and U49801 (N_49801,N_46123,N_47795);
nor U49802 (N_49802,N_46147,N_46469);
and U49803 (N_49803,N_46676,N_47267);
and U49804 (N_49804,N_46878,N_47259);
or U49805 (N_49805,N_47848,N_46352);
xor U49806 (N_49806,N_47656,N_47495);
nor U49807 (N_49807,N_47618,N_47064);
nand U49808 (N_49808,N_46756,N_47233);
nand U49809 (N_49809,N_47207,N_47218);
nor U49810 (N_49810,N_46535,N_46116);
and U49811 (N_49811,N_47971,N_46100);
and U49812 (N_49812,N_46363,N_46078);
xor U49813 (N_49813,N_46964,N_47269);
nand U49814 (N_49814,N_46865,N_47309);
nand U49815 (N_49815,N_46937,N_47380);
and U49816 (N_49816,N_47439,N_46658);
nand U49817 (N_49817,N_47139,N_46484);
or U49818 (N_49818,N_46339,N_47945);
nor U49819 (N_49819,N_46278,N_47256);
or U49820 (N_49820,N_46570,N_47886);
xor U49821 (N_49821,N_46205,N_47708);
nor U49822 (N_49822,N_46799,N_47780);
and U49823 (N_49823,N_47797,N_46099);
nor U49824 (N_49824,N_47311,N_46128);
or U49825 (N_49825,N_46925,N_46879);
and U49826 (N_49826,N_47048,N_47892);
and U49827 (N_49827,N_46297,N_46301);
or U49828 (N_49828,N_46538,N_47206);
and U49829 (N_49829,N_46683,N_47478);
or U49830 (N_49830,N_47950,N_46520);
nor U49831 (N_49831,N_47018,N_47790);
and U49832 (N_49832,N_47162,N_47275);
and U49833 (N_49833,N_46747,N_46137);
and U49834 (N_49834,N_46939,N_47866);
nor U49835 (N_49835,N_47150,N_46283);
or U49836 (N_49836,N_46346,N_46312);
xnor U49837 (N_49837,N_47254,N_46852);
and U49838 (N_49838,N_47131,N_47863);
or U49839 (N_49839,N_47306,N_47403);
and U49840 (N_49840,N_47739,N_46642);
xnor U49841 (N_49841,N_46662,N_47633);
and U49842 (N_49842,N_47326,N_46253);
xnor U49843 (N_49843,N_46629,N_47216);
nand U49844 (N_49844,N_46359,N_47824);
nor U49845 (N_49845,N_47080,N_47316);
xnor U49846 (N_49846,N_46523,N_47153);
or U49847 (N_49847,N_46490,N_47725);
nand U49848 (N_49848,N_47072,N_46757);
nand U49849 (N_49849,N_46776,N_46286);
and U49850 (N_49850,N_47887,N_46321);
and U49851 (N_49851,N_46204,N_47289);
nor U49852 (N_49852,N_47353,N_46919);
nand U49853 (N_49853,N_47096,N_47326);
nor U49854 (N_49854,N_46119,N_46456);
nand U49855 (N_49855,N_47014,N_47838);
or U49856 (N_49856,N_47441,N_47382);
nand U49857 (N_49857,N_47796,N_46219);
nand U49858 (N_49858,N_47087,N_46992);
or U49859 (N_49859,N_47398,N_46810);
nand U49860 (N_49860,N_47379,N_46563);
nor U49861 (N_49861,N_46728,N_46410);
nand U49862 (N_49862,N_46506,N_46158);
xnor U49863 (N_49863,N_47353,N_46255);
nand U49864 (N_49864,N_47068,N_47454);
and U49865 (N_49865,N_47013,N_47752);
nand U49866 (N_49866,N_46528,N_47298);
nand U49867 (N_49867,N_47524,N_46439);
and U49868 (N_49868,N_46747,N_46455);
and U49869 (N_49869,N_47559,N_47105);
or U49870 (N_49870,N_46384,N_46865);
nand U49871 (N_49871,N_47639,N_47409);
and U49872 (N_49872,N_46887,N_46647);
nand U49873 (N_49873,N_47205,N_47512);
and U49874 (N_49874,N_46968,N_47493);
nor U49875 (N_49875,N_46509,N_46821);
nand U49876 (N_49876,N_47995,N_46109);
nor U49877 (N_49877,N_47390,N_47063);
or U49878 (N_49878,N_47192,N_46203);
nand U49879 (N_49879,N_46654,N_46546);
or U49880 (N_49880,N_47780,N_47365);
and U49881 (N_49881,N_46234,N_46144);
or U49882 (N_49882,N_47095,N_47157);
nand U49883 (N_49883,N_46826,N_46754);
and U49884 (N_49884,N_47450,N_46167);
nand U49885 (N_49885,N_47051,N_47868);
nand U49886 (N_49886,N_47361,N_46846);
and U49887 (N_49887,N_47186,N_47128);
and U49888 (N_49888,N_46331,N_46178);
or U49889 (N_49889,N_47751,N_46033);
nor U49890 (N_49890,N_46689,N_46112);
or U49891 (N_49891,N_47609,N_46078);
and U49892 (N_49892,N_47638,N_47889);
or U49893 (N_49893,N_47312,N_47518);
and U49894 (N_49894,N_47996,N_47790);
nand U49895 (N_49895,N_47996,N_46767);
and U49896 (N_49896,N_47710,N_47396);
nor U49897 (N_49897,N_46092,N_46658);
nor U49898 (N_49898,N_47938,N_47175);
nand U49899 (N_49899,N_47570,N_46788);
and U49900 (N_49900,N_47301,N_46303);
and U49901 (N_49901,N_47867,N_47795);
nand U49902 (N_49902,N_46040,N_47131);
and U49903 (N_49903,N_47124,N_46258);
nand U49904 (N_49904,N_46215,N_47582);
and U49905 (N_49905,N_47616,N_47851);
nor U49906 (N_49906,N_46330,N_46056);
or U49907 (N_49907,N_46770,N_46219);
or U49908 (N_49908,N_46184,N_46086);
nor U49909 (N_49909,N_46612,N_47498);
and U49910 (N_49910,N_47142,N_46083);
and U49911 (N_49911,N_47082,N_46805);
or U49912 (N_49912,N_47023,N_47555);
nand U49913 (N_49913,N_46711,N_46332);
nor U49914 (N_49914,N_47064,N_46762);
nor U49915 (N_49915,N_47908,N_46745);
and U49916 (N_49916,N_46977,N_47137);
nand U49917 (N_49917,N_47988,N_47631);
and U49918 (N_49918,N_46666,N_46273);
nand U49919 (N_49919,N_46725,N_47985);
or U49920 (N_49920,N_46832,N_46107);
nand U49921 (N_49921,N_46023,N_47545);
nand U49922 (N_49922,N_47514,N_46755);
or U49923 (N_49923,N_47912,N_46488);
nand U49924 (N_49924,N_46341,N_47677);
and U49925 (N_49925,N_47133,N_46946);
and U49926 (N_49926,N_46888,N_47760);
nand U49927 (N_49927,N_47228,N_46040);
nand U49928 (N_49928,N_47467,N_46682);
nor U49929 (N_49929,N_47095,N_46688);
xnor U49930 (N_49930,N_46172,N_47687);
or U49931 (N_49931,N_46659,N_47494);
and U49932 (N_49932,N_47043,N_47129);
nand U49933 (N_49933,N_46841,N_46935);
nand U49934 (N_49934,N_47941,N_47601);
and U49935 (N_49935,N_46698,N_47724);
nor U49936 (N_49936,N_47944,N_46473);
and U49937 (N_49937,N_47017,N_47316);
nand U49938 (N_49938,N_47710,N_46813);
nand U49939 (N_49939,N_47549,N_46977);
or U49940 (N_49940,N_46940,N_47248);
or U49941 (N_49941,N_47353,N_46602);
and U49942 (N_49942,N_46640,N_46309);
nand U49943 (N_49943,N_46234,N_47960);
or U49944 (N_49944,N_46003,N_46944);
nor U49945 (N_49945,N_47028,N_47946);
nor U49946 (N_49946,N_47773,N_47152);
or U49947 (N_49947,N_46195,N_47418);
nor U49948 (N_49948,N_47730,N_47760);
xor U49949 (N_49949,N_46954,N_46844);
nor U49950 (N_49950,N_47858,N_47127);
nand U49951 (N_49951,N_46953,N_46535);
nor U49952 (N_49952,N_47968,N_46511);
nor U49953 (N_49953,N_47700,N_47464);
or U49954 (N_49954,N_47330,N_46614);
nor U49955 (N_49955,N_47957,N_46599);
and U49956 (N_49956,N_46164,N_47314);
and U49957 (N_49957,N_47102,N_47223);
and U49958 (N_49958,N_46961,N_46409);
nor U49959 (N_49959,N_47742,N_47117);
nand U49960 (N_49960,N_47517,N_47096);
nand U49961 (N_49961,N_46165,N_46750);
nand U49962 (N_49962,N_47697,N_46383);
nand U49963 (N_49963,N_47822,N_47397);
nand U49964 (N_49964,N_47939,N_47059);
nor U49965 (N_49965,N_47116,N_47633);
or U49966 (N_49966,N_46368,N_47524);
or U49967 (N_49967,N_47402,N_46971);
nand U49968 (N_49968,N_47659,N_47510);
or U49969 (N_49969,N_47642,N_46158);
nand U49970 (N_49970,N_47941,N_46216);
or U49971 (N_49971,N_46544,N_46285);
and U49972 (N_49972,N_46670,N_46938);
nand U49973 (N_49973,N_46590,N_46632);
nor U49974 (N_49974,N_46687,N_46763);
nor U49975 (N_49975,N_46344,N_46245);
and U49976 (N_49976,N_46288,N_47392);
or U49977 (N_49977,N_46950,N_47503);
and U49978 (N_49978,N_46142,N_47328);
nand U49979 (N_49979,N_47539,N_47782);
nor U49980 (N_49980,N_47469,N_46801);
nor U49981 (N_49981,N_47229,N_47753);
and U49982 (N_49982,N_46316,N_46833);
nor U49983 (N_49983,N_47114,N_47436);
or U49984 (N_49984,N_46078,N_47608);
or U49985 (N_49985,N_46822,N_47995);
and U49986 (N_49986,N_46182,N_46184);
and U49987 (N_49987,N_47786,N_46644);
xor U49988 (N_49988,N_47567,N_46659);
nor U49989 (N_49989,N_47573,N_46948);
and U49990 (N_49990,N_46044,N_46791);
xor U49991 (N_49991,N_47970,N_47821);
and U49992 (N_49992,N_47430,N_47343);
nor U49993 (N_49993,N_47334,N_47567);
and U49994 (N_49994,N_47413,N_46805);
nand U49995 (N_49995,N_47620,N_46117);
or U49996 (N_49996,N_47116,N_46973);
xnor U49997 (N_49997,N_47744,N_46778);
or U49998 (N_49998,N_47101,N_46400);
nand U49999 (N_49999,N_47433,N_47765);
nand UO_0 (O_0,N_49553,N_49996);
nand UO_1 (O_1,N_48059,N_48733);
or UO_2 (O_2,N_48251,N_48812);
or UO_3 (O_3,N_48875,N_49486);
or UO_4 (O_4,N_49800,N_48963);
and UO_5 (O_5,N_48917,N_48809);
or UO_6 (O_6,N_49763,N_48602);
or UO_7 (O_7,N_48062,N_48404);
nor UO_8 (O_8,N_48315,N_48317);
nand UO_9 (O_9,N_48137,N_49739);
nor UO_10 (O_10,N_49610,N_48111);
or UO_11 (O_11,N_48167,N_48632);
nand UO_12 (O_12,N_48598,N_49213);
or UO_13 (O_13,N_48813,N_48369);
nand UO_14 (O_14,N_49359,N_49161);
xor UO_15 (O_15,N_48792,N_48780);
and UO_16 (O_16,N_49226,N_49958);
nand UO_17 (O_17,N_48740,N_48328);
and UO_18 (O_18,N_48377,N_48676);
nand UO_19 (O_19,N_48810,N_48991);
and UO_20 (O_20,N_48063,N_49258);
or UO_21 (O_21,N_49232,N_48634);
and UO_22 (O_22,N_48175,N_49372);
or UO_23 (O_23,N_49050,N_48020);
and UO_24 (O_24,N_49519,N_49592);
or UO_25 (O_25,N_48594,N_49263);
nor UO_26 (O_26,N_48070,N_49555);
nand UO_27 (O_27,N_48470,N_48372);
nand UO_28 (O_28,N_49734,N_49939);
nor UO_29 (O_29,N_49749,N_48435);
or UO_30 (O_30,N_48698,N_49582);
and UO_31 (O_31,N_48086,N_49973);
and UO_32 (O_32,N_49950,N_49709);
nor UO_33 (O_33,N_49275,N_49712);
nand UO_34 (O_34,N_49398,N_49572);
and UO_35 (O_35,N_48541,N_49145);
nand UO_36 (O_36,N_49025,N_48308);
or UO_37 (O_37,N_48544,N_48845);
or UO_38 (O_38,N_48010,N_48718);
nand UO_39 (O_39,N_48233,N_49037);
and UO_40 (O_40,N_48143,N_49424);
nor UO_41 (O_41,N_48411,N_48546);
and UO_42 (O_42,N_48262,N_48774);
nor UO_43 (O_43,N_48030,N_48280);
or UO_44 (O_44,N_48914,N_49838);
nand UO_45 (O_45,N_48322,N_49351);
nor UO_46 (O_46,N_48507,N_49696);
or UO_47 (O_47,N_48343,N_48336);
nor UO_48 (O_48,N_48305,N_49735);
and UO_49 (O_49,N_48007,N_48359);
nor UO_50 (O_50,N_48680,N_49986);
and UO_51 (O_51,N_49971,N_49860);
nand UO_52 (O_52,N_49403,N_48713);
nor UO_53 (O_53,N_48422,N_49629);
or UO_54 (O_54,N_48569,N_49741);
nand UO_55 (O_55,N_49779,N_48552);
or UO_56 (O_56,N_49787,N_48656);
nand UO_57 (O_57,N_49501,N_49068);
nand UO_58 (O_58,N_48088,N_49512);
nand UO_59 (O_59,N_49984,N_49464);
or UO_60 (O_60,N_48094,N_48858);
and UO_61 (O_61,N_48442,N_48169);
or UO_62 (O_62,N_48884,N_48702);
nor UO_63 (O_63,N_48313,N_48110);
nand UO_64 (O_64,N_48530,N_49777);
or UO_65 (O_65,N_48661,N_48784);
or UO_66 (O_66,N_48974,N_48856);
and UO_67 (O_67,N_48686,N_49943);
nand UO_68 (O_68,N_48432,N_49071);
or UO_69 (O_69,N_49142,N_49184);
nand UO_70 (O_70,N_49294,N_49962);
nand UO_71 (O_71,N_49388,N_49172);
nor UO_72 (O_72,N_49328,N_48923);
nand UO_73 (O_73,N_48739,N_48332);
nand UO_74 (O_74,N_49931,N_48868);
nor UO_75 (O_75,N_48482,N_49626);
or UO_76 (O_76,N_48877,N_49008);
or UO_77 (O_77,N_48467,N_49586);
nand UO_78 (O_78,N_48076,N_48558);
and UO_79 (O_79,N_48590,N_48842);
or UO_80 (O_80,N_49558,N_49535);
and UO_81 (O_81,N_48453,N_49446);
or UO_82 (O_82,N_48985,N_49768);
nor UO_83 (O_83,N_49300,N_48023);
nand UO_84 (O_84,N_48256,N_49603);
nand UO_85 (O_85,N_48937,N_48350);
and UO_86 (O_86,N_49652,N_49339);
nand UO_87 (O_87,N_49277,N_49547);
or UO_88 (O_88,N_49571,N_49422);
nand UO_89 (O_89,N_49459,N_49659);
or UO_90 (O_90,N_49759,N_49577);
nor UO_91 (O_91,N_48365,N_48243);
and UO_92 (O_92,N_49549,N_48260);
or UO_93 (O_93,N_48289,N_49761);
nand UO_94 (O_94,N_48014,N_49385);
or UO_95 (O_95,N_49011,N_48886);
and UO_96 (O_96,N_49764,N_48640);
xnor UO_97 (O_97,N_49925,N_48438);
or UO_98 (O_98,N_48954,N_48840);
and UO_99 (O_99,N_48794,N_49615);
and UO_100 (O_100,N_49301,N_49742);
nand UO_101 (O_101,N_49278,N_48491);
or UO_102 (O_102,N_48978,N_48597);
and UO_103 (O_103,N_49798,N_49990);
and UO_104 (O_104,N_48093,N_48203);
nor UO_105 (O_105,N_48098,N_48050);
or UO_106 (O_106,N_49307,N_49831);
or UO_107 (O_107,N_49695,N_48074);
or UO_108 (O_108,N_48879,N_49835);
nand UO_109 (O_109,N_48120,N_49094);
and UO_110 (O_110,N_48814,N_48907);
nor UO_111 (O_111,N_49312,N_48611);
or UO_112 (O_112,N_49518,N_49905);
nor UO_113 (O_113,N_48198,N_49408);
nand UO_114 (O_114,N_48890,N_48061);
nor UO_115 (O_115,N_49253,N_49671);
and UO_116 (O_116,N_49873,N_49108);
nand UO_117 (O_117,N_48752,N_48090);
and UO_118 (O_118,N_48789,N_49368);
nand UO_119 (O_119,N_48997,N_48874);
and UO_120 (O_120,N_48642,N_49751);
nand UO_121 (O_121,N_49323,N_48224);
nand UO_122 (O_122,N_48389,N_48839);
or UO_123 (O_123,N_48992,N_48754);
nand UO_124 (O_124,N_49542,N_49635);
nand UO_125 (O_125,N_49125,N_49225);
and UO_126 (O_126,N_48103,N_48893);
or UO_127 (O_127,N_48679,N_49425);
nor UO_128 (O_128,N_49098,N_48184);
or UO_129 (O_129,N_49684,N_49358);
or UO_130 (O_130,N_48002,N_49076);
nand UO_131 (O_131,N_49435,N_48475);
nand UO_132 (O_132,N_48310,N_48374);
nand UO_133 (O_133,N_48176,N_49233);
nor UO_134 (O_134,N_48926,N_49087);
and UO_135 (O_135,N_48547,N_48827);
and UO_136 (O_136,N_48105,N_48196);
nand UO_137 (O_137,N_48454,N_48246);
nor UO_138 (O_138,N_48832,N_48102);
nand UO_139 (O_139,N_49042,N_49812);
nand UO_140 (O_140,N_49324,N_49165);
nor UO_141 (O_141,N_48881,N_49139);
and UO_142 (O_142,N_48863,N_48019);
nand UO_143 (O_143,N_48747,N_48969);
or UO_144 (O_144,N_48456,N_49148);
nor UO_145 (O_145,N_48637,N_48696);
and UO_146 (O_146,N_48371,N_49663);
nand UO_147 (O_147,N_49389,N_48068);
nor UO_148 (O_148,N_48263,N_48721);
nor UO_149 (O_149,N_48553,N_49951);
xnor UO_150 (O_150,N_49336,N_48716);
or UO_151 (O_151,N_48302,N_49641);
nor UO_152 (O_152,N_49477,N_48849);
nand UO_153 (O_153,N_48542,N_49539);
nand UO_154 (O_154,N_49752,N_49140);
and UO_155 (O_155,N_48887,N_48771);
or UO_156 (O_156,N_49428,N_49030);
nand UO_157 (O_157,N_48555,N_49299);
nor UO_158 (O_158,N_49178,N_48892);
nand UO_159 (O_159,N_48614,N_48587);
nor UO_160 (O_160,N_48517,N_49264);
nor UO_161 (O_161,N_49183,N_48882);
or UO_162 (O_162,N_48770,N_48354);
nand UO_163 (O_163,N_49437,N_48071);
nand UO_164 (O_164,N_49250,N_48357);
nand UO_165 (O_165,N_49997,N_49401);
nor UO_166 (O_166,N_48259,N_49304);
or UO_167 (O_167,N_49999,N_49821);
nor UO_168 (O_168,N_49096,N_49854);
and UO_169 (O_169,N_49255,N_49272);
nand UO_170 (O_170,N_48622,N_49045);
nand UO_171 (O_171,N_49005,N_49107);
nand UO_172 (O_172,N_48218,N_48474);
and UO_173 (O_173,N_48029,N_49186);
nand UO_174 (O_174,N_48975,N_49180);
nor UO_175 (O_175,N_48114,N_48912);
and UO_176 (O_176,N_49719,N_48757);
or UO_177 (O_177,N_49693,N_49536);
nand UO_178 (O_178,N_49772,N_49384);
nand UO_179 (O_179,N_48215,N_49634);
and UO_180 (O_180,N_49793,N_48725);
nand UO_181 (O_181,N_48635,N_48930);
or UO_182 (O_182,N_49920,N_49816);
nor UO_183 (O_183,N_49740,N_49160);
and UO_184 (O_184,N_49820,N_48678);
or UO_185 (O_185,N_49416,N_48013);
nand UO_186 (O_186,N_49157,N_48782);
nand UO_187 (O_187,N_49611,N_49718);
nor UO_188 (O_188,N_49521,N_48621);
nor UO_189 (O_189,N_49009,N_49884);
and UO_190 (O_190,N_48825,N_49297);
nor UO_191 (O_191,N_49972,N_48970);
nor UO_192 (O_192,N_48156,N_48484);
nor UO_193 (O_193,N_48641,N_48488);
nand UO_194 (O_194,N_49061,N_48869);
nor UO_195 (O_195,N_49445,N_49090);
nand UO_196 (O_196,N_48683,N_49033);
or UO_197 (O_197,N_49292,N_48759);
nor UO_198 (O_198,N_48101,N_49126);
and UO_199 (O_199,N_48603,N_49904);
or UO_200 (O_200,N_48387,N_48582);
nor UO_201 (O_201,N_49998,N_49940);
or UO_202 (O_202,N_49482,N_49474);
nand UO_203 (O_203,N_49640,N_48142);
or UO_204 (O_204,N_48091,N_49782);
nor UO_205 (O_205,N_48490,N_48714);
and UO_206 (O_206,N_48146,N_48081);
and UO_207 (O_207,N_49646,N_49612);
and UO_208 (O_208,N_49580,N_48349);
nor UO_209 (O_209,N_49922,N_49326);
nor UO_210 (O_210,N_48031,N_48045);
xor UO_211 (O_211,N_48675,N_49914);
or UO_212 (O_212,N_48950,N_48769);
and UO_213 (O_213,N_48419,N_48445);
and UO_214 (O_214,N_49386,N_49906);
nor UO_215 (O_215,N_49863,N_48178);
and UO_216 (O_216,N_48563,N_49792);
and UO_217 (O_217,N_48133,N_48457);
and UO_218 (O_218,N_49318,N_49209);
and UO_219 (O_219,N_48100,N_49370);
nand UO_220 (O_220,N_48735,N_49607);
nor UO_221 (O_221,N_49097,N_49072);
and UO_222 (O_222,N_48051,N_49155);
or UO_223 (O_223,N_48828,N_49716);
xor UO_224 (O_224,N_49639,N_48451);
nor UO_225 (O_225,N_48551,N_48870);
nand UO_226 (O_226,N_48724,N_48901);
or UO_227 (O_227,N_49419,N_49715);
nand UO_228 (O_228,N_49618,N_49442);
or UO_229 (O_229,N_48841,N_49799);
or UO_230 (O_230,N_49644,N_49010);
nand UO_231 (O_231,N_48158,N_48520);
nor UO_232 (O_232,N_49624,N_48528);
nor UO_233 (O_233,N_48807,N_48727);
nor UO_234 (O_234,N_49393,N_48297);
or UO_235 (O_235,N_49217,N_48557);
nand UO_236 (O_236,N_48258,N_49185);
nand UO_237 (O_237,N_49658,N_48987);
nand UO_238 (O_238,N_48743,N_48538);
and UO_239 (O_239,N_48053,N_49620);
nand UO_240 (O_240,N_49974,N_49462);
or UO_241 (O_241,N_48660,N_48647);
nor UO_242 (O_242,N_49192,N_48666);
and UO_243 (O_243,N_49954,N_48229);
and UO_244 (O_244,N_48899,N_48205);
xnor UO_245 (O_245,N_49282,N_48596);
nand UO_246 (O_246,N_48952,N_49012);
nor UO_247 (O_247,N_48423,N_48136);
nand UO_248 (O_248,N_49786,N_48428);
nand UO_249 (O_249,N_48788,N_49808);
nor UO_250 (O_250,N_48591,N_48844);
or UO_251 (O_251,N_49944,N_49202);
and UO_252 (O_252,N_49016,N_49447);
or UO_253 (O_253,N_48140,N_49177);
or UO_254 (O_254,N_48921,N_48441);
xnor UO_255 (O_255,N_48292,N_48933);
and UO_256 (O_256,N_49948,N_49475);
and UO_257 (O_257,N_48024,N_49632);
nand UO_258 (O_258,N_49724,N_49058);
and UO_259 (O_259,N_49429,N_49167);
and UO_260 (O_260,N_49348,N_48697);
nand UO_261 (O_261,N_49001,N_49055);
nor UO_262 (O_262,N_49814,N_49083);
nand UO_263 (O_263,N_49805,N_49934);
nor UO_264 (O_264,N_48729,N_48961);
and UO_265 (O_265,N_48193,N_49044);
nand UO_266 (O_266,N_49002,N_49861);
or UO_267 (O_267,N_49756,N_48296);
and UO_268 (O_268,N_48157,N_48535);
or UO_269 (O_269,N_49387,N_48608);
nor UO_270 (O_270,N_48499,N_49247);
or UO_271 (O_271,N_48250,N_49622);
nor UO_272 (O_272,N_49551,N_49667);
or UO_273 (O_273,N_49077,N_48511);
or UO_274 (O_274,N_48046,N_49762);
nor UO_275 (O_275,N_48469,N_48909);
nor UO_276 (O_276,N_49063,N_49162);
nand UO_277 (O_277,N_48537,N_49967);
or UO_278 (O_278,N_48798,N_48394);
nand UO_279 (O_279,N_48278,N_48935);
nand UO_280 (O_280,N_49414,N_48505);
nand UO_281 (O_281,N_48385,N_48548);
and UO_282 (O_282,N_49850,N_48461);
nor UO_283 (O_283,N_48958,N_48414);
and UO_284 (O_284,N_48577,N_48004);
nand UO_285 (O_285,N_49891,N_48763);
nor UO_286 (O_286,N_49830,N_49885);
and UO_287 (O_287,N_48211,N_49164);
nand UO_288 (O_288,N_49809,N_49856);
and UO_289 (O_289,N_49991,N_49054);
nand UO_290 (O_290,N_48944,N_48312);
and UO_291 (O_291,N_48352,N_49917);
nor UO_292 (O_292,N_49034,N_48915);
and UO_293 (O_293,N_49257,N_48630);
nand UO_294 (O_294,N_49606,N_49849);
or UO_295 (O_295,N_49362,N_48035);
and UO_296 (O_296,N_49106,N_48615);
or UO_297 (O_297,N_49598,N_49173);
and UO_298 (O_298,N_48271,N_48896);
nor UO_299 (O_299,N_48397,N_49600);
nand UO_300 (O_300,N_49817,N_49691);
and UO_301 (O_301,N_49352,N_49911);
nor UO_302 (O_302,N_48465,N_49137);
and UO_303 (O_303,N_48040,N_48973);
and UO_304 (O_304,N_49395,N_49952);
nor UO_305 (O_305,N_49579,N_49495);
nor UO_306 (O_306,N_49074,N_48130);
nand UO_307 (O_307,N_49841,N_48464);
nand UO_308 (O_308,N_49758,N_49375);
or UO_309 (O_309,N_48108,N_49754);
and UO_310 (O_310,N_48138,N_49857);
nor UO_311 (O_311,N_49427,N_48818);
and UO_312 (O_312,N_49554,N_48638);
nand UO_313 (O_313,N_49811,N_49886);
or UO_314 (O_314,N_48709,N_49478);
and UO_315 (O_315,N_48715,N_48982);
and UO_316 (O_316,N_48391,N_48938);
nand UO_317 (O_317,N_48329,N_49287);
and UO_318 (O_318,N_48304,N_48787);
nand UO_319 (O_319,N_49169,N_49597);
nor UO_320 (O_320,N_49774,N_48363);
nand UO_321 (O_321,N_49665,N_48965);
nor UO_322 (O_322,N_49866,N_49086);
and UO_323 (O_323,N_49229,N_49660);
and UO_324 (O_324,N_49656,N_48180);
nand UO_325 (O_325,N_48052,N_48960);
nand UO_326 (O_326,N_49621,N_48254);
nand UO_327 (O_327,N_48820,N_49676);
nor UO_328 (O_328,N_48947,N_48286);
nand UO_329 (O_329,N_48823,N_49678);
nor UO_330 (O_330,N_49584,N_49291);
or UO_331 (O_331,N_48144,N_49338);
nand UO_332 (O_332,N_48485,N_49065);
nor UO_333 (O_333,N_48562,N_49095);
nor UO_334 (O_334,N_48522,N_48762);
or UO_335 (O_335,N_49988,N_48850);
and UO_336 (O_336,N_49867,N_48885);
nand UO_337 (O_337,N_48356,N_48346);
nor UO_338 (O_338,N_49785,N_49410);
or UO_339 (O_339,N_48192,N_49770);
and UO_340 (O_340,N_48089,N_48121);
nor UO_341 (O_341,N_48135,N_49059);
or UO_342 (O_342,N_49092,N_48943);
nand UO_343 (O_343,N_49713,N_49175);
and UO_344 (O_344,N_48948,N_48241);
nor UO_345 (O_345,N_49360,N_48496);
and UO_346 (O_346,N_49670,N_48413);
nor UO_347 (O_347,N_48934,N_48309);
or UO_348 (O_348,N_49119,N_48913);
and UO_349 (O_349,N_48204,N_49605);
nand UO_350 (O_350,N_49721,N_49132);
nand UO_351 (O_351,N_48426,N_48689);
or UO_352 (O_352,N_48604,N_49067);
or UO_353 (O_353,N_49921,N_48816);
nor UO_354 (O_354,N_49932,N_48468);
or UO_355 (O_355,N_48447,N_49623);
nor UO_356 (O_356,N_48584,N_48351);
nor UO_357 (O_357,N_48036,N_48168);
nand UO_358 (O_358,N_49546,N_48065);
or UO_359 (O_359,N_49982,N_49134);
and UO_360 (O_360,N_49804,N_49647);
nand UO_361 (O_361,N_48772,N_49527);
nor UO_362 (O_362,N_48449,N_48580);
or UO_363 (O_363,N_49374,N_48480);
nand UO_364 (O_364,N_49440,N_48682);
and UO_365 (O_365,N_48510,N_49200);
or UO_366 (O_366,N_48247,N_49563);
nor UO_367 (O_367,N_49672,N_48731);
and UO_368 (O_368,N_49957,N_48402);
nor UO_369 (O_369,N_48448,N_48172);
and UO_370 (O_370,N_48959,N_49460);
and UO_371 (O_371,N_48131,N_49685);
nor UO_372 (O_372,N_48124,N_49942);
nand UO_373 (O_373,N_49214,N_49513);
or UO_374 (O_374,N_49968,N_48589);
nand UO_375 (O_375,N_49941,N_49454);
and UO_376 (O_376,N_48116,N_48382);
nor UO_377 (O_377,N_48139,N_49468);
nor UO_378 (O_378,N_48430,N_49994);
nor UO_379 (O_379,N_48295,N_49484);
nor UO_380 (O_380,N_49882,N_48236);
and UO_381 (O_381,N_48011,N_49767);
nand UO_382 (O_382,N_49784,N_48655);
or UO_383 (O_383,N_49864,N_49587);
nand UO_384 (O_384,N_48920,N_48189);
nand UO_385 (O_385,N_49955,N_49491);
and UO_386 (O_386,N_49559,N_49382);
or UO_387 (O_387,N_48670,N_49455);
nand UO_388 (O_388,N_48012,N_49568);
nor UO_389 (O_389,N_48099,N_49732);
or UO_390 (O_390,N_49893,N_49201);
and UO_391 (O_391,N_49913,N_49130);
or UO_392 (O_392,N_48472,N_49631);
nor UO_393 (O_393,N_48037,N_48860);
nor UO_394 (O_394,N_48166,N_48182);
nand UO_395 (O_395,N_49488,N_49216);
or UO_396 (O_396,N_48941,N_49923);
and UO_397 (O_397,N_48095,N_49397);
nor UO_398 (O_398,N_48235,N_49953);
nand UO_399 (O_399,N_48344,N_48593);
nor UO_400 (O_400,N_48085,N_49028);
nand UO_401 (O_401,N_48303,N_49279);
nand UO_402 (O_402,N_48900,N_48519);
nor UO_403 (O_403,N_48072,N_48878);
or UO_404 (O_404,N_48216,N_49476);
and UO_405 (O_405,N_48880,N_49969);
nand UO_406 (O_406,N_48160,N_49411);
and UO_407 (O_407,N_48364,N_48155);
or UO_408 (O_408,N_48237,N_49935);
nor UO_409 (O_409,N_48183,N_49507);
or UO_410 (O_410,N_48043,N_49918);
nor UO_411 (O_411,N_49625,N_48612);
xor UO_412 (O_412,N_49066,N_48161);
or UO_413 (O_413,N_49898,N_49039);
nand UO_414 (O_414,N_49760,N_48925);
or UO_415 (O_415,N_49677,N_49823);
and UO_416 (O_416,N_49222,N_49115);
or UO_417 (O_417,N_49723,N_48779);
and UO_418 (O_418,N_48534,N_49285);
xnor UO_419 (O_419,N_49268,N_49506);
or UO_420 (O_420,N_48898,N_49069);
and UO_421 (O_421,N_48373,N_49158);
nand UO_422 (O_422,N_49569,N_49589);
and UO_423 (O_423,N_49824,N_48822);
nor UO_424 (O_424,N_48269,N_49581);
nand UO_425 (O_425,N_48338,N_49230);
and UO_426 (O_426,N_49887,N_48261);
nor UO_427 (O_427,N_49879,N_49977);
xnor UO_428 (O_428,N_48924,N_48625);
nand UO_429 (O_429,N_48749,N_48624);
or UO_430 (O_430,N_49206,N_48654);
or UO_431 (O_431,N_48127,N_48658);
nor UO_432 (O_432,N_48345,N_48831);
or UO_433 (O_433,N_49181,N_48026);
xor UO_434 (O_434,N_49281,N_48703);
nor UO_435 (O_435,N_48358,N_48477);
or UO_436 (O_436,N_48032,N_48122);
and UO_437 (O_437,N_48623,N_48571);
nand UO_438 (O_438,N_49170,N_48060);
or UO_439 (O_439,N_48575,N_49947);
nor UO_440 (O_440,N_49241,N_48222);
nand UO_441 (O_441,N_49528,N_48293);
nor UO_442 (O_442,N_49243,N_48483);
nor UO_443 (O_443,N_49755,N_48576);
nor UO_444 (O_444,N_48202,N_48601);
nand UO_445 (O_445,N_48561,N_49190);
nand UO_446 (O_446,N_49638,N_49057);
xor UO_447 (O_447,N_49807,N_49480);
nand UO_448 (O_448,N_48989,N_49104);
nand UO_449 (O_449,N_48775,N_49515);
or UO_450 (O_450,N_49053,N_48836);
and UO_451 (O_451,N_48034,N_48643);
and UO_452 (O_452,N_49341,N_48055);
nor UO_453 (O_453,N_49650,N_48437);
nor UO_454 (O_454,N_48786,N_49203);
nor UO_455 (O_455,N_48560,N_48790);
nor UO_456 (O_456,N_48949,N_49564);
or UO_457 (O_457,N_49070,N_49084);
and UO_458 (O_458,N_48170,N_49688);
nand UO_459 (O_459,N_49645,N_48618);
and UO_460 (O_460,N_49191,N_48768);
nand UO_461 (O_461,N_48502,N_48527);
or UO_462 (O_462,N_49946,N_49593);
or UO_463 (O_463,N_49750,N_48054);
nand UO_464 (O_464,N_48791,N_49796);
nor UO_465 (O_465,N_49692,N_49706);
nor UO_466 (O_466,N_49727,N_48570);
nor UO_467 (O_467,N_49182,N_49007);
and UO_468 (O_468,N_49035,N_49483);
xor UO_469 (O_469,N_49357,N_49004);
or UO_470 (O_470,N_48817,N_49500);
nand UO_471 (O_471,N_48700,N_48244);
nand UO_472 (O_472,N_49235,N_49109);
and UO_473 (O_473,N_48298,N_48931);
and UO_474 (O_474,N_49510,N_49046);
nand UO_475 (O_475,N_48957,N_48273);
and UO_476 (O_476,N_49556,N_48383);
or UO_477 (O_477,N_49062,N_48330);
or UO_478 (O_478,N_49150,N_48486);
and UO_479 (O_479,N_49080,N_49687);
and UO_480 (O_480,N_48574,N_49633);
nor UO_481 (O_481,N_49079,N_48498);
nor UO_482 (O_482,N_48240,N_49060);
nand UO_483 (O_483,N_49021,N_49674);
xor UO_484 (O_484,N_48766,N_49031);
nand UO_485 (O_485,N_48819,N_49138);
nand UO_486 (O_486,N_49211,N_48946);
nand UO_487 (O_487,N_48573,N_49356);
or UO_488 (O_488,N_49810,N_49493);
nand UO_489 (O_489,N_49228,N_49333);
or UO_490 (O_490,N_48529,N_49859);
and UO_491 (O_491,N_49198,N_48039);
or UO_492 (O_492,N_49701,N_48079);
nor UO_493 (O_493,N_48018,N_49381);
nor UO_494 (O_494,N_49818,N_48471);
nand UO_495 (O_495,N_49273,N_48245);
xnor UO_496 (O_496,N_49993,N_49566);
nand UO_497 (O_497,N_49259,N_48797);
or UO_498 (O_498,N_49284,N_48181);
and UO_499 (O_499,N_48672,N_49526);
nand UO_500 (O_500,N_49089,N_49795);
nand UO_501 (O_501,N_48977,N_48227);
nand UO_502 (O_502,N_49827,N_49319);
xnor UO_503 (O_503,N_48776,N_48639);
or UO_504 (O_504,N_49047,N_49912);
and UO_505 (O_505,N_49964,N_48097);
and UO_506 (O_506,N_48238,N_49858);
or UO_507 (O_507,N_48665,N_49305);
nor UO_508 (O_508,N_49049,N_49985);
or UO_509 (O_509,N_48409,N_49806);
nand UO_510 (O_510,N_49657,N_48866);
and UO_511 (O_511,N_49003,N_49469);
nor UO_512 (O_512,N_48760,N_49788);
and UO_513 (O_513,N_49438,N_49655);
nor UO_514 (O_514,N_49583,N_49205);
nand UO_515 (O_515,N_48523,N_48671);
nor UO_516 (O_516,N_49423,N_49544);
nor UO_517 (O_517,N_49364,N_49680);
and UO_518 (O_518,N_48141,N_48016);
nor UO_519 (O_519,N_48104,N_49240);
nor UO_520 (O_520,N_48609,N_49430);
or UO_521 (O_521,N_49862,N_48347);
nand UO_522 (O_522,N_49270,N_48500);
and UO_523 (O_523,N_49872,N_49743);
nand UO_524 (O_524,N_49373,N_48399);
nor UO_525 (O_525,N_48764,N_49842);
and UO_526 (O_526,N_49899,N_48288);
and UO_527 (O_527,N_49567,N_48585);
and UO_528 (O_528,N_48986,N_48669);
nand UO_529 (O_529,N_49027,N_48277);
and UO_530 (O_530,N_48846,N_49753);
nor UO_531 (O_531,N_49855,N_48325);
or UO_532 (O_532,N_49550,N_49141);
or UO_533 (O_533,N_49113,N_49212);
nor UO_534 (O_534,N_48195,N_48755);
and UO_535 (O_535,N_49619,N_48212);
nor UO_536 (O_536,N_49746,N_49869);
or UO_537 (O_537,N_48199,N_49149);
or UO_538 (O_538,N_48125,N_48478);
or UO_539 (O_539,N_49189,N_48695);
or UO_540 (O_540,N_48164,N_49533);
nor UO_541 (O_541,N_48300,N_49231);
and UO_542 (O_542,N_49714,N_49129);
or UO_543 (O_543,N_49245,N_48777);
or UO_544 (O_544,N_48324,N_48514);
and UO_545 (O_545,N_48540,N_49116);
or UO_546 (O_546,N_48793,N_48190);
or UO_547 (O_547,N_49127,N_48421);
and UO_548 (O_548,N_49836,N_48267);
nor UO_549 (O_549,N_49451,N_48811);
and UO_550 (O_550,N_48028,N_49237);
or UO_551 (O_551,N_49538,N_48765);
nand UO_552 (O_552,N_49215,N_48613);
nor UO_553 (O_553,N_48410,N_49329);
nor UO_554 (O_554,N_48871,N_48804);
or UO_555 (O_555,N_48748,N_49269);
nand UO_556 (O_556,N_48194,N_48022);
or UO_557 (O_557,N_49453,N_49023);
or UO_558 (O_558,N_48069,N_49654);
nor UO_559 (O_559,N_49154,N_48439);
or UO_560 (O_560,N_48084,N_48805);
or UO_561 (O_561,N_49135,N_48290);
or UO_562 (O_562,N_49147,N_49280);
or UO_563 (O_563,N_48526,N_48711);
or UO_564 (O_564,N_49653,N_49418);
or UO_565 (O_565,N_48185,N_48862);
and UO_566 (O_566,N_49219,N_49421);
nand UO_567 (O_567,N_48384,N_48545);
xor UO_568 (O_568,N_48631,N_48567);
nand UO_569 (O_569,N_49794,N_48972);
nor UO_570 (O_570,N_49517,N_48966);
or UO_571 (O_571,N_49846,N_49790);
nor UO_572 (O_572,N_49662,N_49681);
or UO_573 (O_573,N_48283,N_48327);
nand UO_574 (O_574,N_48268,N_49965);
and UO_575 (O_575,N_48588,N_49490);
nand UO_576 (O_576,N_49992,N_48559);
or UO_577 (O_577,N_49578,N_48801);
nand UO_578 (O_578,N_49350,N_49588);
or UO_579 (O_579,N_48824,N_49532);
nand UO_580 (O_580,N_48458,N_49839);
or UO_581 (O_581,N_49342,N_49166);
nor UO_582 (O_582,N_49371,N_49327);
nor UO_583 (O_583,N_48436,N_48493);
or UO_584 (O_584,N_49103,N_49596);
nor UO_585 (O_585,N_48843,N_49874);
nor UO_586 (O_586,N_48208,N_49819);
nand UO_587 (O_587,N_48319,N_48460);
or UO_588 (O_588,N_48440,N_49980);
and UO_589 (O_589,N_48512,N_49473);
nand UO_590 (O_590,N_49575,N_48835);
and UO_591 (O_591,N_49013,N_48368);
and UO_592 (O_592,N_49431,N_48781);
and UO_593 (O_593,N_49888,N_48539);
nor UO_594 (O_594,N_49406,N_49239);
nand UO_595 (O_595,N_49498,N_48953);
and UO_596 (O_596,N_48857,N_49366);
and UO_597 (O_597,N_48504,N_49744);
nor UO_598 (O_598,N_49875,N_48407);
nor UO_599 (O_599,N_48000,N_49343);
nor UO_600 (O_600,N_48285,N_49347);
or UO_601 (O_601,N_49552,N_49697);
or UO_602 (O_602,N_49499,N_48891);
nand UO_603 (O_603,N_48188,N_49668);
nand UO_604 (O_604,N_48566,N_49334);
and UO_605 (O_605,N_49252,N_48684);
nor UO_606 (O_606,N_48006,N_48888);
and UO_607 (O_607,N_49910,N_49355);
nor UO_608 (O_608,N_48653,N_49496);
nor UO_609 (O_609,N_48607,N_49995);
nand UO_610 (O_610,N_48126,N_48064);
and UO_611 (O_611,N_48876,N_49609);
or UO_612 (O_612,N_49531,N_48861);
nand UO_613 (O_613,N_49492,N_48657);
nor UO_614 (O_614,N_49249,N_48424);
and UO_615 (O_615,N_49308,N_49413);
or UO_616 (O_616,N_49745,N_48370);
and UO_617 (O_617,N_49694,N_48177);
and UO_618 (O_618,N_49017,N_48922);
or UO_619 (O_619,N_48979,N_49780);
nand UO_620 (O_620,N_48264,N_48734);
xor UO_621 (O_621,N_48153,N_48080);
or UO_622 (O_622,N_49470,N_49895);
xnor UO_623 (O_623,N_49497,N_49458);
or UO_624 (O_624,N_48940,N_48287);
and UO_625 (O_625,N_49311,N_48854);
nor UO_626 (O_626,N_49293,N_49573);
nor UO_627 (O_627,N_49251,N_48515);
or UO_628 (O_628,N_49729,N_48737);
nand UO_629 (O_629,N_48320,N_49594);
and UO_630 (O_630,N_49174,N_48291);
nor UO_631 (O_631,N_49502,N_49043);
or UO_632 (O_632,N_48600,N_48730);
nand UO_633 (O_633,N_48200,N_49883);
nor UO_634 (O_634,N_49315,N_48281);
or UO_635 (O_635,N_48257,N_48586);
and UO_636 (O_636,N_48223,N_48487);
nand UO_637 (O_637,N_49353,N_48513);
and UO_638 (O_638,N_48400,N_48929);
or UO_639 (O_639,N_49335,N_48651);
or UO_640 (O_640,N_49637,N_48995);
or UO_641 (O_641,N_48406,N_48082);
xnor UO_642 (O_642,N_49396,N_48107);
or UO_643 (O_643,N_49876,N_48848);
and UO_644 (O_644,N_48756,N_48838);
or UO_645 (O_645,N_48710,N_49298);
and UO_646 (O_646,N_49987,N_49244);
nand UO_647 (O_647,N_49267,N_49833);
nand UO_648 (O_648,N_49195,N_49412);
or UO_649 (O_649,N_48207,N_49602);
nor UO_650 (O_650,N_49036,N_48663);
nor UO_651 (O_651,N_48939,N_49121);
nor UO_652 (O_652,N_49933,N_49927);
and UO_653 (O_653,N_49112,N_49199);
or UO_654 (O_654,N_48009,N_48617);
or UO_655 (O_655,N_49524,N_49144);
nand UO_656 (O_656,N_49783,N_48796);
xnor UO_657 (O_657,N_49377,N_48745);
and UO_658 (O_658,N_48549,N_49117);
nor UO_659 (O_659,N_48230,N_48726);
and UO_660 (O_660,N_48691,N_48918);
or UO_661 (O_661,N_48983,N_48837);
or UO_662 (O_662,N_49073,N_48038);
or UO_663 (O_663,N_49907,N_49114);
nor UO_664 (O_664,N_48531,N_48221);
nor UO_665 (O_665,N_48964,N_48503);
nand UO_666 (O_666,N_49390,N_48113);
nand UO_667 (O_667,N_48806,N_49560);
and UO_668 (O_668,N_48412,N_49832);
or UO_669 (O_669,N_48708,N_49325);
nor UO_670 (O_670,N_48025,N_48165);
xnor UO_671 (O_671,N_49574,N_48967);
and UO_672 (O_672,N_49781,N_48228);
and UO_673 (O_673,N_48149,N_49101);
nor UO_674 (O_674,N_49306,N_49664);
nand UO_675 (O_675,N_49345,N_49367);
nand UO_676 (O_676,N_49020,N_49930);
nor UO_677 (O_677,N_48742,N_49890);
nand UO_678 (O_678,N_49908,N_48951);
nand UO_679 (O_679,N_49402,N_49604);
nor UO_680 (O_680,N_49099,N_49757);
and UO_681 (O_681,N_48393,N_49441);
nand UO_682 (O_682,N_48688,N_48645);
and UO_683 (O_683,N_48220,N_49194);
nor UO_684 (O_684,N_48706,N_49029);
nor UO_685 (O_685,N_49591,N_48783);
or UO_686 (O_686,N_48728,N_48629);
or UO_687 (O_687,N_48232,N_49110);
and UO_688 (O_688,N_49516,N_48865);
or UO_689 (O_689,N_49979,N_48785);
nand UO_690 (O_690,N_49426,N_48701);
or UO_691 (O_691,N_49179,N_49153);
or UO_692 (O_692,N_49511,N_49710);
and UO_693 (O_693,N_49679,N_49018);
or UO_694 (O_694,N_49405,N_48276);
or UO_695 (O_695,N_49837,N_48916);
nand UO_696 (O_696,N_49014,N_48392);
and UO_697 (O_697,N_48579,N_48096);
or UO_698 (O_698,N_48362,N_48668);
nor UO_699 (O_699,N_49196,N_49349);
and UO_700 (O_700,N_49537,N_48353);
nand UO_701 (O_701,N_49248,N_48583);
nor UO_702 (O_702,N_48897,N_49344);
and UO_703 (O_703,N_49938,N_48659);
or UO_704 (O_704,N_48873,N_49880);
nand UO_705 (O_705,N_48459,N_48524);
nor UO_706 (O_706,N_49223,N_49828);
and UO_707 (O_707,N_49064,N_49983);
nand UO_708 (O_708,N_49363,N_48027);
and UO_709 (O_709,N_49726,N_48677);
nand UO_710 (O_710,N_49815,N_48056);
and UO_711 (O_711,N_49963,N_49124);
and UO_712 (O_712,N_48401,N_48699);
nand UO_713 (O_713,N_49444,N_48106);
xnor UO_714 (O_714,N_49826,N_48339);
nor UO_715 (O_715,N_49168,N_49522);
nand UO_716 (O_716,N_48521,N_48687);
and UO_717 (O_717,N_48331,N_48648);
nand UO_718 (O_718,N_49093,N_49494);
and UO_719 (O_719,N_48209,N_48518);
nor UO_720 (O_720,N_48750,N_48802);
nand UO_721 (O_721,N_49630,N_48083);
nand UO_722 (O_722,N_48154,N_48556);
and UO_723 (O_723,N_49529,N_48318);
or UO_724 (O_724,N_49000,N_49682);
and UO_725 (O_725,N_48872,N_49848);
and UO_726 (O_726,N_48077,N_49928);
and UO_727 (O_727,N_48375,N_48605);
nand UO_728 (O_728,N_48741,N_48867);
nand UO_729 (O_729,N_48129,N_48800);
nand UO_730 (O_730,N_49978,N_49015);
and UO_731 (O_731,N_49467,N_49262);
and UO_732 (O_732,N_48723,N_48173);
nand UO_733 (O_733,N_49032,N_48910);
nor UO_734 (O_734,N_48851,N_49056);
and UO_735 (O_735,N_48058,N_49585);
or UO_736 (O_736,N_48418,N_49616);
or UO_737 (O_737,N_49224,N_49613);
nor UO_738 (O_738,N_49523,N_49207);
nor UO_739 (O_739,N_49797,N_48693);
or UO_740 (O_740,N_49024,N_48554);
nand UO_741 (O_741,N_48187,N_48214);
nor UO_742 (O_742,N_49590,N_48833);
or UO_743 (O_743,N_49290,N_48415);
or UO_744 (O_744,N_49040,N_48501);
and UO_745 (O_745,N_49407,N_49570);
nand UO_746 (O_746,N_48252,N_48803);
nor UO_747 (O_747,N_48853,N_49617);
or UO_748 (O_748,N_49791,N_48429);
and UO_749 (O_749,N_49322,N_48226);
and UO_750 (O_750,N_48316,N_49261);
and UO_751 (O_751,N_49378,N_49840);
nor UO_752 (O_752,N_48301,N_49242);
or UO_753 (O_753,N_49970,N_48980);
and UO_754 (O_754,N_48444,N_48378);
nor UO_755 (O_755,N_48906,N_49091);
and UO_756 (O_756,N_48619,N_49399);
nand UO_757 (O_757,N_49082,N_49961);
nor UO_758 (O_758,N_49699,N_48466);
or UO_759 (O_759,N_48008,N_48994);
or UO_760 (O_760,N_49903,N_49465);
or UO_761 (O_761,N_49197,N_49088);
or UO_762 (O_762,N_49853,N_49924);
xor UO_763 (O_763,N_49989,N_48396);
nand UO_764 (O_764,N_48627,N_49276);
and UO_765 (O_765,N_49210,N_49321);
nor UO_766 (O_766,N_49380,N_48506);
nand UO_767 (O_767,N_49737,N_49118);
nand UO_768 (O_768,N_48649,N_49220);
and UO_769 (O_769,N_49286,N_49878);
nor UO_770 (O_770,N_49975,N_48911);
or UO_771 (O_771,N_49234,N_48073);
nor UO_772 (O_772,N_48826,N_49471);
nor UO_773 (O_773,N_49822,N_48998);
nand UO_774 (O_774,N_48674,N_49417);
nor UO_775 (O_775,N_48834,N_48633);
nand UO_776 (O_776,N_48495,N_49163);
nor UO_777 (O_777,N_49434,N_49929);
or UO_778 (O_778,N_49956,N_49916);
and UO_779 (O_779,N_48213,N_49265);
and UO_780 (O_780,N_49766,N_49520);
or UO_781 (O_781,N_49936,N_49669);
or UO_782 (O_782,N_49801,N_49960);
xnor UO_783 (O_783,N_48446,N_48306);
nor UO_784 (O_784,N_48489,N_48201);
and UO_785 (O_785,N_48455,N_49711);
or UO_786 (O_786,N_48386,N_49433);
nand UO_787 (O_787,N_48463,N_49379);
nor UO_788 (O_788,N_49627,N_49949);
nand UO_789 (O_789,N_48242,N_49466);
nand UO_790 (O_790,N_49508,N_48048);
and UO_791 (O_791,N_49236,N_48395);
nand UO_792 (O_792,N_48905,N_49728);
nor UO_793 (O_793,N_49019,N_48956);
and UO_794 (O_794,N_49081,N_49509);
nor UO_795 (O_795,N_49136,N_49048);
or UO_796 (O_796,N_49773,N_49120);
or UO_797 (O_797,N_48650,N_48361);
nand UO_798 (O_798,N_48830,N_48606);
nand UO_799 (O_799,N_48962,N_49651);
and UO_800 (O_800,N_49976,N_48075);
and UO_801 (O_801,N_48626,N_48145);
and UO_802 (O_802,N_49673,N_48494);
nand UO_803 (O_803,N_49845,N_48509);
or UO_804 (O_804,N_49376,N_48599);
and UO_805 (O_805,N_48497,N_48942);
nand UO_806 (O_806,N_49851,N_48692);
or UO_807 (O_807,N_49151,N_48274);
and UO_808 (O_808,N_48732,N_48981);
nor UO_809 (O_809,N_49829,N_48206);
and UO_810 (O_810,N_48955,N_48335);
and UO_811 (O_811,N_48847,N_49041);
and UO_812 (O_812,N_48543,N_49541);
nand UO_813 (O_813,N_49813,N_48919);
nor UO_814 (O_814,N_48253,N_48408);
nand UO_815 (O_815,N_48128,N_49100);
or UO_816 (O_816,N_48334,N_49485);
nor UO_817 (O_817,N_49843,N_48720);
or UO_818 (O_818,N_48864,N_48163);
nor UO_819 (O_819,N_48667,N_49661);
or UO_820 (O_820,N_49187,N_48294);
and UO_821 (O_821,N_48425,N_48078);
and UO_822 (O_822,N_49881,N_48829);
and UO_823 (O_823,N_49844,N_48225);
nand UO_824 (O_824,N_48067,N_48799);
nand UO_825 (O_825,N_49227,N_49643);
nand UO_826 (O_826,N_49254,N_49038);
nor UO_827 (O_827,N_48323,N_48017);
and UO_828 (O_828,N_48284,N_48533);
and UO_829 (O_829,N_48255,N_48753);
nand UO_830 (O_830,N_48366,N_48171);
xnor UO_831 (O_831,N_48003,N_48664);
or UO_832 (O_832,N_49332,N_49901);
nor UO_833 (O_833,N_48927,N_48644);
nor UO_834 (O_834,N_49557,N_48744);
nand UO_835 (O_835,N_48685,N_49900);
and UO_836 (O_836,N_49051,N_48360);
and UO_837 (O_837,N_49877,N_49420);
or UO_838 (O_838,N_49266,N_49540);
or UO_839 (O_839,N_49303,N_48266);
nor UO_840 (O_840,N_48492,N_49204);
or UO_841 (O_841,N_48279,N_49152);
or UO_842 (O_842,N_48047,N_49705);
and UO_843 (O_843,N_49937,N_48808);
and UO_844 (O_844,N_48525,N_49525);
xor UO_845 (O_845,N_49725,N_48738);
nand UO_846 (O_846,N_49565,N_48342);
and UO_847 (O_847,N_49256,N_48572);
or UO_848 (O_848,N_48815,N_49449);
or UO_849 (O_849,N_48147,N_49218);
nand UO_850 (O_850,N_49075,N_49897);
or UO_851 (O_851,N_48662,N_49365);
nor UO_852 (O_852,N_48348,N_49847);
and UO_853 (O_853,N_49505,N_48751);
nor UO_854 (O_854,N_49436,N_49503);
xor UO_855 (O_855,N_49026,N_49765);
and UO_856 (O_856,N_48416,N_49283);
nor UO_857 (O_857,N_49769,N_49085);
nor UO_858 (O_858,N_48152,N_49747);
nor UO_859 (O_859,N_48889,N_49834);
or UO_860 (O_860,N_49628,N_48620);
nand UO_861 (O_861,N_49105,N_48719);
nand UO_862 (O_862,N_49868,N_48673);
or UO_863 (O_863,N_48379,N_49776);
and UO_864 (O_864,N_49703,N_49317);
nor UO_865 (O_865,N_48707,N_48115);
nor UO_866 (O_866,N_49450,N_49530);
or UO_867 (O_867,N_48564,N_48005);
nor UO_868 (O_868,N_48239,N_48536);
and UO_869 (O_869,N_49926,N_49052);
xnor UO_870 (O_870,N_49738,N_48646);
nor UO_871 (O_871,N_48381,N_48333);
nor UO_872 (O_872,N_48433,N_48452);
nand UO_873 (O_873,N_48118,N_48936);
nor UO_874 (O_874,N_49354,N_48341);
nand UO_875 (O_875,N_49775,N_48057);
nor UO_876 (O_876,N_49642,N_48712);
or UO_877 (O_877,N_48398,N_49221);
nor UO_878 (O_878,N_49481,N_48092);
or UO_879 (O_879,N_48990,N_48581);
nand UO_880 (O_880,N_49463,N_48042);
or UO_881 (O_881,N_48337,N_48066);
or UO_882 (O_882,N_48134,N_48717);
or UO_883 (O_883,N_49733,N_48636);
nand UO_884 (O_884,N_48307,N_48186);
nand UO_885 (O_885,N_49870,N_48044);
nand UO_886 (O_886,N_49316,N_49981);
nand UO_887 (O_887,N_48903,N_48159);
and UO_888 (O_888,N_48476,N_48736);
and UO_889 (O_889,N_49320,N_48119);
or UO_890 (O_890,N_48417,N_49310);
nand UO_891 (O_891,N_48112,N_48479);
nand UO_892 (O_892,N_48427,N_49078);
or UO_893 (O_893,N_48999,N_48041);
or UO_894 (O_894,N_49748,N_49133);
or UO_895 (O_895,N_48179,N_49369);
nand UO_896 (O_896,N_48380,N_48431);
nor UO_897 (O_897,N_48550,N_48151);
nor UO_898 (O_898,N_49731,N_48758);
nand UO_899 (O_899,N_48001,N_49803);
nor UO_900 (O_900,N_49159,N_49614);
and UO_901 (O_901,N_49006,N_49545);
or UO_902 (O_902,N_48087,N_48565);
nand UO_903 (O_903,N_49176,N_48852);
and UO_904 (O_904,N_49314,N_49309);
nand UO_905 (O_905,N_48109,N_48988);
nor UO_906 (O_906,N_48403,N_48895);
or UO_907 (O_907,N_48270,N_49489);
xor UO_908 (O_908,N_49340,N_49689);
nand UO_909 (O_909,N_48299,N_48462);
or UO_910 (O_910,N_49871,N_48311);
and UO_911 (O_911,N_49409,N_48902);
or UO_912 (O_912,N_48616,N_49608);
or UO_913 (O_913,N_49707,N_49902);
and UO_914 (O_914,N_49156,N_48150);
or UO_915 (O_915,N_48049,N_49122);
nor UO_916 (O_916,N_48578,N_49894);
nor UO_917 (O_917,N_49778,N_48321);
nand UO_918 (O_918,N_48033,N_49274);
nand UO_919 (O_919,N_49648,N_48993);
xnor UO_920 (O_920,N_49457,N_49548);
nand UO_921 (O_921,N_49361,N_48314);
nor UO_922 (O_922,N_48265,N_49698);
nand UO_923 (O_923,N_48996,N_49461);
and UO_924 (O_924,N_49188,N_48148);
nor UO_925 (O_925,N_48722,N_49404);
and UO_926 (O_926,N_49686,N_48976);
nor UO_927 (O_927,N_49852,N_49288);
and UO_928 (O_928,N_49865,N_49128);
nor UO_929 (O_929,N_48773,N_48248);
nor UO_930 (O_930,N_48210,N_48282);
nand UO_931 (O_931,N_48928,N_49131);
nor UO_932 (O_932,N_49432,N_48945);
nand UO_933 (O_933,N_48568,N_48681);
nor UO_934 (O_934,N_48272,N_49452);
nor UO_935 (O_935,N_48367,N_48968);
or UO_936 (O_936,N_49448,N_48904);
nor UO_937 (O_937,N_49337,N_48420);
nor UO_938 (O_938,N_49415,N_48355);
nor UO_939 (O_939,N_49392,N_49720);
nand UO_940 (O_940,N_48197,N_49534);
nor UO_941 (O_941,N_49238,N_48652);
or UO_942 (O_942,N_48690,N_49246);
and UO_943 (O_943,N_48275,N_48021);
and UO_944 (O_944,N_49599,N_49666);
and UO_945 (O_945,N_48434,N_48894);
nor UO_946 (O_946,N_48376,N_49601);
nand UO_947 (O_947,N_48595,N_48234);
and UO_948 (O_948,N_48694,N_49208);
or UO_949 (O_949,N_49802,N_49022);
nor UO_950 (O_950,N_48473,N_48746);
nand UO_951 (O_951,N_49702,N_49171);
nand UO_952 (O_952,N_48015,N_48326);
and UO_953 (O_953,N_48705,N_49479);
and UO_954 (O_954,N_49111,N_49289);
nand UO_955 (O_955,N_49966,N_48610);
xnor UO_956 (O_956,N_49704,N_48984);
or UO_957 (O_957,N_49331,N_48767);
nor UO_958 (O_958,N_49514,N_49959);
and UO_959 (O_959,N_49789,N_48217);
nor UO_960 (O_960,N_48231,N_48859);
and UO_961 (O_961,N_48932,N_48162);
nor UO_962 (O_962,N_49675,N_49439);
and UO_963 (O_963,N_49260,N_48855);
nor UO_964 (O_964,N_48390,N_48117);
nor UO_965 (O_965,N_49771,N_49919);
and UO_966 (O_966,N_48450,N_49896);
nand UO_967 (O_967,N_48191,N_49683);
nand UO_968 (O_968,N_49562,N_48516);
xor UO_969 (O_969,N_49313,N_49296);
or UO_970 (O_970,N_49595,N_48628);
and UO_971 (O_971,N_49690,N_49543);
or UO_972 (O_972,N_49391,N_49636);
and UO_973 (O_973,N_49456,N_49730);
and UO_974 (O_974,N_49193,N_49271);
nor UO_975 (O_975,N_48249,N_49472);
nand UO_976 (O_976,N_49889,N_49945);
and UO_977 (O_977,N_48132,N_49102);
or UO_978 (O_978,N_49400,N_48388);
and UO_979 (O_979,N_48883,N_49302);
nor UO_980 (O_980,N_49892,N_48704);
nand UO_981 (O_981,N_48123,N_48821);
and UO_982 (O_982,N_48795,N_48508);
or UO_983 (O_983,N_48761,N_49825);
nand UO_984 (O_984,N_49722,N_49330);
nand UO_985 (O_985,N_49700,N_49383);
nand UO_986 (O_986,N_48971,N_49443);
nand UO_987 (O_987,N_48405,N_49295);
nand UO_988 (O_988,N_49717,N_49123);
nor UO_989 (O_989,N_48532,N_48443);
and UO_990 (O_990,N_48481,N_49708);
nand UO_991 (O_991,N_48174,N_49504);
nand UO_992 (O_992,N_49394,N_49649);
or UO_993 (O_993,N_48340,N_49146);
and UO_994 (O_994,N_48908,N_49487);
or UO_995 (O_995,N_49909,N_49346);
or UO_996 (O_996,N_49143,N_49576);
and UO_997 (O_997,N_49915,N_48592);
or UO_998 (O_998,N_49736,N_49561);
xnor UO_999 (O_999,N_48219,N_48778);
and UO_1000 (O_1000,N_49883,N_48109);
or UO_1001 (O_1001,N_48632,N_48160);
nand UO_1002 (O_1002,N_48025,N_48356);
or UO_1003 (O_1003,N_48971,N_49328);
nand UO_1004 (O_1004,N_48854,N_49165);
nor UO_1005 (O_1005,N_49218,N_49413);
or UO_1006 (O_1006,N_49065,N_49357);
and UO_1007 (O_1007,N_49204,N_49747);
or UO_1008 (O_1008,N_49435,N_49588);
or UO_1009 (O_1009,N_49871,N_48640);
or UO_1010 (O_1010,N_49922,N_48618);
nor UO_1011 (O_1011,N_48290,N_49144);
nor UO_1012 (O_1012,N_49608,N_48329);
or UO_1013 (O_1013,N_49297,N_49595);
and UO_1014 (O_1014,N_48897,N_49290);
nor UO_1015 (O_1015,N_48450,N_48605);
or UO_1016 (O_1016,N_48730,N_49037);
or UO_1017 (O_1017,N_49997,N_48279);
nand UO_1018 (O_1018,N_48165,N_48107);
nand UO_1019 (O_1019,N_48496,N_48550);
or UO_1020 (O_1020,N_49483,N_48540);
or UO_1021 (O_1021,N_48250,N_49351);
nor UO_1022 (O_1022,N_49240,N_49551);
nand UO_1023 (O_1023,N_49107,N_49489);
nand UO_1024 (O_1024,N_49012,N_48363);
and UO_1025 (O_1025,N_48111,N_48541);
or UO_1026 (O_1026,N_49966,N_49960);
and UO_1027 (O_1027,N_48078,N_49720);
and UO_1028 (O_1028,N_48912,N_49231);
nor UO_1029 (O_1029,N_49060,N_49204);
nand UO_1030 (O_1030,N_48635,N_49179);
nor UO_1031 (O_1031,N_49022,N_48914);
xor UO_1032 (O_1032,N_48650,N_49654);
nand UO_1033 (O_1033,N_49720,N_48071);
nor UO_1034 (O_1034,N_48360,N_49687);
nand UO_1035 (O_1035,N_49343,N_49928);
or UO_1036 (O_1036,N_49490,N_48429);
or UO_1037 (O_1037,N_49550,N_48072);
nor UO_1038 (O_1038,N_49928,N_49235);
or UO_1039 (O_1039,N_49630,N_48280);
or UO_1040 (O_1040,N_48279,N_49156);
or UO_1041 (O_1041,N_49305,N_48973);
and UO_1042 (O_1042,N_49995,N_48097);
and UO_1043 (O_1043,N_49024,N_49799);
and UO_1044 (O_1044,N_48217,N_49977);
nor UO_1045 (O_1045,N_48605,N_48041);
nand UO_1046 (O_1046,N_48867,N_48657);
nand UO_1047 (O_1047,N_48547,N_49214);
and UO_1048 (O_1048,N_49813,N_49691);
nor UO_1049 (O_1049,N_49063,N_49008);
or UO_1050 (O_1050,N_49578,N_49752);
nor UO_1051 (O_1051,N_49471,N_49148);
or UO_1052 (O_1052,N_49652,N_48813);
nand UO_1053 (O_1053,N_49255,N_48889);
nand UO_1054 (O_1054,N_49554,N_48183);
or UO_1055 (O_1055,N_48172,N_48103);
nand UO_1056 (O_1056,N_48216,N_48859);
nand UO_1057 (O_1057,N_48071,N_49245);
nand UO_1058 (O_1058,N_48975,N_49203);
or UO_1059 (O_1059,N_49857,N_48125);
and UO_1060 (O_1060,N_49062,N_48842);
nor UO_1061 (O_1061,N_48874,N_48270);
and UO_1062 (O_1062,N_49102,N_48943);
nor UO_1063 (O_1063,N_49317,N_49279);
nor UO_1064 (O_1064,N_48492,N_49931);
or UO_1065 (O_1065,N_49738,N_48774);
nand UO_1066 (O_1066,N_49171,N_49413);
and UO_1067 (O_1067,N_49033,N_48144);
nor UO_1068 (O_1068,N_49486,N_48606);
or UO_1069 (O_1069,N_48442,N_48935);
and UO_1070 (O_1070,N_49606,N_49960);
or UO_1071 (O_1071,N_49860,N_48168);
or UO_1072 (O_1072,N_49322,N_49084);
nand UO_1073 (O_1073,N_49632,N_49635);
or UO_1074 (O_1074,N_49208,N_49646);
and UO_1075 (O_1075,N_49954,N_49090);
and UO_1076 (O_1076,N_48934,N_49074);
nand UO_1077 (O_1077,N_49416,N_48177);
and UO_1078 (O_1078,N_49229,N_49565);
or UO_1079 (O_1079,N_48229,N_48544);
or UO_1080 (O_1080,N_48828,N_48841);
nor UO_1081 (O_1081,N_48094,N_48390);
or UO_1082 (O_1082,N_48394,N_49384);
and UO_1083 (O_1083,N_49078,N_48913);
or UO_1084 (O_1084,N_49375,N_48434);
nor UO_1085 (O_1085,N_49174,N_49977);
and UO_1086 (O_1086,N_49950,N_48486);
nand UO_1087 (O_1087,N_48216,N_49772);
nor UO_1088 (O_1088,N_49183,N_49883);
nand UO_1089 (O_1089,N_48504,N_48731);
nor UO_1090 (O_1090,N_48412,N_48479);
and UO_1091 (O_1091,N_48317,N_49309);
or UO_1092 (O_1092,N_48297,N_49775);
nand UO_1093 (O_1093,N_48762,N_49703);
and UO_1094 (O_1094,N_49433,N_49051);
or UO_1095 (O_1095,N_49937,N_49565);
or UO_1096 (O_1096,N_48735,N_49378);
or UO_1097 (O_1097,N_49223,N_49735);
or UO_1098 (O_1098,N_49839,N_49401);
nand UO_1099 (O_1099,N_49019,N_49749);
nor UO_1100 (O_1100,N_48587,N_49533);
and UO_1101 (O_1101,N_48109,N_49811);
or UO_1102 (O_1102,N_48798,N_48882);
or UO_1103 (O_1103,N_48710,N_48400);
nand UO_1104 (O_1104,N_49330,N_48991);
nor UO_1105 (O_1105,N_49577,N_48200);
nor UO_1106 (O_1106,N_48515,N_48379);
nand UO_1107 (O_1107,N_48147,N_48819);
or UO_1108 (O_1108,N_49799,N_48804);
and UO_1109 (O_1109,N_48510,N_48022);
nor UO_1110 (O_1110,N_48984,N_48930);
nand UO_1111 (O_1111,N_49281,N_48263);
nand UO_1112 (O_1112,N_48726,N_48190);
or UO_1113 (O_1113,N_49620,N_49612);
and UO_1114 (O_1114,N_49781,N_48525);
nand UO_1115 (O_1115,N_49279,N_48380);
nand UO_1116 (O_1116,N_48385,N_49856);
or UO_1117 (O_1117,N_49523,N_48334);
and UO_1118 (O_1118,N_48282,N_48251);
nor UO_1119 (O_1119,N_49304,N_49174);
and UO_1120 (O_1120,N_49286,N_48110);
nor UO_1121 (O_1121,N_48727,N_48483);
nor UO_1122 (O_1122,N_49742,N_49514);
and UO_1123 (O_1123,N_48293,N_49583);
and UO_1124 (O_1124,N_48760,N_49178);
nand UO_1125 (O_1125,N_48401,N_49999);
nor UO_1126 (O_1126,N_49052,N_49042);
nor UO_1127 (O_1127,N_48297,N_49908);
or UO_1128 (O_1128,N_48067,N_48435);
nor UO_1129 (O_1129,N_48159,N_49441);
and UO_1130 (O_1130,N_49968,N_48226);
nand UO_1131 (O_1131,N_49083,N_49288);
xnor UO_1132 (O_1132,N_49631,N_48430);
or UO_1133 (O_1133,N_48860,N_49038);
nand UO_1134 (O_1134,N_48224,N_48755);
or UO_1135 (O_1135,N_49936,N_49015);
nor UO_1136 (O_1136,N_49559,N_49729);
nor UO_1137 (O_1137,N_48079,N_48224);
nor UO_1138 (O_1138,N_48740,N_49659);
and UO_1139 (O_1139,N_49161,N_48087);
or UO_1140 (O_1140,N_48546,N_49769);
nand UO_1141 (O_1141,N_48788,N_48093);
and UO_1142 (O_1142,N_49680,N_48702);
and UO_1143 (O_1143,N_48091,N_48718);
and UO_1144 (O_1144,N_49666,N_49849);
nor UO_1145 (O_1145,N_48691,N_49808);
and UO_1146 (O_1146,N_48267,N_48848);
nor UO_1147 (O_1147,N_49223,N_49684);
nor UO_1148 (O_1148,N_49290,N_49955);
nor UO_1149 (O_1149,N_49187,N_49066);
and UO_1150 (O_1150,N_48302,N_49106);
nor UO_1151 (O_1151,N_49704,N_49629);
and UO_1152 (O_1152,N_48254,N_49076);
and UO_1153 (O_1153,N_49064,N_48120);
nand UO_1154 (O_1154,N_48018,N_48739);
nor UO_1155 (O_1155,N_49911,N_49389);
and UO_1156 (O_1156,N_48264,N_49202);
nor UO_1157 (O_1157,N_48152,N_49109);
xor UO_1158 (O_1158,N_48194,N_48722);
and UO_1159 (O_1159,N_49429,N_48278);
nand UO_1160 (O_1160,N_48410,N_49838);
nor UO_1161 (O_1161,N_48662,N_48468);
and UO_1162 (O_1162,N_48482,N_49473);
nand UO_1163 (O_1163,N_49462,N_49080);
nor UO_1164 (O_1164,N_49383,N_48263);
nand UO_1165 (O_1165,N_48814,N_48379);
and UO_1166 (O_1166,N_48051,N_48311);
nor UO_1167 (O_1167,N_49206,N_48613);
nand UO_1168 (O_1168,N_48403,N_48779);
xor UO_1169 (O_1169,N_49777,N_48442);
nand UO_1170 (O_1170,N_48572,N_49639);
nor UO_1171 (O_1171,N_49092,N_49295);
nand UO_1172 (O_1172,N_48207,N_49379);
nand UO_1173 (O_1173,N_48404,N_49008);
and UO_1174 (O_1174,N_49023,N_49371);
nor UO_1175 (O_1175,N_49593,N_49863);
or UO_1176 (O_1176,N_48143,N_49107);
and UO_1177 (O_1177,N_49095,N_48470);
nor UO_1178 (O_1178,N_49139,N_48888);
or UO_1179 (O_1179,N_48062,N_48430);
or UO_1180 (O_1180,N_48161,N_49929);
and UO_1181 (O_1181,N_48113,N_49514);
or UO_1182 (O_1182,N_49258,N_49724);
nand UO_1183 (O_1183,N_48151,N_48783);
nand UO_1184 (O_1184,N_49603,N_49737);
or UO_1185 (O_1185,N_49391,N_48153);
nand UO_1186 (O_1186,N_49179,N_49170);
nand UO_1187 (O_1187,N_49844,N_49006);
nand UO_1188 (O_1188,N_48312,N_49154);
nor UO_1189 (O_1189,N_49247,N_48471);
and UO_1190 (O_1190,N_49738,N_48402);
and UO_1191 (O_1191,N_49667,N_49211);
nand UO_1192 (O_1192,N_49969,N_49670);
or UO_1193 (O_1193,N_49604,N_48610);
nand UO_1194 (O_1194,N_48287,N_48749);
nor UO_1195 (O_1195,N_49969,N_49952);
nor UO_1196 (O_1196,N_48200,N_48331);
nor UO_1197 (O_1197,N_49479,N_49865);
nand UO_1198 (O_1198,N_48814,N_49039);
or UO_1199 (O_1199,N_48076,N_48659);
or UO_1200 (O_1200,N_49877,N_49017);
nor UO_1201 (O_1201,N_48057,N_49937);
nor UO_1202 (O_1202,N_49114,N_48179);
nor UO_1203 (O_1203,N_49796,N_48220);
and UO_1204 (O_1204,N_49097,N_49266);
and UO_1205 (O_1205,N_48223,N_48047);
or UO_1206 (O_1206,N_48395,N_48733);
and UO_1207 (O_1207,N_48656,N_48449);
and UO_1208 (O_1208,N_48620,N_49820);
or UO_1209 (O_1209,N_48676,N_48353);
nor UO_1210 (O_1210,N_48166,N_48123);
nor UO_1211 (O_1211,N_48757,N_48077);
nand UO_1212 (O_1212,N_48005,N_49349);
or UO_1213 (O_1213,N_49995,N_48439);
nand UO_1214 (O_1214,N_48222,N_49568);
nor UO_1215 (O_1215,N_48041,N_48610);
xor UO_1216 (O_1216,N_48852,N_49592);
nand UO_1217 (O_1217,N_48737,N_49891);
nor UO_1218 (O_1218,N_48518,N_49550);
nor UO_1219 (O_1219,N_49220,N_49048);
nand UO_1220 (O_1220,N_48347,N_48948);
nor UO_1221 (O_1221,N_49775,N_49109);
nor UO_1222 (O_1222,N_49630,N_48862);
or UO_1223 (O_1223,N_48053,N_49340);
or UO_1224 (O_1224,N_49164,N_48321);
and UO_1225 (O_1225,N_48617,N_49948);
nor UO_1226 (O_1226,N_49776,N_48826);
and UO_1227 (O_1227,N_49766,N_48518);
and UO_1228 (O_1228,N_48426,N_48921);
nor UO_1229 (O_1229,N_48534,N_48528);
nor UO_1230 (O_1230,N_48697,N_48752);
or UO_1231 (O_1231,N_48435,N_49815);
and UO_1232 (O_1232,N_48242,N_48471);
nor UO_1233 (O_1233,N_48676,N_49152);
nor UO_1234 (O_1234,N_48589,N_48236);
and UO_1235 (O_1235,N_49697,N_48346);
nand UO_1236 (O_1236,N_49662,N_48405);
nand UO_1237 (O_1237,N_48962,N_49374);
and UO_1238 (O_1238,N_49593,N_48281);
or UO_1239 (O_1239,N_49177,N_49981);
and UO_1240 (O_1240,N_48981,N_49780);
nand UO_1241 (O_1241,N_48124,N_48791);
or UO_1242 (O_1242,N_49579,N_48846);
and UO_1243 (O_1243,N_49230,N_48039);
nor UO_1244 (O_1244,N_48155,N_49773);
nor UO_1245 (O_1245,N_48294,N_49966);
nor UO_1246 (O_1246,N_49935,N_49380);
nor UO_1247 (O_1247,N_49374,N_49469);
nand UO_1248 (O_1248,N_49700,N_49769);
nand UO_1249 (O_1249,N_49262,N_49935);
and UO_1250 (O_1250,N_48704,N_48021);
nand UO_1251 (O_1251,N_49664,N_48309);
and UO_1252 (O_1252,N_49531,N_49640);
nor UO_1253 (O_1253,N_49868,N_48152);
or UO_1254 (O_1254,N_48356,N_48009);
nand UO_1255 (O_1255,N_49824,N_49642);
and UO_1256 (O_1256,N_49056,N_49422);
or UO_1257 (O_1257,N_48210,N_49959);
or UO_1258 (O_1258,N_48077,N_48015);
or UO_1259 (O_1259,N_48419,N_48750);
and UO_1260 (O_1260,N_48825,N_49161);
or UO_1261 (O_1261,N_48563,N_49766);
nor UO_1262 (O_1262,N_48209,N_49253);
nand UO_1263 (O_1263,N_49750,N_48881);
xnor UO_1264 (O_1264,N_48521,N_49584);
nand UO_1265 (O_1265,N_49900,N_48919);
nand UO_1266 (O_1266,N_49675,N_49134);
nor UO_1267 (O_1267,N_48862,N_48955);
nand UO_1268 (O_1268,N_49384,N_49118);
and UO_1269 (O_1269,N_48040,N_48649);
and UO_1270 (O_1270,N_48095,N_49559);
nand UO_1271 (O_1271,N_48194,N_49789);
xnor UO_1272 (O_1272,N_49875,N_49627);
or UO_1273 (O_1273,N_48647,N_49005);
xnor UO_1274 (O_1274,N_48615,N_48645);
and UO_1275 (O_1275,N_48139,N_48565);
nor UO_1276 (O_1276,N_49625,N_48196);
nor UO_1277 (O_1277,N_49041,N_49193);
and UO_1278 (O_1278,N_48008,N_49935);
nor UO_1279 (O_1279,N_48942,N_49736);
and UO_1280 (O_1280,N_48254,N_49900);
and UO_1281 (O_1281,N_48867,N_48023);
nor UO_1282 (O_1282,N_49389,N_48847);
and UO_1283 (O_1283,N_48845,N_48088);
nor UO_1284 (O_1284,N_48048,N_49716);
nand UO_1285 (O_1285,N_49499,N_48172);
and UO_1286 (O_1286,N_48232,N_48947);
and UO_1287 (O_1287,N_48270,N_49245);
and UO_1288 (O_1288,N_48003,N_48735);
and UO_1289 (O_1289,N_48122,N_49946);
nand UO_1290 (O_1290,N_48318,N_49008);
nor UO_1291 (O_1291,N_49965,N_48078);
or UO_1292 (O_1292,N_49185,N_49485);
and UO_1293 (O_1293,N_49389,N_48353);
nand UO_1294 (O_1294,N_49847,N_49082);
nand UO_1295 (O_1295,N_49132,N_49304);
nor UO_1296 (O_1296,N_48989,N_49563);
nor UO_1297 (O_1297,N_48085,N_49470);
and UO_1298 (O_1298,N_49784,N_49045);
and UO_1299 (O_1299,N_49191,N_48403);
or UO_1300 (O_1300,N_48291,N_49458);
or UO_1301 (O_1301,N_48234,N_48732);
or UO_1302 (O_1302,N_49709,N_48577);
and UO_1303 (O_1303,N_49269,N_49189);
nand UO_1304 (O_1304,N_48596,N_49157);
or UO_1305 (O_1305,N_49212,N_48224);
nand UO_1306 (O_1306,N_48501,N_49991);
or UO_1307 (O_1307,N_49270,N_49875);
nor UO_1308 (O_1308,N_49579,N_48377);
nor UO_1309 (O_1309,N_48515,N_48794);
nor UO_1310 (O_1310,N_49920,N_48164);
and UO_1311 (O_1311,N_48527,N_48430);
nor UO_1312 (O_1312,N_48201,N_49024);
nor UO_1313 (O_1313,N_49761,N_48960);
nor UO_1314 (O_1314,N_49331,N_48652);
nand UO_1315 (O_1315,N_49086,N_49421);
and UO_1316 (O_1316,N_49454,N_49168);
nand UO_1317 (O_1317,N_49436,N_49597);
or UO_1318 (O_1318,N_48630,N_49676);
nor UO_1319 (O_1319,N_48188,N_49346);
nand UO_1320 (O_1320,N_49085,N_49669);
nand UO_1321 (O_1321,N_48920,N_49592);
or UO_1322 (O_1322,N_48624,N_49033);
nor UO_1323 (O_1323,N_49743,N_49351);
and UO_1324 (O_1324,N_49730,N_49510);
and UO_1325 (O_1325,N_48262,N_48507);
nand UO_1326 (O_1326,N_48931,N_49599);
nor UO_1327 (O_1327,N_48937,N_49155);
nand UO_1328 (O_1328,N_48664,N_49886);
nor UO_1329 (O_1329,N_48325,N_48297);
or UO_1330 (O_1330,N_49621,N_49213);
or UO_1331 (O_1331,N_49338,N_49763);
nor UO_1332 (O_1332,N_48565,N_49837);
xor UO_1333 (O_1333,N_49465,N_49888);
or UO_1334 (O_1334,N_48059,N_49586);
nand UO_1335 (O_1335,N_48869,N_48187);
and UO_1336 (O_1336,N_49367,N_49659);
and UO_1337 (O_1337,N_49370,N_49628);
nor UO_1338 (O_1338,N_48537,N_49309);
and UO_1339 (O_1339,N_49239,N_49193);
nor UO_1340 (O_1340,N_49070,N_49351);
nor UO_1341 (O_1341,N_48141,N_49611);
and UO_1342 (O_1342,N_49860,N_48318);
nor UO_1343 (O_1343,N_48025,N_49998);
nor UO_1344 (O_1344,N_49091,N_48583);
nand UO_1345 (O_1345,N_49295,N_48108);
and UO_1346 (O_1346,N_49772,N_48021);
nand UO_1347 (O_1347,N_49035,N_49947);
nor UO_1348 (O_1348,N_48902,N_49786);
and UO_1349 (O_1349,N_48480,N_49955);
and UO_1350 (O_1350,N_49482,N_49531);
nand UO_1351 (O_1351,N_49109,N_49071);
nor UO_1352 (O_1352,N_49176,N_48517);
nand UO_1353 (O_1353,N_48657,N_49028);
nor UO_1354 (O_1354,N_48815,N_48681);
or UO_1355 (O_1355,N_48189,N_48975);
nor UO_1356 (O_1356,N_48827,N_49190);
or UO_1357 (O_1357,N_49032,N_49708);
and UO_1358 (O_1358,N_48484,N_48628);
or UO_1359 (O_1359,N_48527,N_49743);
or UO_1360 (O_1360,N_49942,N_49828);
and UO_1361 (O_1361,N_49669,N_49839);
or UO_1362 (O_1362,N_49932,N_49927);
nand UO_1363 (O_1363,N_48207,N_48463);
nand UO_1364 (O_1364,N_48432,N_49785);
and UO_1365 (O_1365,N_49052,N_48567);
or UO_1366 (O_1366,N_49485,N_49821);
and UO_1367 (O_1367,N_48531,N_49190);
nand UO_1368 (O_1368,N_49766,N_49643);
nor UO_1369 (O_1369,N_49572,N_48669);
nor UO_1370 (O_1370,N_48311,N_49656);
nand UO_1371 (O_1371,N_48696,N_48300);
and UO_1372 (O_1372,N_49705,N_49872);
nor UO_1373 (O_1373,N_49158,N_48323);
nor UO_1374 (O_1374,N_49774,N_48354);
or UO_1375 (O_1375,N_48215,N_49404);
nor UO_1376 (O_1376,N_48396,N_49125);
and UO_1377 (O_1377,N_49031,N_49026);
and UO_1378 (O_1378,N_49087,N_49080);
nor UO_1379 (O_1379,N_48976,N_49881);
nor UO_1380 (O_1380,N_48903,N_48085);
and UO_1381 (O_1381,N_48543,N_48021);
nor UO_1382 (O_1382,N_49301,N_48728);
and UO_1383 (O_1383,N_49815,N_49276);
nor UO_1384 (O_1384,N_49363,N_48263);
and UO_1385 (O_1385,N_49636,N_49464);
and UO_1386 (O_1386,N_48189,N_48074);
nor UO_1387 (O_1387,N_48432,N_49302);
nand UO_1388 (O_1388,N_49859,N_49887);
nor UO_1389 (O_1389,N_49916,N_48546);
or UO_1390 (O_1390,N_49045,N_49875);
nor UO_1391 (O_1391,N_49299,N_49583);
or UO_1392 (O_1392,N_48827,N_48899);
nor UO_1393 (O_1393,N_49063,N_49988);
or UO_1394 (O_1394,N_49926,N_49772);
or UO_1395 (O_1395,N_48356,N_49428);
or UO_1396 (O_1396,N_49167,N_48632);
and UO_1397 (O_1397,N_48142,N_48941);
nor UO_1398 (O_1398,N_49845,N_48357);
nand UO_1399 (O_1399,N_48050,N_49876);
nor UO_1400 (O_1400,N_48628,N_49804);
nand UO_1401 (O_1401,N_48021,N_49441);
and UO_1402 (O_1402,N_48305,N_49211);
or UO_1403 (O_1403,N_48451,N_48834);
and UO_1404 (O_1404,N_48356,N_49586);
xor UO_1405 (O_1405,N_48683,N_49947);
and UO_1406 (O_1406,N_49957,N_49484);
nor UO_1407 (O_1407,N_49631,N_49336);
nor UO_1408 (O_1408,N_49374,N_48900);
and UO_1409 (O_1409,N_48541,N_48154);
or UO_1410 (O_1410,N_48180,N_49131);
or UO_1411 (O_1411,N_49865,N_49207);
nand UO_1412 (O_1412,N_49949,N_48752);
nand UO_1413 (O_1413,N_48875,N_49746);
and UO_1414 (O_1414,N_49011,N_48422);
nand UO_1415 (O_1415,N_49984,N_49897);
and UO_1416 (O_1416,N_48727,N_48460);
nor UO_1417 (O_1417,N_49678,N_49790);
nand UO_1418 (O_1418,N_49965,N_49561);
xor UO_1419 (O_1419,N_49870,N_48692);
or UO_1420 (O_1420,N_48532,N_49416);
nand UO_1421 (O_1421,N_49575,N_49857);
nand UO_1422 (O_1422,N_49473,N_48514);
nand UO_1423 (O_1423,N_48437,N_49042);
and UO_1424 (O_1424,N_48015,N_49851);
nand UO_1425 (O_1425,N_49482,N_49321);
nand UO_1426 (O_1426,N_48746,N_49373);
and UO_1427 (O_1427,N_49405,N_49462);
nor UO_1428 (O_1428,N_49016,N_48956);
nor UO_1429 (O_1429,N_49508,N_48766);
nand UO_1430 (O_1430,N_49510,N_49197);
or UO_1431 (O_1431,N_48864,N_49995);
and UO_1432 (O_1432,N_49960,N_49368);
nand UO_1433 (O_1433,N_49754,N_49599);
and UO_1434 (O_1434,N_48948,N_49169);
nor UO_1435 (O_1435,N_49235,N_48729);
xnor UO_1436 (O_1436,N_48185,N_49830);
nor UO_1437 (O_1437,N_48734,N_49806);
and UO_1438 (O_1438,N_48443,N_48188);
nand UO_1439 (O_1439,N_48828,N_49668);
nor UO_1440 (O_1440,N_49595,N_49319);
or UO_1441 (O_1441,N_49710,N_48137);
nor UO_1442 (O_1442,N_48094,N_49923);
nor UO_1443 (O_1443,N_49250,N_48126);
nor UO_1444 (O_1444,N_49122,N_48951);
and UO_1445 (O_1445,N_49560,N_49157);
and UO_1446 (O_1446,N_49393,N_48830);
nor UO_1447 (O_1447,N_48152,N_49885);
nor UO_1448 (O_1448,N_49019,N_48646);
xnor UO_1449 (O_1449,N_48397,N_49399);
and UO_1450 (O_1450,N_48638,N_49218);
nand UO_1451 (O_1451,N_48298,N_49640);
nand UO_1452 (O_1452,N_48886,N_49660);
nand UO_1453 (O_1453,N_48037,N_49115);
nor UO_1454 (O_1454,N_49247,N_48525);
and UO_1455 (O_1455,N_48897,N_48334);
and UO_1456 (O_1456,N_48452,N_48062);
nand UO_1457 (O_1457,N_49628,N_49793);
and UO_1458 (O_1458,N_48396,N_49718);
nand UO_1459 (O_1459,N_48771,N_48730);
xnor UO_1460 (O_1460,N_48338,N_49139);
and UO_1461 (O_1461,N_49841,N_49578);
and UO_1462 (O_1462,N_48723,N_48128);
or UO_1463 (O_1463,N_49642,N_49940);
and UO_1464 (O_1464,N_49102,N_48340);
and UO_1465 (O_1465,N_48702,N_48066);
and UO_1466 (O_1466,N_48806,N_49485);
nand UO_1467 (O_1467,N_49137,N_49738);
nand UO_1468 (O_1468,N_48079,N_49580);
or UO_1469 (O_1469,N_48912,N_48909);
nand UO_1470 (O_1470,N_49877,N_49662);
nand UO_1471 (O_1471,N_48885,N_48678);
nand UO_1472 (O_1472,N_48658,N_49079);
nor UO_1473 (O_1473,N_48725,N_49128);
nor UO_1474 (O_1474,N_49459,N_49896);
or UO_1475 (O_1475,N_49688,N_48557);
nor UO_1476 (O_1476,N_48759,N_49846);
nand UO_1477 (O_1477,N_49114,N_49767);
and UO_1478 (O_1478,N_48040,N_49006);
nand UO_1479 (O_1479,N_48736,N_49620);
nor UO_1480 (O_1480,N_48869,N_48666);
or UO_1481 (O_1481,N_48620,N_49258);
nand UO_1482 (O_1482,N_48185,N_49340);
and UO_1483 (O_1483,N_49776,N_48828);
or UO_1484 (O_1484,N_49760,N_48004);
nand UO_1485 (O_1485,N_49708,N_48602);
nand UO_1486 (O_1486,N_49854,N_48956);
and UO_1487 (O_1487,N_49537,N_48769);
or UO_1488 (O_1488,N_48019,N_48472);
and UO_1489 (O_1489,N_49782,N_48106);
and UO_1490 (O_1490,N_49567,N_49820);
nor UO_1491 (O_1491,N_48551,N_49977);
nor UO_1492 (O_1492,N_49399,N_49048);
and UO_1493 (O_1493,N_49677,N_48408);
nor UO_1494 (O_1494,N_48010,N_49481);
or UO_1495 (O_1495,N_48038,N_49066);
and UO_1496 (O_1496,N_49496,N_49988);
or UO_1497 (O_1497,N_49587,N_49037);
nand UO_1498 (O_1498,N_48528,N_48938);
xor UO_1499 (O_1499,N_48023,N_48494);
and UO_1500 (O_1500,N_49044,N_48860);
and UO_1501 (O_1501,N_49307,N_48099);
nand UO_1502 (O_1502,N_48584,N_49764);
nand UO_1503 (O_1503,N_48658,N_49140);
nor UO_1504 (O_1504,N_49680,N_49265);
and UO_1505 (O_1505,N_49185,N_48614);
and UO_1506 (O_1506,N_49507,N_49820);
or UO_1507 (O_1507,N_48940,N_49379);
nand UO_1508 (O_1508,N_48627,N_49364);
nand UO_1509 (O_1509,N_49570,N_49009);
nor UO_1510 (O_1510,N_48907,N_49928);
nand UO_1511 (O_1511,N_48886,N_49493);
nand UO_1512 (O_1512,N_48909,N_49113);
nor UO_1513 (O_1513,N_49216,N_48126);
nor UO_1514 (O_1514,N_48551,N_48832);
and UO_1515 (O_1515,N_49909,N_48260);
or UO_1516 (O_1516,N_48953,N_49511);
or UO_1517 (O_1517,N_48758,N_48325);
and UO_1518 (O_1518,N_48881,N_48170);
or UO_1519 (O_1519,N_48454,N_49478);
or UO_1520 (O_1520,N_49650,N_48848);
and UO_1521 (O_1521,N_49382,N_48426);
nand UO_1522 (O_1522,N_48152,N_48730);
or UO_1523 (O_1523,N_49390,N_48765);
or UO_1524 (O_1524,N_49357,N_49304);
nor UO_1525 (O_1525,N_48862,N_49524);
nor UO_1526 (O_1526,N_49220,N_48416);
and UO_1527 (O_1527,N_49642,N_48911);
nor UO_1528 (O_1528,N_48714,N_49347);
nand UO_1529 (O_1529,N_49974,N_48651);
nand UO_1530 (O_1530,N_48475,N_48131);
nand UO_1531 (O_1531,N_49232,N_49427);
nor UO_1532 (O_1532,N_49574,N_48344);
nand UO_1533 (O_1533,N_49968,N_49963);
nor UO_1534 (O_1534,N_48896,N_49844);
or UO_1535 (O_1535,N_48478,N_49740);
nor UO_1536 (O_1536,N_48032,N_48855);
or UO_1537 (O_1537,N_48901,N_49501);
nand UO_1538 (O_1538,N_49464,N_49325);
nor UO_1539 (O_1539,N_48986,N_48976);
nand UO_1540 (O_1540,N_49017,N_48762);
nand UO_1541 (O_1541,N_49261,N_48822);
or UO_1542 (O_1542,N_48960,N_48302);
nor UO_1543 (O_1543,N_49659,N_49498);
and UO_1544 (O_1544,N_49438,N_48147);
or UO_1545 (O_1545,N_48470,N_49657);
nor UO_1546 (O_1546,N_48221,N_48759);
nor UO_1547 (O_1547,N_48453,N_49947);
and UO_1548 (O_1548,N_48192,N_48791);
or UO_1549 (O_1549,N_49250,N_49023);
or UO_1550 (O_1550,N_48534,N_49328);
nand UO_1551 (O_1551,N_49885,N_49433);
nor UO_1552 (O_1552,N_49270,N_48004);
nand UO_1553 (O_1553,N_49966,N_48633);
or UO_1554 (O_1554,N_48683,N_48382);
and UO_1555 (O_1555,N_49657,N_49941);
and UO_1556 (O_1556,N_49143,N_49029);
or UO_1557 (O_1557,N_48934,N_49530);
and UO_1558 (O_1558,N_49472,N_49324);
nand UO_1559 (O_1559,N_48012,N_49210);
nor UO_1560 (O_1560,N_48734,N_48356);
or UO_1561 (O_1561,N_48832,N_49684);
nor UO_1562 (O_1562,N_48384,N_49278);
nand UO_1563 (O_1563,N_48296,N_48817);
and UO_1564 (O_1564,N_48918,N_48937);
nand UO_1565 (O_1565,N_49570,N_48482);
and UO_1566 (O_1566,N_48697,N_49861);
nor UO_1567 (O_1567,N_48561,N_48722);
nand UO_1568 (O_1568,N_48524,N_48788);
and UO_1569 (O_1569,N_48504,N_48040);
and UO_1570 (O_1570,N_48336,N_49594);
nand UO_1571 (O_1571,N_48689,N_49009);
and UO_1572 (O_1572,N_49303,N_49753);
nor UO_1573 (O_1573,N_49437,N_48077);
and UO_1574 (O_1574,N_49067,N_49008);
nand UO_1575 (O_1575,N_49332,N_49938);
nor UO_1576 (O_1576,N_49187,N_49466);
and UO_1577 (O_1577,N_48535,N_48683);
nor UO_1578 (O_1578,N_49512,N_49740);
and UO_1579 (O_1579,N_48555,N_48581);
nand UO_1580 (O_1580,N_48380,N_49968);
nor UO_1581 (O_1581,N_48207,N_49401);
and UO_1582 (O_1582,N_48263,N_49208);
nor UO_1583 (O_1583,N_49001,N_49143);
nor UO_1584 (O_1584,N_48919,N_48415);
or UO_1585 (O_1585,N_49757,N_48209);
or UO_1586 (O_1586,N_48671,N_48329);
nor UO_1587 (O_1587,N_49439,N_49265);
nand UO_1588 (O_1588,N_48924,N_49301);
or UO_1589 (O_1589,N_49080,N_48957);
nor UO_1590 (O_1590,N_49094,N_49076);
nand UO_1591 (O_1591,N_49106,N_48254);
nor UO_1592 (O_1592,N_48296,N_48291);
nor UO_1593 (O_1593,N_48638,N_49976);
nand UO_1594 (O_1594,N_48994,N_49071);
or UO_1595 (O_1595,N_48870,N_49755);
or UO_1596 (O_1596,N_49874,N_48762);
nand UO_1597 (O_1597,N_48973,N_48360);
or UO_1598 (O_1598,N_49263,N_48496);
nor UO_1599 (O_1599,N_48012,N_49030);
nand UO_1600 (O_1600,N_48284,N_48542);
or UO_1601 (O_1601,N_48030,N_49989);
or UO_1602 (O_1602,N_49725,N_48396);
nand UO_1603 (O_1603,N_49222,N_49586);
nor UO_1604 (O_1604,N_48000,N_48078);
nand UO_1605 (O_1605,N_48216,N_48653);
nand UO_1606 (O_1606,N_48590,N_48492);
nor UO_1607 (O_1607,N_48659,N_48752);
and UO_1608 (O_1608,N_48153,N_48875);
nand UO_1609 (O_1609,N_48396,N_49876);
nand UO_1610 (O_1610,N_49879,N_49128);
nor UO_1611 (O_1611,N_48763,N_49814);
nor UO_1612 (O_1612,N_48506,N_48234);
or UO_1613 (O_1613,N_48973,N_48847);
nand UO_1614 (O_1614,N_48771,N_49291);
nand UO_1615 (O_1615,N_48798,N_49935);
or UO_1616 (O_1616,N_49015,N_49636);
xor UO_1617 (O_1617,N_49865,N_48986);
and UO_1618 (O_1618,N_48451,N_48525);
or UO_1619 (O_1619,N_49102,N_49321);
and UO_1620 (O_1620,N_49861,N_49500);
xor UO_1621 (O_1621,N_48880,N_49633);
or UO_1622 (O_1622,N_49587,N_48452);
or UO_1623 (O_1623,N_48241,N_48820);
nor UO_1624 (O_1624,N_49043,N_49948);
nand UO_1625 (O_1625,N_49743,N_49575);
and UO_1626 (O_1626,N_48818,N_49969);
and UO_1627 (O_1627,N_48141,N_49479);
nor UO_1628 (O_1628,N_49684,N_48001);
or UO_1629 (O_1629,N_49356,N_48392);
and UO_1630 (O_1630,N_48809,N_49306);
nand UO_1631 (O_1631,N_48490,N_48940);
and UO_1632 (O_1632,N_49177,N_49401);
or UO_1633 (O_1633,N_48451,N_48791);
and UO_1634 (O_1634,N_48425,N_49574);
nor UO_1635 (O_1635,N_48620,N_49806);
or UO_1636 (O_1636,N_49646,N_49457);
or UO_1637 (O_1637,N_49608,N_48546);
xnor UO_1638 (O_1638,N_48572,N_49236);
nor UO_1639 (O_1639,N_48768,N_48035);
nand UO_1640 (O_1640,N_49440,N_49428);
nor UO_1641 (O_1641,N_48431,N_48353);
and UO_1642 (O_1642,N_48077,N_49220);
nand UO_1643 (O_1643,N_49945,N_49372);
or UO_1644 (O_1644,N_48871,N_49158);
or UO_1645 (O_1645,N_48227,N_48995);
and UO_1646 (O_1646,N_48308,N_48054);
or UO_1647 (O_1647,N_49164,N_49264);
nand UO_1648 (O_1648,N_49284,N_48552);
and UO_1649 (O_1649,N_48720,N_49225);
or UO_1650 (O_1650,N_49630,N_48902);
nand UO_1651 (O_1651,N_48524,N_48931);
nand UO_1652 (O_1652,N_48924,N_49941);
nand UO_1653 (O_1653,N_49709,N_49232);
nor UO_1654 (O_1654,N_49751,N_48932);
nand UO_1655 (O_1655,N_48242,N_48627);
or UO_1656 (O_1656,N_48139,N_48508);
xor UO_1657 (O_1657,N_48924,N_49355);
nor UO_1658 (O_1658,N_48785,N_49641);
nor UO_1659 (O_1659,N_48114,N_48759);
or UO_1660 (O_1660,N_48474,N_48364);
and UO_1661 (O_1661,N_48480,N_48193);
or UO_1662 (O_1662,N_49338,N_48529);
nand UO_1663 (O_1663,N_49586,N_49387);
nor UO_1664 (O_1664,N_49586,N_49819);
or UO_1665 (O_1665,N_49031,N_49260);
nand UO_1666 (O_1666,N_48954,N_48410);
nand UO_1667 (O_1667,N_48805,N_49613);
nand UO_1668 (O_1668,N_49863,N_48733);
nand UO_1669 (O_1669,N_49186,N_48675);
and UO_1670 (O_1670,N_49594,N_49615);
and UO_1671 (O_1671,N_48894,N_49257);
nand UO_1672 (O_1672,N_48845,N_48535);
nor UO_1673 (O_1673,N_49081,N_48143);
and UO_1674 (O_1674,N_49058,N_48307);
nand UO_1675 (O_1675,N_49101,N_48218);
nand UO_1676 (O_1676,N_48501,N_48488);
and UO_1677 (O_1677,N_48546,N_48307);
xnor UO_1678 (O_1678,N_48591,N_49484);
and UO_1679 (O_1679,N_48695,N_49740);
nor UO_1680 (O_1680,N_48495,N_49454);
nor UO_1681 (O_1681,N_48785,N_49564);
or UO_1682 (O_1682,N_48134,N_49489);
nand UO_1683 (O_1683,N_48570,N_48705);
nor UO_1684 (O_1684,N_49225,N_48072);
nand UO_1685 (O_1685,N_49706,N_49376);
nand UO_1686 (O_1686,N_49192,N_49688);
nor UO_1687 (O_1687,N_48510,N_48410);
nand UO_1688 (O_1688,N_49880,N_48863);
nand UO_1689 (O_1689,N_49505,N_49694);
nand UO_1690 (O_1690,N_49209,N_49749);
nand UO_1691 (O_1691,N_48296,N_49726);
and UO_1692 (O_1692,N_48531,N_49985);
or UO_1693 (O_1693,N_48808,N_49948);
nand UO_1694 (O_1694,N_49528,N_48797);
and UO_1695 (O_1695,N_48061,N_49342);
nor UO_1696 (O_1696,N_48772,N_48365);
and UO_1697 (O_1697,N_48041,N_49438);
nor UO_1698 (O_1698,N_49025,N_49503);
or UO_1699 (O_1699,N_49801,N_48390);
nand UO_1700 (O_1700,N_48513,N_49014);
nor UO_1701 (O_1701,N_49846,N_49370);
or UO_1702 (O_1702,N_48153,N_49142);
nand UO_1703 (O_1703,N_49153,N_49677);
nand UO_1704 (O_1704,N_48458,N_48447);
and UO_1705 (O_1705,N_48873,N_49428);
nand UO_1706 (O_1706,N_48212,N_48260);
nor UO_1707 (O_1707,N_48416,N_49811);
nand UO_1708 (O_1708,N_49792,N_48509);
and UO_1709 (O_1709,N_49405,N_48986);
or UO_1710 (O_1710,N_49969,N_49288);
nand UO_1711 (O_1711,N_48338,N_49331);
nand UO_1712 (O_1712,N_49030,N_48125);
nor UO_1713 (O_1713,N_49344,N_49159);
nand UO_1714 (O_1714,N_48986,N_48151);
nand UO_1715 (O_1715,N_48062,N_48020);
nand UO_1716 (O_1716,N_49705,N_49775);
nand UO_1717 (O_1717,N_49944,N_49473);
nor UO_1718 (O_1718,N_48702,N_49317);
nand UO_1719 (O_1719,N_48695,N_49849);
xnor UO_1720 (O_1720,N_48678,N_48418);
or UO_1721 (O_1721,N_49186,N_48180);
nor UO_1722 (O_1722,N_48440,N_49129);
or UO_1723 (O_1723,N_49650,N_48249);
nor UO_1724 (O_1724,N_49958,N_48344);
nand UO_1725 (O_1725,N_48996,N_48997);
nor UO_1726 (O_1726,N_48470,N_49768);
and UO_1727 (O_1727,N_48987,N_48734);
nor UO_1728 (O_1728,N_49310,N_49377);
or UO_1729 (O_1729,N_48285,N_49793);
and UO_1730 (O_1730,N_49681,N_48075);
nor UO_1731 (O_1731,N_49430,N_48896);
or UO_1732 (O_1732,N_49768,N_49481);
or UO_1733 (O_1733,N_48070,N_48888);
nor UO_1734 (O_1734,N_48451,N_48550);
or UO_1735 (O_1735,N_49804,N_48015);
and UO_1736 (O_1736,N_48219,N_49823);
or UO_1737 (O_1737,N_48826,N_48930);
or UO_1738 (O_1738,N_49361,N_49515);
nor UO_1739 (O_1739,N_48591,N_48103);
and UO_1740 (O_1740,N_48491,N_49649);
nor UO_1741 (O_1741,N_48740,N_49746);
and UO_1742 (O_1742,N_49434,N_49791);
nor UO_1743 (O_1743,N_48306,N_48661);
nor UO_1744 (O_1744,N_49281,N_48611);
nand UO_1745 (O_1745,N_48062,N_49880);
or UO_1746 (O_1746,N_49413,N_48587);
nor UO_1747 (O_1747,N_48094,N_49723);
nor UO_1748 (O_1748,N_49803,N_48045);
and UO_1749 (O_1749,N_48128,N_49381);
nand UO_1750 (O_1750,N_48817,N_49501);
nor UO_1751 (O_1751,N_49222,N_49938);
and UO_1752 (O_1752,N_49214,N_49575);
and UO_1753 (O_1753,N_49317,N_48784);
or UO_1754 (O_1754,N_49040,N_49015);
and UO_1755 (O_1755,N_49204,N_49955);
and UO_1756 (O_1756,N_48280,N_49282);
nand UO_1757 (O_1757,N_48717,N_48467);
or UO_1758 (O_1758,N_48951,N_48360);
and UO_1759 (O_1759,N_48978,N_49401);
nand UO_1760 (O_1760,N_49220,N_48009);
nor UO_1761 (O_1761,N_49031,N_49999);
and UO_1762 (O_1762,N_48735,N_49961);
and UO_1763 (O_1763,N_49965,N_48226);
or UO_1764 (O_1764,N_49974,N_48502);
nand UO_1765 (O_1765,N_48448,N_48841);
and UO_1766 (O_1766,N_49979,N_49714);
or UO_1767 (O_1767,N_49365,N_48968);
and UO_1768 (O_1768,N_49802,N_48314);
nor UO_1769 (O_1769,N_49768,N_49141);
and UO_1770 (O_1770,N_48297,N_49012);
nor UO_1771 (O_1771,N_48350,N_49402);
nand UO_1772 (O_1772,N_48837,N_49258);
or UO_1773 (O_1773,N_49694,N_49605);
nor UO_1774 (O_1774,N_49359,N_48345);
and UO_1775 (O_1775,N_49420,N_48131);
or UO_1776 (O_1776,N_49688,N_49857);
and UO_1777 (O_1777,N_48038,N_49337);
or UO_1778 (O_1778,N_49342,N_48758);
and UO_1779 (O_1779,N_48685,N_49553);
nor UO_1780 (O_1780,N_49102,N_48470);
or UO_1781 (O_1781,N_49880,N_48444);
or UO_1782 (O_1782,N_49081,N_49695);
nand UO_1783 (O_1783,N_48920,N_49502);
nor UO_1784 (O_1784,N_49904,N_48233);
nor UO_1785 (O_1785,N_49670,N_48141);
nor UO_1786 (O_1786,N_48566,N_49401);
nand UO_1787 (O_1787,N_49336,N_49748);
nor UO_1788 (O_1788,N_48787,N_48536);
nand UO_1789 (O_1789,N_48776,N_49920);
and UO_1790 (O_1790,N_48744,N_48405);
nor UO_1791 (O_1791,N_48035,N_49182);
and UO_1792 (O_1792,N_49549,N_48391);
or UO_1793 (O_1793,N_49167,N_49493);
xor UO_1794 (O_1794,N_48503,N_49327);
and UO_1795 (O_1795,N_49262,N_49247);
nand UO_1796 (O_1796,N_48950,N_49359);
nand UO_1797 (O_1797,N_48183,N_48704);
and UO_1798 (O_1798,N_49829,N_48480);
and UO_1799 (O_1799,N_48947,N_48967);
or UO_1800 (O_1800,N_49912,N_49377);
and UO_1801 (O_1801,N_49417,N_48439);
nor UO_1802 (O_1802,N_48452,N_48383);
and UO_1803 (O_1803,N_49862,N_49738);
and UO_1804 (O_1804,N_48623,N_48910);
nor UO_1805 (O_1805,N_48028,N_49445);
nand UO_1806 (O_1806,N_48063,N_48378);
nand UO_1807 (O_1807,N_49181,N_49752);
or UO_1808 (O_1808,N_49341,N_48221);
nor UO_1809 (O_1809,N_49501,N_49554);
nor UO_1810 (O_1810,N_48637,N_49107);
nand UO_1811 (O_1811,N_48264,N_48323);
or UO_1812 (O_1812,N_49657,N_49104);
nor UO_1813 (O_1813,N_48378,N_49346);
nor UO_1814 (O_1814,N_49870,N_49785);
nand UO_1815 (O_1815,N_48550,N_48783);
xnor UO_1816 (O_1816,N_49857,N_48267);
or UO_1817 (O_1817,N_49074,N_49311);
nand UO_1818 (O_1818,N_49560,N_48788);
and UO_1819 (O_1819,N_48029,N_49176);
or UO_1820 (O_1820,N_49844,N_48216);
nand UO_1821 (O_1821,N_49111,N_48820);
nor UO_1822 (O_1822,N_48210,N_48582);
nand UO_1823 (O_1823,N_49877,N_49199);
nand UO_1824 (O_1824,N_49573,N_48207);
nor UO_1825 (O_1825,N_49210,N_49823);
nand UO_1826 (O_1826,N_49222,N_49479);
nor UO_1827 (O_1827,N_48139,N_48612);
and UO_1828 (O_1828,N_49129,N_49661);
nor UO_1829 (O_1829,N_48259,N_49117);
nor UO_1830 (O_1830,N_49757,N_49367);
and UO_1831 (O_1831,N_49000,N_49294);
or UO_1832 (O_1832,N_48994,N_48836);
and UO_1833 (O_1833,N_49043,N_49130);
or UO_1834 (O_1834,N_49668,N_49877);
nor UO_1835 (O_1835,N_48441,N_49667);
and UO_1836 (O_1836,N_48548,N_49251);
or UO_1837 (O_1837,N_48392,N_49676);
or UO_1838 (O_1838,N_48781,N_48766);
and UO_1839 (O_1839,N_48340,N_49748);
nor UO_1840 (O_1840,N_48950,N_49354);
and UO_1841 (O_1841,N_49626,N_48670);
nand UO_1842 (O_1842,N_49117,N_49170);
or UO_1843 (O_1843,N_49798,N_49739);
nor UO_1844 (O_1844,N_49770,N_49200);
nand UO_1845 (O_1845,N_48896,N_49239);
nor UO_1846 (O_1846,N_49684,N_48351);
and UO_1847 (O_1847,N_49762,N_48932);
or UO_1848 (O_1848,N_49063,N_49504);
or UO_1849 (O_1849,N_48234,N_49964);
nor UO_1850 (O_1850,N_48162,N_49387);
nand UO_1851 (O_1851,N_49910,N_48807);
nand UO_1852 (O_1852,N_49120,N_49796);
and UO_1853 (O_1853,N_48760,N_49195);
or UO_1854 (O_1854,N_48115,N_49553);
xor UO_1855 (O_1855,N_48198,N_48232);
or UO_1856 (O_1856,N_49792,N_48111);
nor UO_1857 (O_1857,N_48449,N_48914);
nor UO_1858 (O_1858,N_48367,N_49153);
nand UO_1859 (O_1859,N_49191,N_48864);
nor UO_1860 (O_1860,N_49598,N_49089);
and UO_1861 (O_1861,N_49277,N_48943);
nor UO_1862 (O_1862,N_48653,N_48392);
or UO_1863 (O_1863,N_48722,N_48429);
nand UO_1864 (O_1864,N_48465,N_48480);
and UO_1865 (O_1865,N_48543,N_49325);
nand UO_1866 (O_1866,N_49156,N_48056);
and UO_1867 (O_1867,N_48412,N_49683);
and UO_1868 (O_1868,N_48984,N_49345);
or UO_1869 (O_1869,N_48818,N_48727);
nor UO_1870 (O_1870,N_48529,N_48275);
nand UO_1871 (O_1871,N_48120,N_48865);
nand UO_1872 (O_1872,N_48230,N_48437);
nor UO_1873 (O_1873,N_49617,N_49744);
or UO_1874 (O_1874,N_49132,N_48749);
nor UO_1875 (O_1875,N_48856,N_48077);
nand UO_1876 (O_1876,N_49620,N_49267);
and UO_1877 (O_1877,N_48952,N_48675);
xnor UO_1878 (O_1878,N_48153,N_49176);
or UO_1879 (O_1879,N_49525,N_49060);
nand UO_1880 (O_1880,N_48281,N_49087);
and UO_1881 (O_1881,N_48604,N_49593);
nor UO_1882 (O_1882,N_49083,N_48245);
and UO_1883 (O_1883,N_49719,N_49827);
or UO_1884 (O_1884,N_48763,N_49669);
nor UO_1885 (O_1885,N_48237,N_49261);
or UO_1886 (O_1886,N_48536,N_49259);
nor UO_1887 (O_1887,N_48820,N_48265);
nor UO_1888 (O_1888,N_48650,N_48898);
nand UO_1889 (O_1889,N_49751,N_49299);
and UO_1890 (O_1890,N_48634,N_48553);
or UO_1891 (O_1891,N_49681,N_49773);
nand UO_1892 (O_1892,N_49033,N_48756);
nor UO_1893 (O_1893,N_48421,N_49205);
and UO_1894 (O_1894,N_48581,N_49711);
or UO_1895 (O_1895,N_49456,N_49838);
nand UO_1896 (O_1896,N_48460,N_48339);
nand UO_1897 (O_1897,N_48170,N_48132);
and UO_1898 (O_1898,N_48914,N_48698);
or UO_1899 (O_1899,N_49757,N_49623);
and UO_1900 (O_1900,N_48281,N_49377);
nor UO_1901 (O_1901,N_48875,N_48284);
nand UO_1902 (O_1902,N_49199,N_49204);
and UO_1903 (O_1903,N_48887,N_48365);
xor UO_1904 (O_1904,N_49829,N_48172);
nor UO_1905 (O_1905,N_49249,N_49359);
nor UO_1906 (O_1906,N_48890,N_49759);
nor UO_1907 (O_1907,N_49541,N_49885);
nor UO_1908 (O_1908,N_49665,N_48737);
or UO_1909 (O_1909,N_49657,N_49480);
and UO_1910 (O_1910,N_49534,N_49475);
nand UO_1911 (O_1911,N_49128,N_48476);
nand UO_1912 (O_1912,N_49525,N_49736);
or UO_1913 (O_1913,N_49198,N_48806);
or UO_1914 (O_1914,N_48112,N_48705);
and UO_1915 (O_1915,N_48976,N_49742);
nor UO_1916 (O_1916,N_48720,N_48358);
nor UO_1917 (O_1917,N_49274,N_49491);
nand UO_1918 (O_1918,N_48125,N_49182);
and UO_1919 (O_1919,N_48892,N_48871);
nand UO_1920 (O_1920,N_48414,N_48460);
nor UO_1921 (O_1921,N_48948,N_48714);
and UO_1922 (O_1922,N_49405,N_48840);
or UO_1923 (O_1923,N_48906,N_49404);
and UO_1924 (O_1924,N_48697,N_48409);
or UO_1925 (O_1925,N_49801,N_49604);
nor UO_1926 (O_1926,N_49841,N_48136);
and UO_1927 (O_1927,N_49470,N_48042);
and UO_1928 (O_1928,N_49307,N_49892);
nor UO_1929 (O_1929,N_48468,N_49479);
nor UO_1930 (O_1930,N_49173,N_49873);
nor UO_1931 (O_1931,N_48966,N_49876);
and UO_1932 (O_1932,N_49141,N_49339);
nand UO_1933 (O_1933,N_48915,N_48630);
nor UO_1934 (O_1934,N_48202,N_49340);
nor UO_1935 (O_1935,N_48056,N_49358);
nand UO_1936 (O_1936,N_48460,N_49955);
or UO_1937 (O_1937,N_48725,N_49456);
nand UO_1938 (O_1938,N_48708,N_48252);
nor UO_1939 (O_1939,N_48773,N_49423);
or UO_1940 (O_1940,N_48864,N_49625);
nor UO_1941 (O_1941,N_49972,N_49141);
nor UO_1942 (O_1942,N_49277,N_49568);
nand UO_1943 (O_1943,N_49040,N_49899);
nand UO_1944 (O_1944,N_49011,N_49831);
or UO_1945 (O_1945,N_49705,N_48118);
xor UO_1946 (O_1946,N_49481,N_48680);
and UO_1947 (O_1947,N_48091,N_49974);
nand UO_1948 (O_1948,N_49316,N_49234);
and UO_1949 (O_1949,N_49270,N_49221);
nand UO_1950 (O_1950,N_49266,N_48252);
nand UO_1951 (O_1951,N_48299,N_49417);
and UO_1952 (O_1952,N_48370,N_48659);
nor UO_1953 (O_1953,N_48265,N_49491);
nand UO_1954 (O_1954,N_48386,N_49284);
and UO_1955 (O_1955,N_48069,N_49290);
or UO_1956 (O_1956,N_48897,N_48105);
or UO_1957 (O_1957,N_48745,N_49363);
nand UO_1958 (O_1958,N_48607,N_48006);
xnor UO_1959 (O_1959,N_49017,N_48984);
nand UO_1960 (O_1960,N_49223,N_48925);
nand UO_1961 (O_1961,N_49115,N_48451);
nor UO_1962 (O_1962,N_49363,N_48695);
nand UO_1963 (O_1963,N_49887,N_49133);
nand UO_1964 (O_1964,N_49752,N_49338);
and UO_1965 (O_1965,N_48043,N_49745);
or UO_1966 (O_1966,N_48680,N_49726);
or UO_1967 (O_1967,N_49325,N_48374);
and UO_1968 (O_1968,N_49258,N_49824);
nor UO_1969 (O_1969,N_49386,N_49369);
nor UO_1970 (O_1970,N_49796,N_48055);
and UO_1971 (O_1971,N_49709,N_49133);
or UO_1972 (O_1972,N_48467,N_49048);
or UO_1973 (O_1973,N_49665,N_48026);
nor UO_1974 (O_1974,N_49018,N_49849);
or UO_1975 (O_1975,N_49977,N_49774);
or UO_1976 (O_1976,N_49486,N_48827);
nand UO_1977 (O_1977,N_48860,N_49662);
nor UO_1978 (O_1978,N_49008,N_49310);
and UO_1979 (O_1979,N_49980,N_48716);
nor UO_1980 (O_1980,N_49371,N_49607);
and UO_1981 (O_1981,N_48239,N_48285);
or UO_1982 (O_1982,N_48877,N_49477);
nor UO_1983 (O_1983,N_48101,N_49101);
and UO_1984 (O_1984,N_49004,N_48566);
nand UO_1985 (O_1985,N_48805,N_49723);
and UO_1986 (O_1986,N_49039,N_48464);
or UO_1987 (O_1987,N_48990,N_48242);
nor UO_1988 (O_1988,N_49968,N_49422);
nor UO_1989 (O_1989,N_49911,N_48157);
or UO_1990 (O_1990,N_48500,N_48161);
nand UO_1991 (O_1991,N_48030,N_48357);
nand UO_1992 (O_1992,N_48433,N_49623);
nand UO_1993 (O_1993,N_48744,N_49862);
xor UO_1994 (O_1994,N_49589,N_49330);
and UO_1995 (O_1995,N_48718,N_49168);
nor UO_1996 (O_1996,N_49030,N_48174);
or UO_1997 (O_1997,N_49415,N_49526);
and UO_1998 (O_1998,N_48658,N_49052);
or UO_1999 (O_1999,N_48904,N_49401);
or UO_2000 (O_2000,N_48541,N_48372);
nor UO_2001 (O_2001,N_48672,N_49173);
or UO_2002 (O_2002,N_49848,N_48091);
or UO_2003 (O_2003,N_49275,N_49247);
and UO_2004 (O_2004,N_48082,N_49238);
nor UO_2005 (O_2005,N_48388,N_48826);
nor UO_2006 (O_2006,N_49719,N_49807);
and UO_2007 (O_2007,N_48791,N_49123);
nor UO_2008 (O_2008,N_49880,N_48974);
nor UO_2009 (O_2009,N_49298,N_48567);
nand UO_2010 (O_2010,N_49977,N_49543);
nand UO_2011 (O_2011,N_48523,N_49151);
nor UO_2012 (O_2012,N_49676,N_48472);
nor UO_2013 (O_2013,N_48827,N_49627);
and UO_2014 (O_2014,N_49228,N_48622);
nor UO_2015 (O_2015,N_48983,N_48594);
nand UO_2016 (O_2016,N_48833,N_49383);
or UO_2017 (O_2017,N_48190,N_49794);
nor UO_2018 (O_2018,N_49449,N_49604);
and UO_2019 (O_2019,N_49974,N_49973);
nor UO_2020 (O_2020,N_48952,N_49324);
nor UO_2021 (O_2021,N_49890,N_49981);
nand UO_2022 (O_2022,N_48640,N_49791);
or UO_2023 (O_2023,N_48013,N_48361);
or UO_2024 (O_2024,N_48266,N_48073);
nor UO_2025 (O_2025,N_49872,N_48960);
nor UO_2026 (O_2026,N_48313,N_49090);
nor UO_2027 (O_2027,N_49634,N_48805);
xnor UO_2028 (O_2028,N_49704,N_48455);
nor UO_2029 (O_2029,N_48797,N_49315);
xor UO_2030 (O_2030,N_49734,N_49219);
nand UO_2031 (O_2031,N_49398,N_49416);
nand UO_2032 (O_2032,N_49128,N_49260);
and UO_2033 (O_2033,N_48481,N_48579);
nand UO_2034 (O_2034,N_49307,N_48578);
nand UO_2035 (O_2035,N_48036,N_48605);
and UO_2036 (O_2036,N_49028,N_49112);
nor UO_2037 (O_2037,N_48509,N_49605);
or UO_2038 (O_2038,N_48049,N_49922);
and UO_2039 (O_2039,N_49676,N_48347);
or UO_2040 (O_2040,N_49737,N_48936);
and UO_2041 (O_2041,N_48547,N_49366);
and UO_2042 (O_2042,N_49263,N_49544);
or UO_2043 (O_2043,N_48642,N_48035);
or UO_2044 (O_2044,N_49661,N_48459);
nand UO_2045 (O_2045,N_49571,N_48916);
or UO_2046 (O_2046,N_49864,N_49233);
and UO_2047 (O_2047,N_48981,N_48583);
and UO_2048 (O_2048,N_48400,N_48128);
and UO_2049 (O_2049,N_49335,N_49824);
and UO_2050 (O_2050,N_49274,N_49820);
nand UO_2051 (O_2051,N_49857,N_48566);
nor UO_2052 (O_2052,N_48760,N_49228);
and UO_2053 (O_2053,N_49821,N_48436);
nand UO_2054 (O_2054,N_49453,N_48562);
and UO_2055 (O_2055,N_49138,N_48079);
and UO_2056 (O_2056,N_48868,N_49422);
xor UO_2057 (O_2057,N_49537,N_48023);
or UO_2058 (O_2058,N_48618,N_48719);
nor UO_2059 (O_2059,N_48154,N_49574);
nor UO_2060 (O_2060,N_48803,N_49629);
or UO_2061 (O_2061,N_48849,N_48237);
or UO_2062 (O_2062,N_49646,N_49849);
or UO_2063 (O_2063,N_49014,N_48153);
nor UO_2064 (O_2064,N_48590,N_49734);
nand UO_2065 (O_2065,N_49529,N_49148);
or UO_2066 (O_2066,N_49337,N_48330);
or UO_2067 (O_2067,N_49196,N_49119);
nand UO_2068 (O_2068,N_49092,N_48963);
or UO_2069 (O_2069,N_49534,N_48714);
or UO_2070 (O_2070,N_48554,N_49109);
or UO_2071 (O_2071,N_48054,N_49743);
and UO_2072 (O_2072,N_49998,N_49651);
nor UO_2073 (O_2073,N_49351,N_48016);
or UO_2074 (O_2074,N_49636,N_49969);
and UO_2075 (O_2075,N_49157,N_49679);
nor UO_2076 (O_2076,N_48270,N_49973);
and UO_2077 (O_2077,N_49831,N_48079);
nor UO_2078 (O_2078,N_49587,N_49660);
nand UO_2079 (O_2079,N_49766,N_49614);
and UO_2080 (O_2080,N_49686,N_48241);
and UO_2081 (O_2081,N_48135,N_49117);
nand UO_2082 (O_2082,N_48678,N_48482);
nor UO_2083 (O_2083,N_49961,N_49003);
and UO_2084 (O_2084,N_49364,N_49076);
nor UO_2085 (O_2085,N_48847,N_48365);
nand UO_2086 (O_2086,N_49843,N_48182);
and UO_2087 (O_2087,N_49309,N_48002);
nor UO_2088 (O_2088,N_49308,N_49948);
or UO_2089 (O_2089,N_49679,N_49982);
nor UO_2090 (O_2090,N_49842,N_48919);
nand UO_2091 (O_2091,N_49516,N_48134);
nor UO_2092 (O_2092,N_48963,N_48472);
nor UO_2093 (O_2093,N_49166,N_48655);
or UO_2094 (O_2094,N_49240,N_48642);
and UO_2095 (O_2095,N_49100,N_49196);
nor UO_2096 (O_2096,N_48939,N_49494);
and UO_2097 (O_2097,N_49548,N_48127);
or UO_2098 (O_2098,N_49297,N_48514);
nor UO_2099 (O_2099,N_49866,N_49525);
and UO_2100 (O_2100,N_49452,N_48320);
and UO_2101 (O_2101,N_49366,N_49292);
xnor UO_2102 (O_2102,N_49856,N_49763);
and UO_2103 (O_2103,N_48270,N_48316);
or UO_2104 (O_2104,N_49601,N_48749);
and UO_2105 (O_2105,N_49039,N_49484);
nand UO_2106 (O_2106,N_48529,N_48846);
or UO_2107 (O_2107,N_49337,N_48116);
nor UO_2108 (O_2108,N_49487,N_49910);
nor UO_2109 (O_2109,N_48570,N_49509);
or UO_2110 (O_2110,N_49621,N_49638);
xor UO_2111 (O_2111,N_49591,N_49812);
and UO_2112 (O_2112,N_49563,N_49306);
or UO_2113 (O_2113,N_49739,N_49117);
nand UO_2114 (O_2114,N_49011,N_49184);
or UO_2115 (O_2115,N_49689,N_49371);
nor UO_2116 (O_2116,N_49136,N_49013);
nand UO_2117 (O_2117,N_48313,N_49724);
nand UO_2118 (O_2118,N_48402,N_48881);
and UO_2119 (O_2119,N_48721,N_49813);
and UO_2120 (O_2120,N_49086,N_49290);
or UO_2121 (O_2121,N_49744,N_48259);
nor UO_2122 (O_2122,N_49998,N_49026);
or UO_2123 (O_2123,N_48291,N_48379);
nor UO_2124 (O_2124,N_48947,N_49312);
and UO_2125 (O_2125,N_49081,N_48705);
and UO_2126 (O_2126,N_48570,N_49566);
and UO_2127 (O_2127,N_48457,N_49408);
or UO_2128 (O_2128,N_48860,N_49437);
and UO_2129 (O_2129,N_48850,N_49342);
nand UO_2130 (O_2130,N_48775,N_48202);
nor UO_2131 (O_2131,N_49414,N_48934);
nor UO_2132 (O_2132,N_48623,N_48933);
or UO_2133 (O_2133,N_48820,N_49833);
nand UO_2134 (O_2134,N_48400,N_48121);
nand UO_2135 (O_2135,N_49681,N_48382);
nand UO_2136 (O_2136,N_49182,N_49594);
nor UO_2137 (O_2137,N_48126,N_48315);
nand UO_2138 (O_2138,N_48086,N_49848);
nor UO_2139 (O_2139,N_48510,N_49659);
and UO_2140 (O_2140,N_49592,N_49093);
nand UO_2141 (O_2141,N_48108,N_48744);
or UO_2142 (O_2142,N_48583,N_49556);
or UO_2143 (O_2143,N_48756,N_48382);
or UO_2144 (O_2144,N_49712,N_48044);
nor UO_2145 (O_2145,N_48952,N_48705);
or UO_2146 (O_2146,N_49514,N_49802);
or UO_2147 (O_2147,N_48931,N_48383);
and UO_2148 (O_2148,N_49112,N_48008);
nand UO_2149 (O_2149,N_49084,N_48606);
or UO_2150 (O_2150,N_49660,N_48966);
or UO_2151 (O_2151,N_48679,N_48838);
nor UO_2152 (O_2152,N_49691,N_49510);
and UO_2153 (O_2153,N_49353,N_48521);
nand UO_2154 (O_2154,N_48784,N_48856);
nand UO_2155 (O_2155,N_49136,N_48922);
xor UO_2156 (O_2156,N_49352,N_49424);
or UO_2157 (O_2157,N_49273,N_48268);
nand UO_2158 (O_2158,N_48166,N_48484);
and UO_2159 (O_2159,N_48475,N_48630);
and UO_2160 (O_2160,N_48028,N_49730);
nor UO_2161 (O_2161,N_49729,N_49446);
nand UO_2162 (O_2162,N_49410,N_48118);
and UO_2163 (O_2163,N_49412,N_48673);
nor UO_2164 (O_2164,N_49481,N_48347);
and UO_2165 (O_2165,N_48409,N_48650);
or UO_2166 (O_2166,N_49720,N_48111);
or UO_2167 (O_2167,N_48553,N_48900);
nand UO_2168 (O_2168,N_48858,N_49345);
and UO_2169 (O_2169,N_49923,N_48600);
or UO_2170 (O_2170,N_48993,N_48084);
and UO_2171 (O_2171,N_48628,N_48943);
or UO_2172 (O_2172,N_48644,N_48858);
nand UO_2173 (O_2173,N_48467,N_49848);
and UO_2174 (O_2174,N_48487,N_48560);
nor UO_2175 (O_2175,N_48028,N_48063);
nand UO_2176 (O_2176,N_48041,N_49485);
nor UO_2177 (O_2177,N_49882,N_48521);
nand UO_2178 (O_2178,N_48770,N_49290);
and UO_2179 (O_2179,N_48208,N_48258);
nor UO_2180 (O_2180,N_48635,N_48978);
or UO_2181 (O_2181,N_49027,N_49526);
and UO_2182 (O_2182,N_48059,N_49149);
nand UO_2183 (O_2183,N_49386,N_48858);
nand UO_2184 (O_2184,N_48946,N_49503);
nor UO_2185 (O_2185,N_48295,N_48177);
nand UO_2186 (O_2186,N_48173,N_49284);
and UO_2187 (O_2187,N_49141,N_49671);
nor UO_2188 (O_2188,N_48683,N_49757);
and UO_2189 (O_2189,N_49931,N_48080);
nand UO_2190 (O_2190,N_49729,N_48303);
xor UO_2191 (O_2191,N_49262,N_48890);
or UO_2192 (O_2192,N_48818,N_48700);
nand UO_2193 (O_2193,N_49382,N_49426);
or UO_2194 (O_2194,N_49513,N_48274);
nand UO_2195 (O_2195,N_49069,N_49031);
or UO_2196 (O_2196,N_49943,N_48295);
and UO_2197 (O_2197,N_49984,N_49055);
nor UO_2198 (O_2198,N_49691,N_48807);
nor UO_2199 (O_2199,N_48276,N_49656);
and UO_2200 (O_2200,N_49699,N_48499);
nand UO_2201 (O_2201,N_48836,N_48231);
nor UO_2202 (O_2202,N_48529,N_49221);
nor UO_2203 (O_2203,N_48623,N_48224);
nand UO_2204 (O_2204,N_48630,N_48586);
or UO_2205 (O_2205,N_49068,N_49867);
and UO_2206 (O_2206,N_49631,N_49013);
and UO_2207 (O_2207,N_48875,N_49097);
nor UO_2208 (O_2208,N_48567,N_49698);
and UO_2209 (O_2209,N_49328,N_49147);
and UO_2210 (O_2210,N_49243,N_48525);
or UO_2211 (O_2211,N_48862,N_49518);
nor UO_2212 (O_2212,N_49393,N_49487);
and UO_2213 (O_2213,N_49915,N_49328);
and UO_2214 (O_2214,N_49049,N_48634);
nor UO_2215 (O_2215,N_48709,N_48529);
or UO_2216 (O_2216,N_48025,N_48223);
and UO_2217 (O_2217,N_48231,N_48393);
or UO_2218 (O_2218,N_48824,N_49676);
nand UO_2219 (O_2219,N_48374,N_49367);
nand UO_2220 (O_2220,N_49085,N_49117);
nand UO_2221 (O_2221,N_48781,N_49619);
nand UO_2222 (O_2222,N_48263,N_48369);
or UO_2223 (O_2223,N_48327,N_48913);
nor UO_2224 (O_2224,N_48233,N_48610);
nor UO_2225 (O_2225,N_49936,N_48651);
nor UO_2226 (O_2226,N_48588,N_48813);
and UO_2227 (O_2227,N_49157,N_48515);
nor UO_2228 (O_2228,N_49205,N_48925);
or UO_2229 (O_2229,N_48870,N_48968);
nand UO_2230 (O_2230,N_49818,N_49312);
nand UO_2231 (O_2231,N_49312,N_49336);
and UO_2232 (O_2232,N_48775,N_48364);
and UO_2233 (O_2233,N_49983,N_49095);
nand UO_2234 (O_2234,N_48250,N_48754);
nand UO_2235 (O_2235,N_49609,N_49237);
nand UO_2236 (O_2236,N_48575,N_48177);
nand UO_2237 (O_2237,N_48729,N_49546);
and UO_2238 (O_2238,N_49919,N_48187);
and UO_2239 (O_2239,N_48806,N_49467);
and UO_2240 (O_2240,N_49729,N_49259);
xor UO_2241 (O_2241,N_48878,N_48075);
nand UO_2242 (O_2242,N_48239,N_48040);
nor UO_2243 (O_2243,N_49842,N_49870);
nand UO_2244 (O_2244,N_48177,N_49518);
nor UO_2245 (O_2245,N_48161,N_49785);
and UO_2246 (O_2246,N_49891,N_49804);
nand UO_2247 (O_2247,N_49840,N_48998);
or UO_2248 (O_2248,N_49155,N_49729);
and UO_2249 (O_2249,N_48009,N_49460);
and UO_2250 (O_2250,N_49221,N_49693);
nor UO_2251 (O_2251,N_48606,N_49665);
and UO_2252 (O_2252,N_49898,N_49527);
or UO_2253 (O_2253,N_48979,N_48974);
and UO_2254 (O_2254,N_49865,N_48660);
or UO_2255 (O_2255,N_48877,N_49051);
and UO_2256 (O_2256,N_48232,N_49232);
or UO_2257 (O_2257,N_49078,N_49098);
and UO_2258 (O_2258,N_49816,N_48998);
xnor UO_2259 (O_2259,N_49449,N_48224);
or UO_2260 (O_2260,N_48533,N_49063);
or UO_2261 (O_2261,N_48176,N_48262);
nor UO_2262 (O_2262,N_49698,N_49993);
and UO_2263 (O_2263,N_49774,N_48773);
and UO_2264 (O_2264,N_48528,N_48892);
nor UO_2265 (O_2265,N_48286,N_48270);
and UO_2266 (O_2266,N_49500,N_48963);
nand UO_2267 (O_2267,N_49977,N_49894);
nor UO_2268 (O_2268,N_49801,N_49359);
nand UO_2269 (O_2269,N_48710,N_49983);
xor UO_2270 (O_2270,N_49557,N_48239);
or UO_2271 (O_2271,N_48067,N_48901);
or UO_2272 (O_2272,N_49591,N_48614);
and UO_2273 (O_2273,N_48085,N_49855);
nor UO_2274 (O_2274,N_49585,N_48612);
nand UO_2275 (O_2275,N_49880,N_48440);
and UO_2276 (O_2276,N_48440,N_49126);
and UO_2277 (O_2277,N_49106,N_49955);
xnor UO_2278 (O_2278,N_48514,N_48663);
nor UO_2279 (O_2279,N_48020,N_49413);
or UO_2280 (O_2280,N_48822,N_48483);
and UO_2281 (O_2281,N_48265,N_49708);
or UO_2282 (O_2282,N_48445,N_48234);
or UO_2283 (O_2283,N_49435,N_49594);
or UO_2284 (O_2284,N_48437,N_48954);
and UO_2285 (O_2285,N_48148,N_48064);
or UO_2286 (O_2286,N_49750,N_49153);
nand UO_2287 (O_2287,N_49478,N_49522);
and UO_2288 (O_2288,N_48045,N_48122);
or UO_2289 (O_2289,N_48434,N_49274);
nand UO_2290 (O_2290,N_49247,N_49175);
or UO_2291 (O_2291,N_49004,N_49362);
nor UO_2292 (O_2292,N_48531,N_49203);
nor UO_2293 (O_2293,N_48511,N_49792);
nor UO_2294 (O_2294,N_49684,N_48617);
or UO_2295 (O_2295,N_48530,N_49566);
nand UO_2296 (O_2296,N_49731,N_48740);
nand UO_2297 (O_2297,N_48820,N_49335);
or UO_2298 (O_2298,N_48195,N_49324);
or UO_2299 (O_2299,N_49493,N_49716);
or UO_2300 (O_2300,N_49050,N_48295);
nand UO_2301 (O_2301,N_48424,N_48612);
nand UO_2302 (O_2302,N_48080,N_49930);
and UO_2303 (O_2303,N_49253,N_49350);
or UO_2304 (O_2304,N_48304,N_48754);
nor UO_2305 (O_2305,N_48453,N_48587);
nor UO_2306 (O_2306,N_49325,N_48475);
nor UO_2307 (O_2307,N_48246,N_49502);
nor UO_2308 (O_2308,N_49463,N_49681);
or UO_2309 (O_2309,N_49277,N_49522);
xnor UO_2310 (O_2310,N_48867,N_49511);
or UO_2311 (O_2311,N_49592,N_48710);
nand UO_2312 (O_2312,N_49451,N_48915);
xor UO_2313 (O_2313,N_48237,N_48394);
xnor UO_2314 (O_2314,N_48950,N_49935);
or UO_2315 (O_2315,N_48288,N_49261);
nor UO_2316 (O_2316,N_49652,N_49750);
nor UO_2317 (O_2317,N_48435,N_48014);
nor UO_2318 (O_2318,N_48965,N_49153);
xnor UO_2319 (O_2319,N_48883,N_49209);
nand UO_2320 (O_2320,N_48469,N_48735);
and UO_2321 (O_2321,N_48592,N_48111);
nand UO_2322 (O_2322,N_49115,N_49952);
and UO_2323 (O_2323,N_48272,N_48313);
nand UO_2324 (O_2324,N_49370,N_48287);
nand UO_2325 (O_2325,N_49932,N_49461);
nand UO_2326 (O_2326,N_49558,N_48163);
or UO_2327 (O_2327,N_49678,N_49042);
nor UO_2328 (O_2328,N_48804,N_49079);
xor UO_2329 (O_2329,N_48343,N_48697);
nor UO_2330 (O_2330,N_48781,N_49819);
and UO_2331 (O_2331,N_49214,N_49389);
nor UO_2332 (O_2332,N_48044,N_49096);
and UO_2333 (O_2333,N_49958,N_48696);
nor UO_2334 (O_2334,N_48874,N_48437);
nor UO_2335 (O_2335,N_48481,N_48419);
nor UO_2336 (O_2336,N_49669,N_49066);
nand UO_2337 (O_2337,N_49443,N_49081);
or UO_2338 (O_2338,N_48639,N_49811);
nor UO_2339 (O_2339,N_49734,N_49432);
nand UO_2340 (O_2340,N_49264,N_48029);
nor UO_2341 (O_2341,N_49331,N_48603);
nor UO_2342 (O_2342,N_49000,N_49888);
nand UO_2343 (O_2343,N_48901,N_48293);
nor UO_2344 (O_2344,N_49503,N_48853);
nor UO_2345 (O_2345,N_49993,N_48548);
or UO_2346 (O_2346,N_49957,N_49548);
nor UO_2347 (O_2347,N_48512,N_48943);
nor UO_2348 (O_2348,N_49849,N_48235);
nand UO_2349 (O_2349,N_48114,N_48372);
nor UO_2350 (O_2350,N_48459,N_48009);
or UO_2351 (O_2351,N_49180,N_48507);
nor UO_2352 (O_2352,N_49272,N_48101);
nor UO_2353 (O_2353,N_48675,N_48851);
xor UO_2354 (O_2354,N_49391,N_48298);
and UO_2355 (O_2355,N_48765,N_48554);
or UO_2356 (O_2356,N_49671,N_48852);
or UO_2357 (O_2357,N_49341,N_48551);
nor UO_2358 (O_2358,N_48745,N_49745);
and UO_2359 (O_2359,N_48505,N_48588);
nor UO_2360 (O_2360,N_48933,N_48389);
or UO_2361 (O_2361,N_49040,N_49082);
nor UO_2362 (O_2362,N_49861,N_49075);
nor UO_2363 (O_2363,N_49635,N_49758);
nor UO_2364 (O_2364,N_49802,N_49140);
and UO_2365 (O_2365,N_48416,N_48747);
or UO_2366 (O_2366,N_48737,N_49979);
or UO_2367 (O_2367,N_49484,N_48618);
or UO_2368 (O_2368,N_48160,N_48017);
nand UO_2369 (O_2369,N_49764,N_48781);
and UO_2370 (O_2370,N_48227,N_48178);
and UO_2371 (O_2371,N_49583,N_49917);
nand UO_2372 (O_2372,N_49772,N_49817);
nand UO_2373 (O_2373,N_49895,N_48996);
nor UO_2374 (O_2374,N_48845,N_49944);
or UO_2375 (O_2375,N_49153,N_49672);
nor UO_2376 (O_2376,N_48202,N_48837);
nand UO_2377 (O_2377,N_48210,N_48436);
or UO_2378 (O_2378,N_49798,N_49212);
nand UO_2379 (O_2379,N_49695,N_49918);
or UO_2380 (O_2380,N_48100,N_48805);
nand UO_2381 (O_2381,N_49565,N_49735);
nand UO_2382 (O_2382,N_48907,N_48458);
nor UO_2383 (O_2383,N_48078,N_49281);
and UO_2384 (O_2384,N_49028,N_48528);
xnor UO_2385 (O_2385,N_48176,N_49412);
and UO_2386 (O_2386,N_48207,N_48791);
or UO_2387 (O_2387,N_48354,N_48539);
or UO_2388 (O_2388,N_48730,N_48764);
nor UO_2389 (O_2389,N_48478,N_49202);
or UO_2390 (O_2390,N_48029,N_48216);
nand UO_2391 (O_2391,N_48080,N_49316);
and UO_2392 (O_2392,N_48407,N_49044);
and UO_2393 (O_2393,N_49788,N_48376);
or UO_2394 (O_2394,N_49026,N_49852);
nor UO_2395 (O_2395,N_48612,N_49413);
nor UO_2396 (O_2396,N_48909,N_49586);
and UO_2397 (O_2397,N_48826,N_49967);
nand UO_2398 (O_2398,N_48743,N_48253);
or UO_2399 (O_2399,N_49428,N_48747);
or UO_2400 (O_2400,N_49295,N_48577);
and UO_2401 (O_2401,N_48155,N_48011);
or UO_2402 (O_2402,N_48044,N_49856);
and UO_2403 (O_2403,N_48672,N_49824);
nand UO_2404 (O_2404,N_48079,N_48495);
nor UO_2405 (O_2405,N_49290,N_48826);
and UO_2406 (O_2406,N_49814,N_48940);
and UO_2407 (O_2407,N_49917,N_48181);
nor UO_2408 (O_2408,N_48242,N_49549);
and UO_2409 (O_2409,N_49306,N_48807);
nor UO_2410 (O_2410,N_48812,N_48947);
or UO_2411 (O_2411,N_48243,N_49183);
and UO_2412 (O_2412,N_48553,N_49157);
and UO_2413 (O_2413,N_48212,N_48435);
and UO_2414 (O_2414,N_48089,N_48864);
nand UO_2415 (O_2415,N_48851,N_49243);
or UO_2416 (O_2416,N_48640,N_48597);
or UO_2417 (O_2417,N_48824,N_49787);
or UO_2418 (O_2418,N_48879,N_49842);
nor UO_2419 (O_2419,N_48430,N_48652);
nand UO_2420 (O_2420,N_49544,N_48299);
nand UO_2421 (O_2421,N_48643,N_49322);
nand UO_2422 (O_2422,N_49019,N_49174);
and UO_2423 (O_2423,N_49748,N_49206);
nor UO_2424 (O_2424,N_48617,N_49283);
or UO_2425 (O_2425,N_49960,N_49763);
nand UO_2426 (O_2426,N_48448,N_48871);
nor UO_2427 (O_2427,N_49154,N_48741);
or UO_2428 (O_2428,N_49634,N_49097);
nand UO_2429 (O_2429,N_48384,N_49031);
or UO_2430 (O_2430,N_49891,N_48195);
and UO_2431 (O_2431,N_48070,N_48573);
or UO_2432 (O_2432,N_48437,N_49502);
or UO_2433 (O_2433,N_48027,N_49807);
and UO_2434 (O_2434,N_49038,N_49744);
nand UO_2435 (O_2435,N_48307,N_49790);
nand UO_2436 (O_2436,N_48109,N_49157);
nand UO_2437 (O_2437,N_48943,N_48897);
nand UO_2438 (O_2438,N_48044,N_48917);
or UO_2439 (O_2439,N_48029,N_48816);
nand UO_2440 (O_2440,N_48514,N_48516);
or UO_2441 (O_2441,N_49573,N_49178);
xnor UO_2442 (O_2442,N_49989,N_49841);
nand UO_2443 (O_2443,N_49865,N_49183);
and UO_2444 (O_2444,N_48284,N_48818);
nand UO_2445 (O_2445,N_49868,N_48512);
nor UO_2446 (O_2446,N_49441,N_49342);
nand UO_2447 (O_2447,N_48352,N_49634);
or UO_2448 (O_2448,N_48880,N_48175);
or UO_2449 (O_2449,N_48834,N_49992);
nor UO_2450 (O_2450,N_48614,N_49186);
and UO_2451 (O_2451,N_49697,N_48532);
nand UO_2452 (O_2452,N_48126,N_49395);
nor UO_2453 (O_2453,N_49010,N_48485);
nand UO_2454 (O_2454,N_49984,N_48509);
and UO_2455 (O_2455,N_48780,N_48111);
nor UO_2456 (O_2456,N_48941,N_48042);
nor UO_2457 (O_2457,N_49188,N_49779);
and UO_2458 (O_2458,N_48979,N_49064);
and UO_2459 (O_2459,N_48391,N_49768);
and UO_2460 (O_2460,N_48228,N_48175);
and UO_2461 (O_2461,N_48997,N_49629);
or UO_2462 (O_2462,N_48948,N_49559);
or UO_2463 (O_2463,N_48793,N_49556);
and UO_2464 (O_2464,N_49619,N_49164);
or UO_2465 (O_2465,N_48594,N_49291);
and UO_2466 (O_2466,N_48257,N_49614);
nor UO_2467 (O_2467,N_49664,N_49317);
nand UO_2468 (O_2468,N_49088,N_48601);
and UO_2469 (O_2469,N_48284,N_49844);
or UO_2470 (O_2470,N_49742,N_49090);
or UO_2471 (O_2471,N_49973,N_48862);
nor UO_2472 (O_2472,N_49068,N_49725);
nand UO_2473 (O_2473,N_49480,N_48569);
nor UO_2474 (O_2474,N_49074,N_48805);
nand UO_2475 (O_2475,N_49028,N_48848);
or UO_2476 (O_2476,N_48190,N_48492);
or UO_2477 (O_2477,N_48572,N_48150);
nand UO_2478 (O_2478,N_49578,N_48199);
nand UO_2479 (O_2479,N_48120,N_49460);
or UO_2480 (O_2480,N_48582,N_48264);
or UO_2481 (O_2481,N_49067,N_48148);
nand UO_2482 (O_2482,N_49416,N_48286);
nand UO_2483 (O_2483,N_49004,N_48128);
nor UO_2484 (O_2484,N_48433,N_49468);
nor UO_2485 (O_2485,N_49004,N_48146);
or UO_2486 (O_2486,N_49782,N_49270);
or UO_2487 (O_2487,N_49246,N_49458);
nor UO_2488 (O_2488,N_49442,N_48432);
nor UO_2489 (O_2489,N_49807,N_49283);
nand UO_2490 (O_2490,N_48594,N_49460);
nand UO_2491 (O_2491,N_49350,N_49234);
nand UO_2492 (O_2492,N_49204,N_48176);
nor UO_2493 (O_2493,N_48385,N_49772);
and UO_2494 (O_2494,N_48158,N_48264);
nor UO_2495 (O_2495,N_48741,N_48394);
nor UO_2496 (O_2496,N_48102,N_49841);
nor UO_2497 (O_2497,N_48770,N_48439);
nor UO_2498 (O_2498,N_49578,N_48418);
xnor UO_2499 (O_2499,N_49402,N_48946);
or UO_2500 (O_2500,N_49353,N_48149);
and UO_2501 (O_2501,N_48731,N_49870);
and UO_2502 (O_2502,N_49677,N_49941);
nor UO_2503 (O_2503,N_49802,N_49075);
and UO_2504 (O_2504,N_49851,N_48565);
or UO_2505 (O_2505,N_48929,N_49875);
nor UO_2506 (O_2506,N_48455,N_48616);
and UO_2507 (O_2507,N_48111,N_48591);
and UO_2508 (O_2508,N_49185,N_49203);
nor UO_2509 (O_2509,N_48920,N_49832);
or UO_2510 (O_2510,N_48079,N_49958);
nand UO_2511 (O_2511,N_48104,N_48997);
and UO_2512 (O_2512,N_49341,N_49809);
nor UO_2513 (O_2513,N_48086,N_49649);
nand UO_2514 (O_2514,N_49133,N_49554);
nand UO_2515 (O_2515,N_48430,N_48897);
and UO_2516 (O_2516,N_49382,N_49716);
or UO_2517 (O_2517,N_49523,N_49251);
or UO_2518 (O_2518,N_48174,N_49947);
or UO_2519 (O_2519,N_49359,N_49546);
nand UO_2520 (O_2520,N_49713,N_48164);
or UO_2521 (O_2521,N_49042,N_49053);
nor UO_2522 (O_2522,N_48905,N_48827);
and UO_2523 (O_2523,N_48939,N_48322);
nor UO_2524 (O_2524,N_48138,N_48084);
xor UO_2525 (O_2525,N_49811,N_48190);
nand UO_2526 (O_2526,N_48676,N_48315);
and UO_2527 (O_2527,N_48374,N_49895);
or UO_2528 (O_2528,N_49190,N_49282);
nor UO_2529 (O_2529,N_49152,N_48053);
or UO_2530 (O_2530,N_48243,N_49479);
nor UO_2531 (O_2531,N_48159,N_49177);
nor UO_2532 (O_2532,N_49466,N_49130);
and UO_2533 (O_2533,N_49329,N_48705);
nand UO_2534 (O_2534,N_49287,N_49465);
or UO_2535 (O_2535,N_48057,N_48981);
nand UO_2536 (O_2536,N_49446,N_49180);
nand UO_2537 (O_2537,N_49196,N_49094);
nor UO_2538 (O_2538,N_48854,N_48957);
and UO_2539 (O_2539,N_49623,N_49374);
nand UO_2540 (O_2540,N_49202,N_48814);
nand UO_2541 (O_2541,N_49830,N_49339);
or UO_2542 (O_2542,N_48667,N_49940);
nand UO_2543 (O_2543,N_49168,N_48335);
or UO_2544 (O_2544,N_49009,N_49127);
or UO_2545 (O_2545,N_48082,N_49613);
nand UO_2546 (O_2546,N_48736,N_48698);
and UO_2547 (O_2547,N_49918,N_49787);
and UO_2548 (O_2548,N_48665,N_48317);
nor UO_2549 (O_2549,N_49322,N_49895);
nor UO_2550 (O_2550,N_48378,N_49093);
and UO_2551 (O_2551,N_49866,N_49765);
and UO_2552 (O_2552,N_49337,N_49427);
nor UO_2553 (O_2553,N_49456,N_48044);
nand UO_2554 (O_2554,N_49446,N_48678);
or UO_2555 (O_2555,N_49821,N_48342);
or UO_2556 (O_2556,N_48800,N_49914);
nand UO_2557 (O_2557,N_48763,N_49106);
and UO_2558 (O_2558,N_48593,N_49562);
nand UO_2559 (O_2559,N_48347,N_48555);
nand UO_2560 (O_2560,N_49481,N_49103);
nand UO_2561 (O_2561,N_49560,N_49250);
and UO_2562 (O_2562,N_48220,N_49940);
and UO_2563 (O_2563,N_49367,N_48017);
and UO_2564 (O_2564,N_49221,N_49809);
or UO_2565 (O_2565,N_49251,N_49071);
and UO_2566 (O_2566,N_49123,N_49605);
or UO_2567 (O_2567,N_48337,N_48438);
or UO_2568 (O_2568,N_49763,N_49974);
or UO_2569 (O_2569,N_48735,N_49359);
and UO_2570 (O_2570,N_48485,N_48634);
and UO_2571 (O_2571,N_48313,N_48301);
and UO_2572 (O_2572,N_48906,N_48220);
or UO_2573 (O_2573,N_48177,N_48409);
or UO_2574 (O_2574,N_49885,N_49839);
nand UO_2575 (O_2575,N_48456,N_48100);
and UO_2576 (O_2576,N_48406,N_48518);
or UO_2577 (O_2577,N_49852,N_48469);
and UO_2578 (O_2578,N_49518,N_49739);
nor UO_2579 (O_2579,N_49971,N_48642);
nor UO_2580 (O_2580,N_49048,N_49812);
and UO_2581 (O_2581,N_48083,N_49275);
or UO_2582 (O_2582,N_49915,N_49626);
and UO_2583 (O_2583,N_48598,N_48081);
nor UO_2584 (O_2584,N_49851,N_48621);
nand UO_2585 (O_2585,N_49621,N_49427);
and UO_2586 (O_2586,N_49937,N_48225);
nand UO_2587 (O_2587,N_48781,N_49229);
and UO_2588 (O_2588,N_48340,N_48993);
and UO_2589 (O_2589,N_48375,N_49841);
or UO_2590 (O_2590,N_48512,N_48493);
or UO_2591 (O_2591,N_49520,N_49282);
and UO_2592 (O_2592,N_49465,N_48125);
or UO_2593 (O_2593,N_48661,N_48222);
nand UO_2594 (O_2594,N_49076,N_48133);
nor UO_2595 (O_2595,N_48721,N_48052);
nor UO_2596 (O_2596,N_49063,N_49083);
and UO_2597 (O_2597,N_49602,N_49629);
and UO_2598 (O_2598,N_48582,N_48838);
nor UO_2599 (O_2599,N_48409,N_48482);
nand UO_2600 (O_2600,N_49442,N_49801);
or UO_2601 (O_2601,N_48233,N_48265);
or UO_2602 (O_2602,N_48562,N_48321);
and UO_2603 (O_2603,N_48386,N_48364);
xor UO_2604 (O_2604,N_49701,N_48478);
or UO_2605 (O_2605,N_48845,N_49045);
nor UO_2606 (O_2606,N_49998,N_49967);
nand UO_2607 (O_2607,N_49444,N_48694);
or UO_2608 (O_2608,N_49779,N_48773);
and UO_2609 (O_2609,N_48607,N_49048);
and UO_2610 (O_2610,N_49501,N_48734);
and UO_2611 (O_2611,N_49941,N_48241);
or UO_2612 (O_2612,N_49846,N_48377);
nand UO_2613 (O_2613,N_49155,N_49862);
nand UO_2614 (O_2614,N_49497,N_48411);
nand UO_2615 (O_2615,N_49819,N_49769);
or UO_2616 (O_2616,N_48098,N_48836);
and UO_2617 (O_2617,N_49098,N_49344);
nand UO_2618 (O_2618,N_49624,N_49198);
nor UO_2619 (O_2619,N_49871,N_49248);
xor UO_2620 (O_2620,N_48551,N_48335);
nand UO_2621 (O_2621,N_49126,N_49467);
and UO_2622 (O_2622,N_48272,N_49243);
nor UO_2623 (O_2623,N_49107,N_48504);
nor UO_2624 (O_2624,N_48960,N_49519);
nor UO_2625 (O_2625,N_48640,N_48641);
nand UO_2626 (O_2626,N_49892,N_49816);
nand UO_2627 (O_2627,N_49329,N_49063);
and UO_2628 (O_2628,N_49840,N_48776);
nor UO_2629 (O_2629,N_49293,N_49616);
or UO_2630 (O_2630,N_49982,N_49742);
or UO_2631 (O_2631,N_48490,N_48561);
or UO_2632 (O_2632,N_49651,N_49658);
or UO_2633 (O_2633,N_49488,N_48606);
or UO_2634 (O_2634,N_49486,N_48689);
nor UO_2635 (O_2635,N_48127,N_48895);
and UO_2636 (O_2636,N_49748,N_48349);
and UO_2637 (O_2637,N_49514,N_49753);
and UO_2638 (O_2638,N_49334,N_49426);
and UO_2639 (O_2639,N_49089,N_48244);
nor UO_2640 (O_2640,N_48115,N_48307);
or UO_2641 (O_2641,N_49793,N_49644);
nor UO_2642 (O_2642,N_49880,N_49980);
nand UO_2643 (O_2643,N_48527,N_49984);
nand UO_2644 (O_2644,N_49772,N_49438);
or UO_2645 (O_2645,N_49452,N_49711);
nor UO_2646 (O_2646,N_48551,N_48309);
nand UO_2647 (O_2647,N_49861,N_48943);
nand UO_2648 (O_2648,N_49636,N_49075);
and UO_2649 (O_2649,N_49756,N_49171);
nor UO_2650 (O_2650,N_48911,N_49389);
nor UO_2651 (O_2651,N_49368,N_49358);
and UO_2652 (O_2652,N_48507,N_48315);
nor UO_2653 (O_2653,N_49984,N_48561);
nor UO_2654 (O_2654,N_49016,N_49769);
and UO_2655 (O_2655,N_49550,N_49731);
nand UO_2656 (O_2656,N_48617,N_48027);
and UO_2657 (O_2657,N_48712,N_49824);
nand UO_2658 (O_2658,N_48448,N_48238);
or UO_2659 (O_2659,N_49473,N_49529);
nand UO_2660 (O_2660,N_49569,N_48485);
nor UO_2661 (O_2661,N_48953,N_48543);
nor UO_2662 (O_2662,N_48981,N_48833);
nor UO_2663 (O_2663,N_49518,N_48987);
nand UO_2664 (O_2664,N_48881,N_48940);
or UO_2665 (O_2665,N_48876,N_48473);
xnor UO_2666 (O_2666,N_49816,N_49993);
or UO_2667 (O_2667,N_48043,N_48559);
or UO_2668 (O_2668,N_48157,N_48870);
or UO_2669 (O_2669,N_49677,N_48845);
nand UO_2670 (O_2670,N_49889,N_49626);
or UO_2671 (O_2671,N_49119,N_49225);
or UO_2672 (O_2672,N_48410,N_48739);
nor UO_2673 (O_2673,N_49439,N_48757);
and UO_2674 (O_2674,N_49593,N_49285);
or UO_2675 (O_2675,N_48523,N_49892);
nor UO_2676 (O_2676,N_49733,N_49879);
nor UO_2677 (O_2677,N_48116,N_48372);
nand UO_2678 (O_2678,N_48144,N_49304);
nand UO_2679 (O_2679,N_48512,N_48552);
and UO_2680 (O_2680,N_49147,N_48322);
xor UO_2681 (O_2681,N_49877,N_49720);
and UO_2682 (O_2682,N_49552,N_49953);
nor UO_2683 (O_2683,N_48655,N_48521);
or UO_2684 (O_2684,N_49032,N_48600);
xnor UO_2685 (O_2685,N_49681,N_48543);
nand UO_2686 (O_2686,N_48444,N_48998);
nand UO_2687 (O_2687,N_48967,N_48526);
or UO_2688 (O_2688,N_49793,N_48155);
and UO_2689 (O_2689,N_48686,N_49465);
nand UO_2690 (O_2690,N_49095,N_48760);
or UO_2691 (O_2691,N_49273,N_48165);
nor UO_2692 (O_2692,N_48774,N_48906);
or UO_2693 (O_2693,N_49828,N_49567);
nand UO_2694 (O_2694,N_49421,N_48335);
nor UO_2695 (O_2695,N_49562,N_49565);
or UO_2696 (O_2696,N_48564,N_48853);
and UO_2697 (O_2697,N_49142,N_48810);
or UO_2698 (O_2698,N_49022,N_49284);
nand UO_2699 (O_2699,N_49785,N_48398);
nor UO_2700 (O_2700,N_49131,N_49804);
or UO_2701 (O_2701,N_49602,N_49426);
nor UO_2702 (O_2702,N_48986,N_49560);
and UO_2703 (O_2703,N_49366,N_48553);
nor UO_2704 (O_2704,N_49469,N_49558);
nor UO_2705 (O_2705,N_48805,N_48980);
or UO_2706 (O_2706,N_49662,N_49029);
and UO_2707 (O_2707,N_49779,N_49025);
and UO_2708 (O_2708,N_49456,N_48106);
nand UO_2709 (O_2709,N_49166,N_49569);
nand UO_2710 (O_2710,N_49523,N_49629);
nand UO_2711 (O_2711,N_48200,N_49964);
nor UO_2712 (O_2712,N_49198,N_49054);
or UO_2713 (O_2713,N_48899,N_48874);
or UO_2714 (O_2714,N_48809,N_48104);
and UO_2715 (O_2715,N_49631,N_48799);
nand UO_2716 (O_2716,N_49256,N_48331);
and UO_2717 (O_2717,N_49590,N_49885);
nor UO_2718 (O_2718,N_48426,N_49774);
and UO_2719 (O_2719,N_48484,N_49066);
and UO_2720 (O_2720,N_49534,N_48222);
xnor UO_2721 (O_2721,N_49155,N_48056);
or UO_2722 (O_2722,N_49157,N_48244);
or UO_2723 (O_2723,N_48153,N_49898);
or UO_2724 (O_2724,N_49469,N_48365);
nor UO_2725 (O_2725,N_48723,N_48609);
or UO_2726 (O_2726,N_49797,N_49686);
nor UO_2727 (O_2727,N_49966,N_48721);
nand UO_2728 (O_2728,N_49146,N_48626);
nand UO_2729 (O_2729,N_48272,N_49423);
nor UO_2730 (O_2730,N_48085,N_49499);
or UO_2731 (O_2731,N_49680,N_48123);
and UO_2732 (O_2732,N_48129,N_48152);
xor UO_2733 (O_2733,N_49972,N_49150);
and UO_2734 (O_2734,N_48918,N_48163);
nor UO_2735 (O_2735,N_49433,N_49091);
and UO_2736 (O_2736,N_49620,N_48358);
or UO_2737 (O_2737,N_49186,N_49552);
nand UO_2738 (O_2738,N_48799,N_49832);
xor UO_2739 (O_2739,N_48482,N_48985);
nor UO_2740 (O_2740,N_49280,N_48448);
and UO_2741 (O_2741,N_49770,N_49031);
or UO_2742 (O_2742,N_49636,N_48774);
and UO_2743 (O_2743,N_48148,N_49248);
nor UO_2744 (O_2744,N_48138,N_49980);
nand UO_2745 (O_2745,N_48737,N_49967);
nand UO_2746 (O_2746,N_49538,N_48475);
and UO_2747 (O_2747,N_48471,N_48930);
and UO_2748 (O_2748,N_48761,N_48704);
nand UO_2749 (O_2749,N_48661,N_48549);
and UO_2750 (O_2750,N_48698,N_49511);
and UO_2751 (O_2751,N_49758,N_49955);
or UO_2752 (O_2752,N_49720,N_48249);
or UO_2753 (O_2753,N_49728,N_49508);
nor UO_2754 (O_2754,N_49696,N_49311);
nand UO_2755 (O_2755,N_48318,N_49253);
xnor UO_2756 (O_2756,N_49654,N_48916);
or UO_2757 (O_2757,N_48882,N_48675);
nand UO_2758 (O_2758,N_48199,N_49461);
or UO_2759 (O_2759,N_49167,N_48361);
nand UO_2760 (O_2760,N_49753,N_49117);
or UO_2761 (O_2761,N_49860,N_48417);
nand UO_2762 (O_2762,N_48417,N_48222);
nor UO_2763 (O_2763,N_49629,N_49470);
and UO_2764 (O_2764,N_49386,N_49365);
or UO_2765 (O_2765,N_49229,N_49194);
nor UO_2766 (O_2766,N_48421,N_49385);
nor UO_2767 (O_2767,N_48018,N_49889);
or UO_2768 (O_2768,N_49920,N_49481);
nand UO_2769 (O_2769,N_49106,N_48235);
and UO_2770 (O_2770,N_49008,N_48928);
nand UO_2771 (O_2771,N_49420,N_49991);
nand UO_2772 (O_2772,N_49271,N_49968);
or UO_2773 (O_2773,N_49740,N_49652);
or UO_2774 (O_2774,N_48458,N_49884);
or UO_2775 (O_2775,N_49839,N_49133);
nor UO_2776 (O_2776,N_49515,N_48325);
nand UO_2777 (O_2777,N_49242,N_48612);
xor UO_2778 (O_2778,N_48461,N_49560);
and UO_2779 (O_2779,N_48869,N_49616);
nor UO_2780 (O_2780,N_48669,N_48292);
nand UO_2781 (O_2781,N_49151,N_48771);
or UO_2782 (O_2782,N_49756,N_48633);
or UO_2783 (O_2783,N_49252,N_49807);
and UO_2784 (O_2784,N_49602,N_49845);
xor UO_2785 (O_2785,N_49304,N_49810);
or UO_2786 (O_2786,N_49372,N_49287);
nand UO_2787 (O_2787,N_49356,N_48186);
and UO_2788 (O_2788,N_48531,N_49513);
or UO_2789 (O_2789,N_49736,N_48292);
or UO_2790 (O_2790,N_48406,N_48645);
and UO_2791 (O_2791,N_49166,N_48113);
and UO_2792 (O_2792,N_49086,N_49383);
nand UO_2793 (O_2793,N_49187,N_48169);
nand UO_2794 (O_2794,N_49979,N_48419);
nor UO_2795 (O_2795,N_48890,N_49802);
or UO_2796 (O_2796,N_48752,N_49714);
nor UO_2797 (O_2797,N_49316,N_48188);
nor UO_2798 (O_2798,N_48980,N_49248);
nor UO_2799 (O_2799,N_49971,N_48610);
or UO_2800 (O_2800,N_48306,N_48184);
or UO_2801 (O_2801,N_49335,N_48196);
nor UO_2802 (O_2802,N_48882,N_49684);
and UO_2803 (O_2803,N_49262,N_48001);
and UO_2804 (O_2804,N_48696,N_49357);
or UO_2805 (O_2805,N_48384,N_49538);
and UO_2806 (O_2806,N_48008,N_48388);
nand UO_2807 (O_2807,N_49870,N_48304);
or UO_2808 (O_2808,N_48602,N_48990);
and UO_2809 (O_2809,N_49768,N_48220);
nor UO_2810 (O_2810,N_49127,N_49586);
and UO_2811 (O_2811,N_48597,N_49008);
nor UO_2812 (O_2812,N_48950,N_48621);
or UO_2813 (O_2813,N_48525,N_48873);
nor UO_2814 (O_2814,N_48223,N_49739);
or UO_2815 (O_2815,N_48285,N_48737);
nand UO_2816 (O_2816,N_49026,N_48103);
or UO_2817 (O_2817,N_48409,N_49731);
xnor UO_2818 (O_2818,N_49612,N_49006);
and UO_2819 (O_2819,N_49788,N_48499);
or UO_2820 (O_2820,N_49120,N_48832);
nor UO_2821 (O_2821,N_49044,N_49825);
or UO_2822 (O_2822,N_48425,N_49963);
or UO_2823 (O_2823,N_49820,N_49565);
nor UO_2824 (O_2824,N_49121,N_48462);
and UO_2825 (O_2825,N_48776,N_48669);
and UO_2826 (O_2826,N_48140,N_48098);
or UO_2827 (O_2827,N_48866,N_49366);
nand UO_2828 (O_2828,N_48483,N_48076);
or UO_2829 (O_2829,N_49368,N_48622);
nand UO_2830 (O_2830,N_49932,N_49933);
xnor UO_2831 (O_2831,N_49077,N_49111);
or UO_2832 (O_2832,N_48132,N_48585);
nor UO_2833 (O_2833,N_49809,N_49664);
nand UO_2834 (O_2834,N_49542,N_49069);
nand UO_2835 (O_2835,N_49308,N_48012);
or UO_2836 (O_2836,N_48951,N_49117);
or UO_2837 (O_2837,N_49190,N_49049);
nand UO_2838 (O_2838,N_49849,N_48523);
nor UO_2839 (O_2839,N_48427,N_49855);
or UO_2840 (O_2840,N_49723,N_49541);
and UO_2841 (O_2841,N_49570,N_49536);
nor UO_2842 (O_2842,N_48366,N_49175);
and UO_2843 (O_2843,N_49400,N_48480);
or UO_2844 (O_2844,N_49535,N_48966);
or UO_2845 (O_2845,N_49291,N_49362);
nor UO_2846 (O_2846,N_49355,N_48440);
nor UO_2847 (O_2847,N_48758,N_49464);
or UO_2848 (O_2848,N_49535,N_49172);
or UO_2849 (O_2849,N_49610,N_49182);
or UO_2850 (O_2850,N_48539,N_49625);
nor UO_2851 (O_2851,N_48097,N_49215);
nand UO_2852 (O_2852,N_49584,N_48184);
and UO_2853 (O_2853,N_48629,N_49251);
or UO_2854 (O_2854,N_48748,N_48520);
nand UO_2855 (O_2855,N_49924,N_48558);
and UO_2856 (O_2856,N_49803,N_48168);
nand UO_2857 (O_2857,N_48104,N_48196);
xor UO_2858 (O_2858,N_48479,N_48489);
nor UO_2859 (O_2859,N_48981,N_49086);
nand UO_2860 (O_2860,N_49017,N_48526);
nand UO_2861 (O_2861,N_49607,N_48440);
and UO_2862 (O_2862,N_48376,N_48413);
nand UO_2863 (O_2863,N_49513,N_48726);
or UO_2864 (O_2864,N_48445,N_49194);
nor UO_2865 (O_2865,N_48056,N_49801);
nand UO_2866 (O_2866,N_49662,N_49701);
and UO_2867 (O_2867,N_48188,N_49472);
and UO_2868 (O_2868,N_49603,N_48349);
nand UO_2869 (O_2869,N_49072,N_49974);
and UO_2870 (O_2870,N_48701,N_48741);
or UO_2871 (O_2871,N_48283,N_48795);
and UO_2872 (O_2872,N_48427,N_48817);
or UO_2873 (O_2873,N_48072,N_48036);
or UO_2874 (O_2874,N_48898,N_49278);
or UO_2875 (O_2875,N_49947,N_49739);
or UO_2876 (O_2876,N_49220,N_48963);
or UO_2877 (O_2877,N_49262,N_48773);
nand UO_2878 (O_2878,N_49918,N_48780);
nand UO_2879 (O_2879,N_48189,N_49452);
or UO_2880 (O_2880,N_48075,N_49982);
nand UO_2881 (O_2881,N_48159,N_49577);
or UO_2882 (O_2882,N_48991,N_49005);
and UO_2883 (O_2883,N_48638,N_48549);
nor UO_2884 (O_2884,N_49841,N_48520);
or UO_2885 (O_2885,N_49247,N_48790);
or UO_2886 (O_2886,N_48665,N_48149);
nor UO_2887 (O_2887,N_49745,N_49325);
or UO_2888 (O_2888,N_49353,N_49127);
and UO_2889 (O_2889,N_49055,N_48398);
nor UO_2890 (O_2890,N_49673,N_48211);
nor UO_2891 (O_2891,N_49151,N_49801);
nand UO_2892 (O_2892,N_48158,N_49415);
and UO_2893 (O_2893,N_49081,N_49712);
nor UO_2894 (O_2894,N_48451,N_49878);
nor UO_2895 (O_2895,N_49421,N_48032);
or UO_2896 (O_2896,N_48909,N_49619);
xnor UO_2897 (O_2897,N_48444,N_48879);
and UO_2898 (O_2898,N_49503,N_49615);
or UO_2899 (O_2899,N_48871,N_48558);
nand UO_2900 (O_2900,N_48981,N_49606);
or UO_2901 (O_2901,N_48097,N_48465);
and UO_2902 (O_2902,N_49314,N_49127);
nand UO_2903 (O_2903,N_49988,N_48028);
or UO_2904 (O_2904,N_49097,N_49194);
nor UO_2905 (O_2905,N_48811,N_49259);
and UO_2906 (O_2906,N_48731,N_49077);
and UO_2907 (O_2907,N_48237,N_48757);
nor UO_2908 (O_2908,N_49266,N_49319);
and UO_2909 (O_2909,N_49017,N_49150);
nor UO_2910 (O_2910,N_48001,N_49477);
or UO_2911 (O_2911,N_49694,N_49925);
and UO_2912 (O_2912,N_48618,N_49275);
or UO_2913 (O_2913,N_48982,N_49828);
and UO_2914 (O_2914,N_49735,N_49432);
nand UO_2915 (O_2915,N_49381,N_49075);
nand UO_2916 (O_2916,N_49335,N_49356);
nand UO_2917 (O_2917,N_49377,N_49879);
nor UO_2918 (O_2918,N_49467,N_49107);
nand UO_2919 (O_2919,N_48097,N_48702);
and UO_2920 (O_2920,N_48792,N_48768);
nand UO_2921 (O_2921,N_49055,N_49277);
nand UO_2922 (O_2922,N_49561,N_49975);
nand UO_2923 (O_2923,N_48544,N_48302);
nor UO_2924 (O_2924,N_49750,N_48698);
nor UO_2925 (O_2925,N_49334,N_48305);
or UO_2926 (O_2926,N_48623,N_48633);
or UO_2927 (O_2927,N_49947,N_48338);
nor UO_2928 (O_2928,N_48395,N_48114);
or UO_2929 (O_2929,N_48614,N_49628);
and UO_2930 (O_2930,N_48146,N_49299);
nor UO_2931 (O_2931,N_48194,N_49347);
or UO_2932 (O_2932,N_48231,N_49937);
nand UO_2933 (O_2933,N_48250,N_48265);
or UO_2934 (O_2934,N_48882,N_48494);
nor UO_2935 (O_2935,N_48658,N_48927);
nor UO_2936 (O_2936,N_49342,N_48980);
and UO_2937 (O_2937,N_49223,N_48507);
or UO_2938 (O_2938,N_48403,N_49236);
nor UO_2939 (O_2939,N_49590,N_48039);
nand UO_2940 (O_2940,N_48242,N_49080);
xor UO_2941 (O_2941,N_49633,N_49148);
nor UO_2942 (O_2942,N_49599,N_49881);
and UO_2943 (O_2943,N_48443,N_49429);
nor UO_2944 (O_2944,N_48277,N_49232);
and UO_2945 (O_2945,N_49246,N_49572);
or UO_2946 (O_2946,N_48907,N_49593);
nor UO_2947 (O_2947,N_48037,N_48047);
and UO_2948 (O_2948,N_48059,N_48866);
or UO_2949 (O_2949,N_49099,N_48137);
nor UO_2950 (O_2950,N_48208,N_48402);
and UO_2951 (O_2951,N_48744,N_49027);
or UO_2952 (O_2952,N_49864,N_49600);
nand UO_2953 (O_2953,N_49949,N_49964);
nor UO_2954 (O_2954,N_49973,N_48157);
nand UO_2955 (O_2955,N_48981,N_49446);
or UO_2956 (O_2956,N_48409,N_49982);
and UO_2957 (O_2957,N_48651,N_48720);
and UO_2958 (O_2958,N_48698,N_48102);
nor UO_2959 (O_2959,N_49979,N_49990);
nor UO_2960 (O_2960,N_49799,N_48745);
nand UO_2961 (O_2961,N_48743,N_49852);
and UO_2962 (O_2962,N_49695,N_49156);
xnor UO_2963 (O_2963,N_49049,N_48149);
or UO_2964 (O_2964,N_48006,N_49369);
or UO_2965 (O_2965,N_48050,N_49934);
or UO_2966 (O_2966,N_49583,N_48069);
nor UO_2967 (O_2967,N_48621,N_49678);
nand UO_2968 (O_2968,N_49901,N_48441);
nand UO_2969 (O_2969,N_48123,N_49954);
and UO_2970 (O_2970,N_49223,N_48587);
nand UO_2971 (O_2971,N_48915,N_49709);
nor UO_2972 (O_2972,N_49803,N_48999);
and UO_2973 (O_2973,N_48218,N_49856);
or UO_2974 (O_2974,N_49966,N_48879);
or UO_2975 (O_2975,N_49800,N_48952);
nand UO_2976 (O_2976,N_49710,N_48815);
nor UO_2977 (O_2977,N_48801,N_48683);
and UO_2978 (O_2978,N_49876,N_49221);
or UO_2979 (O_2979,N_49012,N_49315);
nor UO_2980 (O_2980,N_48374,N_49879);
nand UO_2981 (O_2981,N_48988,N_49238);
or UO_2982 (O_2982,N_49436,N_48350);
nor UO_2983 (O_2983,N_49309,N_48706);
nor UO_2984 (O_2984,N_48413,N_48763);
or UO_2985 (O_2985,N_48435,N_48736);
xor UO_2986 (O_2986,N_48562,N_49721);
nor UO_2987 (O_2987,N_49466,N_49125);
or UO_2988 (O_2988,N_49284,N_48910);
or UO_2989 (O_2989,N_48734,N_49261);
nor UO_2990 (O_2990,N_48211,N_48139);
nand UO_2991 (O_2991,N_48949,N_48552);
nand UO_2992 (O_2992,N_48563,N_49447);
nor UO_2993 (O_2993,N_49516,N_49150);
nor UO_2994 (O_2994,N_48897,N_48747);
nor UO_2995 (O_2995,N_49558,N_49482);
nor UO_2996 (O_2996,N_49612,N_49776);
or UO_2997 (O_2997,N_48241,N_49342);
nor UO_2998 (O_2998,N_49681,N_49781);
or UO_2999 (O_2999,N_49872,N_49423);
nor UO_3000 (O_3000,N_48480,N_48342);
and UO_3001 (O_3001,N_48169,N_49889);
and UO_3002 (O_3002,N_49428,N_48655);
and UO_3003 (O_3003,N_48376,N_49007);
nor UO_3004 (O_3004,N_48461,N_48289);
nand UO_3005 (O_3005,N_49450,N_49012);
nand UO_3006 (O_3006,N_48273,N_49680);
nor UO_3007 (O_3007,N_49601,N_48386);
xnor UO_3008 (O_3008,N_49807,N_49766);
nand UO_3009 (O_3009,N_48305,N_48737);
nor UO_3010 (O_3010,N_49063,N_49218);
or UO_3011 (O_3011,N_49311,N_49575);
nor UO_3012 (O_3012,N_49016,N_49612);
nor UO_3013 (O_3013,N_48720,N_48012);
nor UO_3014 (O_3014,N_49715,N_48256);
or UO_3015 (O_3015,N_48978,N_48222);
or UO_3016 (O_3016,N_49312,N_49719);
and UO_3017 (O_3017,N_49232,N_49478);
or UO_3018 (O_3018,N_48506,N_49841);
nand UO_3019 (O_3019,N_49444,N_49538);
nor UO_3020 (O_3020,N_48704,N_49150);
and UO_3021 (O_3021,N_48996,N_49660);
and UO_3022 (O_3022,N_48042,N_49132);
and UO_3023 (O_3023,N_49468,N_48905);
nor UO_3024 (O_3024,N_48593,N_49460);
nand UO_3025 (O_3025,N_48623,N_48565);
or UO_3026 (O_3026,N_49412,N_49797);
and UO_3027 (O_3027,N_48247,N_48365);
or UO_3028 (O_3028,N_49810,N_49556);
nand UO_3029 (O_3029,N_48497,N_48163);
and UO_3030 (O_3030,N_48693,N_49193);
and UO_3031 (O_3031,N_49481,N_48223);
nand UO_3032 (O_3032,N_48018,N_48097);
and UO_3033 (O_3033,N_49426,N_48375);
or UO_3034 (O_3034,N_48800,N_48450);
and UO_3035 (O_3035,N_48299,N_49521);
nand UO_3036 (O_3036,N_48888,N_49814);
nor UO_3037 (O_3037,N_48136,N_49006);
nand UO_3038 (O_3038,N_49506,N_49668);
and UO_3039 (O_3039,N_48279,N_48739);
nor UO_3040 (O_3040,N_49868,N_48511);
or UO_3041 (O_3041,N_48536,N_49464);
nand UO_3042 (O_3042,N_49090,N_49592);
nand UO_3043 (O_3043,N_48337,N_49601);
or UO_3044 (O_3044,N_49300,N_48494);
nor UO_3045 (O_3045,N_48577,N_49708);
and UO_3046 (O_3046,N_49522,N_48821);
nand UO_3047 (O_3047,N_49146,N_48047);
nand UO_3048 (O_3048,N_49108,N_49680);
and UO_3049 (O_3049,N_49161,N_49343);
nand UO_3050 (O_3050,N_49621,N_48729);
and UO_3051 (O_3051,N_49172,N_48045);
nand UO_3052 (O_3052,N_49292,N_49383);
or UO_3053 (O_3053,N_48291,N_48971);
and UO_3054 (O_3054,N_49456,N_48526);
or UO_3055 (O_3055,N_48058,N_48942);
nand UO_3056 (O_3056,N_48957,N_48402);
or UO_3057 (O_3057,N_48393,N_48416);
nor UO_3058 (O_3058,N_48701,N_48926);
nor UO_3059 (O_3059,N_49025,N_49596);
or UO_3060 (O_3060,N_48487,N_48450);
or UO_3061 (O_3061,N_49001,N_48337);
or UO_3062 (O_3062,N_48852,N_49142);
or UO_3063 (O_3063,N_49341,N_48083);
or UO_3064 (O_3064,N_48290,N_49498);
nand UO_3065 (O_3065,N_48312,N_48041);
or UO_3066 (O_3066,N_48393,N_48978);
nand UO_3067 (O_3067,N_48781,N_49520);
or UO_3068 (O_3068,N_48660,N_49697);
nor UO_3069 (O_3069,N_49121,N_48875);
and UO_3070 (O_3070,N_49859,N_48895);
nand UO_3071 (O_3071,N_48026,N_49589);
and UO_3072 (O_3072,N_48673,N_48118);
nand UO_3073 (O_3073,N_48881,N_49961);
and UO_3074 (O_3074,N_49540,N_48012);
and UO_3075 (O_3075,N_48418,N_48894);
and UO_3076 (O_3076,N_49462,N_49280);
nor UO_3077 (O_3077,N_49706,N_48604);
nor UO_3078 (O_3078,N_48745,N_49762);
and UO_3079 (O_3079,N_49797,N_48999);
nor UO_3080 (O_3080,N_49736,N_49761);
nand UO_3081 (O_3081,N_49678,N_49348);
and UO_3082 (O_3082,N_49213,N_49134);
nand UO_3083 (O_3083,N_48913,N_49759);
or UO_3084 (O_3084,N_48012,N_48577);
nand UO_3085 (O_3085,N_49822,N_48014);
or UO_3086 (O_3086,N_49984,N_48386);
and UO_3087 (O_3087,N_48478,N_49115);
nor UO_3088 (O_3088,N_49888,N_48567);
and UO_3089 (O_3089,N_49047,N_48154);
nor UO_3090 (O_3090,N_49267,N_48677);
and UO_3091 (O_3091,N_48752,N_48121);
and UO_3092 (O_3092,N_49202,N_49851);
nor UO_3093 (O_3093,N_49335,N_49120);
nor UO_3094 (O_3094,N_48400,N_49272);
nand UO_3095 (O_3095,N_49864,N_48942);
or UO_3096 (O_3096,N_48207,N_48971);
or UO_3097 (O_3097,N_49708,N_48412);
or UO_3098 (O_3098,N_48451,N_49903);
and UO_3099 (O_3099,N_49285,N_49435);
or UO_3100 (O_3100,N_48641,N_48098);
nor UO_3101 (O_3101,N_48674,N_49253);
nand UO_3102 (O_3102,N_48946,N_48113);
nor UO_3103 (O_3103,N_49533,N_48590);
nand UO_3104 (O_3104,N_48371,N_48121);
xnor UO_3105 (O_3105,N_48790,N_49861);
or UO_3106 (O_3106,N_49175,N_49307);
and UO_3107 (O_3107,N_49816,N_48020);
nor UO_3108 (O_3108,N_49047,N_49481);
nor UO_3109 (O_3109,N_48886,N_48959);
nand UO_3110 (O_3110,N_49058,N_49694);
and UO_3111 (O_3111,N_48490,N_48344);
nor UO_3112 (O_3112,N_48079,N_49805);
nor UO_3113 (O_3113,N_49924,N_48012);
and UO_3114 (O_3114,N_48578,N_48187);
or UO_3115 (O_3115,N_49452,N_49748);
nand UO_3116 (O_3116,N_49417,N_49274);
nand UO_3117 (O_3117,N_48329,N_48129);
or UO_3118 (O_3118,N_48619,N_48068);
and UO_3119 (O_3119,N_49179,N_49638);
nor UO_3120 (O_3120,N_48146,N_49033);
and UO_3121 (O_3121,N_49711,N_49042);
nand UO_3122 (O_3122,N_48214,N_49007);
xor UO_3123 (O_3123,N_48714,N_48373);
and UO_3124 (O_3124,N_48554,N_49411);
or UO_3125 (O_3125,N_48824,N_49970);
and UO_3126 (O_3126,N_48806,N_48730);
or UO_3127 (O_3127,N_49171,N_48656);
nand UO_3128 (O_3128,N_48485,N_49035);
nor UO_3129 (O_3129,N_48592,N_49815);
nor UO_3130 (O_3130,N_49223,N_49435);
xor UO_3131 (O_3131,N_49836,N_49474);
or UO_3132 (O_3132,N_48831,N_49825);
or UO_3133 (O_3133,N_48018,N_48769);
or UO_3134 (O_3134,N_49687,N_49328);
and UO_3135 (O_3135,N_49473,N_49371);
or UO_3136 (O_3136,N_48793,N_49366);
or UO_3137 (O_3137,N_49863,N_49691);
and UO_3138 (O_3138,N_49337,N_48768);
nand UO_3139 (O_3139,N_48222,N_49466);
nor UO_3140 (O_3140,N_49527,N_49107);
and UO_3141 (O_3141,N_48028,N_49774);
nor UO_3142 (O_3142,N_49256,N_49569);
and UO_3143 (O_3143,N_49175,N_48603);
xor UO_3144 (O_3144,N_48290,N_49121);
nor UO_3145 (O_3145,N_48812,N_48492);
nor UO_3146 (O_3146,N_49858,N_49035);
nor UO_3147 (O_3147,N_48776,N_48024);
or UO_3148 (O_3148,N_49770,N_48967);
nand UO_3149 (O_3149,N_49292,N_48990);
nand UO_3150 (O_3150,N_49224,N_49699);
nand UO_3151 (O_3151,N_48815,N_49528);
or UO_3152 (O_3152,N_48807,N_48856);
or UO_3153 (O_3153,N_49329,N_48192);
nor UO_3154 (O_3154,N_48762,N_48148);
nor UO_3155 (O_3155,N_48274,N_48858);
or UO_3156 (O_3156,N_48503,N_49469);
nor UO_3157 (O_3157,N_48144,N_49263);
and UO_3158 (O_3158,N_49027,N_49262);
or UO_3159 (O_3159,N_49147,N_48623);
nor UO_3160 (O_3160,N_48982,N_49750);
or UO_3161 (O_3161,N_48530,N_48122);
nor UO_3162 (O_3162,N_48344,N_49297);
nor UO_3163 (O_3163,N_48962,N_48911);
and UO_3164 (O_3164,N_49843,N_49696);
or UO_3165 (O_3165,N_48996,N_49874);
or UO_3166 (O_3166,N_49743,N_49838);
nand UO_3167 (O_3167,N_48290,N_48681);
and UO_3168 (O_3168,N_48688,N_49256);
or UO_3169 (O_3169,N_49523,N_48586);
nand UO_3170 (O_3170,N_49340,N_48856);
or UO_3171 (O_3171,N_49600,N_49909);
and UO_3172 (O_3172,N_49219,N_49439);
and UO_3173 (O_3173,N_48489,N_49651);
and UO_3174 (O_3174,N_48181,N_49233);
nor UO_3175 (O_3175,N_49831,N_48990);
and UO_3176 (O_3176,N_48421,N_49163);
or UO_3177 (O_3177,N_48306,N_48498);
or UO_3178 (O_3178,N_49755,N_49010);
nor UO_3179 (O_3179,N_48845,N_48532);
nor UO_3180 (O_3180,N_48947,N_48838);
and UO_3181 (O_3181,N_49695,N_48554);
xnor UO_3182 (O_3182,N_49461,N_48074);
nor UO_3183 (O_3183,N_48982,N_49083);
and UO_3184 (O_3184,N_49190,N_48695);
and UO_3185 (O_3185,N_49486,N_49942);
nor UO_3186 (O_3186,N_48506,N_48635);
and UO_3187 (O_3187,N_48190,N_48616);
or UO_3188 (O_3188,N_49552,N_48889);
or UO_3189 (O_3189,N_49270,N_48168);
nand UO_3190 (O_3190,N_49730,N_48276);
nand UO_3191 (O_3191,N_48096,N_48589);
and UO_3192 (O_3192,N_48909,N_48158);
nor UO_3193 (O_3193,N_48672,N_48563);
or UO_3194 (O_3194,N_48263,N_48885);
nor UO_3195 (O_3195,N_48771,N_49706);
nor UO_3196 (O_3196,N_48160,N_48108);
or UO_3197 (O_3197,N_48154,N_49073);
and UO_3198 (O_3198,N_48727,N_48212);
nor UO_3199 (O_3199,N_48342,N_49948);
nand UO_3200 (O_3200,N_48405,N_48224);
and UO_3201 (O_3201,N_48484,N_49674);
nor UO_3202 (O_3202,N_49310,N_49781);
nand UO_3203 (O_3203,N_48512,N_49213);
nand UO_3204 (O_3204,N_49550,N_48496);
nor UO_3205 (O_3205,N_48661,N_48418);
nand UO_3206 (O_3206,N_48674,N_49838);
or UO_3207 (O_3207,N_49140,N_48131);
nor UO_3208 (O_3208,N_49221,N_48565);
xnor UO_3209 (O_3209,N_48987,N_48448);
nor UO_3210 (O_3210,N_49298,N_49511);
nand UO_3211 (O_3211,N_49366,N_48969);
nand UO_3212 (O_3212,N_49471,N_48037);
nor UO_3213 (O_3213,N_49001,N_49881);
and UO_3214 (O_3214,N_48763,N_49512);
and UO_3215 (O_3215,N_48877,N_48858);
nor UO_3216 (O_3216,N_48953,N_49330);
and UO_3217 (O_3217,N_49317,N_48044);
nor UO_3218 (O_3218,N_49535,N_48953);
or UO_3219 (O_3219,N_48357,N_48489);
or UO_3220 (O_3220,N_48746,N_48969);
nor UO_3221 (O_3221,N_49507,N_48577);
or UO_3222 (O_3222,N_48266,N_48124);
or UO_3223 (O_3223,N_49614,N_49098);
or UO_3224 (O_3224,N_49014,N_48114);
nor UO_3225 (O_3225,N_49137,N_48270);
or UO_3226 (O_3226,N_48133,N_48037);
or UO_3227 (O_3227,N_48357,N_48355);
and UO_3228 (O_3228,N_49071,N_48444);
nand UO_3229 (O_3229,N_49542,N_49761);
or UO_3230 (O_3230,N_49944,N_49781);
and UO_3231 (O_3231,N_48362,N_49142);
and UO_3232 (O_3232,N_48861,N_49973);
or UO_3233 (O_3233,N_49414,N_49432);
and UO_3234 (O_3234,N_49756,N_48327);
nand UO_3235 (O_3235,N_49833,N_49913);
and UO_3236 (O_3236,N_48210,N_48947);
or UO_3237 (O_3237,N_48142,N_48426);
nand UO_3238 (O_3238,N_48565,N_49529);
and UO_3239 (O_3239,N_49347,N_48383);
and UO_3240 (O_3240,N_49939,N_49843);
and UO_3241 (O_3241,N_48401,N_49670);
nor UO_3242 (O_3242,N_48650,N_49371);
nor UO_3243 (O_3243,N_48882,N_48883);
nor UO_3244 (O_3244,N_49515,N_49252);
and UO_3245 (O_3245,N_48545,N_48770);
nand UO_3246 (O_3246,N_49891,N_48709);
nand UO_3247 (O_3247,N_48038,N_49849);
and UO_3248 (O_3248,N_48912,N_49988);
nor UO_3249 (O_3249,N_48747,N_48503);
or UO_3250 (O_3250,N_49270,N_48518);
and UO_3251 (O_3251,N_48358,N_48050);
nand UO_3252 (O_3252,N_48036,N_48602);
nor UO_3253 (O_3253,N_49572,N_48901);
or UO_3254 (O_3254,N_49644,N_49850);
nand UO_3255 (O_3255,N_49256,N_49979);
nor UO_3256 (O_3256,N_49197,N_48217);
and UO_3257 (O_3257,N_48368,N_49405);
nor UO_3258 (O_3258,N_48273,N_49898);
nand UO_3259 (O_3259,N_48965,N_48640);
xnor UO_3260 (O_3260,N_49010,N_49006);
nor UO_3261 (O_3261,N_48817,N_49663);
and UO_3262 (O_3262,N_48102,N_49425);
nor UO_3263 (O_3263,N_48434,N_49087);
and UO_3264 (O_3264,N_48072,N_49853);
nand UO_3265 (O_3265,N_48144,N_49621);
or UO_3266 (O_3266,N_48310,N_49542);
nand UO_3267 (O_3267,N_48100,N_49235);
xnor UO_3268 (O_3268,N_48400,N_48451);
and UO_3269 (O_3269,N_48834,N_49201);
or UO_3270 (O_3270,N_48024,N_48299);
nand UO_3271 (O_3271,N_49843,N_49094);
nor UO_3272 (O_3272,N_49144,N_49482);
nand UO_3273 (O_3273,N_49710,N_48621);
nand UO_3274 (O_3274,N_49810,N_49803);
or UO_3275 (O_3275,N_48179,N_48231);
or UO_3276 (O_3276,N_49629,N_48137);
nor UO_3277 (O_3277,N_48319,N_49916);
nor UO_3278 (O_3278,N_48471,N_48280);
nand UO_3279 (O_3279,N_48972,N_48079);
nor UO_3280 (O_3280,N_48610,N_48718);
nand UO_3281 (O_3281,N_48627,N_48391);
nand UO_3282 (O_3282,N_48731,N_48906);
and UO_3283 (O_3283,N_48550,N_49843);
nand UO_3284 (O_3284,N_49927,N_49415);
or UO_3285 (O_3285,N_49154,N_48421);
nand UO_3286 (O_3286,N_48798,N_49077);
or UO_3287 (O_3287,N_48387,N_49408);
nand UO_3288 (O_3288,N_48992,N_49588);
or UO_3289 (O_3289,N_49105,N_48917);
or UO_3290 (O_3290,N_48000,N_48773);
nor UO_3291 (O_3291,N_48541,N_49192);
xor UO_3292 (O_3292,N_49285,N_48814);
nor UO_3293 (O_3293,N_49531,N_49019);
nor UO_3294 (O_3294,N_48022,N_48698);
nand UO_3295 (O_3295,N_49903,N_48047);
nand UO_3296 (O_3296,N_48383,N_49372);
or UO_3297 (O_3297,N_49930,N_48679);
nor UO_3298 (O_3298,N_49350,N_48484);
nor UO_3299 (O_3299,N_49152,N_48117);
nand UO_3300 (O_3300,N_48184,N_49525);
nor UO_3301 (O_3301,N_48629,N_49529);
or UO_3302 (O_3302,N_49144,N_48574);
nand UO_3303 (O_3303,N_49679,N_48786);
or UO_3304 (O_3304,N_48235,N_48084);
and UO_3305 (O_3305,N_49022,N_49473);
nor UO_3306 (O_3306,N_49834,N_48729);
or UO_3307 (O_3307,N_48493,N_49433);
nor UO_3308 (O_3308,N_49752,N_48896);
or UO_3309 (O_3309,N_49995,N_48032);
nor UO_3310 (O_3310,N_48383,N_48188);
nand UO_3311 (O_3311,N_49043,N_49035);
and UO_3312 (O_3312,N_49379,N_49027);
nand UO_3313 (O_3313,N_48423,N_48742);
and UO_3314 (O_3314,N_49028,N_48136);
nand UO_3315 (O_3315,N_49646,N_48249);
or UO_3316 (O_3316,N_48978,N_48911);
nor UO_3317 (O_3317,N_49710,N_48761);
and UO_3318 (O_3318,N_48133,N_48114);
or UO_3319 (O_3319,N_49232,N_48134);
xor UO_3320 (O_3320,N_48067,N_49576);
and UO_3321 (O_3321,N_48918,N_49209);
nor UO_3322 (O_3322,N_48763,N_49400);
and UO_3323 (O_3323,N_48379,N_48959);
or UO_3324 (O_3324,N_48929,N_49986);
or UO_3325 (O_3325,N_49715,N_49706);
nor UO_3326 (O_3326,N_49952,N_48518);
nand UO_3327 (O_3327,N_48127,N_48264);
xor UO_3328 (O_3328,N_49431,N_48181);
and UO_3329 (O_3329,N_48705,N_48560);
and UO_3330 (O_3330,N_49365,N_48007);
or UO_3331 (O_3331,N_48878,N_49857);
nor UO_3332 (O_3332,N_49781,N_49235);
and UO_3333 (O_3333,N_49943,N_48462);
and UO_3334 (O_3334,N_48411,N_49666);
nand UO_3335 (O_3335,N_49091,N_49843);
nand UO_3336 (O_3336,N_49746,N_49573);
nand UO_3337 (O_3337,N_48307,N_48076);
xor UO_3338 (O_3338,N_48764,N_48964);
or UO_3339 (O_3339,N_48806,N_48141);
or UO_3340 (O_3340,N_48093,N_48938);
nand UO_3341 (O_3341,N_49198,N_49139);
or UO_3342 (O_3342,N_48676,N_49339);
or UO_3343 (O_3343,N_49236,N_48009);
nor UO_3344 (O_3344,N_48107,N_48582);
or UO_3345 (O_3345,N_49381,N_48997);
or UO_3346 (O_3346,N_48943,N_48164);
nor UO_3347 (O_3347,N_48522,N_49730);
or UO_3348 (O_3348,N_49398,N_48184);
nor UO_3349 (O_3349,N_48116,N_49391);
nor UO_3350 (O_3350,N_49514,N_48979);
nor UO_3351 (O_3351,N_49702,N_49297);
and UO_3352 (O_3352,N_49868,N_49796);
and UO_3353 (O_3353,N_48620,N_49139);
nor UO_3354 (O_3354,N_49073,N_49895);
nor UO_3355 (O_3355,N_48889,N_48945);
or UO_3356 (O_3356,N_49457,N_49015);
and UO_3357 (O_3357,N_49183,N_48902);
nor UO_3358 (O_3358,N_49801,N_48272);
and UO_3359 (O_3359,N_49487,N_48452);
or UO_3360 (O_3360,N_48819,N_49809);
or UO_3361 (O_3361,N_48867,N_48037);
or UO_3362 (O_3362,N_48542,N_48142);
and UO_3363 (O_3363,N_48752,N_48019);
and UO_3364 (O_3364,N_48151,N_48749);
nor UO_3365 (O_3365,N_48384,N_49883);
and UO_3366 (O_3366,N_48931,N_49514);
nand UO_3367 (O_3367,N_49996,N_49268);
or UO_3368 (O_3368,N_48859,N_49190);
and UO_3369 (O_3369,N_48395,N_48819);
nand UO_3370 (O_3370,N_48065,N_49041);
or UO_3371 (O_3371,N_48288,N_49048);
or UO_3372 (O_3372,N_49974,N_49863);
nand UO_3373 (O_3373,N_48457,N_48587);
or UO_3374 (O_3374,N_48269,N_48495);
and UO_3375 (O_3375,N_49247,N_48488);
and UO_3376 (O_3376,N_49214,N_49956);
nor UO_3377 (O_3377,N_48382,N_49410);
nand UO_3378 (O_3378,N_48136,N_49235);
nor UO_3379 (O_3379,N_48613,N_48275);
and UO_3380 (O_3380,N_49923,N_48662);
or UO_3381 (O_3381,N_49834,N_49252);
nand UO_3382 (O_3382,N_49977,N_48501);
and UO_3383 (O_3383,N_49507,N_48366);
or UO_3384 (O_3384,N_48051,N_48224);
nor UO_3385 (O_3385,N_48591,N_49306);
nor UO_3386 (O_3386,N_49991,N_49965);
nand UO_3387 (O_3387,N_49170,N_48749);
nand UO_3388 (O_3388,N_49656,N_48214);
nor UO_3389 (O_3389,N_48821,N_48538);
or UO_3390 (O_3390,N_48367,N_49225);
and UO_3391 (O_3391,N_48758,N_49146);
nand UO_3392 (O_3392,N_49726,N_49247);
nand UO_3393 (O_3393,N_48251,N_49504);
nor UO_3394 (O_3394,N_49236,N_49112);
nor UO_3395 (O_3395,N_49750,N_49229);
nor UO_3396 (O_3396,N_48534,N_49778);
or UO_3397 (O_3397,N_48121,N_48764);
nand UO_3398 (O_3398,N_48157,N_48209);
nor UO_3399 (O_3399,N_48706,N_48127);
and UO_3400 (O_3400,N_49594,N_49675);
or UO_3401 (O_3401,N_49673,N_49491);
nand UO_3402 (O_3402,N_49492,N_48739);
and UO_3403 (O_3403,N_49203,N_48413);
nand UO_3404 (O_3404,N_49795,N_49103);
nand UO_3405 (O_3405,N_49302,N_49880);
nand UO_3406 (O_3406,N_49648,N_49523);
and UO_3407 (O_3407,N_49544,N_48896);
and UO_3408 (O_3408,N_49564,N_49545);
or UO_3409 (O_3409,N_49506,N_48468);
xnor UO_3410 (O_3410,N_48907,N_48669);
nor UO_3411 (O_3411,N_49361,N_49626);
nor UO_3412 (O_3412,N_49201,N_49244);
nand UO_3413 (O_3413,N_48981,N_48497);
and UO_3414 (O_3414,N_48198,N_49555);
or UO_3415 (O_3415,N_49940,N_49460);
and UO_3416 (O_3416,N_48845,N_48763);
nor UO_3417 (O_3417,N_48025,N_49446);
or UO_3418 (O_3418,N_48832,N_49428);
nor UO_3419 (O_3419,N_49179,N_49426);
nand UO_3420 (O_3420,N_49741,N_49716);
nand UO_3421 (O_3421,N_48610,N_48565);
and UO_3422 (O_3422,N_49369,N_48228);
or UO_3423 (O_3423,N_49847,N_49739);
and UO_3424 (O_3424,N_48160,N_48154);
nand UO_3425 (O_3425,N_48825,N_49475);
nor UO_3426 (O_3426,N_49774,N_48648);
nand UO_3427 (O_3427,N_49628,N_48930);
or UO_3428 (O_3428,N_48909,N_48633);
or UO_3429 (O_3429,N_48728,N_48921);
and UO_3430 (O_3430,N_48832,N_48127);
nor UO_3431 (O_3431,N_48120,N_48543);
nor UO_3432 (O_3432,N_48646,N_49497);
or UO_3433 (O_3433,N_49869,N_49528);
and UO_3434 (O_3434,N_48877,N_48843);
or UO_3435 (O_3435,N_49691,N_49846);
nand UO_3436 (O_3436,N_48447,N_48517);
or UO_3437 (O_3437,N_49557,N_48266);
nand UO_3438 (O_3438,N_49471,N_49122);
and UO_3439 (O_3439,N_49818,N_49406);
and UO_3440 (O_3440,N_49678,N_49494);
nand UO_3441 (O_3441,N_48688,N_48774);
or UO_3442 (O_3442,N_49548,N_48910);
nand UO_3443 (O_3443,N_49404,N_48810);
nor UO_3444 (O_3444,N_48488,N_48835);
or UO_3445 (O_3445,N_48997,N_48666);
nor UO_3446 (O_3446,N_49886,N_49578);
or UO_3447 (O_3447,N_49792,N_49532);
xnor UO_3448 (O_3448,N_49245,N_49037);
nand UO_3449 (O_3449,N_49952,N_48681);
and UO_3450 (O_3450,N_48610,N_48265);
and UO_3451 (O_3451,N_48728,N_48548);
nand UO_3452 (O_3452,N_49266,N_49955);
nor UO_3453 (O_3453,N_49204,N_49397);
and UO_3454 (O_3454,N_49616,N_49934);
or UO_3455 (O_3455,N_48175,N_49338);
and UO_3456 (O_3456,N_49945,N_48279);
or UO_3457 (O_3457,N_48876,N_49412);
nand UO_3458 (O_3458,N_48212,N_48426);
or UO_3459 (O_3459,N_49088,N_48532);
nand UO_3460 (O_3460,N_49140,N_48876);
and UO_3461 (O_3461,N_49154,N_49628);
nor UO_3462 (O_3462,N_48262,N_48271);
nor UO_3463 (O_3463,N_49456,N_48525);
nand UO_3464 (O_3464,N_48143,N_49016);
and UO_3465 (O_3465,N_48589,N_48366);
and UO_3466 (O_3466,N_48991,N_48952);
and UO_3467 (O_3467,N_48613,N_48068);
or UO_3468 (O_3468,N_49145,N_48797);
nand UO_3469 (O_3469,N_48369,N_48663);
nand UO_3470 (O_3470,N_48338,N_48835);
or UO_3471 (O_3471,N_49413,N_49459);
nor UO_3472 (O_3472,N_49084,N_49596);
nand UO_3473 (O_3473,N_49054,N_48877);
nor UO_3474 (O_3474,N_48906,N_48249);
and UO_3475 (O_3475,N_48664,N_48232);
nand UO_3476 (O_3476,N_49428,N_48651);
and UO_3477 (O_3477,N_48782,N_48299);
and UO_3478 (O_3478,N_48269,N_48493);
nand UO_3479 (O_3479,N_49557,N_49033);
or UO_3480 (O_3480,N_48374,N_49238);
nor UO_3481 (O_3481,N_48329,N_49430);
nand UO_3482 (O_3482,N_49976,N_48412);
and UO_3483 (O_3483,N_48030,N_48225);
nand UO_3484 (O_3484,N_48200,N_48521);
nor UO_3485 (O_3485,N_49823,N_49306);
nand UO_3486 (O_3486,N_49822,N_48498);
and UO_3487 (O_3487,N_49417,N_49383);
or UO_3488 (O_3488,N_49675,N_48964);
and UO_3489 (O_3489,N_48948,N_48960);
nand UO_3490 (O_3490,N_49877,N_48516);
nor UO_3491 (O_3491,N_48137,N_48039);
and UO_3492 (O_3492,N_48842,N_48928);
nor UO_3493 (O_3493,N_49253,N_48859);
nor UO_3494 (O_3494,N_49445,N_48640);
nor UO_3495 (O_3495,N_48631,N_49223);
or UO_3496 (O_3496,N_48920,N_49052);
nor UO_3497 (O_3497,N_49056,N_48977);
or UO_3498 (O_3498,N_49720,N_48948);
and UO_3499 (O_3499,N_48147,N_48766);
nor UO_3500 (O_3500,N_48977,N_49479);
or UO_3501 (O_3501,N_48185,N_48681);
nor UO_3502 (O_3502,N_49508,N_48525);
nor UO_3503 (O_3503,N_49717,N_48394);
or UO_3504 (O_3504,N_48738,N_48842);
nor UO_3505 (O_3505,N_48641,N_49891);
xnor UO_3506 (O_3506,N_48276,N_48650);
nand UO_3507 (O_3507,N_48670,N_49069);
or UO_3508 (O_3508,N_49276,N_48146);
and UO_3509 (O_3509,N_49789,N_48885);
nand UO_3510 (O_3510,N_49258,N_48082);
and UO_3511 (O_3511,N_49171,N_48296);
nand UO_3512 (O_3512,N_49765,N_49304);
and UO_3513 (O_3513,N_49868,N_48442);
or UO_3514 (O_3514,N_48522,N_48649);
nor UO_3515 (O_3515,N_49233,N_48946);
or UO_3516 (O_3516,N_49619,N_49351);
and UO_3517 (O_3517,N_49971,N_49210);
nor UO_3518 (O_3518,N_48943,N_48484);
xor UO_3519 (O_3519,N_49069,N_48510);
nand UO_3520 (O_3520,N_49248,N_49416);
nor UO_3521 (O_3521,N_49344,N_49742);
and UO_3522 (O_3522,N_49171,N_48080);
and UO_3523 (O_3523,N_49207,N_48761);
nand UO_3524 (O_3524,N_48642,N_48745);
nor UO_3525 (O_3525,N_49256,N_49596);
and UO_3526 (O_3526,N_49645,N_48349);
nor UO_3527 (O_3527,N_49871,N_49905);
and UO_3528 (O_3528,N_48074,N_49674);
nor UO_3529 (O_3529,N_49486,N_49374);
and UO_3530 (O_3530,N_48666,N_48546);
nand UO_3531 (O_3531,N_48573,N_49822);
nand UO_3532 (O_3532,N_49644,N_49243);
xor UO_3533 (O_3533,N_48264,N_48915);
or UO_3534 (O_3534,N_48461,N_49327);
nor UO_3535 (O_3535,N_48039,N_48387);
nand UO_3536 (O_3536,N_48523,N_48997);
nor UO_3537 (O_3537,N_49962,N_48986);
or UO_3538 (O_3538,N_49489,N_48745);
or UO_3539 (O_3539,N_49551,N_49510);
nor UO_3540 (O_3540,N_49445,N_49457);
nand UO_3541 (O_3541,N_48214,N_49957);
nor UO_3542 (O_3542,N_49169,N_49127);
or UO_3543 (O_3543,N_49692,N_48408);
nand UO_3544 (O_3544,N_49879,N_48476);
nor UO_3545 (O_3545,N_48231,N_48726);
nand UO_3546 (O_3546,N_49387,N_49480);
nor UO_3547 (O_3547,N_48026,N_49359);
or UO_3548 (O_3548,N_49847,N_49897);
and UO_3549 (O_3549,N_49608,N_49638);
and UO_3550 (O_3550,N_49603,N_48923);
nand UO_3551 (O_3551,N_48070,N_49496);
nand UO_3552 (O_3552,N_49965,N_48606);
nand UO_3553 (O_3553,N_49202,N_49470);
and UO_3554 (O_3554,N_49886,N_48395);
nor UO_3555 (O_3555,N_48524,N_48169);
and UO_3556 (O_3556,N_48692,N_49849);
nand UO_3557 (O_3557,N_49599,N_48916);
xnor UO_3558 (O_3558,N_48233,N_49566);
nand UO_3559 (O_3559,N_48037,N_48769);
nand UO_3560 (O_3560,N_48159,N_49329);
or UO_3561 (O_3561,N_48479,N_48682);
and UO_3562 (O_3562,N_49317,N_49509);
nor UO_3563 (O_3563,N_49018,N_49649);
or UO_3564 (O_3564,N_48009,N_49070);
nor UO_3565 (O_3565,N_48467,N_48524);
or UO_3566 (O_3566,N_48777,N_48229);
and UO_3567 (O_3567,N_48102,N_48209);
or UO_3568 (O_3568,N_49193,N_49435);
or UO_3569 (O_3569,N_49423,N_49097);
or UO_3570 (O_3570,N_48797,N_48474);
and UO_3571 (O_3571,N_49875,N_48162);
or UO_3572 (O_3572,N_49187,N_49975);
nor UO_3573 (O_3573,N_48211,N_48243);
nor UO_3574 (O_3574,N_49818,N_49036);
nand UO_3575 (O_3575,N_48045,N_49907);
and UO_3576 (O_3576,N_49293,N_49110);
and UO_3577 (O_3577,N_48461,N_49576);
nor UO_3578 (O_3578,N_49690,N_49807);
nor UO_3579 (O_3579,N_49390,N_48039);
nor UO_3580 (O_3580,N_48269,N_49639);
nand UO_3581 (O_3581,N_48669,N_48668);
nor UO_3582 (O_3582,N_48024,N_48038);
nor UO_3583 (O_3583,N_49939,N_49240);
and UO_3584 (O_3584,N_48981,N_48277);
nor UO_3585 (O_3585,N_48929,N_49762);
nor UO_3586 (O_3586,N_48477,N_48061);
nor UO_3587 (O_3587,N_48811,N_49561);
or UO_3588 (O_3588,N_49869,N_48061);
nand UO_3589 (O_3589,N_48752,N_48245);
nand UO_3590 (O_3590,N_49331,N_48859);
or UO_3591 (O_3591,N_49034,N_49785);
or UO_3592 (O_3592,N_48787,N_49736);
and UO_3593 (O_3593,N_49484,N_48874);
and UO_3594 (O_3594,N_48313,N_49484);
nor UO_3595 (O_3595,N_48190,N_48499);
and UO_3596 (O_3596,N_49213,N_48856);
or UO_3597 (O_3597,N_49946,N_48077);
or UO_3598 (O_3598,N_48045,N_48438);
nor UO_3599 (O_3599,N_48322,N_48093);
nor UO_3600 (O_3600,N_49200,N_48045);
nand UO_3601 (O_3601,N_49528,N_48929);
nor UO_3602 (O_3602,N_48828,N_48046);
or UO_3603 (O_3603,N_48682,N_49408);
nor UO_3604 (O_3604,N_48000,N_48465);
or UO_3605 (O_3605,N_49914,N_48303);
and UO_3606 (O_3606,N_49212,N_49709);
nor UO_3607 (O_3607,N_48036,N_48863);
nor UO_3608 (O_3608,N_48674,N_49998);
or UO_3609 (O_3609,N_48553,N_49966);
nor UO_3610 (O_3610,N_48108,N_49647);
nor UO_3611 (O_3611,N_48472,N_48759);
or UO_3612 (O_3612,N_49004,N_48599);
and UO_3613 (O_3613,N_49553,N_48250);
xor UO_3614 (O_3614,N_48170,N_49564);
or UO_3615 (O_3615,N_49168,N_49347);
nand UO_3616 (O_3616,N_49762,N_49314);
or UO_3617 (O_3617,N_49051,N_48816);
nor UO_3618 (O_3618,N_48020,N_48045);
and UO_3619 (O_3619,N_49594,N_48388);
nand UO_3620 (O_3620,N_49974,N_49335);
and UO_3621 (O_3621,N_48418,N_49375);
or UO_3622 (O_3622,N_48719,N_48468);
or UO_3623 (O_3623,N_48550,N_49234);
nand UO_3624 (O_3624,N_49505,N_49579);
and UO_3625 (O_3625,N_49731,N_48551);
and UO_3626 (O_3626,N_49878,N_48959);
nor UO_3627 (O_3627,N_48118,N_49528);
nand UO_3628 (O_3628,N_49566,N_49338);
or UO_3629 (O_3629,N_49346,N_48736);
nor UO_3630 (O_3630,N_49692,N_49386);
nand UO_3631 (O_3631,N_49771,N_49322);
nand UO_3632 (O_3632,N_48179,N_49294);
or UO_3633 (O_3633,N_48491,N_48020);
nand UO_3634 (O_3634,N_49689,N_49874);
nand UO_3635 (O_3635,N_48126,N_49884);
or UO_3636 (O_3636,N_48190,N_48517);
or UO_3637 (O_3637,N_48660,N_49471);
and UO_3638 (O_3638,N_48953,N_49229);
or UO_3639 (O_3639,N_49419,N_48944);
nor UO_3640 (O_3640,N_49857,N_48842);
and UO_3641 (O_3641,N_49272,N_48939);
or UO_3642 (O_3642,N_49986,N_48041);
and UO_3643 (O_3643,N_48370,N_48152);
nor UO_3644 (O_3644,N_48837,N_49726);
nand UO_3645 (O_3645,N_48190,N_48977);
and UO_3646 (O_3646,N_49272,N_48971);
nand UO_3647 (O_3647,N_49491,N_49227);
nand UO_3648 (O_3648,N_49416,N_49110);
nand UO_3649 (O_3649,N_48329,N_48428);
or UO_3650 (O_3650,N_48975,N_49750);
xor UO_3651 (O_3651,N_49814,N_49886);
nor UO_3652 (O_3652,N_48206,N_49651);
or UO_3653 (O_3653,N_49296,N_49691);
nand UO_3654 (O_3654,N_48412,N_48771);
nor UO_3655 (O_3655,N_48192,N_48232);
nand UO_3656 (O_3656,N_48399,N_48772);
nor UO_3657 (O_3657,N_49474,N_49945);
and UO_3658 (O_3658,N_49827,N_48929);
or UO_3659 (O_3659,N_49443,N_49638);
or UO_3660 (O_3660,N_49531,N_48880);
nor UO_3661 (O_3661,N_49479,N_49496);
or UO_3662 (O_3662,N_48147,N_49798);
nor UO_3663 (O_3663,N_48276,N_48127);
nor UO_3664 (O_3664,N_48241,N_48221);
nand UO_3665 (O_3665,N_48346,N_48954);
and UO_3666 (O_3666,N_49099,N_48749);
or UO_3667 (O_3667,N_49874,N_49228);
xnor UO_3668 (O_3668,N_48440,N_48130);
or UO_3669 (O_3669,N_48690,N_49466);
and UO_3670 (O_3670,N_48366,N_48062);
and UO_3671 (O_3671,N_49429,N_48833);
nor UO_3672 (O_3672,N_49251,N_49473);
nand UO_3673 (O_3673,N_49272,N_48898);
nor UO_3674 (O_3674,N_49827,N_49984);
nor UO_3675 (O_3675,N_49573,N_49763);
and UO_3676 (O_3676,N_48906,N_49371);
or UO_3677 (O_3677,N_48570,N_49100);
or UO_3678 (O_3678,N_49682,N_48414);
nand UO_3679 (O_3679,N_48257,N_49983);
and UO_3680 (O_3680,N_49207,N_49279);
nor UO_3681 (O_3681,N_48337,N_49110);
xnor UO_3682 (O_3682,N_48776,N_49681);
nand UO_3683 (O_3683,N_49633,N_49866);
nor UO_3684 (O_3684,N_49206,N_49687);
and UO_3685 (O_3685,N_49185,N_49317);
nand UO_3686 (O_3686,N_49124,N_49885);
xor UO_3687 (O_3687,N_49599,N_49879);
and UO_3688 (O_3688,N_49152,N_49077);
or UO_3689 (O_3689,N_48464,N_48608);
nand UO_3690 (O_3690,N_48646,N_48225);
and UO_3691 (O_3691,N_49320,N_49125);
and UO_3692 (O_3692,N_48395,N_48969);
nor UO_3693 (O_3693,N_49648,N_49644);
and UO_3694 (O_3694,N_49729,N_49998);
and UO_3695 (O_3695,N_49790,N_48543);
xnor UO_3696 (O_3696,N_49884,N_48620);
and UO_3697 (O_3697,N_48240,N_48292);
nor UO_3698 (O_3698,N_48782,N_49772);
nor UO_3699 (O_3699,N_48621,N_48103);
nor UO_3700 (O_3700,N_49803,N_48461);
or UO_3701 (O_3701,N_49211,N_49247);
nor UO_3702 (O_3702,N_48697,N_49483);
nor UO_3703 (O_3703,N_48314,N_49401);
and UO_3704 (O_3704,N_49729,N_49642);
or UO_3705 (O_3705,N_49190,N_48372);
nand UO_3706 (O_3706,N_49626,N_48938);
or UO_3707 (O_3707,N_48555,N_49404);
xor UO_3708 (O_3708,N_48935,N_49921);
or UO_3709 (O_3709,N_49276,N_49560);
or UO_3710 (O_3710,N_48227,N_49523);
or UO_3711 (O_3711,N_49121,N_49225);
and UO_3712 (O_3712,N_49496,N_48417);
nand UO_3713 (O_3713,N_49919,N_48605);
nand UO_3714 (O_3714,N_48477,N_49451);
or UO_3715 (O_3715,N_48594,N_49894);
nor UO_3716 (O_3716,N_49670,N_48313);
or UO_3717 (O_3717,N_49328,N_48814);
nor UO_3718 (O_3718,N_48143,N_48067);
and UO_3719 (O_3719,N_49921,N_49036);
and UO_3720 (O_3720,N_49110,N_48603);
nand UO_3721 (O_3721,N_48706,N_48829);
nor UO_3722 (O_3722,N_48707,N_48213);
or UO_3723 (O_3723,N_48531,N_48103);
and UO_3724 (O_3724,N_48805,N_48682);
or UO_3725 (O_3725,N_49318,N_49393);
xor UO_3726 (O_3726,N_49902,N_48501);
nand UO_3727 (O_3727,N_49303,N_48177);
nand UO_3728 (O_3728,N_48292,N_49077);
and UO_3729 (O_3729,N_49411,N_49014);
or UO_3730 (O_3730,N_49069,N_48270);
nor UO_3731 (O_3731,N_48146,N_49864);
nand UO_3732 (O_3732,N_49483,N_48104);
nor UO_3733 (O_3733,N_48213,N_49711);
nand UO_3734 (O_3734,N_49355,N_49713);
nor UO_3735 (O_3735,N_48080,N_49284);
and UO_3736 (O_3736,N_49376,N_49294);
and UO_3737 (O_3737,N_49723,N_49033);
or UO_3738 (O_3738,N_49923,N_49425);
nand UO_3739 (O_3739,N_49462,N_48132);
and UO_3740 (O_3740,N_49686,N_49401);
nor UO_3741 (O_3741,N_48544,N_48699);
nand UO_3742 (O_3742,N_49689,N_48033);
or UO_3743 (O_3743,N_49113,N_49355);
and UO_3744 (O_3744,N_48409,N_49659);
and UO_3745 (O_3745,N_49187,N_49819);
xor UO_3746 (O_3746,N_48066,N_49940);
nand UO_3747 (O_3747,N_49550,N_48600);
or UO_3748 (O_3748,N_49880,N_49016);
and UO_3749 (O_3749,N_49899,N_48033);
and UO_3750 (O_3750,N_48142,N_49809);
nand UO_3751 (O_3751,N_49312,N_49542);
or UO_3752 (O_3752,N_49255,N_49435);
nor UO_3753 (O_3753,N_48051,N_49422);
or UO_3754 (O_3754,N_48085,N_49839);
nor UO_3755 (O_3755,N_49002,N_49480);
and UO_3756 (O_3756,N_48840,N_49509);
or UO_3757 (O_3757,N_48693,N_49159);
xnor UO_3758 (O_3758,N_48105,N_49446);
nor UO_3759 (O_3759,N_49972,N_49706);
nor UO_3760 (O_3760,N_49310,N_48605);
and UO_3761 (O_3761,N_48024,N_49995);
xnor UO_3762 (O_3762,N_48752,N_49897);
or UO_3763 (O_3763,N_48583,N_48463);
nor UO_3764 (O_3764,N_49216,N_49363);
and UO_3765 (O_3765,N_49452,N_48640);
nor UO_3766 (O_3766,N_49130,N_49410);
and UO_3767 (O_3767,N_49479,N_48296);
nor UO_3768 (O_3768,N_49966,N_48119);
and UO_3769 (O_3769,N_48034,N_48554);
or UO_3770 (O_3770,N_48414,N_48984);
nor UO_3771 (O_3771,N_49667,N_48578);
nand UO_3772 (O_3772,N_49035,N_48368);
or UO_3773 (O_3773,N_49836,N_48546);
and UO_3774 (O_3774,N_48045,N_49793);
nand UO_3775 (O_3775,N_48871,N_49906);
nand UO_3776 (O_3776,N_49674,N_48221);
and UO_3777 (O_3777,N_48792,N_49126);
or UO_3778 (O_3778,N_49112,N_48281);
and UO_3779 (O_3779,N_48650,N_49727);
and UO_3780 (O_3780,N_48763,N_48145);
or UO_3781 (O_3781,N_48630,N_49797);
nor UO_3782 (O_3782,N_48792,N_48724);
or UO_3783 (O_3783,N_48930,N_49921);
nand UO_3784 (O_3784,N_49174,N_49793);
and UO_3785 (O_3785,N_49182,N_48851);
and UO_3786 (O_3786,N_48538,N_49315);
nand UO_3787 (O_3787,N_48692,N_49344);
nand UO_3788 (O_3788,N_49671,N_48117);
nand UO_3789 (O_3789,N_49428,N_49051);
nor UO_3790 (O_3790,N_48758,N_48656);
nor UO_3791 (O_3791,N_49489,N_49323);
nand UO_3792 (O_3792,N_48613,N_49813);
nor UO_3793 (O_3793,N_48757,N_48596);
nor UO_3794 (O_3794,N_49738,N_49122);
or UO_3795 (O_3795,N_48474,N_48685);
and UO_3796 (O_3796,N_49164,N_49882);
and UO_3797 (O_3797,N_49913,N_48541);
nor UO_3798 (O_3798,N_49674,N_48432);
nor UO_3799 (O_3799,N_48723,N_48165);
nand UO_3800 (O_3800,N_48404,N_48796);
and UO_3801 (O_3801,N_49547,N_49064);
and UO_3802 (O_3802,N_49197,N_48367);
or UO_3803 (O_3803,N_48111,N_48860);
or UO_3804 (O_3804,N_48893,N_49540);
nor UO_3805 (O_3805,N_49907,N_49768);
nand UO_3806 (O_3806,N_49084,N_49588);
or UO_3807 (O_3807,N_48708,N_48209);
and UO_3808 (O_3808,N_49304,N_49952);
nand UO_3809 (O_3809,N_49538,N_48077);
nand UO_3810 (O_3810,N_48789,N_48338);
nand UO_3811 (O_3811,N_48978,N_48563);
or UO_3812 (O_3812,N_49193,N_48110);
and UO_3813 (O_3813,N_48823,N_48081);
nor UO_3814 (O_3814,N_49717,N_49818);
or UO_3815 (O_3815,N_49983,N_49577);
nand UO_3816 (O_3816,N_48215,N_49917);
or UO_3817 (O_3817,N_49257,N_48879);
nor UO_3818 (O_3818,N_49258,N_48161);
nor UO_3819 (O_3819,N_49070,N_49542);
and UO_3820 (O_3820,N_48695,N_49936);
nand UO_3821 (O_3821,N_48351,N_49151);
nand UO_3822 (O_3822,N_48166,N_48996);
and UO_3823 (O_3823,N_48935,N_48422);
and UO_3824 (O_3824,N_48834,N_49046);
nor UO_3825 (O_3825,N_49921,N_49696);
nand UO_3826 (O_3826,N_49169,N_49438);
nand UO_3827 (O_3827,N_49174,N_49299);
nor UO_3828 (O_3828,N_48804,N_48392);
and UO_3829 (O_3829,N_49734,N_49010);
and UO_3830 (O_3830,N_48982,N_49404);
and UO_3831 (O_3831,N_49299,N_48107);
nand UO_3832 (O_3832,N_48856,N_49888);
nor UO_3833 (O_3833,N_48395,N_48158);
and UO_3834 (O_3834,N_48779,N_49451);
nor UO_3835 (O_3835,N_49618,N_48593);
nor UO_3836 (O_3836,N_49109,N_48640);
nand UO_3837 (O_3837,N_48505,N_48517);
or UO_3838 (O_3838,N_49669,N_49364);
nand UO_3839 (O_3839,N_48883,N_48139);
or UO_3840 (O_3840,N_48584,N_49771);
and UO_3841 (O_3841,N_48658,N_48406);
or UO_3842 (O_3842,N_48508,N_49728);
and UO_3843 (O_3843,N_49189,N_48200);
or UO_3844 (O_3844,N_49845,N_49818);
nand UO_3845 (O_3845,N_48630,N_49075);
nand UO_3846 (O_3846,N_49004,N_49249);
and UO_3847 (O_3847,N_48688,N_49065);
nor UO_3848 (O_3848,N_48426,N_48482);
and UO_3849 (O_3849,N_49346,N_48123);
and UO_3850 (O_3850,N_48238,N_48887);
and UO_3851 (O_3851,N_48501,N_49358);
and UO_3852 (O_3852,N_49387,N_49632);
nand UO_3853 (O_3853,N_49820,N_49930);
or UO_3854 (O_3854,N_49472,N_49055);
or UO_3855 (O_3855,N_49251,N_48190);
nand UO_3856 (O_3856,N_49972,N_49502);
nand UO_3857 (O_3857,N_48467,N_49513);
nand UO_3858 (O_3858,N_49940,N_49760);
or UO_3859 (O_3859,N_48246,N_49477);
nor UO_3860 (O_3860,N_48950,N_49165);
or UO_3861 (O_3861,N_48605,N_48591);
nand UO_3862 (O_3862,N_49640,N_49224);
or UO_3863 (O_3863,N_48144,N_48954);
nand UO_3864 (O_3864,N_48917,N_48562);
and UO_3865 (O_3865,N_49721,N_48419);
nor UO_3866 (O_3866,N_48084,N_49623);
nand UO_3867 (O_3867,N_49014,N_48925);
and UO_3868 (O_3868,N_49264,N_48200);
nand UO_3869 (O_3869,N_49834,N_48161);
and UO_3870 (O_3870,N_49395,N_48476);
and UO_3871 (O_3871,N_49076,N_48277);
nand UO_3872 (O_3872,N_48841,N_49846);
nand UO_3873 (O_3873,N_48912,N_49695);
or UO_3874 (O_3874,N_48108,N_48575);
or UO_3875 (O_3875,N_49205,N_48368);
nor UO_3876 (O_3876,N_49732,N_48427);
and UO_3877 (O_3877,N_48809,N_49246);
nand UO_3878 (O_3878,N_49069,N_49294);
nand UO_3879 (O_3879,N_48055,N_49438);
nand UO_3880 (O_3880,N_48343,N_49774);
nor UO_3881 (O_3881,N_48106,N_48073);
nand UO_3882 (O_3882,N_49275,N_49967);
and UO_3883 (O_3883,N_49871,N_49988);
and UO_3884 (O_3884,N_49949,N_49691);
nand UO_3885 (O_3885,N_49858,N_48583);
and UO_3886 (O_3886,N_49789,N_48631);
nand UO_3887 (O_3887,N_49436,N_48197);
and UO_3888 (O_3888,N_49054,N_49192);
and UO_3889 (O_3889,N_49209,N_49072);
and UO_3890 (O_3890,N_48440,N_48129);
or UO_3891 (O_3891,N_48598,N_49740);
nand UO_3892 (O_3892,N_49171,N_49443);
nor UO_3893 (O_3893,N_48578,N_48459);
nor UO_3894 (O_3894,N_48350,N_49615);
or UO_3895 (O_3895,N_49211,N_48762);
and UO_3896 (O_3896,N_49193,N_48810);
or UO_3897 (O_3897,N_49145,N_49560);
and UO_3898 (O_3898,N_49082,N_49551);
nor UO_3899 (O_3899,N_48551,N_48263);
and UO_3900 (O_3900,N_49186,N_48410);
or UO_3901 (O_3901,N_48244,N_49069);
or UO_3902 (O_3902,N_49736,N_49176);
nand UO_3903 (O_3903,N_49698,N_48189);
or UO_3904 (O_3904,N_48164,N_49552);
and UO_3905 (O_3905,N_49838,N_49899);
and UO_3906 (O_3906,N_49465,N_49456);
or UO_3907 (O_3907,N_48128,N_48278);
nand UO_3908 (O_3908,N_49789,N_48808);
nand UO_3909 (O_3909,N_49193,N_49826);
nand UO_3910 (O_3910,N_48278,N_48448);
and UO_3911 (O_3911,N_48247,N_49811);
or UO_3912 (O_3912,N_48073,N_49187);
nand UO_3913 (O_3913,N_48404,N_48387);
and UO_3914 (O_3914,N_49838,N_49880);
nor UO_3915 (O_3915,N_48089,N_49276);
nand UO_3916 (O_3916,N_49306,N_48017);
or UO_3917 (O_3917,N_49045,N_49258);
nand UO_3918 (O_3918,N_48958,N_49660);
or UO_3919 (O_3919,N_48900,N_48322);
and UO_3920 (O_3920,N_49180,N_49123);
nor UO_3921 (O_3921,N_48159,N_48018);
and UO_3922 (O_3922,N_49388,N_48781);
or UO_3923 (O_3923,N_49884,N_48587);
or UO_3924 (O_3924,N_48672,N_49558);
or UO_3925 (O_3925,N_48834,N_49698);
and UO_3926 (O_3926,N_48961,N_49498);
and UO_3927 (O_3927,N_49795,N_49974);
nor UO_3928 (O_3928,N_49087,N_49499);
nor UO_3929 (O_3929,N_49385,N_49003);
or UO_3930 (O_3930,N_49317,N_49425);
nor UO_3931 (O_3931,N_49488,N_49178);
nand UO_3932 (O_3932,N_48605,N_49579);
nor UO_3933 (O_3933,N_48138,N_49220);
or UO_3934 (O_3934,N_48970,N_49099);
and UO_3935 (O_3935,N_49835,N_49813);
nand UO_3936 (O_3936,N_48006,N_49839);
nor UO_3937 (O_3937,N_48452,N_48103);
nor UO_3938 (O_3938,N_48280,N_49764);
xnor UO_3939 (O_3939,N_49270,N_48746);
nand UO_3940 (O_3940,N_49633,N_49098);
nor UO_3941 (O_3941,N_48916,N_48299);
nand UO_3942 (O_3942,N_49857,N_49435);
and UO_3943 (O_3943,N_49669,N_48214);
or UO_3944 (O_3944,N_49746,N_49694);
or UO_3945 (O_3945,N_49287,N_49259);
xor UO_3946 (O_3946,N_48440,N_49789);
and UO_3947 (O_3947,N_48060,N_49251);
nand UO_3948 (O_3948,N_49941,N_48020);
nand UO_3949 (O_3949,N_49581,N_49855);
nor UO_3950 (O_3950,N_48128,N_49016);
nor UO_3951 (O_3951,N_49505,N_49752);
or UO_3952 (O_3952,N_48370,N_49249);
nand UO_3953 (O_3953,N_49453,N_48829);
nor UO_3954 (O_3954,N_48206,N_48180);
nand UO_3955 (O_3955,N_49320,N_48376);
xnor UO_3956 (O_3956,N_49384,N_49009);
nor UO_3957 (O_3957,N_48806,N_49584);
or UO_3958 (O_3958,N_49077,N_48289);
nand UO_3959 (O_3959,N_49297,N_49528);
nor UO_3960 (O_3960,N_48784,N_48027);
or UO_3961 (O_3961,N_48309,N_49808);
nand UO_3962 (O_3962,N_48793,N_49311);
nand UO_3963 (O_3963,N_49386,N_49203);
nand UO_3964 (O_3964,N_48806,N_49804);
and UO_3965 (O_3965,N_48155,N_48350);
or UO_3966 (O_3966,N_48629,N_49317);
and UO_3967 (O_3967,N_48636,N_48862);
or UO_3968 (O_3968,N_48973,N_49583);
or UO_3969 (O_3969,N_49084,N_49355);
nand UO_3970 (O_3970,N_48555,N_48730);
or UO_3971 (O_3971,N_49414,N_49212);
xor UO_3972 (O_3972,N_49037,N_48998);
nor UO_3973 (O_3973,N_49893,N_49462);
or UO_3974 (O_3974,N_48203,N_49826);
nand UO_3975 (O_3975,N_49082,N_48645);
or UO_3976 (O_3976,N_49424,N_49626);
and UO_3977 (O_3977,N_48226,N_48720);
or UO_3978 (O_3978,N_48785,N_48149);
nor UO_3979 (O_3979,N_48468,N_49437);
or UO_3980 (O_3980,N_48441,N_48149);
or UO_3981 (O_3981,N_49420,N_48077);
or UO_3982 (O_3982,N_48121,N_48535);
nor UO_3983 (O_3983,N_48611,N_48883);
nor UO_3984 (O_3984,N_48029,N_48144);
or UO_3985 (O_3985,N_48904,N_49961);
or UO_3986 (O_3986,N_49172,N_49470);
and UO_3987 (O_3987,N_49923,N_49492);
nand UO_3988 (O_3988,N_48487,N_49684);
nor UO_3989 (O_3989,N_48133,N_48759);
nand UO_3990 (O_3990,N_48796,N_49488);
nand UO_3991 (O_3991,N_48173,N_48487);
or UO_3992 (O_3992,N_48406,N_48548);
nor UO_3993 (O_3993,N_49404,N_48306);
nor UO_3994 (O_3994,N_48739,N_48400);
or UO_3995 (O_3995,N_48589,N_48804);
and UO_3996 (O_3996,N_49830,N_49291);
xor UO_3997 (O_3997,N_49510,N_48988);
or UO_3998 (O_3998,N_49089,N_48282);
nand UO_3999 (O_3999,N_49040,N_48451);
nor UO_4000 (O_4000,N_48495,N_48395);
nand UO_4001 (O_4001,N_48825,N_49398);
or UO_4002 (O_4002,N_48078,N_48370);
nor UO_4003 (O_4003,N_48963,N_48917);
and UO_4004 (O_4004,N_49167,N_49224);
nor UO_4005 (O_4005,N_49406,N_48728);
or UO_4006 (O_4006,N_48062,N_48546);
nor UO_4007 (O_4007,N_49401,N_49907);
nand UO_4008 (O_4008,N_48485,N_49262);
and UO_4009 (O_4009,N_48243,N_48986);
nand UO_4010 (O_4010,N_48450,N_48410);
or UO_4011 (O_4011,N_49306,N_49329);
nand UO_4012 (O_4012,N_49839,N_49508);
nand UO_4013 (O_4013,N_49723,N_49714);
and UO_4014 (O_4014,N_49638,N_48165);
nand UO_4015 (O_4015,N_49695,N_49202);
nor UO_4016 (O_4016,N_49542,N_48240);
nand UO_4017 (O_4017,N_49888,N_48811);
or UO_4018 (O_4018,N_48134,N_49863);
nand UO_4019 (O_4019,N_48025,N_48728);
and UO_4020 (O_4020,N_48113,N_49077);
xnor UO_4021 (O_4021,N_49737,N_49643);
nor UO_4022 (O_4022,N_49822,N_49614);
and UO_4023 (O_4023,N_48425,N_48065);
xnor UO_4024 (O_4024,N_49672,N_49490);
or UO_4025 (O_4025,N_48563,N_48634);
and UO_4026 (O_4026,N_49397,N_48643);
nor UO_4027 (O_4027,N_49688,N_48271);
or UO_4028 (O_4028,N_49915,N_48301);
nand UO_4029 (O_4029,N_49655,N_49005);
nand UO_4030 (O_4030,N_48508,N_49989);
or UO_4031 (O_4031,N_48161,N_49025);
nor UO_4032 (O_4032,N_48954,N_48663);
xnor UO_4033 (O_4033,N_49421,N_49707);
and UO_4034 (O_4034,N_48217,N_48232);
and UO_4035 (O_4035,N_48532,N_48488);
nand UO_4036 (O_4036,N_48319,N_48980);
nand UO_4037 (O_4037,N_48608,N_49880);
nand UO_4038 (O_4038,N_48247,N_48827);
and UO_4039 (O_4039,N_49207,N_49546);
xor UO_4040 (O_4040,N_48235,N_49303);
nand UO_4041 (O_4041,N_48907,N_49271);
and UO_4042 (O_4042,N_48191,N_49864);
nor UO_4043 (O_4043,N_49555,N_48351);
nand UO_4044 (O_4044,N_49639,N_49185);
nor UO_4045 (O_4045,N_48025,N_48161);
nor UO_4046 (O_4046,N_49697,N_49532);
nor UO_4047 (O_4047,N_48898,N_49488);
and UO_4048 (O_4048,N_48628,N_48518);
nand UO_4049 (O_4049,N_48441,N_49023);
and UO_4050 (O_4050,N_48514,N_48706);
or UO_4051 (O_4051,N_48228,N_49116);
and UO_4052 (O_4052,N_49135,N_48194);
nand UO_4053 (O_4053,N_49803,N_49062);
nand UO_4054 (O_4054,N_49608,N_48703);
nand UO_4055 (O_4055,N_49045,N_48353);
and UO_4056 (O_4056,N_48866,N_48501);
nor UO_4057 (O_4057,N_49683,N_49689);
or UO_4058 (O_4058,N_49787,N_48493);
or UO_4059 (O_4059,N_48633,N_49525);
or UO_4060 (O_4060,N_49667,N_48919);
and UO_4061 (O_4061,N_48982,N_49772);
nor UO_4062 (O_4062,N_48631,N_48557);
and UO_4063 (O_4063,N_48229,N_49977);
nor UO_4064 (O_4064,N_49577,N_49478);
and UO_4065 (O_4065,N_49338,N_48200);
and UO_4066 (O_4066,N_48846,N_48117);
nor UO_4067 (O_4067,N_48539,N_48766);
and UO_4068 (O_4068,N_49965,N_48202);
or UO_4069 (O_4069,N_49747,N_48455);
nand UO_4070 (O_4070,N_48315,N_48439);
and UO_4071 (O_4071,N_49132,N_48085);
nor UO_4072 (O_4072,N_48615,N_48194);
nor UO_4073 (O_4073,N_49723,N_48064);
and UO_4074 (O_4074,N_48330,N_48229);
nor UO_4075 (O_4075,N_49959,N_49116);
and UO_4076 (O_4076,N_48626,N_48601);
nor UO_4077 (O_4077,N_48743,N_49941);
or UO_4078 (O_4078,N_48745,N_48196);
and UO_4079 (O_4079,N_48155,N_48716);
and UO_4080 (O_4080,N_48350,N_48930);
nor UO_4081 (O_4081,N_49420,N_49251);
or UO_4082 (O_4082,N_48689,N_48433);
nand UO_4083 (O_4083,N_49601,N_49511);
or UO_4084 (O_4084,N_48960,N_49076);
and UO_4085 (O_4085,N_49074,N_48534);
and UO_4086 (O_4086,N_49399,N_48517);
and UO_4087 (O_4087,N_49463,N_48141);
or UO_4088 (O_4088,N_49469,N_48827);
nand UO_4089 (O_4089,N_49927,N_49855);
nor UO_4090 (O_4090,N_49978,N_49289);
and UO_4091 (O_4091,N_48569,N_49876);
xor UO_4092 (O_4092,N_49323,N_49867);
nand UO_4093 (O_4093,N_49659,N_48603);
and UO_4094 (O_4094,N_48558,N_48649);
nor UO_4095 (O_4095,N_49320,N_49511);
or UO_4096 (O_4096,N_49952,N_48398);
nor UO_4097 (O_4097,N_49705,N_48144);
xnor UO_4098 (O_4098,N_48241,N_49490);
or UO_4099 (O_4099,N_48016,N_48401);
or UO_4100 (O_4100,N_49274,N_48699);
or UO_4101 (O_4101,N_48625,N_48280);
or UO_4102 (O_4102,N_49845,N_48141);
nor UO_4103 (O_4103,N_49363,N_48889);
nor UO_4104 (O_4104,N_48215,N_49918);
and UO_4105 (O_4105,N_49156,N_49859);
and UO_4106 (O_4106,N_48885,N_48283);
and UO_4107 (O_4107,N_48123,N_49077);
or UO_4108 (O_4108,N_49585,N_48016);
and UO_4109 (O_4109,N_49717,N_48154);
nand UO_4110 (O_4110,N_49405,N_49440);
nor UO_4111 (O_4111,N_49404,N_49479);
and UO_4112 (O_4112,N_48712,N_49341);
nor UO_4113 (O_4113,N_48096,N_49591);
and UO_4114 (O_4114,N_49931,N_49094);
and UO_4115 (O_4115,N_49152,N_48509);
or UO_4116 (O_4116,N_48600,N_48376);
nand UO_4117 (O_4117,N_49744,N_48139);
nor UO_4118 (O_4118,N_49362,N_48555);
and UO_4119 (O_4119,N_48354,N_49973);
or UO_4120 (O_4120,N_49017,N_48042);
xnor UO_4121 (O_4121,N_48767,N_48484);
nand UO_4122 (O_4122,N_48462,N_49804);
nor UO_4123 (O_4123,N_49374,N_48119);
or UO_4124 (O_4124,N_49651,N_48837);
nand UO_4125 (O_4125,N_49962,N_48852);
nor UO_4126 (O_4126,N_49285,N_48553);
and UO_4127 (O_4127,N_48412,N_49330);
nor UO_4128 (O_4128,N_49909,N_49195);
nor UO_4129 (O_4129,N_49066,N_49763);
or UO_4130 (O_4130,N_48671,N_48388);
nand UO_4131 (O_4131,N_48721,N_48407);
xor UO_4132 (O_4132,N_48364,N_49671);
nand UO_4133 (O_4133,N_49752,N_48871);
nand UO_4134 (O_4134,N_48270,N_49108);
nand UO_4135 (O_4135,N_48906,N_49082);
or UO_4136 (O_4136,N_48205,N_48124);
nor UO_4137 (O_4137,N_49133,N_48047);
nor UO_4138 (O_4138,N_49743,N_49750);
and UO_4139 (O_4139,N_49170,N_49722);
or UO_4140 (O_4140,N_49416,N_48984);
nand UO_4141 (O_4141,N_48013,N_48988);
nand UO_4142 (O_4142,N_49428,N_49495);
nand UO_4143 (O_4143,N_48908,N_49181);
xnor UO_4144 (O_4144,N_49634,N_48866);
nand UO_4145 (O_4145,N_48050,N_48938);
nor UO_4146 (O_4146,N_49607,N_49524);
or UO_4147 (O_4147,N_49924,N_48010);
nor UO_4148 (O_4148,N_48100,N_48865);
and UO_4149 (O_4149,N_49454,N_49656);
nand UO_4150 (O_4150,N_49153,N_49665);
nor UO_4151 (O_4151,N_49228,N_49941);
nand UO_4152 (O_4152,N_49422,N_48102);
or UO_4153 (O_4153,N_49169,N_49810);
nor UO_4154 (O_4154,N_49507,N_49700);
xor UO_4155 (O_4155,N_48543,N_48160);
and UO_4156 (O_4156,N_49954,N_49641);
and UO_4157 (O_4157,N_49631,N_49363);
and UO_4158 (O_4158,N_49317,N_48973);
nor UO_4159 (O_4159,N_49988,N_49183);
nand UO_4160 (O_4160,N_48588,N_48674);
and UO_4161 (O_4161,N_49000,N_48452);
or UO_4162 (O_4162,N_49441,N_48541);
nor UO_4163 (O_4163,N_49787,N_49773);
or UO_4164 (O_4164,N_49939,N_49181);
or UO_4165 (O_4165,N_49495,N_48083);
and UO_4166 (O_4166,N_48676,N_49758);
and UO_4167 (O_4167,N_48235,N_48618);
nand UO_4168 (O_4168,N_49157,N_48573);
nor UO_4169 (O_4169,N_49622,N_49882);
and UO_4170 (O_4170,N_48427,N_49796);
nand UO_4171 (O_4171,N_48066,N_49054);
nor UO_4172 (O_4172,N_48566,N_49715);
and UO_4173 (O_4173,N_49652,N_49289);
or UO_4174 (O_4174,N_49146,N_49754);
xnor UO_4175 (O_4175,N_48244,N_48626);
or UO_4176 (O_4176,N_49243,N_48213);
nor UO_4177 (O_4177,N_49270,N_48761);
nand UO_4178 (O_4178,N_49989,N_48600);
nor UO_4179 (O_4179,N_48030,N_48172);
and UO_4180 (O_4180,N_49926,N_48097);
nand UO_4181 (O_4181,N_48153,N_48776);
nor UO_4182 (O_4182,N_48961,N_48553);
and UO_4183 (O_4183,N_49936,N_49486);
and UO_4184 (O_4184,N_49787,N_49791);
nor UO_4185 (O_4185,N_48818,N_48419);
nor UO_4186 (O_4186,N_48444,N_49813);
and UO_4187 (O_4187,N_48741,N_48817);
and UO_4188 (O_4188,N_48043,N_48478);
and UO_4189 (O_4189,N_48686,N_48175);
and UO_4190 (O_4190,N_48727,N_48073);
and UO_4191 (O_4191,N_48561,N_49266);
or UO_4192 (O_4192,N_48805,N_49469);
nor UO_4193 (O_4193,N_48131,N_48860);
nor UO_4194 (O_4194,N_48042,N_49637);
and UO_4195 (O_4195,N_49238,N_49777);
nand UO_4196 (O_4196,N_49282,N_49669);
nor UO_4197 (O_4197,N_48082,N_49761);
or UO_4198 (O_4198,N_49710,N_49157);
and UO_4199 (O_4199,N_48884,N_49412);
nand UO_4200 (O_4200,N_49203,N_49567);
nor UO_4201 (O_4201,N_49490,N_49422);
or UO_4202 (O_4202,N_48907,N_48939);
nand UO_4203 (O_4203,N_49540,N_48937);
nor UO_4204 (O_4204,N_48174,N_49218);
nor UO_4205 (O_4205,N_49223,N_48782);
and UO_4206 (O_4206,N_49036,N_48620);
nand UO_4207 (O_4207,N_49533,N_49027);
nor UO_4208 (O_4208,N_49812,N_48770);
nand UO_4209 (O_4209,N_49496,N_49289);
nor UO_4210 (O_4210,N_48398,N_49851);
nand UO_4211 (O_4211,N_49778,N_49963);
nand UO_4212 (O_4212,N_49850,N_49544);
nand UO_4213 (O_4213,N_49781,N_48713);
nand UO_4214 (O_4214,N_49079,N_49395);
and UO_4215 (O_4215,N_49287,N_49189);
or UO_4216 (O_4216,N_48212,N_48408);
nand UO_4217 (O_4217,N_49614,N_48412);
and UO_4218 (O_4218,N_48018,N_49262);
nor UO_4219 (O_4219,N_48360,N_49928);
and UO_4220 (O_4220,N_49154,N_48592);
or UO_4221 (O_4221,N_49349,N_48485);
nor UO_4222 (O_4222,N_49290,N_48169);
nor UO_4223 (O_4223,N_49202,N_48619);
nand UO_4224 (O_4224,N_49839,N_48501);
or UO_4225 (O_4225,N_48634,N_49581);
and UO_4226 (O_4226,N_48067,N_48053);
nand UO_4227 (O_4227,N_48452,N_48557);
or UO_4228 (O_4228,N_49560,N_49291);
nand UO_4229 (O_4229,N_49058,N_48766);
xor UO_4230 (O_4230,N_49341,N_49488);
nor UO_4231 (O_4231,N_49511,N_48508);
and UO_4232 (O_4232,N_49469,N_48061);
or UO_4233 (O_4233,N_48888,N_48733);
nand UO_4234 (O_4234,N_48894,N_49880);
nand UO_4235 (O_4235,N_48793,N_48288);
nor UO_4236 (O_4236,N_49216,N_49532);
or UO_4237 (O_4237,N_48939,N_48419);
and UO_4238 (O_4238,N_49102,N_48929);
and UO_4239 (O_4239,N_48552,N_48198);
nand UO_4240 (O_4240,N_49706,N_48007);
nand UO_4241 (O_4241,N_48598,N_48991);
or UO_4242 (O_4242,N_49217,N_49931);
nand UO_4243 (O_4243,N_48837,N_49449);
nand UO_4244 (O_4244,N_49034,N_49899);
and UO_4245 (O_4245,N_48828,N_49896);
nand UO_4246 (O_4246,N_48848,N_48058);
or UO_4247 (O_4247,N_49665,N_49892);
nand UO_4248 (O_4248,N_48265,N_48811);
nand UO_4249 (O_4249,N_49113,N_49316);
nand UO_4250 (O_4250,N_49479,N_49347);
or UO_4251 (O_4251,N_48969,N_48284);
and UO_4252 (O_4252,N_48447,N_49062);
and UO_4253 (O_4253,N_48374,N_49516);
or UO_4254 (O_4254,N_48276,N_49594);
nand UO_4255 (O_4255,N_49759,N_48510);
and UO_4256 (O_4256,N_48953,N_49080);
and UO_4257 (O_4257,N_49635,N_49752);
and UO_4258 (O_4258,N_48392,N_48728);
nor UO_4259 (O_4259,N_48794,N_48944);
and UO_4260 (O_4260,N_48906,N_49670);
nand UO_4261 (O_4261,N_48796,N_48942);
and UO_4262 (O_4262,N_48926,N_48599);
or UO_4263 (O_4263,N_49831,N_48688);
and UO_4264 (O_4264,N_48437,N_48486);
nand UO_4265 (O_4265,N_49263,N_48688);
nor UO_4266 (O_4266,N_49866,N_48408);
nor UO_4267 (O_4267,N_49771,N_49144);
nand UO_4268 (O_4268,N_48964,N_49410);
or UO_4269 (O_4269,N_48246,N_49157);
nor UO_4270 (O_4270,N_48781,N_48383);
nand UO_4271 (O_4271,N_48189,N_49666);
or UO_4272 (O_4272,N_49166,N_48961);
nand UO_4273 (O_4273,N_49239,N_48016);
and UO_4274 (O_4274,N_48362,N_48853);
and UO_4275 (O_4275,N_49481,N_48760);
nand UO_4276 (O_4276,N_49506,N_48082);
and UO_4277 (O_4277,N_49087,N_48575);
nand UO_4278 (O_4278,N_49068,N_48860);
nor UO_4279 (O_4279,N_49484,N_49046);
or UO_4280 (O_4280,N_49954,N_49966);
nor UO_4281 (O_4281,N_49882,N_49448);
and UO_4282 (O_4282,N_48497,N_49669);
nor UO_4283 (O_4283,N_49895,N_48069);
and UO_4284 (O_4284,N_48546,N_48711);
or UO_4285 (O_4285,N_48860,N_48500);
nor UO_4286 (O_4286,N_49188,N_49372);
or UO_4287 (O_4287,N_49329,N_48887);
or UO_4288 (O_4288,N_48703,N_49888);
nand UO_4289 (O_4289,N_48577,N_49472);
or UO_4290 (O_4290,N_49083,N_49946);
and UO_4291 (O_4291,N_49860,N_48010);
or UO_4292 (O_4292,N_49966,N_49538);
and UO_4293 (O_4293,N_49882,N_48924);
nand UO_4294 (O_4294,N_49843,N_49446);
nor UO_4295 (O_4295,N_48864,N_48565);
and UO_4296 (O_4296,N_49564,N_49201);
nor UO_4297 (O_4297,N_48000,N_49884);
nand UO_4298 (O_4298,N_48748,N_49905);
or UO_4299 (O_4299,N_48703,N_49901);
nor UO_4300 (O_4300,N_48202,N_49567);
nor UO_4301 (O_4301,N_48688,N_49715);
nand UO_4302 (O_4302,N_49774,N_48812);
xnor UO_4303 (O_4303,N_48232,N_48481);
and UO_4304 (O_4304,N_49230,N_48088);
nand UO_4305 (O_4305,N_48814,N_49487);
or UO_4306 (O_4306,N_49283,N_48587);
or UO_4307 (O_4307,N_49468,N_49551);
and UO_4308 (O_4308,N_48300,N_49164);
nor UO_4309 (O_4309,N_49936,N_49540);
or UO_4310 (O_4310,N_49685,N_48955);
and UO_4311 (O_4311,N_48266,N_49813);
or UO_4312 (O_4312,N_49122,N_48582);
nor UO_4313 (O_4313,N_48182,N_49901);
and UO_4314 (O_4314,N_48573,N_48950);
and UO_4315 (O_4315,N_49579,N_48355);
nand UO_4316 (O_4316,N_49148,N_48322);
and UO_4317 (O_4317,N_49257,N_48828);
or UO_4318 (O_4318,N_49291,N_48465);
nand UO_4319 (O_4319,N_49170,N_48868);
nand UO_4320 (O_4320,N_48004,N_49484);
nor UO_4321 (O_4321,N_48176,N_48030);
nand UO_4322 (O_4322,N_49232,N_48846);
nor UO_4323 (O_4323,N_49530,N_49792);
and UO_4324 (O_4324,N_49791,N_49013);
and UO_4325 (O_4325,N_49548,N_49293);
nor UO_4326 (O_4326,N_49804,N_49310);
nand UO_4327 (O_4327,N_49132,N_49330);
nand UO_4328 (O_4328,N_48496,N_48455);
or UO_4329 (O_4329,N_48957,N_48073);
and UO_4330 (O_4330,N_48700,N_48297);
or UO_4331 (O_4331,N_48166,N_49776);
and UO_4332 (O_4332,N_48736,N_48571);
and UO_4333 (O_4333,N_49114,N_48455);
and UO_4334 (O_4334,N_48087,N_48256);
and UO_4335 (O_4335,N_48609,N_48789);
or UO_4336 (O_4336,N_49525,N_48435);
nand UO_4337 (O_4337,N_49852,N_48422);
and UO_4338 (O_4338,N_49022,N_48728);
nand UO_4339 (O_4339,N_48937,N_48244);
or UO_4340 (O_4340,N_49009,N_49369);
nor UO_4341 (O_4341,N_49519,N_49254);
nor UO_4342 (O_4342,N_48707,N_49246);
nand UO_4343 (O_4343,N_48680,N_49503);
or UO_4344 (O_4344,N_49982,N_49237);
and UO_4345 (O_4345,N_48819,N_49530);
nor UO_4346 (O_4346,N_49466,N_48908);
nor UO_4347 (O_4347,N_49969,N_48091);
nand UO_4348 (O_4348,N_48128,N_48920);
xnor UO_4349 (O_4349,N_48372,N_48145);
or UO_4350 (O_4350,N_49184,N_49718);
or UO_4351 (O_4351,N_48296,N_49497);
or UO_4352 (O_4352,N_49037,N_49457);
or UO_4353 (O_4353,N_49351,N_48063);
or UO_4354 (O_4354,N_48055,N_48421);
and UO_4355 (O_4355,N_49023,N_49617);
nor UO_4356 (O_4356,N_48461,N_48388);
or UO_4357 (O_4357,N_48033,N_48116);
or UO_4358 (O_4358,N_48524,N_48062);
nand UO_4359 (O_4359,N_48856,N_48389);
and UO_4360 (O_4360,N_48566,N_48553);
nand UO_4361 (O_4361,N_48635,N_49209);
and UO_4362 (O_4362,N_48764,N_48813);
nand UO_4363 (O_4363,N_48471,N_48261);
xnor UO_4364 (O_4364,N_49380,N_48721);
nand UO_4365 (O_4365,N_48489,N_48130);
or UO_4366 (O_4366,N_48739,N_48192);
nand UO_4367 (O_4367,N_48820,N_48274);
nor UO_4368 (O_4368,N_49226,N_49881);
or UO_4369 (O_4369,N_48284,N_49935);
nand UO_4370 (O_4370,N_48523,N_49979);
nand UO_4371 (O_4371,N_48152,N_49611);
and UO_4372 (O_4372,N_49728,N_48106);
or UO_4373 (O_4373,N_49931,N_49427);
or UO_4374 (O_4374,N_49883,N_48181);
and UO_4375 (O_4375,N_48303,N_48121);
nor UO_4376 (O_4376,N_48795,N_49196);
and UO_4377 (O_4377,N_48644,N_49064);
nor UO_4378 (O_4378,N_48777,N_48558);
and UO_4379 (O_4379,N_48316,N_48575);
nand UO_4380 (O_4380,N_48838,N_49685);
and UO_4381 (O_4381,N_49169,N_48081);
nor UO_4382 (O_4382,N_48476,N_48000);
and UO_4383 (O_4383,N_49439,N_49405);
nor UO_4384 (O_4384,N_48777,N_49499);
nor UO_4385 (O_4385,N_48949,N_48561);
or UO_4386 (O_4386,N_48436,N_49462);
nand UO_4387 (O_4387,N_48740,N_49831);
or UO_4388 (O_4388,N_49000,N_48289);
nor UO_4389 (O_4389,N_49153,N_48510);
nand UO_4390 (O_4390,N_48537,N_49666);
or UO_4391 (O_4391,N_49257,N_49495);
nand UO_4392 (O_4392,N_49572,N_49653);
nand UO_4393 (O_4393,N_48466,N_49159);
nand UO_4394 (O_4394,N_49683,N_48953);
or UO_4395 (O_4395,N_49233,N_49682);
xor UO_4396 (O_4396,N_49180,N_49637);
nand UO_4397 (O_4397,N_49113,N_48687);
or UO_4398 (O_4398,N_49028,N_49472);
nand UO_4399 (O_4399,N_48290,N_48234);
nand UO_4400 (O_4400,N_48636,N_48791);
nor UO_4401 (O_4401,N_49624,N_49610);
nor UO_4402 (O_4402,N_49381,N_48632);
nand UO_4403 (O_4403,N_48651,N_48958);
and UO_4404 (O_4404,N_48147,N_48719);
or UO_4405 (O_4405,N_48124,N_49754);
and UO_4406 (O_4406,N_49144,N_49917);
nand UO_4407 (O_4407,N_48971,N_49813);
and UO_4408 (O_4408,N_49714,N_48670);
nor UO_4409 (O_4409,N_48848,N_49424);
nor UO_4410 (O_4410,N_49716,N_48388);
and UO_4411 (O_4411,N_48881,N_49529);
nor UO_4412 (O_4412,N_49715,N_48861);
and UO_4413 (O_4413,N_48685,N_49136);
or UO_4414 (O_4414,N_48219,N_49100);
and UO_4415 (O_4415,N_48939,N_49123);
nand UO_4416 (O_4416,N_49628,N_48700);
and UO_4417 (O_4417,N_48273,N_49325);
nand UO_4418 (O_4418,N_49663,N_49525);
and UO_4419 (O_4419,N_49480,N_48963);
nor UO_4420 (O_4420,N_48452,N_48286);
and UO_4421 (O_4421,N_49152,N_48058);
nand UO_4422 (O_4422,N_48662,N_49130);
or UO_4423 (O_4423,N_49430,N_49327);
or UO_4424 (O_4424,N_49120,N_48671);
and UO_4425 (O_4425,N_48782,N_49723);
nor UO_4426 (O_4426,N_49367,N_48401);
nand UO_4427 (O_4427,N_49690,N_49427);
or UO_4428 (O_4428,N_49837,N_49342);
nor UO_4429 (O_4429,N_49300,N_49783);
and UO_4430 (O_4430,N_48776,N_49700);
nand UO_4431 (O_4431,N_49680,N_49113);
nand UO_4432 (O_4432,N_48802,N_49799);
or UO_4433 (O_4433,N_49726,N_48775);
nand UO_4434 (O_4434,N_49748,N_48343);
nor UO_4435 (O_4435,N_49037,N_48892);
nor UO_4436 (O_4436,N_48904,N_49427);
or UO_4437 (O_4437,N_49633,N_48503);
nor UO_4438 (O_4438,N_48875,N_49476);
nand UO_4439 (O_4439,N_48041,N_49370);
and UO_4440 (O_4440,N_49500,N_48047);
nand UO_4441 (O_4441,N_48714,N_49474);
nand UO_4442 (O_4442,N_48482,N_49955);
and UO_4443 (O_4443,N_49259,N_49082);
nand UO_4444 (O_4444,N_48801,N_49714);
nand UO_4445 (O_4445,N_49351,N_48834);
and UO_4446 (O_4446,N_49127,N_49027);
or UO_4447 (O_4447,N_49023,N_48888);
and UO_4448 (O_4448,N_48342,N_49687);
nor UO_4449 (O_4449,N_49766,N_48666);
or UO_4450 (O_4450,N_49152,N_49685);
nand UO_4451 (O_4451,N_48348,N_48739);
nand UO_4452 (O_4452,N_48083,N_49847);
nor UO_4453 (O_4453,N_48365,N_49789);
nand UO_4454 (O_4454,N_48391,N_48711);
and UO_4455 (O_4455,N_49645,N_49986);
and UO_4456 (O_4456,N_49368,N_49353);
or UO_4457 (O_4457,N_48050,N_48865);
or UO_4458 (O_4458,N_49689,N_49214);
or UO_4459 (O_4459,N_49907,N_49551);
and UO_4460 (O_4460,N_48570,N_49915);
or UO_4461 (O_4461,N_48443,N_48454);
and UO_4462 (O_4462,N_49506,N_48256);
and UO_4463 (O_4463,N_49471,N_49659);
and UO_4464 (O_4464,N_48337,N_49245);
and UO_4465 (O_4465,N_48866,N_49900);
nor UO_4466 (O_4466,N_49171,N_48257);
and UO_4467 (O_4467,N_48612,N_48356);
nor UO_4468 (O_4468,N_48159,N_48777);
nand UO_4469 (O_4469,N_48796,N_49644);
nand UO_4470 (O_4470,N_48208,N_49154);
nor UO_4471 (O_4471,N_48451,N_48038);
nor UO_4472 (O_4472,N_49535,N_48203);
xnor UO_4473 (O_4473,N_49688,N_49235);
or UO_4474 (O_4474,N_48115,N_49893);
and UO_4475 (O_4475,N_48469,N_48336);
and UO_4476 (O_4476,N_48310,N_49058);
and UO_4477 (O_4477,N_48018,N_48080);
and UO_4478 (O_4478,N_48176,N_48895);
and UO_4479 (O_4479,N_48239,N_49561);
nor UO_4480 (O_4480,N_49835,N_49558);
nand UO_4481 (O_4481,N_49386,N_49487);
and UO_4482 (O_4482,N_49702,N_49078);
nor UO_4483 (O_4483,N_49599,N_49978);
or UO_4484 (O_4484,N_49908,N_49393);
xor UO_4485 (O_4485,N_49594,N_48790);
nand UO_4486 (O_4486,N_49320,N_49560);
nand UO_4487 (O_4487,N_48357,N_48747);
and UO_4488 (O_4488,N_49298,N_49336);
nand UO_4489 (O_4489,N_48281,N_48392);
nand UO_4490 (O_4490,N_49269,N_49890);
nand UO_4491 (O_4491,N_49097,N_48418);
nor UO_4492 (O_4492,N_49211,N_48957);
or UO_4493 (O_4493,N_48075,N_48078);
nor UO_4494 (O_4494,N_49735,N_48761);
or UO_4495 (O_4495,N_49833,N_49883);
or UO_4496 (O_4496,N_48929,N_48563);
and UO_4497 (O_4497,N_48476,N_49732);
nand UO_4498 (O_4498,N_48474,N_48181);
nand UO_4499 (O_4499,N_49893,N_49542);
and UO_4500 (O_4500,N_49803,N_49842);
or UO_4501 (O_4501,N_49862,N_48197);
and UO_4502 (O_4502,N_49199,N_48269);
and UO_4503 (O_4503,N_49630,N_49727);
nand UO_4504 (O_4504,N_49944,N_48426);
nand UO_4505 (O_4505,N_48741,N_49649);
nor UO_4506 (O_4506,N_49285,N_49373);
nand UO_4507 (O_4507,N_49680,N_48745);
nand UO_4508 (O_4508,N_48810,N_48119);
nor UO_4509 (O_4509,N_48046,N_49244);
or UO_4510 (O_4510,N_48067,N_48971);
nor UO_4511 (O_4511,N_48018,N_49732);
nand UO_4512 (O_4512,N_48791,N_48727);
nand UO_4513 (O_4513,N_48790,N_48625);
or UO_4514 (O_4514,N_49035,N_49160);
and UO_4515 (O_4515,N_49083,N_48554);
nand UO_4516 (O_4516,N_48142,N_49400);
or UO_4517 (O_4517,N_48367,N_49565);
or UO_4518 (O_4518,N_48841,N_48559);
and UO_4519 (O_4519,N_48431,N_49185);
nor UO_4520 (O_4520,N_48108,N_49441);
nor UO_4521 (O_4521,N_49876,N_49975);
and UO_4522 (O_4522,N_49285,N_49492);
nor UO_4523 (O_4523,N_49742,N_49498);
nand UO_4524 (O_4524,N_49695,N_48937);
nor UO_4525 (O_4525,N_49073,N_49236);
nor UO_4526 (O_4526,N_49608,N_49775);
nor UO_4527 (O_4527,N_48421,N_48414);
nor UO_4528 (O_4528,N_48864,N_48704);
nor UO_4529 (O_4529,N_49772,N_49994);
nor UO_4530 (O_4530,N_49606,N_49311);
nand UO_4531 (O_4531,N_49537,N_49641);
or UO_4532 (O_4532,N_48280,N_49651);
and UO_4533 (O_4533,N_49651,N_49715);
or UO_4534 (O_4534,N_48215,N_49596);
nor UO_4535 (O_4535,N_49896,N_49182);
or UO_4536 (O_4536,N_49997,N_49827);
nand UO_4537 (O_4537,N_48812,N_49871);
nor UO_4538 (O_4538,N_49287,N_48794);
and UO_4539 (O_4539,N_48943,N_49925);
nand UO_4540 (O_4540,N_49977,N_49645);
and UO_4541 (O_4541,N_49721,N_49467);
or UO_4542 (O_4542,N_49432,N_48192);
nor UO_4543 (O_4543,N_49264,N_48863);
and UO_4544 (O_4544,N_49161,N_48111);
nand UO_4545 (O_4545,N_49062,N_48916);
nand UO_4546 (O_4546,N_49596,N_48672);
and UO_4547 (O_4547,N_48888,N_49192);
and UO_4548 (O_4548,N_49907,N_48049);
nor UO_4549 (O_4549,N_48049,N_48700);
and UO_4550 (O_4550,N_48548,N_49581);
nand UO_4551 (O_4551,N_49061,N_48687);
and UO_4552 (O_4552,N_49995,N_48030);
nor UO_4553 (O_4553,N_49850,N_49167);
and UO_4554 (O_4554,N_49106,N_48811);
and UO_4555 (O_4555,N_48841,N_49595);
xor UO_4556 (O_4556,N_49254,N_49193);
xor UO_4557 (O_4557,N_48394,N_48203);
nand UO_4558 (O_4558,N_48875,N_49794);
xor UO_4559 (O_4559,N_49151,N_48659);
nor UO_4560 (O_4560,N_49891,N_48328);
nor UO_4561 (O_4561,N_48702,N_48887);
nor UO_4562 (O_4562,N_48127,N_48702);
nand UO_4563 (O_4563,N_48536,N_49649);
nor UO_4564 (O_4564,N_48807,N_49451);
nor UO_4565 (O_4565,N_49371,N_48958);
or UO_4566 (O_4566,N_48985,N_49667);
or UO_4567 (O_4567,N_49813,N_48303);
nor UO_4568 (O_4568,N_49829,N_48005);
or UO_4569 (O_4569,N_49579,N_48071);
nor UO_4570 (O_4570,N_48214,N_49522);
nor UO_4571 (O_4571,N_48161,N_49870);
or UO_4572 (O_4572,N_49975,N_48571);
or UO_4573 (O_4573,N_48102,N_49563);
and UO_4574 (O_4574,N_49035,N_48200);
nand UO_4575 (O_4575,N_49379,N_49810);
or UO_4576 (O_4576,N_48922,N_48018);
nor UO_4577 (O_4577,N_49643,N_49188);
nor UO_4578 (O_4578,N_49731,N_49818);
nand UO_4579 (O_4579,N_49870,N_48589);
nand UO_4580 (O_4580,N_48873,N_48640);
or UO_4581 (O_4581,N_49425,N_49640);
nand UO_4582 (O_4582,N_49109,N_49288);
and UO_4583 (O_4583,N_48653,N_49130);
nand UO_4584 (O_4584,N_48264,N_48139);
nor UO_4585 (O_4585,N_49408,N_48313);
and UO_4586 (O_4586,N_49591,N_49068);
or UO_4587 (O_4587,N_48896,N_49568);
or UO_4588 (O_4588,N_48887,N_48349);
or UO_4589 (O_4589,N_48176,N_49509);
and UO_4590 (O_4590,N_48532,N_48260);
nand UO_4591 (O_4591,N_49206,N_48015);
nand UO_4592 (O_4592,N_48081,N_49108);
or UO_4593 (O_4593,N_48136,N_48626);
or UO_4594 (O_4594,N_48618,N_49200);
or UO_4595 (O_4595,N_48500,N_49347);
and UO_4596 (O_4596,N_48687,N_48004);
nor UO_4597 (O_4597,N_48399,N_49809);
or UO_4598 (O_4598,N_49556,N_49420);
or UO_4599 (O_4599,N_48253,N_49266);
or UO_4600 (O_4600,N_49377,N_49904);
or UO_4601 (O_4601,N_48421,N_49528);
or UO_4602 (O_4602,N_48781,N_48692);
or UO_4603 (O_4603,N_49731,N_48947);
and UO_4604 (O_4604,N_48048,N_48510);
or UO_4605 (O_4605,N_48242,N_49250);
or UO_4606 (O_4606,N_48232,N_48694);
nor UO_4607 (O_4607,N_48390,N_48191);
and UO_4608 (O_4608,N_48778,N_49394);
nand UO_4609 (O_4609,N_48984,N_48977);
nand UO_4610 (O_4610,N_49745,N_48909);
xor UO_4611 (O_4611,N_48723,N_49510);
xor UO_4612 (O_4612,N_49561,N_48687);
or UO_4613 (O_4613,N_48835,N_48666);
or UO_4614 (O_4614,N_49554,N_48006);
or UO_4615 (O_4615,N_49330,N_49968);
and UO_4616 (O_4616,N_49744,N_49654);
nand UO_4617 (O_4617,N_49919,N_49634);
nand UO_4618 (O_4618,N_48759,N_49349);
nand UO_4619 (O_4619,N_49085,N_49653);
nor UO_4620 (O_4620,N_48557,N_48497);
and UO_4621 (O_4621,N_48842,N_49121);
nor UO_4622 (O_4622,N_49655,N_48075);
nor UO_4623 (O_4623,N_48489,N_48114);
and UO_4624 (O_4624,N_49292,N_48458);
nand UO_4625 (O_4625,N_48497,N_49904);
xnor UO_4626 (O_4626,N_49267,N_48119);
nand UO_4627 (O_4627,N_48017,N_49678);
nand UO_4628 (O_4628,N_49763,N_49445);
and UO_4629 (O_4629,N_48587,N_49124);
nand UO_4630 (O_4630,N_49155,N_49997);
or UO_4631 (O_4631,N_49633,N_48885);
nand UO_4632 (O_4632,N_49401,N_48655);
and UO_4633 (O_4633,N_49738,N_49969);
nor UO_4634 (O_4634,N_48077,N_49921);
and UO_4635 (O_4635,N_48853,N_48587);
nand UO_4636 (O_4636,N_48343,N_48404);
or UO_4637 (O_4637,N_49538,N_49521);
or UO_4638 (O_4638,N_48772,N_49163);
nand UO_4639 (O_4639,N_49407,N_48545);
nor UO_4640 (O_4640,N_48509,N_49289);
and UO_4641 (O_4641,N_49311,N_48100);
nand UO_4642 (O_4642,N_49773,N_49054);
xor UO_4643 (O_4643,N_48775,N_48404);
or UO_4644 (O_4644,N_48408,N_49291);
and UO_4645 (O_4645,N_48461,N_49802);
nor UO_4646 (O_4646,N_49811,N_49773);
or UO_4647 (O_4647,N_49740,N_49950);
nand UO_4648 (O_4648,N_49329,N_49344);
and UO_4649 (O_4649,N_49089,N_48045);
and UO_4650 (O_4650,N_49709,N_48179);
and UO_4651 (O_4651,N_48113,N_48077);
and UO_4652 (O_4652,N_49437,N_49153);
and UO_4653 (O_4653,N_49538,N_49875);
and UO_4654 (O_4654,N_49338,N_48399);
or UO_4655 (O_4655,N_49223,N_49886);
nor UO_4656 (O_4656,N_49304,N_48567);
and UO_4657 (O_4657,N_49365,N_48576);
nor UO_4658 (O_4658,N_49892,N_49497);
or UO_4659 (O_4659,N_48147,N_49992);
nor UO_4660 (O_4660,N_48006,N_49504);
nor UO_4661 (O_4661,N_48428,N_48049);
or UO_4662 (O_4662,N_49637,N_49077);
nor UO_4663 (O_4663,N_49403,N_49420);
or UO_4664 (O_4664,N_49026,N_48603);
nand UO_4665 (O_4665,N_48646,N_49000);
nor UO_4666 (O_4666,N_48297,N_48341);
and UO_4667 (O_4667,N_48973,N_49162);
or UO_4668 (O_4668,N_48021,N_48771);
nand UO_4669 (O_4669,N_48370,N_49228);
nor UO_4670 (O_4670,N_49166,N_48156);
nor UO_4671 (O_4671,N_49553,N_49687);
nand UO_4672 (O_4672,N_48663,N_48420);
or UO_4673 (O_4673,N_48774,N_49746);
or UO_4674 (O_4674,N_48765,N_48433);
nor UO_4675 (O_4675,N_49470,N_49025);
and UO_4676 (O_4676,N_49448,N_49824);
and UO_4677 (O_4677,N_48534,N_48192);
and UO_4678 (O_4678,N_48478,N_48609);
and UO_4679 (O_4679,N_49404,N_48590);
or UO_4680 (O_4680,N_49635,N_48889);
or UO_4681 (O_4681,N_49298,N_49308);
nand UO_4682 (O_4682,N_49330,N_48134);
nand UO_4683 (O_4683,N_49844,N_48816);
xnor UO_4684 (O_4684,N_48392,N_48428);
or UO_4685 (O_4685,N_49643,N_49030);
nor UO_4686 (O_4686,N_48560,N_49066);
or UO_4687 (O_4687,N_49465,N_49347);
nand UO_4688 (O_4688,N_48412,N_48297);
nor UO_4689 (O_4689,N_49866,N_49418);
and UO_4690 (O_4690,N_49468,N_48014);
nor UO_4691 (O_4691,N_49575,N_48400);
or UO_4692 (O_4692,N_48374,N_49451);
and UO_4693 (O_4693,N_48011,N_48986);
and UO_4694 (O_4694,N_48659,N_48572);
nor UO_4695 (O_4695,N_49687,N_48163);
nand UO_4696 (O_4696,N_48133,N_48752);
and UO_4697 (O_4697,N_49505,N_49617);
nand UO_4698 (O_4698,N_49331,N_49955);
or UO_4699 (O_4699,N_48815,N_49361);
nor UO_4700 (O_4700,N_48272,N_48823);
or UO_4701 (O_4701,N_48658,N_48723);
nor UO_4702 (O_4702,N_49206,N_48880);
nand UO_4703 (O_4703,N_48739,N_49559);
nand UO_4704 (O_4704,N_48541,N_48835);
and UO_4705 (O_4705,N_49263,N_49339);
and UO_4706 (O_4706,N_48230,N_49646);
or UO_4707 (O_4707,N_49067,N_49426);
or UO_4708 (O_4708,N_48070,N_48822);
nand UO_4709 (O_4709,N_49489,N_49510);
or UO_4710 (O_4710,N_48463,N_49072);
or UO_4711 (O_4711,N_48423,N_48051);
nor UO_4712 (O_4712,N_49700,N_48798);
xnor UO_4713 (O_4713,N_49029,N_49730);
nor UO_4714 (O_4714,N_48507,N_48722);
and UO_4715 (O_4715,N_49989,N_48223);
nor UO_4716 (O_4716,N_49537,N_49698);
and UO_4717 (O_4717,N_49953,N_48651);
and UO_4718 (O_4718,N_48386,N_49337);
nor UO_4719 (O_4719,N_48604,N_48529);
and UO_4720 (O_4720,N_48432,N_49718);
or UO_4721 (O_4721,N_48984,N_48937);
and UO_4722 (O_4722,N_48849,N_49170);
or UO_4723 (O_4723,N_48876,N_49683);
xnor UO_4724 (O_4724,N_49057,N_48908);
or UO_4725 (O_4725,N_48792,N_48242);
nor UO_4726 (O_4726,N_48549,N_49694);
or UO_4727 (O_4727,N_49637,N_48614);
nor UO_4728 (O_4728,N_49970,N_49343);
nand UO_4729 (O_4729,N_49872,N_48702);
nand UO_4730 (O_4730,N_49271,N_49040);
or UO_4731 (O_4731,N_48440,N_48182);
or UO_4732 (O_4732,N_48408,N_48198);
nor UO_4733 (O_4733,N_49679,N_49709);
nor UO_4734 (O_4734,N_48330,N_48651);
nand UO_4735 (O_4735,N_48555,N_49290);
xnor UO_4736 (O_4736,N_48470,N_49565);
or UO_4737 (O_4737,N_48511,N_48756);
nand UO_4738 (O_4738,N_49719,N_49869);
and UO_4739 (O_4739,N_48696,N_48568);
nand UO_4740 (O_4740,N_48615,N_49139);
nor UO_4741 (O_4741,N_49442,N_49789);
nand UO_4742 (O_4742,N_48464,N_48108);
and UO_4743 (O_4743,N_49557,N_48667);
nand UO_4744 (O_4744,N_48027,N_48404);
nor UO_4745 (O_4745,N_49370,N_49771);
or UO_4746 (O_4746,N_49822,N_49141);
nor UO_4747 (O_4747,N_48041,N_48148);
or UO_4748 (O_4748,N_48659,N_48942);
and UO_4749 (O_4749,N_49547,N_48385);
nand UO_4750 (O_4750,N_49823,N_49529);
nor UO_4751 (O_4751,N_49238,N_49716);
nor UO_4752 (O_4752,N_49340,N_48502);
nor UO_4753 (O_4753,N_48179,N_48884);
nand UO_4754 (O_4754,N_48243,N_48322);
or UO_4755 (O_4755,N_48161,N_48180);
and UO_4756 (O_4756,N_49838,N_49070);
or UO_4757 (O_4757,N_49473,N_48010);
and UO_4758 (O_4758,N_49448,N_48027);
nand UO_4759 (O_4759,N_48366,N_48600);
nor UO_4760 (O_4760,N_49913,N_49291);
nor UO_4761 (O_4761,N_49122,N_49292);
nand UO_4762 (O_4762,N_48315,N_49709);
nor UO_4763 (O_4763,N_49893,N_48987);
nand UO_4764 (O_4764,N_48538,N_48333);
nor UO_4765 (O_4765,N_49113,N_48410);
and UO_4766 (O_4766,N_49287,N_49404);
nand UO_4767 (O_4767,N_48399,N_48655);
nor UO_4768 (O_4768,N_49456,N_49425);
nand UO_4769 (O_4769,N_48140,N_49881);
nor UO_4770 (O_4770,N_49486,N_48361);
and UO_4771 (O_4771,N_49432,N_49077);
and UO_4772 (O_4772,N_49357,N_49942);
and UO_4773 (O_4773,N_49194,N_49340);
nand UO_4774 (O_4774,N_48547,N_49496);
nand UO_4775 (O_4775,N_48646,N_49113);
or UO_4776 (O_4776,N_49480,N_48204);
and UO_4777 (O_4777,N_48985,N_49865);
and UO_4778 (O_4778,N_49431,N_49015);
nand UO_4779 (O_4779,N_49188,N_48870);
nor UO_4780 (O_4780,N_49342,N_49365);
or UO_4781 (O_4781,N_49060,N_49956);
and UO_4782 (O_4782,N_48473,N_48403);
nand UO_4783 (O_4783,N_48941,N_48880);
nand UO_4784 (O_4784,N_48279,N_49596);
nand UO_4785 (O_4785,N_48017,N_49209);
or UO_4786 (O_4786,N_49937,N_49609);
or UO_4787 (O_4787,N_48354,N_48261);
and UO_4788 (O_4788,N_48025,N_48787);
nor UO_4789 (O_4789,N_48167,N_49860);
and UO_4790 (O_4790,N_48276,N_49832);
nor UO_4791 (O_4791,N_48873,N_49398);
and UO_4792 (O_4792,N_49458,N_49968);
nand UO_4793 (O_4793,N_49656,N_48483);
and UO_4794 (O_4794,N_48341,N_49894);
nor UO_4795 (O_4795,N_49181,N_48357);
nor UO_4796 (O_4796,N_48940,N_48149);
or UO_4797 (O_4797,N_49692,N_49819);
and UO_4798 (O_4798,N_49582,N_48792);
nor UO_4799 (O_4799,N_48840,N_48206);
or UO_4800 (O_4800,N_49768,N_49566);
nand UO_4801 (O_4801,N_49760,N_49884);
or UO_4802 (O_4802,N_49383,N_49861);
or UO_4803 (O_4803,N_48776,N_49733);
and UO_4804 (O_4804,N_49582,N_48287);
or UO_4805 (O_4805,N_49818,N_48076);
nor UO_4806 (O_4806,N_48654,N_48288);
and UO_4807 (O_4807,N_48846,N_49186);
and UO_4808 (O_4808,N_48272,N_48123);
nand UO_4809 (O_4809,N_48860,N_48419);
nor UO_4810 (O_4810,N_49850,N_48604);
nor UO_4811 (O_4811,N_48683,N_49328);
and UO_4812 (O_4812,N_48477,N_49670);
nand UO_4813 (O_4813,N_49889,N_49776);
or UO_4814 (O_4814,N_49614,N_48999);
nand UO_4815 (O_4815,N_48974,N_49362);
and UO_4816 (O_4816,N_48768,N_49241);
nand UO_4817 (O_4817,N_49662,N_48885);
nor UO_4818 (O_4818,N_49416,N_48388);
nand UO_4819 (O_4819,N_49477,N_49844);
or UO_4820 (O_4820,N_48277,N_48597);
and UO_4821 (O_4821,N_48254,N_49211);
nor UO_4822 (O_4822,N_48732,N_48379);
nand UO_4823 (O_4823,N_48293,N_48636);
or UO_4824 (O_4824,N_48140,N_49650);
or UO_4825 (O_4825,N_48242,N_48892);
nand UO_4826 (O_4826,N_49904,N_49309);
nor UO_4827 (O_4827,N_49252,N_49778);
nor UO_4828 (O_4828,N_48873,N_48978);
and UO_4829 (O_4829,N_49776,N_48564);
nand UO_4830 (O_4830,N_48463,N_49751);
and UO_4831 (O_4831,N_48299,N_48737);
and UO_4832 (O_4832,N_48519,N_49173);
or UO_4833 (O_4833,N_48721,N_49173);
nor UO_4834 (O_4834,N_49583,N_49179);
and UO_4835 (O_4835,N_49165,N_48077);
and UO_4836 (O_4836,N_49297,N_48391);
and UO_4837 (O_4837,N_49611,N_48303);
or UO_4838 (O_4838,N_49426,N_48867);
nand UO_4839 (O_4839,N_49312,N_49675);
or UO_4840 (O_4840,N_48722,N_49495);
and UO_4841 (O_4841,N_48739,N_48030);
nor UO_4842 (O_4842,N_48725,N_48257);
nand UO_4843 (O_4843,N_48167,N_48719);
and UO_4844 (O_4844,N_49788,N_48362);
or UO_4845 (O_4845,N_49145,N_49033);
nand UO_4846 (O_4846,N_49271,N_49943);
nor UO_4847 (O_4847,N_49276,N_48204);
or UO_4848 (O_4848,N_48934,N_49263);
and UO_4849 (O_4849,N_48570,N_49606);
nor UO_4850 (O_4850,N_49453,N_48455);
and UO_4851 (O_4851,N_49388,N_49355);
and UO_4852 (O_4852,N_49844,N_48350);
nor UO_4853 (O_4853,N_48955,N_48095);
and UO_4854 (O_4854,N_49358,N_49610);
and UO_4855 (O_4855,N_49787,N_49794);
nor UO_4856 (O_4856,N_49515,N_48425);
nor UO_4857 (O_4857,N_48499,N_49214);
nor UO_4858 (O_4858,N_49779,N_49252);
nor UO_4859 (O_4859,N_48954,N_49609);
nand UO_4860 (O_4860,N_48459,N_49783);
or UO_4861 (O_4861,N_49785,N_49715);
nand UO_4862 (O_4862,N_48451,N_49388);
or UO_4863 (O_4863,N_49780,N_49250);
or UO_4864 (O_4864,N_49730,N_49567);
nor UO_4865 (O_4865,N_49831,N_48687);
nor UO_4866 (O_4866,N_49634,N_48861);
or UO_4867 (O_4867,N_49828,N_48196);
nand UO_4868 (O_4868,N_48002,N_49632);
nor UO_4869 (O_4869,N_49476,N_49234);
nor UO_4870 (O_4870,N_49757,N_48874);
or UO_4871 (O_4871,N_48967,N_48080);
nand UO_4872 (O_4872,N_48205,N_49794);
and UO_4873 (O_4873,N_48023,N_49608);
nor UO_4874 (O_4874,N_49020,N_49037);
nor UO_4875 (O_4875,N_48005,N_49786);
nand UO_4876 (O_4876,N_49245,N_49179);
nand UO_4877 (O_4877,N_49780,N_48925);
nand UO_4878 (O_4878,N_49528,N_48226);
and UO_4879 (O_4879,N_48086,N_48511);
nand UO_4880 (O_4880,N_48013,N_49232);
nor UO_4881 (O_4881,N_49663,N_48728);
nand UO_4882 (O_4882,N_49140,N_49358);
nor UO_4883 (O_4883,N_48872,N_48593);
nand UO_4884 (O_4884,N_49819,N_49471);
nand UO_4885 (O_4885,N_49134,N_48730);
or UO_4886 (O_4886,N_48131,N_49854);
nand UO_4887 (O_4887,N_49548,N_48886);
nor UO_4888 (O_4888,N_49527,N_48608);
nand UO_4889 (O_4889,N_49288,N_48241);
nand UO_4890 (O_4890,N_49083,N_49734);
or UO_4891 (O_4891,N_49304,N_48076);
nor UO_4892 (O_4892,N_48778,N_49241);
nor UO_4893 (O_4893,N_48944,N_48565);
and UO_4894 (O_4894,N_49979,N_49437);
and UO_4895 (O_4895,N_48752,N_49452);
nand UO_4896 (O_4896,N_48962,N_49828);
nand UO_4897 (O_4897,N_49149,N_49190);
and UO_4898 (O_4898,N_48598,N_49238);
nor UO_4899 (O_4899,N_49572,N_49719);
nor UO_4900 (O_4900,N_49231,N_49050);
and UO_4901 (O_4901,N_49537,N_49904);
xnor UO_4902 (O_4902,N_48880,N_48644);
nor UO_4903 (O_4903,N_49499,N_48614);
or UO_4904 (O_4904,N_49114,N_48410);
and UO_4905 (O_4905,N_48758,N_48158);
and UO_4906 (O_4906,N_48497,N_49051);
nor UO_4907 (O_4907,N_48176,N_48177);
and UO_4908 (O_4908,N_49496,N_48382);
or UO_4909 (O_4909,N_48096,N_49549);
and UO_4910 (O_4910,N_48166,N_49892);
or UO_4911 (O_4911,N_48334,N_49421);
or UO_4912 (O_4912,N_49893,N_48142);
nor UO_4913 (O_4913,N_49092,N_49746);
and UO_4914 (O_4914,N_49754,N_49906);
nand UO_4915 (O_4915,N_48446,N_48431);
and UO_4916 (O_4916,N_48501,N_49832);
or UO_4917 (O_4917,N_48716,N_48386);
nand UO_4918 (O_4918,N_49491,N_48602);
and UO_4919 (O_4919,N_48716,N_48552);
nor UO_4920 (O_4920,N_48269,N_49695);
nor UO_4921 (O_4921,N_48273,N_48252);
nand UO_4922 (O_4922,N_48289,N_49381);
nand UO_4923 (O_4923,N_48531,N_49623);
nand UO_4924 (O_4924,N_48963,N_48460);
nor UO_4925 (O_4925,N_49511,N_49121);
nor UO_4926 (O_4926,N_48308,N_48060);
or UO_4927 (O_4927,N_49476,N_49815);
nand UO_4928 (O_4928,N_49794,N_49599);
nand UO_4929 (O_4929,N_49808,N_48519);
and UO_4930 (O_4930,N_48285,N_48859);
nand UO_4931 (O_4931,N_48992,N_49367);
xnor UO_4932 (O_4932,N_48124,N_48587);
nor UO_4933 (O_4933,N_48633,N_49919);
or UO_4934 (O_4934,N_49716,N_49512);
and UO_4935 (O_4935,N_48225,N_48003);
nor UO_4936 (O_4936,N_49096,N_49775);
nor UO_4937 (O_4937,N_49157,N_49898);
and UO_4938 (O_4938,N_49684,N_48590);
nand UO_4939 (O_4939,N_48359,N_48690);
or UO_4940 (O_4940,N_49511,N_49032);
and UO_4941 (O_4941,N_48509,N_49832);
or UO_4942 (O_4942,N_48094,N_49781);
and UO_4943 (O_4943,N_49182,N_49431);
xnor UO_4944 (O_4944,N_49930,N_49559);
or UO_4945 (O_4945,N_48920,N_49075);
and UO_4946 (O_4946,N_49202,N_49110);
and UO_4947 (O_4947,N_48384,N_49584);
and UO_4948 (O_4948,N_49727,N_49953);
or UO_4949 (O_4949,N_48367,N_49043);
or UO_4950 (O_4950,N_48992,N_48327);
nand UO_4951 (O_4951,N_49568,N_49492);
and UO_4952 (O_4952,N_48433,N_49828);
nor UO_4953 (O_4953,N_48021,N_48697);
or UO_4954 (O_4954,N_49361,N_49320);
and UO_4955 (O_4955,N_48659,N_48432);
and UO_4956 (O_4956,N_49836,N_48211);
nor UO_4957 (O_4957,N_48250,N_49526);
or UO_4958 (O_4958,N_49614,N_48480);
and UO_4959 (O_4959,N_48178,N_48257);
nand UO_4960 (O_4960,N_48619,N_48413);
or UO_4961 (O_4961,N_49318,N_48730);
or UO_4962 (O_4962,N_48926,N_49299);
or UO_4963 (O_4963,N_48940,N_48604);
nand UO_4964 (O_4964,N_48708,N_49660);
nor UO_4965 (O_4965,N_48956,N_49122);
or UO_4966 (O_4966,N_48198,N_48929);
xnor UO_4967 (O_4967,N_49304,N_48447);
nor UO_4968 (O_4968,N_48689,N_49008);
nor UO_4969 (O_4969,N_48207,N_49284);
nand UO_4970 (O_4970,N_48907,N_49637);
and UO_4971 (O_4971,N_48239,N_49660);
nor UO_4972 (O_4972,N_48434,N_49335);
and UO_4973 (O_4973,N_49027,N_48688);
nand UO_4974 (O_4974,N_49644,N_49179);
and UO_4975 (O_4975,N_48216,N_48994);
or UO_4976 (O_4976,N_49688,N_48785);
nand UO_4977 (O_4977,N_49364,N_48173);
nor UO_4978 (O_4978,N_49195,N_48108);
and UO_4979 (O_4979,N_49962,N_49094);
and UO_4980 (O_4980,N_48695,N_49899);
nand UO_4981 (O_4981,N_48758,N_48635);
nor UO_4982 (O_4982,N_48420,N_49369);
nor UO_4983 (O_4983,N_48955,N_49414);
or UO_4984 (O_4984,N_49123,N_48860);
nand UO_4985 (O_4985,N_49433,N_48820);
or UO_4986 (O_4986,N_49198,N_49667);
and UO_4987 (O_4987,N_49113,N_49034);
and UO_4988 (O_4988,N_49329,N_49198);
nor UO_4989 (O_4989,N_49084,N_48473);
or UO_4990 (O_4990,N_49400,N_49498);
nand UO_4991 (O_4991,N_49847,N_49700);
nor UO_4992 (O_4992,N_48062,N_49568);
nor UO_4993 (O_4993,N_48953,N_49819);
xnor UO_4994 (O_4994,N_49582,N_49693);
or UO_4995 (O_4995,N_49702,N_48465);
or UO_4996 (O_4996,N_49517,N_48543);
and UO_4997 (O_4997,N_48613,N_48014);
nand UO_4998 (O_4998,N_48484,N_48316);
nor UO_4999 (O_4999,N_48189,N_48704);
endmodule