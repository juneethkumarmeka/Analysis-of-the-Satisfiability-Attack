module basic_1000_10000_1500_10_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_421,In_471);
or U1 (N_1,In_279,In_142);
or U2 (N_2,In_633,In_475);
and U3 (N_3,In_379,In_606);
xor U4 (N_4,In_392,In_349);
and U5 (N_5,In_191,In_99);
or U6 (N_6,In_424,In_187);
xor U7 (N_7,In_954,In_505);
or U8 (N_8,In_667,In_709);
and U9 (N_9,In_708,In_931);
or U10 (N_10,In_464,In_453);
and U11 (N_11,In_998,In_530);
and U12 (N_12,In_696,In_79);
or U13 (N_13,In_964,In_718);
or U14 (N_14,In_157,In_582);
and U15 (N_15,In_200,In_752);
nand U16 (N_16,In_12,In_771);
and U17 (N_17,In_875,In_972);
or U18 (N_18,In_827,In_647);
or U19 (N_19,In_252,In_271);
and U20 (N_20,In_975,In_436);
nand U21 (N_21,In_49,In_994);
nand U22 (N_22,In_591,In_60);
nor U23 (N_23,In_676,In_618);
nor U24 (N_24,In_461,In_634);
nand U25 (N_25,In_761,In_323);
nor U26 (N_26,In_171,In_312);
nand U27 (N_27,In_319,In_820);
and U28 (N_28,In_892,In_380);
nand U29 (N_29,In_8,In_318);
nor U30 (N_30,In_898,In_432);
nor U31 (N_31,In_384,In_899);
or U32 (N_32,In_679,In_258);
or U33 (N_33,In_427,In_304);
nor U34 (N_34,In_592,In_517);
or U35 (N_35,In_443,In_145);
nand U36 (N_36,In_388,In_241);
nor U37 (N_37,In_498,In_366);
and U38 (N_38,In_948,In_814);
and U39 (N_39,In_439,In_22);
and U40 (N_40,In_617,In_91);
or U41 (N_41,In_212,In_872);
and U42 (N_42,In_149,In_494);
and U43 (N_43,In_455,In_558);
nor U44 (N_44,In_857,In_999);
nor U45 (N_45,In_393,In_952);
nand U46 (N_46,In_37,In_275);
or U47 (N_47,In_514,In_0);
or U48 (N_48,In_425,In_57);
and U49 (N_49,In_949,In_929);
nor U50 (N_50,In_309,In_557);
and U51 (N_51,In_819,In_614);
nand U52 (N_52,In_886,In_354);
nand U53 (N_53,In_501,In_404);
nand U54 (N_54,In_325,In_563);
nor U55 (N_55,In_382,In_732);
nor U56 (N_56,In_358,In_347);
nor U57 (N_57,In_877,In_273);
or U58 (N_58,In_903,In_835);
nand U59 (N_59,In_504,In_214);
or U60 (N_60,In_155,In_265);
nor U61 (N_61,In_56,In_226);
nor U62 (N_62,In_654,In_598);
nor U63 (N_63,In_109,In_509);
nor U64 (N_64,In_562,In_518);
or U65 (N_65,In_719,In_564);
and U66 (N_66,In_763,In_102);
or U67 (N_67,In_81,In_694);
and U68 (N_68,In_525,In_869);
nand U69 (N_69,In_210,In_127);
or U70 (N_70,In_734,In_181);
nand U71 (N_71,In_327,In_589);
or U72 (N_72,In_405,In_477);
and U73 (N_73,In_105,In_45);
and U74 (N_74,In_278,In_905);
nand U75 (N_75,In_277,In_217);
and U76 (N_76,In_925,In_174);
and U77 (N_77,In_411,In_78);
nor U78 (N_78,In_153,In_300);
nand U79 (N_79,In_507,In_788);
nand U80 (N_80,In_288,In_516);
or U81 (N_81,In_396,In_729);
and U82 (N_82,In_726,In_996);
or U83 (N_83,In_860,In_699);
nor U84 (N_84,In_790,In_14);
nand U85 (N_85,In_840,In_923);
or U86 (N_86,In_772,In_355);
and U87 (N_87,In_635,In_986);
nand U88 (N_88,In_283,In_714);
nor U89 (N_89,In_307,In_337);
and U90 (N_90,In_574,In_64);
and U91 (N_91,In_743,In_576);
nor U92 (N_92,In_966,In_561);
or U93 (N_93,In_566,In_549);
or U94 (N_94,In_813,In_104);
nand U95 (N_95,In_13,In_551);
or U96 (N_96,In_737,In_39);
and U97 (N_97,In_403,In_496);
or U98 (N_98,In_433,In_850);
and U99 (N_99,In_976,In_141);
nor U100 (N_100,In_243,In_34);
nor U101 (N_101,In_410,In_851);
nor U102 (N_102,In_855,In_467);
xnor U103 (N_103,In_513,In_926);
nor U104 (N_104,In_920,In_764);
and U105 (N_105,In_208,In_622);
and U106 (N_106,In_276,In_867);
nand U107 (N_107,In_150,In_779);
nor U108 (N_108,In_386,In_299);
and U109 (N_109,In_417,In_987);
or U110 (N_110,In_267,In_639);
nor U111 (N_111,In_579,In_538);
nand U112 (N_112,In_569,In_871);
xor U113 (N_113,In_612,In_712);
or U114 (N_114,In_293,In_281);
nand U115 (N_115,In_967,In_470);
nor U116 (N_116,In_428,In_520);
nand U117 (N_117,In_342,In_984);
nand U118 (N_118,In_842,In_286);
and U119 (N_119,In_703,In_673);
nand U120 (N_120,In_691,In_817);
nor U121 (N_121,In_919,In_824);
or U122 (N_122,In_655,In_810);
nor U123 (N_123,In_503,In_768);
or U124 (N_124,In_641,In_414);
nor U125 (N_125,In_27,In_314);
nor U126 (N_126,In_995,In_130);
nor U127 (N_127,In_936,In_448);
nor U128 (N_128,In_462,In_648);
xor U129 (N_129,In_154,In_701);
and U130 (N_130,In_492,In_236);
or U131 (N_131,In_692,In_683);
and U132 (N_132,In_610,In_222);
or U133 (N_133,In_483,In_339);
or U134 (N_134,In_77,In_670);
or U135 (N_135,In_733,In_990);
nor U136 (N_136,In_962,In_693);
nor U137 (N_137,In_391,In_945);
nand U138 (N_138,In_435,In_515);
nor U139 (N_139,In_854,In_266);
and U140 (N_140,In_922,In_572);
or U141 (N_141,In_251,In_874);
nand U142 (N_142,In_913,In_653);
and U143 (N_143,In_660,In_666);
and U144 (N_144,In_5,In_237);
and U145 (N_145,In_893,In_837);
xor U146 (N_146,In_158,In_284);
nand U147 (N_147,In_6,In_782);
and U148 (N_148,In_548,In_166);
and U149 (N_149,In_628,In_108);
or U150 (N_150,In_303,In_664);
xor U151 (N_151,In_578,In_184);
nand U152 (N_152,In_583,In_4);
nor U153 (N_153,In_651,In_378);
and U154 (N_154,In_727,In_754);
nor U155 (N_155,In_451,In_649);
nand U156 (N_156,In_374,In_787);
nor U157 (N_157,In_642,In_545);
nand U158 (N_158,In_121,In_400);
xor U159 (N_159,In_637,In_848);
and U160 (N_160,In_242,In_740);
nand U161 (N_161,In_480,In_211);
nand U162 (N_162,In_92,In_491);
and U163 (N_163,In_459,In_983);
nand U164 (N_164,In_844,In_554);
and U165 (N_165,In_678,In_390);
nand U166 (N_166,In_107,In_904);
and U167 (N_167,In_381,In_112);
nand U168 (N_168,In_136,In_981);
xnor U169 (N_169,In_408,In_24);
nor U170 (N_170,In_113,In_257);
nand U171 (N_171,In_434,In_484);
or U172 (N_172,In_725,In_625);
and U173 (N_173,In_399,In_430);
and U174 (N_174,In_807,In_993);
or U175 (N_175,In_82,In_129);
nor U176 (N_176,In_956,In_262);
nor U177 (N_177,In_270,In_873);
nand U178 (N_178,In_769,In_26);
or U179 (N_179,In_9,In_608);
or U180 (N_180,In_3,In_254);
or U181 (N_181,In_47,In_826);
nor U182 (N_182,In_440,In_974);
nand U183 (N_183,In_539,In_600);
and U184 (N_184,In_613,In_61);
or U185 (N_185,In_684,In_225);
nor U186 (N_186,In_593,In_23);
or U187 (N_187,In_992,In_881);
and U188 (N_188,In_846,In_602);
or U189 (N_189,In_555,In_44);
nand U190 (N_190,In_720,In_746);
nor U191 (N_191,In_802,In_192);
nand U192 (N_192,In_700,In_728);
and U193 (N_193,In_889,In_415);
or U194 (N_194,In_117,In_10);
and U195 (N_195,In_294,In_918);
and U196 (N_196,In_785,In_409);
and U197 (N_197,In_295,In_134);
nand U198 (N_198,In_19,In_182);
nand U199 (N_199,In_175,In_84);
and U200 (N_200,In_88,In_698);
nand U201 (N_201,In_958,In_937);
or U202 (N_202,In_989,In_685);
nand U203 (N_203,In_41,In_316);
and U204 (N_204,In_54,In_33);
nand U205 (N_205,In_512,In_624);
nand U206 (N_206,In_706,In_97);
or U207 (N_207,In_103,In_710);
and U208 (N_208,In_702,In_83);
or U209 (N_209,In_80,In_759);
and U210 (N_210,In_959,In_152);
and U211 (N_211,In_841,In_407);
nand U212 (N_212,In_261,In_385);
and U213 (N_213,In_422,In_148);
and U214 (N_214,In_206,In_970);
and U215 (N_215,In_343,In_452);
nor U216 (N_216,In_586,In_196);
nor U217 (N_217,In_527,In_997);
and U218 (N_218,In_526,In_308);
and U219 (N_219,In_124,In_739);
nor U220 (N_220,In_784,In_264);
nor U221 (N_221,In_370,In_674);
and U222 (N_222,In_645,In_528);
and U223 (N_223,In_32,In_575);
and U224 (N_224,In_292,In_297);
and U225 (N_225,In_173,In_863);
and U226 (N_226,In_968,In_845);
or U227 (N_227,In_28,In_159);
xor U228 (N_228,In_868,In_495);
nand U229 (N_229,In_547,In_511);
and U230 (N_230,In_951,In_162);
or U231 (N_231,In_268,In_786);
nor U232 (N_232,In_862,In_114);
xnor U233 (N_233,In_71,In_991);
nor U234 (N_234,In_603,In_172);
nand U235 (N_235,In_963,In_798);
and U236 (N_236,In_357,In_531);
or U237 (N_237,In_128,In_256);
nor U238 (N_238,In_38,In_194);
nand U239 (N_239,In_481,In_53);
or U240 (N_240,In_878,In_541);
nor U241 (N_241,In_429,In_506);
and U242 (N_242,In_140,In_177);
nor U243 (N_243,In_466,In_67);
and U244 (N_244,In_794,In_935);
nor U245 (N_245,In_359,In_486);
nand U246 (N_246,In_247,In_816);
nand U247 (N_247,In_132,In_915);
and U248 (N_248,In_960,In_879);
and U249 (N_249,In_675,In_147);
and U250 (N_250,In_260,In_59);
or U251 (N_251,In_943,In_218);
nand U252 (N_252,In_442,In_63);
and U253 (N_253,In_890,In_285);
xor U254 (N_254,In_444,In_536);
and U255 (N_255,In_738,In_317);
nor U256 (N_256,In_490,In_465);
and U257 (N_257,In_885,In_950);
and U258 (N_258,In_809,In_800);
nand U259 (N_259,In_336,In_902);
nor U260 (N_260,In_601,In_197);
and U261 (N_261,In_735,In_185);
or U262 (N_262,In_362,In_361);
xnor U263 (N_263,In_111,In_135);
nand U264 (N_264,In_2,In_830);
nand U265 (N_265,In_646,In_398);
and U266 (N_266,In_86,In_626);
and U267 (N_267,In_305,In_401);
nor U268 (N_268,In_681,In_30);
and U269 (N_269,In_927,In_487);
and U270 (N_270,In_352,In_544);
and U271 (N_271,In_240,In_219);
or U272 (N_272,In_156,In_521);
nand U273 (N_273,In_532,In_630);
or U274 (N_274,In_395,In_818);
and U275 (N_275,In_472,In_246);
or U276 (N_276,In_632,In_324);
and U277 (N_277,In_20,In_372);
nor U278 (N_278,In_456,In_650);
and U279 (N_279,In_668,In_540);
and U280 (N_280,In_62,In_493);
and U281 (N_281,In_238,In_722);
and U282 (N_282,In_638,In_988);
nand U283 (N_283,In_447,In_231);
or U284 (N_284,In_631,In_94);
nand U285 (N_285,In_468,In_944);
nand U286 (N_286,In_368,In_289);
or U287 (N_287,In_912,In_757);
and U288 (N_288,In_619,In_330);
nand U289 (N_289,In_812,In_916);
nor U290 (N_290,In_640,In_463);
or U291 (N_291,In_940,In_406);
nor U292 (N_292,In_235,In_657);
nor U293 (N_293,In_263,In_418);
nand U294 (N_294,In_365,In_957);
nor U295 (N_295,In_143,In_793);
nand U296 (N_296,In_856,In_865);
nor U297 (N_297,In_350,In_914);
nand U298 (N_298,In_315,In_93);
or U299 (N_299,In_707,In_985);
nor U300 (N_300,In_351,In_338);
nor U301 (N_301,In_165,In_804);
or U302 (N_302,In_901,In_203);
and U303 (N_303,In_377,In_170);
or U304 (N_304,In_423,In_239);
or U305 (N_305,In_228,In_120);
and U306 (N_306,In_721,In_609);
or U307 (N_307,In_715,In_806);
xnor U308 (N_308,In_230,In_450);
nand U309 (N_309,In_965,In_560);
and U310 (N_310,In_753,In_705);
or U311 (N_311,In_412,In_133);
nor U312 (N_312,In_119,In_449);
nor U313 (N_313,In_607,In_774);
and U314 (N_314,In_934,In_758);
nor U315 (N_315,In_616,In_190);
nor U316 (N_316,In_933,In_596);
and U317 (N_317,In_783,In_580);
and U318 (N_318,In_95,In_473);
and U319 (N_319,In_125,In_205);
and U320 (N_320,In_831,In_280);
or U321 (N_321,In_98,In_438);
nor U322 (N_322,In_864,In_302);
nor U323 (N_323,In_777,In_402);
nand U324 (N_324,In_776,In_595);
and U325 (N_325,In_924,In_478);
and U326 (N_326,In_322,In_792);
nand U327 (N_327,In_216,In_887);
and U328 (N_328,In_751,In_144);
or U329 (N_329,In_745,In_204);
nor U330 (N_330,In_310,In_65);
xnor U331 (N_331,In_978,In_849);
nor U332 (N_332,In_106,In_195);
nand U333 (N_333,In_55,In_233);
nor U334 (N_334,In_202,In_479);
nand U335 (N_335,In_89,In_224);
or U336 (N_336,In_559,In_568);
nor U337 (N_337,In_389,In_394);
or U338 (N_338,In_454,In_604);
nand U339 (N_339,In_229,In_234);
and U340 (N_340,In_510,In_223);
nand U341 (N_341,In_870,In_522);
xor U342 (N_342,In_852,In_48);
nand U343 (N_343,In_193,In_894);
nor U344 (N_344,In_340,In_533);
or U345 (N_345,In_335,In_419);
or U346 (N_346,In_320,In_942);
nand U347 (N_347,In_791,In_847);
nand U348 (N_348,In_115,In_326);
and U349 (N_349,In_489,In_888);
and U350 (N_350,In_420,In_90);
or U351 (N_351,In_373,In_571);
xnor U352 (N_352,In_884,In_543);
and U353 (N_353,In_573,In_762);
xnor U354 (N_354,In_755,In_704);
nand U355 (N_355,In_973,In_137);
nand U356 (N_356,In_68,In_534);
nand U357 (N_357,In_749,In_348);
or U358 (N_358,In_979,In_163);
and U359 (N_359,In_446,In_717);
or U360 (N_360,In_311,In_662);
and U361 (N_361,In_524,In_587);
nand U362 (N_362,In_244,In_167);
nand U363 (N_363,In_383,In_553);
nor U364 (N_364,In_680,In_584);
nor U365 (N_365,In_31,In_766);
or U366 (N_366,In_169,In_87);
nand U367 (N_367,In_535,In_883);
nor U368 (N_368,In_151,In_866);
nand U369 (N_369,In_25,In_341);
nand U370 (N_370,In_1,In_801);
and U371 (N_371,In_938,In_756);
nor U372 (N_372,In_74,In_485);
nand U373 (N_373,In_101,In_35);
and U374 (N_374,In_209,In_72);
and U375 (N_375,In_76,In_66);
or U376 (N_376,In_828,In_669);
nand U377 (N_377,In_360,In_656);
or U378 (N_378,In_861,In_227);
and U379 (N_379,In_274,In_760);
and U380 (N_380,In_565,In_376);
or U381 (N_381,In_808,In_689);
and U382 (N_382,In_953,In_253);
and U383 (N_383,In_843,In_895);
and U384 (N_384,In_971,In_821);
or U385 (N_385,In_930,In_96);
and U386 (N_386,In_682,In_482);
and U387 (N_387,In_773,In_838);
nor U388 (N_388,In_296,In_353);
or U389 (N_389,In_900,In_550);
and U390 (N_390,In_795,In_387);
or U391 (N_391,In_75,In_588);
nand U392 (N_392,In_859,In_825);
nor U393 (N_393,In_908,In_146);
xnor U394 (N_394,In_687,In_939);
nor U395 (N_395,In_906,In_476);
or U396 (N_396,In_179,In_329);
nand U397 (N_397,In_441,In_546);
nor U398 (N_398,In_741,In_43);
and U399 (N_399,In_724,In_331);
and U400 (N_400,In_711,In_597);
nand U401 (N_401,In_747,In_803);
and U402 (N_402,In_176,In_138);
or U403 (N_403,In_85,In_909);
and U404 (N_404,In_858,In_652);
and U405 (N_405,In_697,In_36);
nand U406 (N_406,In_805,In_189);
or U407 (N_407,In_921,In_585);
and U408 (N_408,In_291,In_232);
nand U409 (N_409,In_977,In_928);
and U410 (N_410,In_11,In_917);
nor U411 (N_411,In_627,In_853);
and U412 (N_412,In_397,In_269);
nor U413 (N_413,In_876,In_42);
nor U414 (N_414,In_832,In_413);
and U415 (N_415,In_488,In_199);
or U416 (N_416,In_896,In_164);
nand U417 (N_417,In_426,In_58);
or U418 (N_418,In_474,In_248);
xor U419 (N_419,In_69,In_122);
nand U420 (N_420,In_567,In_690);
or U421 (N_421,In_213,In_183);
and U422 (N_422,In_552,In_781);
nor U423 (N_423,In_911,In_100);
nor U424 (N_424,In_332,In_537);
nor U425 (N_425,In_829,In_178);
nand U426 (N_426,In_910,In_519);
or U427 (N_427,In_730,In_52);
nand U428 (N_428,In_502,In_364);
and U429 (N_429,In_542,In_731);
nand U430 (N_430,In_523,In_961);
or U431 (N_431,In_416,In_123);
nor U432 (N_432,In_529,In_298);
nor U433 (N_433,In_797,In_767);
nor U434 (N_434,In_605,In_198);
and U435 (N_435,In_29,In_328);
nor U436 (N_436,In_369,In_775);
nand U437 (N_437,In_367,In_445);
xor U438 (N_438,In_671,In_833);
nor U439 (N_439,In_659,In_880);
and U440 (N_440,In_834,In_180);
xnor U441 (N_441,In_118,In_126);
and U442 (N_442,In_139,In_131);
nor U443 (N_443,In_723,In_643);
or U444 (N_444,In_161,In_250);
and U445 (N_445,In_932,In_629);
nor U446 (N_446,In_290,In_882);
or U447 (N_447,In_437,In_255);
nand U448 (N_448,In_16,In_375);
and U449 (N_449,In_168,In_306);
nand U450 (N_450,In_644,In_249);
nor U451 (N_451,In_70,In_508);
nand U452 (N_452,In_811,In_946);
nand U453 (N_453,In_982,In_658);
nand U454 (N_454,In_891,In_695);
nor U455 (N_455,In_259,In_941);
nand U456 (N_456,In_663,In_713);
and U457 (N_457,In_497,In_313);
and U458 (N_458,In_577,In_599);
or U459 (N_459,In_796,In_21);
and U460 (N_460,In_50,In_371);
and U461 (N_461,In_748,In_980);
nor U462 (N_462,In_73,In_188);
and U463 (N_463,In_346,In_661);
nor U464 (N_464,In_686,In_18);
nand U465 (N_465,In_839,In_815);
and U466 (N_466,In_556,In_590);
nand U467 (N_467,In_363,In_40);
nor U468 (N_468,In_907,In_7);
and U469 (N_469,In_611,In_51);
and U470 (N_470,In_160,In_744);
nand U471 (N_471,In_822,In_799);
nand U472 (N_472,In_594,In_688);
or U473 (N_473,In_969,In_301);
or U474 (N_474,In_615,In_186);
nand U475 (N_475,In_344,In_469);
nand U476 (N_476,In_742,In_823);
and U477 (N_477,In_620,In_457);
nor U478 (N_478,In_623,In_220);
and U479 (N_479,In_778,In_716);
nand U480 (N_480,In_272,In_207);
nand U481 (N_481,In_46,In_110);
and U482 (N_482,In_345,In_581);
or U483 (N_483,In_897,In_215);
nand U484 (N_484,In_500,In_955);
xnor U485 (N_485,In_947,In_672);
and U486 (N_486,In_334,In_621);
nor U487 (N_487,In_836,In_333);
and U488 (N_488,In_770,In_789);
nor U489 (N_489,In_201,In_17);
and U490 (N_490,In_570,In_665);
nor U491 (N_491,In_499,In_282);
nand U492 (N_492,In_458,In_750);
nor U493 (N_493,In_780,In_356);
nor U494 (N_494,In_431,In_221);
and U495 (N_495,In_287,In_245);
and U496 (N_496,In_321,In_765);
or U497 (N_497,In_736,In_677);
and U498 (N_498,In_460,In_15);
and U499 (N_499,In_116,In_636);
nand U500 (N_500,In_480,In_579);
and U501 (N_501,In_683,In_163);
nand U502 (N_502,In_520,In_795);
and U503 (N_503,In_639,In_608);
or U504 (N_504,In_263,In_502);
and U505 (N_505,In_556,In_13);
nor U506 (N_506,In_197,In_904);
and U507 (N_507,In_476,In_307);
nor U508 (N_508,In_167,In_320);
nand U509 (N_509,In_127,In_444);
nor U510 (N_510,In_348,In_752);
nand U511 (N_511,In_690,In_14);
or U512 (N_512,In_461,In_860);
or U513 (N_513,In_425,In_98);
or U514 (N_514,In_39,In_614);
nor U515 (N_515,In_977,In_853);
and U516 (N_516,In_171,In_349);
or U517 (N_517,In_866,In_973);
nor U518 (N_518,In_894,In_636);
and U519 (N_519,In_586,In_216);
nor U520 (N_520,In_760,In_895);
and U521 (N_521,In_966,In_673);
or U522 (N_522,In_505,In_806);
nand U523 (N_523,In_837,In_187);
and U524 (N_524,In_897,In_579);
and U525 (N_525,In_669,In_484);
and U526 (N_526,In_405,In_901);
and U527 (N_527,In_69,In_374);
and U528 (N_528,In_738,In_774);
nand U529 (N_529,In_177,In_616);
and U530 (N_530,In_661,In_815);
or U531 (N_531,In_357,In_402);
and U532 (N_532,In_855,In_867);
and U533 (N_533,In_473,In_579);
nor U534 (N_534,In_85,In_984);
nand U535 (N_535,In_370,In_967);
nor U536 (N_536,In_258,In_714);
nand U537 (N_537,In_255,In_337);
or U538 (N_538,In_154,In_663);
and U539 (N_539,In_131,In_432);
nor U540 (N_540,In_45,In_385);
nor U541 (N_541,In_985,In_714);
and U542 (N_542,In_329,In_11);
and U543 (N_543,In_227,In_358);
nor U544 (N_544,In_540,In_605);
or U545 (N_545,In_47,In_703);
or U546 (N_546,In_787,In_372);
or U547 (N_547,In_789,In_374);
nor U548 (N_548,In_446,In_109);
nand U549 (N_549,In_293,In_45);
and U550 (N_550,In_959,In_395);
and U551 (N_551,In_481,In_645);
or U552 (N_552,In_507,In_137);
and U553 (N_553,In_377,In_993);
and U554 (N_554,In_198,In_427);
nand U555 (N_555,In_29,In_518);
nand U556 (N_556,In_791,In_414);
or U557 (N_557,In_809,In_979);
and U558 (N_558,In_709,In_759);
nor U559 (N_559,In_377,In_816);
or U560 (N_560,In_693,In_478);
and U561 (N_561,In_504,In_935);
nor U562 (N_562,In_390,In_593);
xor U563 (N_563,In_816,In_75);
nor U564 (N_564,In_202,In_841);
nor U565 (N_565,In_174,In_587);
nor U566 (N_566,In_308,In_985);
or U567 (N_567,In_53,In_709);
nand U568 (N_568,In_118,In_674);
and U569 (N_569,In_753,In_804);
xor U570 (N_570,In_91,In_321);
and U571 (N_571,In_261,In_599);
nor U572 (N_572,In_152,In_285);
and U573 (N_573,In_73,In_460);
and U574 (N_574,In_155,In_939);
nor U575 (N_575,In_155,In_170);
nor U576 (N_576,In_102,In_359);
or U577 (N_577,In_894,In_577);
and U578 (N_578,In_702,In_148);
nor U579 (N_579,In_393,In_946);
and U580 (N_580,In_80,In_579);
and U581 (N_581,In_208,In_76);
or U582 (N_582,In_894,In_472);
nand U583 (N_583,In_705,In_307);
nand U584 (N_584,In_835,In_965);
and U585 (N_585,In_193,In_438);
nand U586 (N_586,In_378,In_528);
and U587 (N_587,In_195,In_437);
nand U588 (N_588,In_431,In_947);
nand U589 (N_589,In_348,In_160);
or U590 (N_590,In_707,In_179);
nor U591 (N_591,In_643,In_542);
and U592 (N_592,In_786,In_142);
nor U593 (N_593,In_560,In_428);
nor U594 (N_594,In_162,In_481);
nand U595 (N_595,In_746,In_185);
nor U596 (N_596,In_239,In_47);
nand U597 (N_597,In_813,In_382);
nor U598 (N_598,In_594,In_340);
nand U599 (N_599,In_222,In_601);
and U600 (N_600,In_531,In_922);
or U601 (N_601,In_898,In_22);
and U602 (N_602,In_44,In_106);
or U603 (N_603,In_545,In_754);
nor U604 (N_604,In_621,In_371);
nand U605 (N_605,In_277,In_126);
nor U606 (N_606,In_768,In_178);
and U607 (N_607,In_527,In_959);
nand U608 (N_608,In_596,In_440);
or U609 (N_609,In_433,In_92);
nand U610 (N_610,In_221,In_460);
or U611 (N_611,In_12,In_744);
nor U612 (N_612,In_119,In_191);
nor U613 (N_613,In_137,In_970);
nand U614 (N_614,In_692,In_279);
nor U615 (N_615,In_729,In_754);
or U616 (N_616,In_65,In_725);
nand U617 (N_617,In_277,In_308);
nand U618 (N_618,In_25,In_350);
nand U619 (N_619,In_145,In_614);
nor U620 (N_620,In_480,In_46);
or U621 (N_621,In_309,In_116);
and U622 (N_622,In_196,In_855);
and U623 (N_623,In_749,In_978);
nor U624 (N_624,In_642,In_578);
or U625 (N_625,In_612,In_529);
or U626 (N_626,In_203,In_805);
or U627 (N_627,In_176,In_994);
and U628 (N_628,In_79,In_711);
xor U629 (N_629,In_739,In_136);
and U630 (N_630,In_355,In_575);
nand U631 (N_631,In_925,In_61);
and U632 (N_632,In_790,In_197);
nor U633 (N_633,In_457,In_856);
nand U634 (N_634,In_901,In_5);
nand U635 (N_635,In_674,In_216);
and U636 (N_636,In_894,In_219);
nand U637 (N_637,In_650,In_436);
or U638 (N_638,In_759,In_204);
and U639 (N_639,In_64,In_109);
nor U640 (N_640,In_0,In_512);
and U641 (N_641,In_14,In_833);
nor U642 (N_642,In_636,In_821);
nand U643 (N_643,In_899,In_956);
xor U644 (N_644,In_869,In_251);
and U645 (N_645,In_254,In_930);
and U646 (N_646,In_379,In_797);
and U647 (N_647,In_894,In_98);
nor U648 (N_648,In_409,In_350);
nor U649 (N_649,In_808,In_993);
nor U650 (N_650,In_843,In_423);
and U651 (N_651,In_256,In_104);
nor U652 (N_652,In_70,In_958);
and U653 (N_653,In_416,In_411);
and U654 (N_654,In_236,In_751);
or U655 (N_655,In_540,In_63);
and U656 (N_656,In_990,In_412);
or U657 (N_657,In_279,In_178);
nor U658 (N_658,In_326,In_26);
nor U659 (N_659,In_369,In_461);
and U660 (N_660,In_997,In_514);
or U661 (N_661,In_553,In_534);
or U662 (N_662,In_44,In_751);
or U663 (N_663,In_152,In_292);
nand U664 (N_664,In_188,In_92);
nor U665 (N_665,In_957,In_728);
and U666 (N_666,In_182,In_189);
xor U667 (N_667,In_974,In_918);
and U668 (N_668,In_76,In_660);
nand U669 (N_669,In_418,In_892);
nor U670 (N_670,In_305,In_717);
and U671 (N_671,In_473,In_940);
xor U672 (N_672,In_745,In_798);
nand U673 (N_673,In_551,In_217);
or U674 (N_674,In_812,In_692);
nor U675 (N_675,In_146,In_458);
and U676 (N_676,In_153,In_485);
nor U677 (N_677,In_719,In_470);
nor U678 (N_678,In_41,In_65);
or U679 (N_679,In_200,In_196);
or U680 (N_680,In_324,In_46);
and U681 (N_681,In_810,In_190);
or U682 (N_682,In_9,In_25);
nand U683 (N_683,In_572,In_746);
nand U684 (N_684,In_435,In_82);
and U685 (N_685,In_872,In_948);
or U686 (N_686,In_60,In_891);
nor U687 (N_687,In_964,In_402);
nand U688 (N_688,In_826,In_936);
nand U689 (N_689,In_562,In_252);
or U690 (N_690,In_653,In_341);
or U691 (N_691,In_656,In_233);
nand U692 (N_692,In_515,In_988);
or U693 (N_693,In_820,In_20);
nand U694 (N_694,In_452,In_949);
nand U695 (N_695,In_965,In_362);
nand U696 (N_696,In_244,In_155);
xnor U697 (N_697,In_165,In_918);
or U698 (N_698,In_573,In_214);
or U699 (N_699,In_853,In_494);
nor U700 (N_700,In_588,In_479);
and U701 (N_701,In_154,In_413);
and U702 (N_702,In_681,In_232);
or U703 (N_703,In_843,In_158);
and U704 (N_704,In_134,In_241);
or U705 (N_705,In_171,In_997);
and U706 (N_706,In_203,In_300);
and U707 (N_707,In_372,In_238);
nand U708 (N_708,In_434,In_416);
and U709 (N_709,In_866,In_55);
nor U710 (N_710,In_894,In_680);
nand U711 (N_711,In_485,In_804);
or U712 (N_712,In_207,In_75);
and U713 (N_713,In_931,In_262);
and U714 (N_714,In_872,In_392);
nor U715 (N_715,In_419,In_752);
and U716 (N_716,In_479,In_145);
xor U717 (N_717,In_71,In_427);
and U718 (N_718,In_232,In_819);
nand U719 (N_719,In_773,In_670);
nand U720 (N_720,In_49,In_538);
nand U721 (N_721,In_150,In_988);
and U722 (N_722,In_188,In_492);
nor U723 (N_723,In_939,In_707);
nand U724 (N_724,In_340,In_583);
or U725 (N_725,In_940,In_809);
nor U726 (N_726,In_589,In_761);
nor U727 (N_727,In_237,In_665);
or U728 (N_728,In_187,In_958);
and U729 (N_729,In_359,In_781);
and U730 (N_730,In_383,In_289);
nor U731 (N_731,In_602,In_750);
nand U732 (N_732,In_392,In_862);
nor U733 (N_733,In_493,In_925);
nand U734 (N_734,In_135,In_649);
nor U735 (N_735,In_379,In_78);
nor U736 (N_736,In_843,In_344);
or U737 (N_737,In_637,In_745);
and U738 (N_738,In_613,In_308);
nand U739 (N_739,In_339,In_35);
or U740 (N_740,In_774,In_60);
and U741 (N_741,In_192,In_6);
nand U742 (N_742,In_237,In_331);
nand U743 (N_743,In_962,In_253);
nand U744 (N_744,In_336,In_792);
and U745 (N_745,In_104,In_433);
or U746 (N_746,In_779,In_329);
xnor U747 (N_747,In_982,In_191);
and U748 (N_748,In_285,In_169);
and U749 (N_749,In_782,In_843);
and U750 (N_750,In_988,In_577);
or U751 (N_751,In_347,In_270);
nor U752 (N_752,In_311,In_43);
nand U753 (N_753,In_321,In_956);
or U754 (N_754,In_148,In_825);
and U755 (N_755,In_770,In_886);
nor U756 (N_756,In_128,In_332);
nor U757 (N_757,In_135,In_554);
and U758 (N_758,In_742,In_411);
and U759 (N_759,In_969,In_249);
or U760 (N_760,In_206,In_864);
nor U761 (N_761,In_390,In_582);
nor U762 (N_762,In_901,In_512);
and U763 (N_763,In_219,In_962);
xor U764 (N_764,In_156,In_63);
nand U765 (N_765,In_873,In_120);
nand U766 (N_766,In_402,In_937);
or U767 (N_767,In_728,In_490);
nor U768 (N_768,In_250,In_463);
and U769 (N_769,In_855,In_687);
nor U770 (N_770,In_610,In_242);
and U771 (N_771,In_471,In_788);
and U772 (N_772,In_97,In_36);
and U773 (N_773,In_632,In_919);
nand U774 (N_774,In_818,In_763);
and U775 (N_775,In_67,In_79);
nand U776 (N_776,In_747,In_420);
nor U777 (N_777,In_893,In_486);
nand U778 (N_778,In_297,In_503);
nor U779 (N_779,In_678,In_477);
or U780 (N_780,In_642,In_128);
or U781 (N_781,In_215,In_312);
and U782 (N_782,In_111,In_318);
or U783 (N_783,In_120,In_983);
nand U784 (N_784,In_569,In_229);
nand U785 (N_785,In_911,In_40);
and U786 (N_786,In_597,In_422);
nor U787 (N_787,In_39,In_226);
or U788 (N_788,In_870,In_865);
or U789 (N_789,In_848,In_781);
nor U790 (N_790,In_150,In_853);
nor U791 (N_791,In_402,In_727);
and U792 (N_792,In_363,In_50);
nand U793 (N_793,In_662,In_135);
nand U794 (N_794,In_110,In_235);
or U795 (N_795,In_966,In_875);
nor U796 (N_796,In_820,In_781);
or U797 (N_797,In_5,In_469);
nor U798 (N_798,In_192,In_39);
nand U799 (N_799,In_333,In_864);
nand U800 (N_800,In_575,In_306);
xor U801 (N_801,In_726,In_125);
nand U802 (N_802,In_16,In_880);
nand U803 (N_803,In_774,In_802);
or U804 (N_804,In_209,In_287);
nor U805 (N_805,In_227,In_58);
nand U806 (N_806,In_693,In_660);
or U807 (N_807,In_638,In_388);
nand U808 (N_808,In_309,In_318);
and U809 (N_809,In_499,In_762);
nor U810 (N_810,In_906,In_78);
nor U811 (N_811,In_534,In_456);
nor U812 (N_812,In_169,In_673);
and U813 (N_813,In_632,In_286);
or U814 (N_814,In_24,In_419);
nor U815 (N_815,In_688,In_206);
nand U816 (N_816,In_151,In_99);
nor U817 (N_817,In_108,In_204);
nor U818 (N_818,In_956,In_117);
xnor U819 (N_819,In_116,In_983);
and U820 (N_820,In_613,In_862);
or U821 (N_821,In_769,In_134);
xor U822 (N_822,In_683,In_177);
nor U823 (N_823,In_391,In_211);
nor U824 (N_824,In_104,In_366);
nor U825 (N_825,In_466,In_248);
nor U826 (N_826,In_772,In_683);
nand U827 (N_827,In_175,In_928);
or U828 (N_828,In_983,In_725);
and U829 (N_829,In_984,In_865);
and U830 (N_830,In_267,In_22);
nand U831 (N_831,In_971,In_399);
nand U832 (N_832,In_88,In_31);
nand U833 (N_833,In_899,In_462);
and U834 (N_834,In_736,In_418);
nor U835 (N_835,In_663,In_880);
nand U836 (N_836,In_78,In_913);
nand U837 (N_837,In_644,In_515);
and U838 (N_838,In_902,In_982);
nor U839 (N_839,In_602,In_719);
and U840 (N_840,In_466,In_852);
nor U841 (N_841,In_861,In_556);
nand U842 (N_842,In_568,In_910);
and U843 (N_843,In_134,In_338);
nand U844 (N_844,In_422,In_627);
nand U845 (N_845,In_73,In_18);
nand U846 (N_846,In_565,In_511);
and U847 (N_847,In_491,In_186);
nor U848 (N_848,In_797,In_864);
or U849 (N_849,In_559,In_851);
nor U850 (N_850,In_440,In_818);
and U851 (N_851,In_782,In_127);
or U852 (N_852,In_99,In_482);
or U853 (N_853,In_962,In_123);
or U854 (N_854,In_581,In_759);
and U855 (N_855,In_855,In_980);
nand U856 (N_856,In_166,In_692);
nand U857 (N_857,In_60,In_379);
nand U858 (N_858,In_288,In_557);
nand U859 (N_859,In_522,In_187);
and U860 (N_860,In_220,In_327);
nand U861 (N_861,In_383,In_15);
nand U862 (N_862,In_671,In_784);
nor U863 (N_863,In_593,In_884);
or U864 (N_864,In_510,In_514);
nand U865 (N_865,In_989,In_796);
nor U866 (N_866,In_37,In_65);
nand U867 (N_867,In_906,In_703);
or U868 (N_868,In_476,In_900);
nand U869 (N_869,In_645,In_122);
or U870 (N_870,In_615,In_297);
xnor U871 (N_871,In_824,In_560);
nand U872 (N_872,In_510,In_758);
nand U873 (N_873,In_94,In_986);
or U874 (N_874,In_821,In_449);
and U875 (N_875,In_801,In_298);
nand U876 (N_876,In_556,In_174);
nand U877 (N_877,In_292,In_875);
and U878 (N_878,In_381,In_719);
nor U879 (N_879,In_529,In_528);
and U880 (N_880,In_60,In_755);
and U881 (N_881,In_755,In_542);
or U882 (N_882,In_34,In_91);
nand U883 (N_883,In_953,In_493);
nand U884 (N_884,In_498,In_8);
nor U885 (N_885,In_808,In_140);
and U886 (N_886,In_621,In_957);
xor U887 (N_887,In_516,In_374);
or U888 (N_888,In_993,In_443);
and U889 (N_889,In_301,In_203);
nor U890 (N_890,In_823,In_918);
nor U891 (N_891,In_108,In_465);
and U892 (N_892,In_347,In_873);
or U893 (N_893,In_967,In_616);
and U894 (N_894,In_432,In_424);
nand U895 (N_895,In_206,In_597);
nand U896 (N_896,In_569,In_972);
nand U897 (N_897,In_261,In_913);
and U898 (N_898,In_389,In_593);
nand U899 (N_899,In_552,In_461);
nand U900 (N_900,In_164,In_790);
nand U901 (N_901,In_736,In_334);
or U902 (N_902,In_334,In_754);
and U903 (N_903,In_936,In_696);
nand U904 (N_904,In_729,In_571);
and U905 (N_905,In_812,In_546);
nor U906 (N_906,In_551,In_799);
or U907 (N_907,In_772,In_590);
nor U908 (N_908,In_205,In_937);
or U909 (N_909,In_39,In_504);
or U910 (N_910,In_325,In_761);
nor U911 (N_911,In_888,In_80);
or U912 (N_912,In_996,In_7);
nand U913 (N_913,In_817,In_736);
nand U914 (N_914,In_129,In_703);
nand U915 (N_915,In_109,In_499);
nand U916 (N_916,In_568,In_19);
nor U917 (N_917,In_690,In_681);
and U918 (N_918,In_286,In_234);
or U919 (N_919,In_163,In_60);
nor U920 (N_920,In_64,In_555);
nor U921 (N_921,In_271,In_90);
and U922 (N_922,In_133,In_190);
nand U923 (N_923,In_97,In_112);
nand U924 (N_924,In_108,In_557);
nand U925 (N_925,In_364,In_35);
and U926 (N_926,In_131,In_569);
nor U927 (N_927,In_544,In_906);
nand U928 (N_928,In_618,In_360);
nor U929 (N_929,In_798,In_359);
and U930 (N_930,In_183,In_459);
and U931 (N_931,In_457,In_843);
or U932 (N_932,In_325,In_33);
nand U933 (N_933,In_390,In_736);
xnor U934 (N_934,In_238,In_740);
nor U935 (N_935,In_777,In_707);
nand U936 (N_936,In_793,In_931);
or U937 (N_937,In_704,In_699);
nor U938 (N_938,In_91,In_434);
nor U939 (N_939,In_188,In_312);
nor U940 (N_940,In_231,In_905);
or U941 (N_941,In_846,In_500);
nand U942 (N_942,In_296,In_200);
nor U943 (N_943,In_872,In_743);
or U944 (N_944,In_206,In_844);
and U945 (N_945,In_427,In_70);
and U946 (N_946,In_299,In_313);
or U947 (N_947,In_944,In_343);
xnor U948 (N_948,In_536,In_71);
or U949 (N_949,In_3,In_923);
nor U950 (N_950,In_527,In_851);
nor U951 (N_951,In_777,In_584);
and U952 (N_952,In_877,In_623);
nand U953 (N_953,In_745,In_840);
nand U954 (N_954,In_184,In_846);
nor U955 (N_955,In_852,In_713);
nand U956 (N_956,In_727,In_845);
nand U957 (N_957,In_602,In_99);
or U958 (N_958,In_500,In_629);
or U959 (N_959,In_1,In_469);
or U960 (N_960,In_865,In_557);
nand U961 (N_961,In_801,In_837);
nand U962 (N_962,In_511,In_363);
and U963 (N_963,In_656,In_636);
or U964 (N_964,In_907,In_860);
nor U965 (N_965,In_479,In_742);
and U966 (N_966,In_787,In_857);
nand U967 (N_967,In_219,In_842);
and U968 (N_968,In_601,In_356);
xor U969 (N_969,In_438,In_137);
or U970 (N_970,In_20,In_314);
nand U971 (N_971,In_288,In_901);
nand U972 (N_972,In_694,In_877);
and U973 (N_973,In_767,In_691);
nand U974 (N_974,In_486,In_849);
nand U975 (N_975,In_177,In_224);
or U976 (N_976,In_854,In_111);
or U977 (N_977,In_458,In_38);
nand U978 (N_978,In_49,In_78);
or U979 (N_979,In_340,In_289);
nand U980 (N_980,In_270,In_390);
nor U981 (N_981,In_805,In_105);
nor U982 (N_982,In_136,In_473);
or U983 (N_983,In_714,In_543);
nand U984 (N_984,In_836,In_693);
and U985 (N_985,In_761,In_687);
or U986 (N_986,In_94,In_149);
nand U987 (N_987,In_499,In_455);
nor U988 (N_988,In_146,In_993);
nor U989 (N_989,In_739,In_435);
nor U990 (N_990,In_745,In_847);
nor U991 (N_991,In_534,In_231);
or U992 (N_992,In_76,In_380);
or U993 (N_993,In_368,In_816);
or U994 (N_994,In_247,In_173);
or U995 (N_995,In_131,In_457);
nand U996 (N_996,In_556,In_468);
and U997 (N_997,In_789,In_757);
nand U998 (N_998,In_392,In_724);
nor U999 (N_999,In_999,In_826);
nor U1000 (N_1000,N_69,N_871);
and U1001 (N_1001,N_428,N_357);
nand U1002 (N_1002,N_302,N_445);
and U1003 (N_1003,N_405,N_762);
nor U1004 (N_1004,N_543,N_306);
and U1005 (N_1005,N_728,N_168);
nand U1006 (N_1006,N_855,N_316);
nand U1007 (N_1007,N_459,N_845);
or U1008 (N_1008,N_456,N_644);
and U1009 (N_1009,N_551,N_438);
nand U1010 (N_1010,N_144,N_174);
and U1011 (N_1011,N_145,N_641);
or U1012 (N_1012,N_476,N_392);
nor U1013 (N_1013,N_881,N_536);
or U1014 (N_1014,N_196,N_679);
and U1015 (N_1015,N_495,N_265);
or U1016 (N_1016,N_336,N_92);
and U1017 (N_1017,N_226,N_654);
and U1018 (N_1018,N_53,N_124);
nor U1019 (N_1019,N_149,N_88);
or U1020 (N_1020,N_841,N_81);
and U1021 (N_1021,N_709,N_540);
nor U1022 (N_1022,N_458,N_947);
or U1023 (N_1023,N_719,N_868);
nand U1024 (N_1024,N_194,N_991);
nor U1025 (N_1025,N_922,N_110);
or U1026 (N_1026,N_751,N_776);
nand U1027 (N_1027,N_492,N_975);
or U1028 (N_1028,N_250,N_322);
nand U1029 (N_1029,N_32,N_470);
nor U1030 (N_1030,N_840,N_127);
and U1031 (N_1031,N_851,N_400);
or U1032 (N_1032,N_234,N_489);
or U1033 (N_1033,N_285,N_299);
or U1034 (N_1034,N_598,N_972);
nor U1035 (N_1035,N_443,N_878);
nand U1036 (N_1036,N_1,N_687);
nor U1037 (N_1037,N_605,N_839);
nand U1038 (N_1038,N_921,N_488);
nand U1039 (N_1039,N_510,N_201);
or U1040 (N_1040,N_589,N_673);
nor U1041 (N_1041,N_457,N_227);
xor U1042 (N_1042,N_882,N_100);
or U1043 (N_1043,N_827,N_918);
nor U1044 (N_1044,N_67,N_943);
and U1045 (N_1045,N_232,N_38);
xnor U1046 (N_1046,N_786,N_600);
or U1047 (N_1047,N_782,N_650);
or U1048 (N_1048,N_792,N_122);
or U1049 (N_1049,N_515,N_266);
xnor U1050 (N_1050,N_318,N_622);
nand U1051 (N_1051,N_633,N_118);
nand U1052 (N_1052,N_615,N_61);
nand U1053 (N_1053,N_531,N_404);
nand U1054 (N_1054,N_970,N_214);
or U1055 (N_1055,N_572,N_460);
or U1056 (N_1056,N_158,N_397);
nand U1057 (N_1057,N_288,N_101);
xnor U1058 (N_1058,N_765,N_399);
nor U1059 (N_1059,N_80,N_703);
nand U1060 (N_1060,N_13,N_575);
nand U1061 (N_1061,N_235,N_678);
nor U1062 (N_1062,N_321,N_542);
or U1063 (N_1063,N_933,N_512);
or U1064 (N_1064,N_983,N_668);
nor U1065 (N_1065,N_718,N_793);
nor U1066 (N_1066,N_468,N_927);
nor U1067 (N_1067,N_995,N_653);
nor U1068 (N_1068,N_570,N_51);
nor U1069 (N_1069,N_899,N_451);
nor U1070 (N_1070,N_97,N_329);
nor U1071 (N_1071,N_906,N_857);
nand U1072 (N_1072,N_330,N_325);
and U1073 (N_1073,N_638,N_340);
or U1074 (N_1074,N_375,N_346);
or U1075 (N_1075,N_130,N_629);
and U1076 (N_1076,N_212,N_382);
nor U1077 (N_1077,N_713,N_213);
nor U1078 (N_1078,N_463,N_772);
nand U1079 (N_1079,N_305,N_619);
nand U1080 (N_1080,N_754,N_953);
nor U1081 (N_1081,N_467,N_643);
and U1082 (N_1082,N_362,N_537);
and U1083 (N_1083,N_780,N_612);
nand U1084 (N_1084,N_656,N_17);
and U1085 (N_1085,N_828,N_592);
nor U1086 (N_1086,N_702,N_788);
nand U1087 (N_1087,N_422,N_221);
or U1088 (N_1088,N_509,N_395);
nor U1089 (N_1089,N_816,N_850);
nand U1090 (N_1090,N_18,N_96);
nand U1091 (N_1091,N_402,N_87);
nor U1092 (N_1092,N_401,N_34);
nand U1093 (N_1093,N_313,N_108);
or U1094 (N_1094,N_834,N_370);
or U1095 (N_1095,N_126,N_603);
nor U1096 (N_1096,N_291,N_939);
or U1097 (N_1097,N_339,N_490);
nor U1098 (N_1098,N_717,N_189);
xnor U1099 (N_1099,N_270,N_930);
and U1100 (N_1100,N_160,N_867);
or U1101 (N_1101,N_117,N_987);
nor U1102 (N_1102,N_71,N_70);
nor U1103 (N_1103,N_699,N_215);
or U1104 (N_1104,N_90,N_72);
or U1105 (N_1105,N_573,N_19);
or U1106 (N_1106,N_7,N_833);
and U1107 (N_1107,N_353,N_990);
or U1108 (N_1108,N_611,N_989);
or U1109 (N_1109,N_279,N_799);
xor U1110 (N_1110,N_480,N_271);
nor U1111 (N_1111,N_91,N_301);
and U1112 (N_1112,N_435,N_294);
or U1113 (N_1113,N_154,N_686);
nor U1114 (N_1114,N_932,N_550);
nand U1115 (N_1115,N_333,N_43);
nand U1116 (N_1116,N_711,N_278);
or U1117 (N_1117,N_585,N_31);
nand U1118 (N_1118,N_159,N_712);
or U1119 (N_1119,N_197,N_599);
nor U1120 (N_1120,N_511,N_387);
and U1121 (N_1121,N_167,N_920);
xor U1122 (N_1122,N_95,N_426);
and U1123 (N_1123,N_390,N_56);
and U1124 (N_1124,N_162,N_5);
and U1125 (N_1125,N_556,N_916);
nand U1126 (N_1126,N_548,N_716);
and U1127 (N_1127,N_809,N_513);
and U1128 (N_1128,N_350,N_580);
and U1129 (N_1129,N_693,N_264);
nor U1130 (N_1130,N_450,N_566);
nor U1131 (N_1131,N_787,N_647);
nand U1132 (N_1132,N_186,N_631);
nand U1133 (N_1133,N_231,N_873);
nor U1134 (N_1134,N_637,N_273);
and U1135 (N_1135,N_262,N_103);
and U1136 (N_1136,N_913,N_961);
or U1137 (N_1137,N_836,N_398);
nand U1138 (N_1138,N_888,N_247);
and U1139 (N_1139,N_134,N_147);
nor U1140 (N_1140,N_645,N_892);
and U1141 (N_1141,N_132,N_946);
nand U1142 (N_1142,N_623,N_574);
or U1143 (N_1143,N_307,N_113);
nor U1144 (N_1144,N_85,N_874);
and U1145 (N_1145,N_671,N_576);
xor U1146 (N_1146,N_284,N_926);
or U1147 (N_1147,N_140,N_198);
nor U1148 (N_1148,N_430,N_44);
and U1149 (N_1149,N_50,N_176);
and U1150 (N_1150,N_449,N_937);
or U1151 (N_1151,N_242,N_204);
and U1152 (N_1152,N_706,N_859);
nand U1153 (N_1153,N_484,N_852);
and U1154 (N_1154,N_314,N_311);
and U1155 (N_1155,N_727,N_406);
nand U1156 (N_1156,N_666,N_384);
nand U1157 (N_1157,N_224,N_903);
or U1158 (N_1158,N_994,N_199);
nor U1159 (N_1159,N_944,N_758);
and U1160 (N_1160,N_800,N_976);
and U1161 (N_1161,N_843,N_334);
nor U1162 (N_1162,N_900,N_94);
nor U1163 (N_1163,N_41,N_487);
nand U1164 (N_1164,N_137,N_68);
and U1165 (N_1165,N_378,N_896);
and U1166 (N_1166,N_564,N_496);
and U1167 (N_1167,N_343,N_829);
nor U1168 (N_1168,N_30,N_997);
nand U1169 (N_1169,N_355,N_486);
or U1170 (N_1170,N_440,N_965);
or U1171 (N_1171,N_689,N_697);
or U1172 (N_1172,N_909,N_373);
and U1173 (N_1173,N_520,N_142);
or U1174 (N_1174,N_465,N_823);
nand U1175 (N_1175,N_614,N_606);
nor U1176 (N_1176,N_905,N_931);
and U1177 (N_1177,N_519,N_664);
or U1178 (N_1178,N_309,N_907);
nand U1179 (N_1179,N_919,N_218);
and U1180 (N_1180,N_82,N_889);
and U1181 (N_1181,N_796,N_177);
and U1182 (N_1182,N_10,N_791);
or U1183 (N_1183,N_323,N_532);
and U1184 (N_1184,N_26,N_195);
xnor U1185 (N_1185,N_77,N_523);
and U1186 (N_1186,N_182,N_741);
nand U1187 (N_1187,N_750,N_794);
or U1188 (N_1188,N_720,N_152);
or U1189 (N_1189,N_27,N_846);
nand U1190 (N_1190,N_724,N_534);
nor U1191 (N_1191,N_55,N_674);
or U1192 (N_1192,N_261,N_587);
and U1193 (N_1193,N_832,N_58);
and U1194 (N_1194,N_86,N_295);
nor U1195 (N_1195,N_958,N_24);
nand U1196 (N_1196,N_917,N_950);
nand U1197 (N_1197,N_66,N_277);
nor U1198 (N_1198,N_442,N_815);
xnor U1199 (N_1199,N_973,N_683);
or U1200 (N_1200,N_814,N_856);
or U1201 (N_1201,N_191,N_607);
or U1202 (N_1202,N_811,N_139);
and U1203 (N_1203,N_848,N_183);
or U1204 (N_1204,N_745,N_230);
nor U1205 (N_1205,N_640,N_769);
and U1206 (N_1206,N_483,N_415);
or U1207 (N_1207,N_744,N_854);
and U1208 (N_1208,N_381,N_303);
nand U1209 (N_1209,N_36,N_114);
or U1210 (N_1210,N_16,N_865);
and U1211 (N_1211,N_942,N_696);
or U1212 (N_1212,N_354,N_659);
or U1213 (N_1213,N_363,N_698);
nor U1214 (N_1214,N_388,N_651);
nor U1215 (N_1215,N_393,N_684);
nand U1216 (N_1216,N_57,N_173);
and U1217 (N_1217,N_692,N_42);
xnor U1218 (N_1218,N_286,N_726);
or U1219 (N_1219,N_352,N_785);
nor U1220 (N_1220,N_968,N_842);
nand U1221 (N_1221,N_813,N_8);
and U1222 (N_1222,N_984,N_898);
and U1223 (N_1223,N_447,N_617);
nand U1224 (N_1224,N_368,N_327);
and U1225 (N_1225,N_151,N_268);
nand U1226 (N_1226,N_773,N_675);
nand U1227 (N_1227,N_634,N_437);
or U1228 (N_1228,N_672,N_967);
or U1229 (N_1229,N_337,N_418);
nand U1230 (N_1230,N_347,N_798);
nand U1231 (N_1231,N_642,N_568);
and U1232 (N_1232,N_148,N_948);
nand U1233 (N_1233,N_396,N_131);
or U1234 (N_1234,N_209,N_715);
or U1235 (N_1235,N_150,N_365);
nor U1236 (N_1236,N_190,N_880);
nand U1237 (N_1237,N_552,N_102);
nand U1238 (N_1238,N_872,N_45);
or U1239 (N_1239,N_136,N_680);
xnor U1240 (N_1240,N_344,N_662);
and U1241 (N_1241,N_98,N_359);
nand U1242 (N_1242,N_563,N_240);
and U1243 (N_1243,N_924,N_915);
or U1244 (N_1244,N_251,N_14);
nand U1245 (N_1245,N_665,N_471);
nor U1246 (N_1246,N_602,N_626);
xnor U1247 (N_1247,N_249,N_554);
or U1248 (N_1248,N_39,N_707);
and U1249 (N_1249,N_328,N_192);
nand U1250 (N_1250,N_421,N_371);
nand U1251 (N_1251,N_826,N_789);
or U1252 (N_1252,N_923,N_748);
nand U1253 (N_1253,N_394,N_407);
nor U1254 (N_1254,N_739,N_992);
nor U1255 (N_1255,N_93,N_47);
or U1256 (N_1256,N_596,N_356);
nor U1257 (N_1257,N_505,N_525);
nor U1258 (N_1258,N_263,N_960);
xor U1259 (N_1259,N_172,N_964);
or U1260 (N_1260,N_755,N_613);
xnor U1261 (N_1261,N_529,N_508);
and U1262 (N_1262,N_770,N_475);
and U1263 (N_1263,N_115,N_372);
or U1264 (N_1264,N_893,N_778);
or U1265 (N_1265,N_819,N_795);
nand U1266 (N_1266,N_389,N_267);
or U1267 (N_1267,N_335,N_481);
or U1268 (N_1268,N_52,N_620);
and U1269 (N_1269,N_446,N_584);
nor U1270 (N_1270,N_743,N_431);
xnor U1271 (N_1271,N_831,N_660);
nor U1272 (N_1272,N_171,N_908);
nand U1273 (N_1273,N_805,N_830);
xnor U1274 (N_1274,N_416,N_287);
or U1275 (N_1275,N_582,N_749);
nor U1276 (N_1276,N_812,N_601);
and U1277 (N_1277,N_507,N_506);
nand U1278 (N_1278,N_763,N_894);
and U1279 (N_1279,N_466,N_364);
nor U1280 (N_1280,N_616,N_590);
or U1281 (N_1281,N_982,N_521);
nor U1282 (N_1282,N_527,N_141);
or U1283 (N_1283,N_89,N_245);
and U1284 (N_1284,N_220,N_414);
and U1285 (N_1285,N_156,N_83);
or U1286 (N_1286,N_822,N_380);
or U1287 (N_1287,N_817,N_559);
nand U1288 (N_1288,N_806,N_635);
nor U1289 (N_1289,N_383,N_586);
nand U1290 (N_1290,N_424,N_569);
or U1291 (N_1291,N_260,N_106);
nor U1292 (N_1292,N_121,N_0);
nand U1293 (N_1293,N_928,N_562);
nor U1294 (N_1294,N_76,N_236);
and U1295 (N_1295,N_593,N_135);
nand U1296 (N_1296,N_479,N_516);
or U1297 (N_1297,N_253,N_835);
or U1298 (N_1298,N_25,N_434);
and U1299 (N_1299,N_317,N_256);
nor U1300 (N_1300,N_54,N_630);
or U1301 (N_1301,N_891,N_175);
nor U1302 (N_1302,N_708,N_169);
nor U1303 (N_1303,N_345,N_376);
and U1304 (N_1304,N_21,N_652);
and U1305 (N_1305,N_412,N_233);
nor U1306 (N_1306,N_632,N_409);
and U1307 (N_1307,N_272,N_771);
and U1308 (N_1308,N_825,N_441);
nor U1309 (N_1309,N_75,N_366);
or U1310 (N_1310,N_700,N_107);
and U1311 (N_1311,N_732,N_723);
or U1312 (N_1312,N_936,N_105);
or U1313 (N_1313,N_99,N_565);
or U1314 (N_1314,N_738,N_956);
or U1315 (N_1315,N_377,N_290);
xnor U1316 (N_1316,N_636,N_897);
nand U1317 (N_1317,N_914,N_292);
nand U1318 (N_1318,N_883,N_462);
or U1319 (N_1319,N_688,N_23);
nor U1320 (N_1320,N_40,N_248);
and U1321 (N_1321,N_500,N_858);
nor U1322 (N_1322,N_608,N_461);
nand U1323 (N_1323,N_863,N_999);
nand U1324 (N_1324,N_977,N_257);
nand U1325 (N_1325,N_497,N_385);
nor U1326 (N_1326,N_818,N_297);
and U1327 (N_1327,N_319,N_704);
or U1328 (N_1328,N_403,N_801);
and U1329 (N_1329,N_133,N_553);
or U1330 (N_1330,N_861,N_109);
or U1331 (N_1331,N_735,N_170);
and U1332 (N_1332,N_747,N_361);
nand U1333 (N_1333,N_955,N_65);
or U1334 (N_1334,N_22,N_60);
or U1335 (N_1335,N_207,N_324);
nor U1336 (N_1336,N_493,N_781);
or U1337 (N_1337,N_996,N_3);
nand U1338 (N_1338,N_351,N_962);
nor U1339 (N_1339,N_369,N_4);
xnor U1340 (N_1340,N_420,N_482);
and U1341 (N_1341,N_15,N_890);
nor U1342 (N_1342,N_119,N_934);
or U1343 (N_1343,N_244,N_208);
nand U1344 (N_1344,N_911,N_649);
nand U1345 (N_1345,N_957,N_941);
or U1346 (N_1346,N_432,N_386);
xor U1347 (N_1347,N_283,N_225);
nor U1348 (N_1348,N_761,N_676);
nand U1349 (N_1349,N_59,N_29);
nor U1350 (N_1350,N_777,N_541);
nand U1351 (N_1351,N_966,N_705);
nor U1352 (N_1352,N_945,N_206);
and U1353 (N_1353,N_963,N_326);
nor U1354 (N_1354,N_320,N_20);
and U1355 (N_1355,N_433,N_84);
nand U1356 (N_1356,N_112,N_11);
or U1357 (N_1357,N_193,N_538);
and U1358 (N_1358,N_222,N_804);
nor U1359 (N_1359,N_904,N_444);
nand U1360 (N_1360,N_558,N_658);
or U1361 (N_1361,N_737,N_165);
or U1362 (N_1362,N_628,N_837);
nor U1363 (N_1363,N_760,N_618);
or U1364 (N_1364,N_312,N_79);
or U1365 (N_1365,N_217,N_238);
nand U1366 (N_1366,N_949,N_978);
or U1367 (N_1367,N_581,N_701);
nor U1368 (N_1368,N_503,N_866);
nor U1369 (N_1369,N_464,N_535);
or U1370 (N_1370,N_498,N_610);
or U1371 (N_1371,N_448,N_875);
or U1372 (N_1372,N_423,N_533);
nand U1373 (N_1373,N_501,N_627);
nand U1374 (N_1374,N_621,N_824);
nor U1375 (N_1375,N_200,N_413);
or U1376 (N_1376,N_986,N_655);
nand U1377 (N_1377,N_969,N_417);
nor U1378 (N_1378,N_239,N_111);
and U1379 (N_1379,N_123,N_935);
nor U1380 (N_1380,N_864,N_869);
nand U1381 (N_1381,N_667,N_821);
and U1382 (N_1382,N_988,N_116);
xor U1383 (N_1383,N_155,N_661);
and U1384 (N_1384,N_847,N_298);
and U1385 (N_1385,N_885,N_849);
nor U1386 (N_1386,N_341,N_571);
nand U1387 (N_1387,N_669,N_408);
or U1388 (N_1388,N_128,N_560);
or U1389 (N_1389,N_491,N_895);
nor U1390 (N_1390,N_379,N_731);
or U1391 (N_1391,N_6,N_591);
or U1392 (N_1392,N_280,N_528);
nand U1393 (N_1393,N_241,N_710);
and U1394 (N_1394,N_539,N_522);
or U1395 (N_1395,N_657,N_682);
and U1396 (N_1396,N_547,N_546);
or U1397 (N_1397,N_721,N_205);
or U1398 (N_1398,N_677,N_243);
and U1399 (N_1399,N_803,N_729);
and U1400 (N_1400,N_853,N_161);
or U1401 (N_1401,N_879,N_959);
or U1402 (N_1402,N_427,N_518);
nand U1403 (N_1403,N_223,N_597);
and U1404 (N_1404,N_951,N_179);
xnor U1405 (N_1405,N_348,N_300);
or U1406 (N_1406,N_64,N_129);
or U1407 (N_1407,N_595,N_742);
or U1408 (N_1408,N_74,N_410);
nor U1409 (N_1409,N_281,N_293);
or U1410 (N_1410,N_419,N_504);
nor U1411 (N_1411,N_544,N_246);
nor U1412 (N_1412,N_734,N_929);
and U1413 (N_1413,N_436,N_624);
nand U1414 (N_1414,N_517,N_358);
nand U1415 (N_1415,N_971,N_940);
nor U1416 (N_1416,N_210,N_808);
and U1417 (N_1417,N_993,N_494);
nand U1418 (N_1418,N_998,N_579);
nor U1419 (N_1419,N_429,N_802);
and U1420 (N_1420,N_910,N_981);
nand U1421 (N_1421,N_545,N_120);
nand U1422 (N_1422,N_764,N_153);
and U1423 (N_1423,N_736,N_255);
or U1424 (N_1424,N_567,N_577);
and U1425 (N_1425,N_877,N_530);
nand U1426 (N_1426,N_391,N_663);
or U1427 (N_1427,N_478,N_695);
and U1428 (N_1428,N_767,N_274);
or U1429 (N_1429,N_766,N_304);
and U1430 (N_1430,N_48,N_746);
and U1431 (N_1431,N_714,N_37);
nand U1432 (N_1432,N_779,N_588);
xor U1433 (N_1433,N_163,N_164);
and U1434 (N_1434,N_331,N_578);
nand U1435 (N_1435,N_775,N_12);
nand U1436 (N_1436,N_876,N_768);
xor U1437 (N_1437,N_73,N_9);
or U1438 (N_1438,N_797,N_887);
and U1439 (N_1439,N_954,N_49);
or U1440 (N_1440,N_925,N_146);
nand U1441 (N_1441,N_374,N_985);
and U1442 (N_1442,N_187,N_157);
and U1443 (N_1443,N_203,N_469);
nor U1444 (N_1444,N_604,N_282);
and U1445 (N_1445,N_360,N_557);
nand U1446 (N_1446,N_725,N_884);
and U1447 (N_1447,N_912,N_807);
nand U1448 (N_1448,N_790,N_514);
nor U1449 (N_1449,N_35,N_28);
and U1450 (N_1450,N_974,N_104);
nor U1451 (N_1451,N_237,N_276);
nand U1452 (N_1452,N_838,N_901);
nand U1453 (N_1453,N_338,N_753);
or U1454 (N_1454,N_180,N_477);
nand U1455 (N_1455,N_33,N_583);
or U1456 (N_1456,N_252,N_499);
nand U1457 (N_1457,N_485,N_774);
and U1458 (N_1458,N_228,N_594);
nor U1459 (N_1459,N_216,N_609);
and U1460 (N_1460,N_125,N_862);
and U1461 (N_1461,N_46,N_902);
or U1462 (N_1462,N_308,N_425);
nand U1463 (N_1463,N_979,N_844);
and U1464 (N_1464,N_202,N_783);
nand U1465 (N_1465,N_63,N_980);
or U1466 (N_1466,N_184,N_860);
and U1467 (N_1467,N_691,N_820);
or U1468 (N_1468,N_78,N_62);
nand U1469 (N_1469,N_2,N_315);
nand U1470 (N_1470,N_269,N_188);
nand U1471 (N_1471,N_526,N_258);
and U1472 (N_1472,N_411,N_452);
nor U1473 (N_1473,N_555,N_646);
nor U1474 (N_1474,N_952,N_648);
nor U1475 (N_1475,N_474,N_757);
and U1476 (N_1476,N_938,N_181);
nand U1477 (N_1477,N_342,N_694);
and U1478 (N_1478,N_759,N_670);
nand U1479 (N_1479,N_524,N_756);
or U1480 (N_1480,N_439,N_289);
nand U1481 (N_1481,N_685,N_502);
nor U1482 (N_1482,N_454,N_455);
nand U1483 (N_1483,N_229,N_211);
nor U1484 (N_1484,N_733,N_639);
and U1485 (N_1485,N_259,N_166);
or U1486 (N_1486,N_219,N_730);
and U1487 (N_1487,N_332,N_810);
nand U1488 (N_1488,N_681,N_349);
and U1489 (N_1489,N_143,N_870);
nor U1490 (N_1490,N_886,N_690);
nor U1491 (N_1491,N_138,N_472);
and U1492 (N_1492,N_275,N_722);
or U1493 (N_1493,N_367,N_752);
or U1494 (N_1494,N_296,N_625);
nand U1495 (N_1495,N_473,N_740);
nand U1496 (N_1496,N_178,N_561);
or U1497 (N_1497,N_185,N_784);
nand U1498 (N_1498,N_453,N_549);
nand U1499 (N_1499,N_310,N_254);
or U1500 (N_1500,N_754,N_422);
nor U1501 (N_1501,N_655,N_636);
nand U1502 (N_1502,N_112,N_192);
nor U1503 (N_1503,N_280,N_952);
nor U1504 (N_1504,N_162,N_502);
and U1505 (N_1505,N_461,N_145);
and U1506 (N_1506,N_944,N_670);
xor U1507 (N_1507,N_868,N_824);
xor U1508 (N_1508,N_515,N_400);
nand U1509 (N_1509,N_811,N_493);
or U1510 (N_1510,N_393,N_179);
or U1511 (N_1511,N_330,N_777);
nor U1512 (N_1512,N_866,N_436);
nor U1513 (N_1513,N_984,N_726);
and U1514 (N_1514,N_333,N_331);
nor U1515 (N_1515,N_405,N_968);
and U1516 (N_1516,N_618,N_5);
nor U1517 (N_1517,N_468,N_627);
nor U1518 (N_1518,N_26,N_879);
nand U1519 (N_1519,N_994,N_998);
or U1520 (N_1520,N_92,N_649);
and U1521 (N_1521,N_831,N_984);
and U1522 (N_1522,N_999,N_50);
and U1523 (N_1523,N_686,N_777);
or U1524 (N_1524,N_322,N_972);
nor U1525 (N_1525,N_726,N_890);
nand U1526 (N_1526,N_823,N_381);
nand U1527 (N_1527,N_494,N_660);
or U1528 (N_1528,N_516,N_25);
or U1529 (N_1529,N_628,N_39);
or U1530 (N_1530,N_188,N_103);
or U1531 (N_1531,N_7,N_918);
and U1532 (N_1532,N_242,N_285);
nand U1533 (N_1533,N_88,N_682);
or U1534 (N_1534,N_987,N_270);
or U1535 (N_1535,N_920,N_509);
nand U1536 (N_1536,N_511,N_275);
nor U1537 (N_1537,N_135,N_971);
nor U1538 (N_1538,N_27,N_960);
or U1539 (N_1539,N_136,N_994);
and U1540 (N_1540,N_284,N_191);
nand U1541 (N_1541,N_926,N_486);
and U1542 (N_1542,N_147,N_350);
and U1543 (N_1543,N_431,N_970);
nand U1544 (N_1544,N_309,N_657);
and U1545 (N_1545,N_941,N_304);
nand U1546 (N_1546,N_702,N_428);
nor U1547 (N_1547,N_494,N_683);
or U1548 (N_1548,N_230,N_957);
or U1549 (N_1549,N_236,N_460);
xor U1550 (N_1550,N_620,N_160);
and U1551 (N_1551,N_145,N_453);
nor U1552 (N_1552,N_514,N_151);
nand U1553 (N_1553,N_347,N_29);
nor U1554 (N_1554,N_930,N_100);
or U1555 (N_1555,N_776,N_813);
or U1556 (N_1556,N_761,N_671);
nand U1557 (N_1557,N_565,N_833);
nand U1558 (N_1558,N_827,N_242);
nor U1559 (N_1559,N_237,N_826);
nand U1560 (N_1560,N_291,N_193);
nand U1561 (N_1561,N_929,N_919);
or U1562 (N_1562,N_640,N_191);
or U1563 (N_1563,N_979,N_109);
nand U1564 (N_1564,N_319,N_995);
or U1565 (N_1565,N_279,N_299);
nand U1566 (N_1566,N_298,N_521);
or U1567 (N_1567,N_188,N_381);
nor U1568 (N_1568,N_375,N_903);
and U1569 (N_1569,N_613,N_743);
or U1570 (N_1570,N_326,N_683);
nand U1571 (N_1571,N_822,N_164);
or U1572 (N_1572,N_144,N_71);
or U1573 (N_1573,N_587,N_595);
nand U1574 (N_1574,N_38,N_937);
nor U1575 (N_1575,N_208,N_432);
nor U1576 (N_1576,N_729,N_628);
or U1577 (N_1577,N_349,N_921);
or U1578 (N_1578,N_754,N_16);
and U1579 (N_1579,N_899,N_831);
nand U1580 (N_1580,N_828,N_7);
nand U1581 (N_1581,N_662,N_228);
or U1582 (N_1582,N_208,N_786);
nor U1583 (N_1583,N_319,N_255);
nand U1584 (N_1584,N_5,N_776);
nor U1585 (N_1585,N_161,N_789);
and U1586 (N_1586,N_223,N_510);
or U1587 (N_1587,N_135,N_964);
and U1588 (N_1588,N_86,N_926);
nor U1589 (N_1589,N_721,N_321);
nor U1590 (N_1590,N_114,N_820);
and U1591 (N_1591,N_744,N_122);
nor U1592 (N_1592,N_295,N_986);
or U1593 (N_1593,N_954,N_917);
nor U1594 (N_1594,N_449,N_504);
nand U1595 (N_1595,N_108,N_271);
xor U1596 (N_1596,N_180,N_637);
nor U1597 (N_1597,N_823,N_962);
xnor U1598 (N_1598,N_431,N_454);
nand U1599 (N_1599,N_316,N_898);
nand U1600 (N_1600,N_159,N_911);
and U1601 (N_1601,N_65,N_439);
or U1602 (N_1602,N_532,N_314);
nand U1603 (N_1603,N_537,N_770);
xnor U1604 (N_1604,N_574,N_989);
or U1605 (N_1605,N_900,N_367);
and U1606 (N_1606,N_334,N_384);
nor U1607 (N_1607,N_10,N_665);
xnor U1608 (N_1608,N_491,N_322);
and U1609 (N_1609,N_599,N_683);
or U1610 (N_1610,N_377,N_560);
and U1611 (N_1611,N_975,N_531);
xnor U1612 (N_1612,N_722,N_453);
or U1613 (N_1613,N_264,N_384);
and U1614 (N_1614,N_562,N_625);
and U1615 (N_1615,N_400,N_117);
nor U1616 (N_1616,N_37,N_459);
nor U1617 (N_1617,N_425,N_981);
xnor U1618 (N_1618,N_760,N_190);
or U1619 (N_1619,N_527,N_852);
nor U1620 (N_1620,N_735,N_825);
and U1621 (N_1621,N_437,N_231);
nand U1622 (N_1622,N_144,N_791);
or U1623 (N_1623,N_985,N_57);
nor U1624 (N_1624,N_293,N_280);
or U1625 (N_1625,N_273,N_53);
nor U1626 (N_1626,N_501,N_98);
or U1627 (N_1627,N_432,N_917);
and U1628 (N_1628,N_482,N_737);
or U1629 (N_1629,N_620,N_196);
nor U1630 (N_1630,N_180,N_54);
nor U1631 (N_1631,N_617,N_904);
nor U1632 (N_1632,N_443,N_208);
nand U1633 (N_1633,N_595,N_634);
or U1634 (N_1634,N_599,N_968);
and U1635 (N_1635,N_90,N_822);
or U1636 (N_1636,N_902,N_483);
nand U1637 (N_1637,N_703,N_800);
nand U1638 (N_1638,N_174,N_772);
nand U1639 (N_1639,N_839,N_543);
nand U1640 (N_1640,N_967,N_447);
nand U1641 (N_1641,N_299,N_709);
or U1642 (N_1642,N_989,N_104);
or U1643 (N_1643,N_956,N_130);
or U1644 (N_1644,N_785,N_502);
nor U1645 (N_1645,N_184,N_395);
and U1646 (N_1646,N_706,N_683);
and U1647 (N_1647,N_684,N_620);
and U1648 (N_1648,N_62,N_25);
nand U1649 (N_1649,N_954,N_510);
or U1650 (N_1650,N_763,N_642);
or U1651 (N_1651,N_775,N_409);
or U1652 (N_1652,N_197,N_356);
and U1653 (N_1653,N_713,N_359);
and U1654 (N_1654,N_476,N_973);
nor U1655 (N_1655,N_898,N_619);
or U1656 (N_1656,N_505,N_57);
nand U1657 (N_1657,N_387,N_607);
and U1658 (N_1658,N_91,N_249);
and U1659 (N_1659,N_24,N_474);
or U1660 (N_1660,N_179,N_217);
nor U1661 (N_1661,N_13,N_925);
nor U1662 (N_1662,N_819,N_897);
or U1663 (N_1663,N_854,N_941);
nor U1664 (N_1664,N_899,N_501);
nand U1665 (N_1665,N_611,N_696);
nor U1666 (N_1666,N_156,N_337);
nand U1667 (N_1667,N_826,N_144);
nand U1668 (N_1668,N_147,N_89);
and U1669 (N_1669,N_522,N_29);
nor U1670 (N_1670,N_965,N_583);
nand U1671 (N_1671,N_396,N_780);
nand U1672 (N_1672,N_321,N_4);
nor U1673 (N_1673,N_457,N_111);
and U1674 (N_1674,N_359,N_960);
or U1675 (N_1675,N_964,N_905);
or U1676 (N_1676,N_878,N_818);
nor U1677 (N_1677,N_8,N_844);
nor U1678 (N_1678,N_442,N_10);
nand U1679 (N_1679,N_71,N_274);
or U1680 (N_1680,N_151,N_419);
nor U1681 (N_1681,N_245,N_552);
nor U1682 (N_1682,N_842,N_298);
and U1683 (N_1683,N_804,N_712);
and U1684 (N_1684,N_639,N_189);
or U1685 (N_1685,N_103,N_181);
and U1686 (N_1686,N_121,N_417);
or U1687 (N_1687,N_594,N_657);
nand U1688 (N_1688,N_939,N_736);
nor U1689 (N_1689,N_86,N_273);
xnor U1690 (N_1690,N_391,N_401);
and U1691 (N_1691,N_344,N_289);
nand U1692 (N_1692,N_371,N_912);
nor U1693 (N_1693,N_790,N_530);
nor U1694 (N_1694,N_641,N_111);
nand U1695 (N_1695,N_904,N_353);
nor U1696 (N_1696,N_997,N_150);
nor U1697 (N_1697,N_224,N_142);
and U1698 (N_1698,N_897,N_882);
nor U1699 (N_1699,N_247,N_171);
nor U1700 (N_1700,N_590,N_413);
or U1701 (N_1701,N_260,N_254);
or U1702 (N_1702,N_519,N_314);
nand U1703 (N_1703,N_812,N_430);
and U1704 (N_1704,N_205,N_43);
nor U1705 (N_1705,N_138,N_302);
nand U1706 (N_1706,N_763,N_616);
or U1707 (N_1707,N_700,N_811);
xor U1708 (N_1708,N_177,N_905);
nand U1709 (N_1709,N_886,N_9);
xnor U1710 (N_1710,N_907,N_490);
nor U1711 (N_1711,N_9,N_946);
nand U1712 (N_1712,N_309,N_139);
nand U1713 (N_1713,N_168,N_926);
nand U1714 (N_1714,N_853,N_0);
nor U1715 (N_1715,N_268,N_865);
or U1716 (N_1716,N_551,N_962);
or U1717 (N_1717,N_192,N_759);
or U1718 (N_1718,N_860,N_308);
nor U1719 (N_1719,N_431,N_374);
nor U1720 (N_1720,N_673,N_10);
nand U1721 (N_1721,N_67,N_202);
or U1722 (N_1722,N_674,N_59);
and U1723 (N_1723,N_373,N_884);
or U1724 (N_1724,N_81,N_571);
and U1725 (N_1725,N_877,N_506);
and U1726 (N_1726,N_465,N_977);
and U1727 (N_1727,N_711,N_161);
or U1728 (N_1728,N_659,N_246);
or U1729 (N_1729,N_617,N_24);
xor U1730 (N_1730,N_1,N_940);
nand U1731 (N_1731,N_770,N_213);
or U1732 (N_1732,N_523,N_200);
nand U1733 (N_1733,N_471,N_204);
nand U1734 (N_1734,N_325,N_547);
or U1735 (N_1735,N_517,N_280);
and U1736 (N_1736,N_728,N_601);
nand U1737 (N_1737,N_173,N_545);
nor U1738 (N_1738,N_723,N_373);
nand U1739 (N_1739,N_847,N_198);
and U1740 (N_1740,N_933,N_273);
nand U1741 (N_1741,N_336,N_602);
and U1742 (N_1742,N_630,N_514);
nand U1743 (N_1743,N_577,N_413);
or U1744 (N_1744,N_120,N_334);
and U1745 (N_1745,N_865,N_127);
nand U1746 (N_1746,N_563,N_616);
or U1747 (N_1747,N_654,N_511);
and U1748 (N_1748,N_239,N_957);
nor U1749 (N_1749,N_139,N_128);
or U1750 (N_1750,N_172,N_730);
nor U1751 (N_1751,N_144,N_269);
or U1752 (N_1752,N_386,N_361);
or U1753 (N_1753,N_842,N_780);
or U1754 (N_1754,N_32,N_654);
or U1755 (N_1755,N_745,N_217);
and U1756 (N_1756,N_777,N_870);
xnor U1757 (N_1757,N_296,N_230);
nor U1758 (N_1758,N_648,N_494);
nand U1759 (N_1759,N_368,N_402);
and U1760 (N_1760,N_47,N_409);
nand U1761 (N_1761,N_964,N_864);
nand U1762 (N_1762,N_716,N_113);
nand U1763 (N_1763,N_463,N_838);
and U1764 (N_1764,N_488,N_899);
xnor U1765 (N_1765,N_497,N_842);
and U1766 (N_1766,N_690,N_246);
xor U1767 (N_1767,N_729,N_285);
nand U1768 (N_1768,N_261,N_454);
and U1769 (N_1769,N_512,N_133);
nand U1770 (N_1770,N_530,N_267);
nor U1771 (N_1771,N_121,N_662);
xnor U1772 (N_1772,N_611,N_615);
and U1773 (N_1773,N_833,N_369);
or U1774 (N_1774,N_271,N_646);
and U1775 (N_1775,N_82,N_483);
or U1776 (N_1776,N_79,N_333);
xor U1777 (N_1777,N_729,N_711);
and U1778 (N_1778,N_292,N_475);
and U1779 (N_1779,N_890,N_940);
and U1780 (N_1780,N_537,N_930);
and U1781 (N_1781,N_470,N_654);
nand U1782 (N_1782,N_760,N_959);
nor U1783 (N_1783,N_345,N_473);
and U1784 (N_1784,N_148,N_515);
nand U1785 (N_1785,N_695,N_266);
nand U1786 (N_1786,N_438,N_945);
and U1787 (N_1787,N_963,N_164);
and U1788 (N_1788,N_947,N_79);
and U1789 (N_1789,N_397,N_748);
nand U1790 (N_1790,N_828,N_629);
and U1791 (N_1791,N_924,N_769);
nand U1792 (N_1792,N_675,N_712);
nor U1793 (N_1793,N_40,N_73);
nand U1794 (N_1794,N_36,N_910);
nor U1795 (N_1795,N_225,N_470);
or U1796 (N_1796,N_722,N_437);
or U1797 (N_1797,N_232,N_379);
or U1798 (N_1798,N_152,N_836);
and U1799 (N_1799,N_536,N_725);
nand U1800 (N_1800,N_347,N_148);
and U1801 (N_1801,N_614,N_340);
or U1802 (N_1802,N_347,N_417);
or U1803 (N_1803,N_344,N_300);
and U1804 (N_1804,N_391,N_730);
nand U1805 (N_1805,N_267,N_872);
nor U1806 (N_1806,N_456,N_309);
or U1807 (N_1807,N_948,N_584);
and U1808 (N_1808,N_490,N_206);
or U1809 (N_1809,N_99,N_911);
or U1810 (N_1810,N_761,N_315);
nor U1811 (N_1811,N_268,N_346);
nand U1812 (N_1812,N_839,N_901);
and U1813 (N_1813,N_624,N_833);
nand U1814 (N_1814,N_298,N_79);
nand U1815 (N_1815,N_583,N_4);
and U1816 (N_1816,N_950,N_109);
or U1817 (N_1817,N_769,N_700);
nor U1818 (N_1818,N_820,N_946);
and U1819 (N_1819,N_852,N_194);
and U1820 (N_1820,N_57,N_397);
nand U1821 (N_1821,N_932,N_446);
and U1822 (N_1822,N_677,N_223);
nand U1823 (N_1823,N_234,N_672);
and U1824 (N_1824,N_613,N_586);
and U1825 (N_1825,N_431,N_395);
nor U1826 (N_1826,N_413,N_57);
nor U1827 (N_1827,N_128,N_216);
nand U1828 (N_1828,N_430,N_52);
or U1829 (N_1829,N_644,N_773);
nor U1830 (N_1830,N_51,N_615);
nand U1831 (N_1831,N_44,N_20);
nor U1832 (N_1832,N_624,N_527);
nand U1833 (N_1833,N_364,N_776);
or U1834 (N_1834,N_539,N_741);
nor U1835 (N_1835,N_617,N_35);
nor U1836 (N_1836,N_437,N_173);
xnor U1837 (N_1837,N_359,N_340);
and U1838 (N_1838,N_788,N_112);
nand U1839 (N_1839,N_354,N_566);
xor U1840 (N_1840,N_696,N_186);
nor U1841 (N_1841,N_187,N_285);
nand U1842 (N_1842,N_279,N_388);
nand U1843 (N_1843,N_604,N_610);
nand U1844 (N_1844,N_378,N_614);
or U1845 (N_1845,N_870,N_620);
and U1846 (N_1846,N_810,N_720);
nand U1847 (N_1847,N_375,N_664);
or U1848 (N_1848,N_816,N_476);
and U1849 (N_1849,N_762,N_915);
or U1850 (N_1850,N_117,N_323);
nor U1851 (N_1851,N_788,N_286);
xor U1852 (N_1852,N_756,N_842);
and U1853 (N_1853,N_701,N_734);
nand U1854 (N_1854,N_366,N_494);
or U1855 (N_1855,N_837,N_826);
nor U1856 (N_1856,N_610,N_575);
or U1857 (N_1857,N_278,N_688);
nor U1858 (N_1858,N_704,N_499);
and U1859 (N_1859,N_240,N_407);
and U1860 (N_1860,N_496,N_849);
and U1861 (N_1861,N_995,N_852);
and U1862 (N_1862,N_324,N_753);
nor U1863 (N_1863,N_487,N_854);
and U1864 (N_1864,N_21,N_645);
xnor U1865 (N_1865,N_684,N_404);
or U1866 (N_1866,N_527,N_410);
nor U1867 (N_1867,N_637,N_26);
nor U1868 (N_1868,N_49,N_581);
or U1869 (N_1869,N_648,N_508);
nor U1870 (N_1870,N_919,N_607);
or U1871 (N_1871,N_11,N_163);
and U1872 (N_1872,N_777,N_801);
nor U1873 (N_1873,N_64,N_706);
nor U1874 (N_1874,N_572,N_354);
nand U1875 (N_1875,N_355,N_206);
and U1876 (N_1876,N_949,N_594);
nor U1877 (N_1877,N_779,N_385);
nand U1878 (N_1878,N_582,N_417);
and U1879 (N_1879,N_155,N_394);
or U1880 (N_1880,N_499,N_369);
nor U1881 (N_1881,N_882,N_213);
nand U1882 (N_1882,N_250,N_164);
or U1883 (N_1883,N_721,N_804);
nor U1884 (N_1884,N_957,N_430);
and U1885 (N_1885,N_244,N_626);
and U1886 (N_1886,N_908,N_486);
nor U1887 (N_1887,N_175,N_808);
nor U1888 (N_1888,N_686,N_442);
nor U1889 (N_1889,N_155,N_654);
or U1890 (N_1890,N_845,N_151);
or U1891 (N_1891,N_346,N_392);
nor U1892 (N_1892,N_980,N_869);
or U1893 (N_1893,N_707,N_995);
or U1894 (N_1894,N_803,N_122);
nor U1895 (N_1895,N_797,N_46);
or U1896 (N_1896,N_756,N_433);
nor U1897 (N_1897,N_445,N_602);
and U1898 (N_1898,N_802,N_845);
nor U1899 (N_1899,N_367,N_855);
or U1900 (N_1900,N_863,N_818);
nand U1901 (N_1901,N_809,N_920);
or U1902 (N_1902,N_608,N_50);
and U1903 (N_1903,N_582,N_624);
nand U1904 (N_1904,N_108,N_810);
or U1905 (N_1905,N_422,N_590);
or U1906 (N_1906,N_272,N_558);
or U1907 (N_1907,N_211,N_990);
nor U1908 (N_1908,N_966,N_571);
and U1909 (N_1909,N_947,N_293);
or U1910 (N_1910,N_836,N_508);
nand U1911 (N_1911,N_358,N_138);
nand U1912 (N_1912,N_78,N_939);
xnor U1913 (N_1913,N_545,N_581);
nand U1914 (N_1914,N_620,N_306);
nor U1915 (N_1915,N_13,N_230);
and U1916 (N_1916,N_456,N_570);
and U1917 (N_1917,N_158,N_845);
and U1918 (N_1918,N_333,N_244);
or U1919 (N_1919,N_340,N_716);
or U1920 (N_1920,N_944,N_216);
nor U1921 (N_1921,N_366,N_668);
nand U1922 (N_1922,N_699,N_807);
and U1923 (N_1923,N_927,N_738);
nor U1924 (N_1924,N_661,N_819);
and U1925 (N_1925,N_227,N_659);
nor U1926 (N_1926,N_764,N_385);
nor U1927 (N_1927,N_957,N_938);
and U1928 (N_1928,N_425,N_785);
nand U1929 (N_1929,N_97,N_126);
or U1930 (N_1930,N_838,N_529);
and U1931 (N_1931,N_470,N_569);
nor U1932 (N_1932,N_89,N_507);
or U1933 (N_1933,N_949,N_465);
nand U1934 (N_1934,N_757,N_581);
or U1935 (N_1935,N_420,N_381);
nor U1936 (N_1936,N_849,N_894);
and U1937 (N_1937,N_36,N_927);
and U1938 (N_1938,N_225,N_614);
and U1939 (N_1939,N_49,N_406);
or U1940 (N_1940,N_250,N_546);
or U1941 (N_1941,N_903,N_757);
nor U1942 (N_1942,N_520,N_545);
and U1943 (N_1943,N_746,N_54);
and U1944 (N_1944,N_989,N_479);
nand U1945 (N_1945,N_442,N_201);
or U1946 (N_1946,N_538,N_726);
nor U1947 (N_1947,N_215,N_879);
nand U1948 (N_1948,N_762,N_394);
nor U1949 (N_1949,N_726,N_91);
nand U1950 (N_1950,N_749,N_549);
nor U1951 (N_1951,N_982,N_60);
nor U1952 (N_1952,N_458,N_351);
nor U1953 (N_1953,N_32,N_319);
nand U1954 (N_1954,N_859,N_52);
nand U1955 (N_1955,N_115,N_174);
and U1956 (N_1956,N_586,N_95);
nor U1957 (N_1957,N_925,N_469);
and U1958 (N_1958,N_280,N_755);
nand U1959 (N_1959,N_962,N_791);
nand U1960 (N_1960,N_861,N_634);
nand U1961 (N_1961,N_425,N_109);
or U1962 (N_1962,N_927,N_91);
or U1963 (N_1963,N_463,N_407);
or U1964 (N_1964,N_945,N_677);
nand U1965 (N_1965,N_422,N_112);
or U1966 (N_1966,N_632,N_188);
nor U1967 (N_1967,N_241,N_999);
xor U1968 (N_1968,N_769,N_414);
or U1969 (N_1969,N_961,N_184);
and U1970 (N_1970,N_932,N_367);
nand U1971 (N_1971,N_894,N_252);
nor U1972 (N_1972,N_63,N_719);
or U1973 (N_1973,N_445,N_412);
nand U1974 (N_1974,N_672,N_988);
or U1975 (N_1975,N_20,N_613);
or U1976 (N_1976,N_433,N_596);
or U1977 (N_1977,N_813,N_534);
or U1978 (N_1978,N_943,N_344);
or U1979 (N_1979,N_984,N_812);
and U1980 (N_1980,N_542,N_583);
nand U1981 (N_1981,N_95,N_929);
and U1982 (N_1982,N_985,N_231);
nor U1983 (N_1983,N_628,N_416);
nand U1984 (N_1984,N_730,N_343);
or U1985 (N_1985,N_886,N_775);
nand U1986 (N_1986,N_375,N_3);
or U1987 (N_1987,N_418,N_718);
or U1988 (N_1988,N_566,N_32);
nand U1989 (N_1989,N_996,N_926);
or U1990 (N_1990,N_225,N_802);
or U1991 (N_1991,N_123,N_77);
and U1992 (N_1992,N_223,N_347);
nor U1993 (N_1993,N_27,N_900);
nor U1994 (N_1994,N_123,N_176);
or U1995 (N_1995,N_916,N_370);
nor U1996 (N_1996,N_513,N_975);
or U1997 (N_1997,N_958,N_303);
nand U1998 (N_1998,N_114,N_10);
nand U1999 (N_1999,N_925,N_150);
or U2000 (N_2000,N_1408,N_1350);
or U2001 (N_2001,N_1638,N_1001);
or U2002 (N_2002,N_1454,N_1251);
and U2003 (N_2003,N_1306,N_1129);
nand U2004 (N_2004,N_1246,N_1403);
nand U2005 (N_2005,N_1154,N_1749);
and U2006 (N_2006,N_1823,N_1139);
and U2007 (N_2007,N_1962,N_1833);
or U2008 (N_2008,N_1472,N_1560);
or U2009 (N_2009,N_1898,N_1554);
and U2010 (N_2010,N_1465,N_1121);
nor U2011 (N_2011,N_1343,N_1031);
or U2012 (N_2012,N_1200,N_1353);
nand U2013 (N_2013,N_1889,N_1789);
nor U2014 (N_2014,N_1960,N_1432);
nor U2015 (N_2015,N_1456,N_1892);
nand U2016 (N_2016,N_1376,N_1046);
and U2017 (N_2017,N_1559,N_1097);
and U2018 (N_2018,N_1014,N_1581);
and U2019 (N_2019,N_1997,N_1304);
nor U2020 (N_2020,N_1618,N_1886);
or U2021 (N_2021,N_1224,N_1307);
or U2022 (N_2022,N_1932,N_1363);
and U2023 (N_2023,N_1631,N_1821);
nor U2024 (N_2024,N_1023,N_1923);
nor U2025 (N_2025,N_1634,N_1217);
nor U2026 (N_2026,N_1378,N_1066);
or U2027 (N_2027,N_1776,N_1924);
nand U2028 (N_2028,N_1077,N_1446);
xnor U2029 (N_2029,N_1564,N_1142);
or U2030 (N_2030,N_1820,N_1054);
nand U2031 (N_2031,N_1042,N_1799);
nand U2032 (N_2032,N_1538,N_1872);
nand U2033 (N_2033,N_1991,N_1484);
nor U2034 (N_2034,N_1106,N_1429);
or U2035 (N_2035,N_1040,N_1173);
or U2036 (N_2036,N_1951,N_1431);
or U2037 (N_2037,N_1727,N_1852);
and U2038 (N_2038,N_1632,N_1393);
nand U2039 (N_2039,N_1164,N_1528);
or U2040 (N_2040,N_1627,N_1779);
nor U2041 (N_2041,N_1233,N_1558);
or U2042 (N_2042,N_1733,N_1642);
nand U2043 (N_2043,N_1483,N_1263);
or U2044 (N_2044,N_1152,N_1518);
nor U2045 (N_2045,N_1838,N_1260);
nand U2046 (N_2046,N_1747,N_1442);
and U2047 (N_2047,N_1404,N_1803);
and U2048 (N_2048,N_1970,N_1658);
and U2049 (N_2049,N_1150,N_1875);
nor U2050 (N_2050,N_1525,N_1989);
nand U2051 (N_2051,N_1676,N_1226);
nor U2052 (N_2052,N_1006,N_1594);
nor U2053 (N_2053,N_1252,N_1880);
or U2054 (N_2054,N_1385,N_1271);
and U2055 (N_2055,N_1178,N_1461);
or U2056 (N_2056,N_1993,N_1422);
nor U2057 (N_2057,N_1878,N_1457);
nand U2058 (N_2058,N_1814,N_1496);
nand U2059 (N_2059,N_1505,N_1187);
nor U2060 (N_2060,N_1689,N_1739);
nor U2061 (N_2061,N_1717,N_1633);
nand U2062 (N_2062,N_1563,N_1711);
nand U2063 (N_2063,N_1433,N_1963);
nand U2064 (N_2064,N_1920,N_1944);
or U2065 (N_2065,N_1375,N_1402);
or U2066 (N_2066,N_1613,N_1839);
nor U2067 (N_2067,N_1131,N_1625);
and U2068 (N_2068,N_1188,N_1024);
nor U2069 (N_2069,N_1844,N_1621);
nor U2070 (N_2070,N_1639,N_1225);
and U2071 (N_2071,N_1215,N_1010);
and U2072 (N_2072,N_1041,N_1980);
or U2073 (N_2073,N_1474,N_1718);
and U2074 (N_2074,N_1987,N_1612);
nand U2075 (N_2075,N_1949,N_1245);
nand U2076 (N_2076,N_1545,N_1888);
or U2077 (N_2077,N_1834,N_1339);
nor U2078 (N_2078,N_1262,N_1128);
or U2079 (N_2079,N_1212,N_1331);
and U2080 (N_2080,N_1975,N_1397);
or U2081 (N_2081,N_1818,N_1981);
nand U2082 (N_2082,N_1922,N_1824);
or U2083 (N_2083,N_1382,N_1421);
and U2084 (N_2084,N_1323,N_1943);
nor U2085 (N_2085,N_1760,N_1035);
or U2086 (N_2086,N_1971,N_1598);
or U2087 (N_2087,N_1259,N_1293);
nor U2088 (N_2088,N_1794,N_1517);
or U2089 (N_2089,N_1601,N_1022);
nand U2090 (N_2090,N_1705,N_1316);
nor U2091 (N_2091,N_1591,N_1276);
nor U2092 (N_2092,N_1478,N_1854);
and U2093 (N_2093,N_1935,N_1462);
nand U2094 (N_2094,N_1440,N_1078);
nor U2095 (N_2095,N_1907,N_1074);
or U2096 (N_2096,N_1085,N_1133);
and U2097 (N_2097,N_1374,N_1241);
or U2098 (N_2098,N_1978,N_1681);
nand U2099 (N_2099,N_1902,N_1752);
nand U2100 (N_2100,N_1651,N_1044);
nand U2101 (N_2101,N_1469,N_1290);
nor U2102 (N_2102,N_1955,N_1851);
and U2103 (N_2103,N_1202,N_1027);
nand U2104 (N_2104,N_1561,N_1018);
nand U2105 (N_2105,N_1855,N_1835);
nor U2106 (N_2106,N_1361,N_1029);
or U2107 (N_2107,N_1798,N_1707);
nand U2108 (N_2108,N_1848,N_1118);
nor U2109 (N_2109,N_1593,N_1566);
nand U2110 (N_2110,N_1012,N_1455);
and U2111 (N_2111,N_1911,N_1864);
nor U2112 (N_2112,N_1901,N_1569);
or U2113 (N_2113,N_1883,N_1900);
nor U2114 (N_2114,N_1265,N_1926);
or U2115 (N_2115,N_1751,N_1736);
nor U2116 (N_2116,N_1495,N_1715);
nand U2117 (N_2117,N_1910,N_1028);
nor U2118 (N_2118,N_1586,N_1572);
and U2119 (N_2119,N_1657,N_1829);
nor U2120 (N_2120,N_1135,N_1624);
nor U2121 (N_2121,N_1573,N_1275);
or U2122 (N_2122,N_1600,N_1415);
and U2123 (N_2123,N_1849,N_1744);
nor U2124 (N_2124,N_1296,N_1994);
or U2125 (N_2125,N_1103,N_1716);
and U2126 (N_2126,N_1510,N_1948);
or U2127 (N_2127,N_1746,N_1666);
and U2128 (N_2128,N_1940,N_1592);
or U2129 (N_2129,N_1753,N_1567);
or U2130 (N_2130,N_1800,N_1430);
nand U2131 (N_2131,N_1201,N_1058);
nor U2132 (N_2132,N_1206,N_1072);
or U2133 (N_2133,N_1614,N_1395);
or U2134 (N_2134,N_1847,N_1207);
nor U2135 (N_2135,N_1804,N_1936);
nand U2136 (N_2136,N_1303,N_1730);
or U2137 (N_2137,N_1856,N_1328);
and U2138 (N_2138,N_1386,N_1368);
or U2139 (N_2139,N_1050,N_1372);
nor U2140 (N_2140,N_1273,N_1391);
nor U2141 (N_2141,N_1211,N_1373);
nand U2142 (N_2142,N_1729,N_1180);
or U2143 (N_2143,N_1623,N_1228);
nor U2144 (N_2144,N_1222,N_1837);
nor U2145 (N_2145,N_1700,N_1933);
or U2146 (N_2146,N_1289,N_1258);
and U2147 (N_2147,N_1861,N_1967);
xor U2148 (N_2148,N_1037,N_1537);
and U2149 (N_2149,N_1846,N_1390);
nor U2150 (N_2150,N_1604,N_1866);
nor U2151 (N_2151,N_1620,N_1370);
and U2152 (N_2152,N_1874,N_1655);
and U2153 (N_2153,N_1519,N_1908);
or U2154 (N_2154,N_1722,N_1611);
or U2155 (N_2155,N_1792,N_1570);
xor U2156 (N_2156,N_1341,N_1702);
nor U2157 (N_2157,N_1137,N_1223);
nor U2158 (N_2158,N_1953,N_1025);
nor U2159 (N_2159,N_1253,N_1919);
or U2160 (N_2160,N_1492,N_1269);
nor U2161 (N_2161,N_1055,N_1915);
and U2162 (N_2162,N_1762,N_1205);
or U2163 (N_2163,N_1310,N_1358);
nand U2164 (N_2164,N_1629,N_1141);
and U2165 (N_2165,N_1644,N_1239);
or U2166 (N_2166,N_1366,N_1785);
and U2167 (N_2167,N_1236,N_1797);
nand U2168 (N_2168,N_1802,N_1190);
and U2169 (N_2169,N_1539,N_1218);
nor U2170 (N_2170,N_1016,N_1931);
or U2171 (N_2171,N_1448,N_1683);
nand U2172 (N_2172,N_1983,N_1556);
and U2173 (N_2173,N_1314,N_1136);
xor U2174 (N_2174,N_1708,N_1551);
and U2175 (N_2175,N_1266,N_1562);
or U2176 (N_2176,N_1487,N_1053);
and U2177 (N_2177,N_1536,N_1870);
and U2178 (N_2178,N_1759,N_1713);
or U2179 (N_2179,N_1979,N_1862);
nor U2180 (N_2180,N_1523,N_1858);
nor U2181 (N_2181,N_1512,N_1111);
nand U2182 (N_2182,N_1688,N_1740);
or U2183 (N_2183,N_1232,N_1966);
or U2184 (N_2184,N_1184,N_1147);
or U2185 (N_2185,N_1685,N_1039);
nand U2186 (N_2186,N_1819,N_1895);
or U2187 (N_2187,N_1256,N_1294);
nor U2188 (N_2188,N_1768,N_1687);
and U2189 (N_2189,N_1489,N_1434);
nand U2190 (N_2190,N_1565,N_1104);
xnor U2191 (N_2191,N_1175,N_1196);
or U2192 (N_2192,N_1941,N_1126);
nand U2193 (N_2193,N_1897,N_1257);
and U2194 (N_2194,N_1764,N_1143);
nor U2195 (N_2195,N_1083,N_1588);
nand U2196 (N_2196,N_1977,N_1105);
nand U2197 (N_2197,N_1669,N_1845);
nor U2198 (N_2198,N_1396,N_1937);
and U2199 (N_2199,N_1065,N_1783);
nor U2200 (N_2200,N_1369,N_1480);
nand U2201 (N_2201,N_1628,N_1805);
nand U2202 (N_2202,N_1925,N_1221);
nor U2203 (N_2203,N_1720,N_1984);
nand U2204 (N_2204,N_1460,N_1243);
or U2205 (N_2205,N_1424,N_1284);
nor U2206 (N_2206,N_1318,N_1299);
or U2207 (N_2207,N_1905,N_1344);
and U2208 (N_2208,N_1507,N_1313);
and U2209 (N_2209,N_1521,N_1287);
and U2210 (N_2210,N_1153,N_1686);
nor U2211 (N_2211,N_1169,N_1504);
or U2212 (N_2212,N_1985,N_1167);
nand U2213 (N_2213,N_1636,N_1511);
nand U2214 (N_2214,N_1815,N_1927);
and U2215 (N_2215,N_1635,N_1494);
or U2216 (N_2216,N_1787,N_1671);
nor U2217 (N_2217,N_1930,N_1362);
nor U2218 (N_2218,N_1876,N_1120);
and U2219 (N_2219,N_1181,N_1399);
nand U2220 (N_2220,N_1697,N_1264);
nand U2221 (N_2221,N_1324,N_1019);
and U2222 (N_2222,N_1615,N_1070);
nor U2223 (N_2223,N_1502,N_1577);
nor U2224 (N_2224,N_1282,N_1379);
or U2225 (N_2225,N_1826,N_1364);
nand U2226 (N_2226,N_1351,N_1807);
nand U2227 (N_2227,N_1295,N_1367);
nand U2228 (N_2228,N_1812,N_1542);
xnor U2229 (N_2229,N_1830,N_1437);
nand U2230 (N_2230,N_1348,N_1738);
and U2231 (N_2231,N_1513,N_1850);
nor U2232 (N_2232,N_1904,N_1360);
and U2233 (N_2233,N_1400,N_1587);
and U2234 (N_2234,N_1912,N_1509);
or U2235 (N_2235,N_1132,N_1485);
nor U2236 (N_2236,N_1842,N_1896);
or U2237 (N_2237,N_1388,N_1235);
and U2238 (N_2238,N_1068,N_1667);
nand U2239 (N_2239,N_1359,N_1801);
nand U2240 (N_2240,N_1300,N_1267);
or U2241 (N_2241,N_1859,N_1109);
nor U2242 (N_2242,N_1832,N_1113);
nor U2243 (N_2243,N_1630,N_1534);
and U2244 (N_2244,N_1772,N_1159);
or U2245 (N_2245,N_1988,N_1192);
or U2246 (N_2246,N_1464,N_1062);
nor U2247 (N_2247,N_1092,N_1813);
or U2248 (N_2248,N_1420,N_1795);
nand U2249 (N_2249,N_1398,N_1721);
or U2250 (N_2250,N_1954,N_1122);
or U2251 (N_2251,N_1654,N_1384);
or U2252 (N_2252,N_1706,N_1516);
and U2253 (N_2253,N_1439,N_1728);
and U2254 (N_2254,N_1426,N_1419);
and U2255 (N_2255,N_1491,N_1547);
or U2256 (N_2256,N_1166,N_1774);
nor U2257 (N_2257,N_1088,N_1352);
nor U2258 (N_2258,N_1034,N_1081);
xor U2259 (N_2259,N_1288,N_1575);
or U2260 (N_2260,N_1679,N_1840);
and U2261 (N_2261,N_1349,N_1755);
and U2262 (N_2262,N_1127,N_1186);
nand U2263 (N_2263,N_1501,N_1191);
nor U2264 (N_2264,N_1336,N_1499);
nor U2265 (N_2265,N_1394,N_1096);
nand U2266 (N_2266,N_1021,N_1475);
nand U2267 (N_2267,N_1580,N_1769);
and U2268 (N_2268,N_1094,N_1436);
or U2269 (N_2269,N_1292,N_1914);
nor U2270 (N_2270,N_1865,N_1605);
nand U2271 (N_2271,N_1778,N_1999);
nand U2272 (N_2272,N_1003,N_1959);
nor U2273 (N_2273,N_1043,N_1882);
nor U2274 (N_2274,N_1274,N_1045);
or U2275 (N_2275,N_1603,N_1757);
nand U2276 (N_2276,N_1737,N_1449);
and U2277 (N_2277,N_1145,N_1441);
or U2278 (N_2278,N_1405,N_1668);
nor U2279 (N_2279,N_1725,N_1409);
nand U2280 (N_2280,N_1986,N_1061);
nor U2281 (N_2281,N_1881,N_1506);
and U2282 (N_2282,N_1766,N_1788);
or U2283 (N_2283,N_1095,N_1330);
nor U2284 (N_2284,N_1112,N_1146);
or U2285 (N_2285,N_1298,N_1057);
and U2286 (N_2286,N_1650,N_1281);
nand U2287 (N_2287,N_1622,N_1087);
and U2288 (N_2288,N_1038,N_1197);
nor U2289 (N_2289,N_1459,N_1584);
and U2290 (N_2290,N_1672,N_1140);
nor U2291 (N_2291,N_1522,N_1945);
or U2292 (N_2292,N_1515,N_1806);
nor U2293 (N_2293,N_1340,N_1108);
nor U2294 (N_2294,N_1007,N_1822);
nor U2295 (N_2295,N_1890,N_1110);
and U2296 (N_2296,N_1756,N_1675);
and U2297 (N_2297,N_1020,N_1860);
and U2298 (N_2298,N_1972,N_1056);
nand U2299 (N_2299,N_1952,N_1950);
nor U2300 (N_2300,N_1148,N_1315);
or U2301 (N_2301,N_1743,N_1790);
nor U2302 (N_2302,N_1219,N_1312);
nor U2303 (N_2303,N_1481,N_1548);
nor U2304 (N_2304,N_1453,N_1445);
and U2305 (N_2305,N_1503,N_1526);
xnor U2306 (N_2306,N_1867,N_1447);
or U2307 (N_2307,N_1242,N_1701);
or U2308 (N_2308,N_1237,N_1013);
nand U2309 (N_2309,N_1982,N_1906);
xor U2310 (N_2310,N_1036,N_1529);
or U2311 (N_2311,N_1745,N_1249);
or U2312 (N_2312,N_1199,N_1115);
nor U2313 (N_2313,N_1231,N_1125);
and U2314 (N_2314,N_1723,N_1338);
and U2315 (N_2315,N_1609,N_1144);
and U2316 (N_2316,N_1387,N_1765);
nor U2317 (N_2317,N_1585,N_1791);
or U2318 (N_2318,N_1064,N_1268);
nor U2319 (N_2319,N_1060,N_1073);
nand U2320 (N_2320,N_1117,N_1377);
nand U2321 (N_2321,N_1048,N_1332);
or U2322 (N_2322,N_1270,N_1786);
nor U2323 (N_2323,N_1011,N_1968);
nor U2324 (N_2324,N_1877,N_1535);
nor U2325 (N_2325,N_1468,N_1508);
nor U2326 (N_2326,N_1810,N_1780);
and U2327 (N_2327,N_1541,N_1008);
nor U2328 (N_2328,N_1283,N_1557);
nand U2329 (N_2329,N_1401,N_1767);
nand U2330 (N_2330,N_1182,N_1894);
nor U2331 (N_2331,N_1413,N_1450);
or U2332 (N_2332,N_1498,N_1607);
or U2333 (N_2333,N_1857,N_1887);
and U2334 (N_2334,N_1724,N_1520);
nand U2335 (N_2335,N_1305,N_1076);
or U2336 (N_2336,N_1356,N_1107);
and U2337 (N_2337,N_1185,N_1544);
or U2338 (N_2338,N_1793,N_1082);
nand U2339 (N_2339,N_1208,N_1712);
or U2340 (N_2340,N_1345,N_1347);
nand U2341 (N_2341,N_1261,N_1909);
and U2342 (N_2342,N_1406,N_1130);
nand U2343 (N_2343,N_1868,N_1086);
or U2344 (N_2344,N_1916,N_1194);
or U2345 (N_2345,N_1354,N_1254);
xor U2346 (N_2346,N_1546,N_1486);
nand U2347 (N_2347,N_1719,N_1781);
nand U2348 (N_2348,N_1162,N_1337);
and U2349 (N_2349,N_1342,N_1663);
or U2350 (N_2350,N_1407,N_1165);
or U2351 (N_2351,N_1903,N_1230);
and U2352 (N_2352,N_1410,N_1100);
nand U2353 (N_2353,N_1665,N_1873);
nand U2354 (N_2354,N_1583,N_1365);
nand U2355 (N_2355,N_1383,N_1831);
nand U2356 (N_2356,N_1051,N_1928);
nand U2357 (N_2357,N_1714,N_1099);
and U2358 (N_2358,N_1423,N_1380);
or U2359 (N_2359,N_1741,N_1451);
and U2360 (N_2360,N_1578,N_1661);
nand U2361 (N_2361,N_1311,N_1158);
nor U2362 (N_2362,N_1549,N_1552);
and U2363 (N_2363,N_1280,N_1255);
nor U2364 (N_2364,N_1240,N_1617);
nor U2365 (N_2365,N_1809,N_1015);
nor U2366 (N_2366,N_1005,N_1698);
nand U2367 (N_2367,N_1335,N_1616);
or U2368 (N_2368,N_1470,N_1673);
nand U2369 (N_2369,N_1428,N_1637);
and U2370 (N_2370,N_1381,N_1091);
and U2371 (N_2371,N_1947,N_1893);
nand U2372 (N_2372,N_1179,N_1550);
nand U2373 (N_2373,N_1033,N_1471);
nor U2374 (N_2374,N_1695,N_1773);
or U2375 (N_2375,N_1116,N_1193);
and U2376 (N_2376,N_1004,N_1684);
nor U2377 (N_2377,N_1956,N_1411);
and U2378 (N_2378,N_1782,N_1836);
and U2379 (N_2379,N_1063,N_1704);
or U2380 (N_2380,N_1319,N_1899);
nand U2381 (N_2381,N_1102,N_1524);
nand U2382 (N_2382,N_1477,N_1589);
and U2383 (N_2383,N_1995,N_1748);
and U2384 (N_2384,N_1841,N_1731);
or U2385 (N_2385,N_1286,N_1216);
nor U2386 (N_2386,N_1879,N_1168);
nand U2387 (N_2387,N_1134,N_1458);
and U2388 (N_2388,N_1238,N_1244);
nor U2389 (N_2389,N_1693,N_1047);
or U2390 (N_2390,N_1418,N_1427);
or U2391 (N_2391,N_1690,N_1101);
nand U2392 (N_2392,N_1827,N_1250);
and U2393 (N_2393,N_1160,N_1079);
nand U2394 (N_2394,N_1843,N_1417);
and U2395 (N_2395,N_1177,N_1530);
or U2396 (N_2396,N_1123,N_1750);
and U2397 (N_2397,N_1579,N_1389);
and U2398 (N_2398,N_1770,N_1302);
nand U2399 (N_2399,N_1692,N_1098);
or U2400 (N_2400,N_1514,N_1229);
nor U2401 (N_2401,N_1998,N_1161);
or U2402 (N_2402,N_1533,N_1853);
or U2403 (N_2403,N_1568,N_1476);
xnor U2404 (N_2404,N_1452,N_1151);
nand U2405 (N_2405,N_1277,N_1149);
nor U2406 (N_2406,N_1754,N_1643);
nor U2407 (N_2407,N_1964,N_1291);
nand U2408 (N_2408,N_1974,N_1195);
or U2409 (N_2409,N_1976,N_1156);
or U2410 (N_2410,N_1002,N_1946);
nand U2411 (N_2411,N_1540,N_1574);
nor U2412 (N_2412,N_1710,N_1597);
nand U2413 (N_2413,N_1080,N_1346);
and U2414 (N_2414,N_1114,N_1863);
nand U2415 (N_2415,N_1334,N_1049);
nand U2416 (N_2416,N_1775,N_1913);
or U2417 (N_2417,N_1326,N_1699);
xor U2418 (N_2418,N_1606,N_1414);
and U2419 (N_2419,N_1957,N_1596);
or U2420 (N_2420,N_1071,N_1412);
nand U2421 (N_2421,N_1308,N_1272);
nand U2422 (N_2422,N_1325,N_1301);
or U2423 (N_2423,N_1248,N_1059);
nand U2424 (N_2424,N_1119,N_1482);
or U2425 (N_2425,N_1828,N_1758);
and U2426 (N_2426,N_1327,N_1884);
or U2427 (N_2427,N_1198,N_1640);
nand U2428 (N_2428,N_1392,N_1320);
nand U2429 (N_2429,N_1210,N_1543);
and U2430 (N_2430,N_1742,N_1734);
or U2431 (N_2431,N_1648,N_1463);
nand U2432 (N_2432,N_1996,N_1234);
nand U2433 (N_2433,N_1816,N_1726);
and U2434 (N_2434,N_1466,N_1576);
and U2435 (N_2435,N_1796,N_1680);
and U2436 (N_2436,N_1204,N_1647);
nand U2437 (N_2437,N_1093,N_1488);
nor U2438 (N_2438,N_1602,N_1333);
nand U2439 (N_2439,N_1652,N_1247);
or U2440 (N_2440,N_1553,N_1934);
nor U2441 (N_2441,N_1732,N_1674);
and U2442 (N_2442,N_1958,N_1473);
nor U2443 (N_2443,N_1026,N_1992);
nor U2444 (N_2444,N_1000,N_1209);
or U2445 (N_2445,N_1662,N_1664);
xor U2446 (N_2446,N_1825,N_1917);
nand U2447 (N_2447,N_1493,N_1084);
nand U2448 (N_2448,N_1531,N_1645);
or U2449 (N_2449,N_1355,N_1694);
or U2450 (N_2450,N_1763,N_1891);
nor U2451 (N_2451,N_1443,N_1297);
or U2452 (N_2452,N_1869,N_1817);
and U2453 (N_2453,N_1075,N_1171);
and U2454 (N_2454,N_1918,N_1961);
nor U2455 (N_2455,N_1490,N_1973);
nand U2456 (N_2456,N_1709,N_1808);
or U2457 (N_2457,N_1599,N_1278);
or U2458 (N_2458,N_1321,N_1641);
and U2459 (N_2459,N_1682,N_1532);
and U2460 (N_2460,N_1582,N_1183);
nor U2461 (N_2461,N_1811,N_1595);
and U2462 (N_2462,N_1571,N_1626);
nor U2463 (N_2463,N_1435,N_1444);
and U2464 (N_2464,N_1220,N_1660);
nor U2465 (N_2465,N_1703,N_1656);
nor U2466 (N_2466,N_1357,N_1214);
or U2467 (N_2467,N_1610,N_1649);
nand U2468 (N_2468,N_1213,N_1138);
or U2469 (N_2469,N_1784,N_1965);
and U2470 (N_2470,N_1309,N_1555);
or U2471 (N_2471,N_1939,N_1329);
nor U2472 (N_2472,N_1317,N_1017);
or U2473 (N_2473,N_1172,N_1157);
nor U2474 (N_2474,N_1942,N_1438);
or U2475 (N_2475,N_1425,N_1069);
nor U2476 (N_2476,N_1590,N_1678);
or U2477 (N_2477,N_1163,N_1990);
nand U2478 (N_2478,N_1170,N_1176);
or U2479 (N_2479,N_1090,N_1691);
or U2480 (N_2480,N_1969,N_1777);
or U2481 (N_2481,N_1527,N_1608);
nand U2482 (N_2482,N_1619,N_1761);
or U2483 (N_2483,N_1871,N_1771);
nand U2484 (N_2484,N_1659,N_1416);
and U2485 (N_2485,N_1670,N_1067);
and U2486 (N_2486,N_1696,N_1646);
nand U2487 (N_2487,N_1371,N_1322);
or U2488 (N_2488,N_1497,N_1279);
and U2489 (N_2489,N_1500,N_1009);
nand U2490 (N_2490,N_1052,N_1124);
nand U2491 (N_2491,N_1929,N_1735);
nand U2492 (N_2492,N_1479,N_1467);
nand U2493 (N_2493,N_1203,N_1938);
or U2494 (N_2494,N_1677,N_1285);
xnor U2495 (N_2495,N_1155,N_1174);
and U2496 (N_2496,N_1089,N_1032);
nand U2497 (N_2497,N_1653,N_1227);
and U2498 (N_2498,N_1030,N_1189);
or U2499 (N_2499,N_1921,N_1885);
or U2500 (N_2500,N_1874,N_1225);
nor U2501 (N_2501,N_1724,N_1494);
nor U2502 (N_2502,N_1391,N_1061);
nor U2503 (N_2503,N_1833,N_1029);
nor U2504 (N_2504,N_1095,N_1164);
and U2505 (N_2505,N_1996,N_1806);
nor U2506 (N_2506,N_1668,N_1040);
or U2507 (N_2507,N_1279,N_1087);
nand U2508 (N_2508,N_1886,N_1061);
xnor U2509 (N_2509,N_1807,N_1501);
or U2510 (N_2510,N_1404,N_1025);
or U2511 (N_2511,N_1713,N_1613);
nor U2512 (N_2512,N_1674,N_1740);
nand U2513 (N_2513,N_1396,N_1421);
and U2514 (N_2514,N_1187,N_1487);
nor U2515 (N_2515,N_1386,N_1284);
or U2516 (N_2516,N_1391,N_1017);
nor U2517 (N_2517,N_1510,N_1164);
nand U2518 (N_2518,N_1913,N_1892);
nor U2519 (N_2519,N_1198,N_1240);
nand U2520 (N_2520,N_1561,N_1895);
or U2521 (N_2521,N_1956,N_1959);
nand U2522 (N_2522,N_1043,N_1438);
and U2523 (N_2523,N_1097,N_1478);
or U2524 (N_2524,N_1990,N_1010);
or U2525 (N_2525,N_1265,N_1229);
nor U2526 (N_2526,N_1133,N_1433);
nor U2527 (N_2527,N_1271,N_1540);
or U2528 (N_2528,N_1652,N_1497);
or U2529 (N_2529,N_1086,N_1303);
nor U2530 (N_2530,N_1271,N_1494);
or U2531 (N_2531,N_1827,N_1739);
xnor U2532 (N_2532,N_1874,N_1344);
nor U2533 (N_2533,N_1725,N_1733);
or U2534 (N_2534,N_1074,N_1683);
or U2535 (N_2535,N_1656,N_1175);
or U2536 (N_2536,N_1509,N_1057);
nand U2537 (N_2537,N_1224,N_1243);
nand U2538 (N_2538,N_1714,N_1319);
nand U2539 (N_2539,N_1198,N_1954);
nor U2540 (N_2540,N_1122,N_1341);
nor U2541 (N_2541,N_1681,N_1760);
nor U2542 (N_2542,N_1149,N_1358);
nor U2543 (N_2543,N_1843,N_1321);
or U2544 (N_2544,N_1891,N_1741);
xnor U2545 (N_2545,N_1331,N_1948);
and U2546 (N_2546,N_1492,N_1135);
nor U2547 (N_2547,N_1230,N_1820);
or U2548 (N_2548,N_1738,N_1146);
nand U2549 (N_2549,N_1668,N_1529);
and U2550 (N_2550,N_1088,N_1481);
or U2551 (N_2551,N_1701,N_1118);
and U2552 (N_2552,N_1391,N_1675);
or U2553 (N_2553,N_1425,N_1308);
nor U2554 (N_2554,N_1168,N_1372);
or U2555 (N_2555,N_1149,N_1116);
and U2556 (N_2556,N_1583,N_1349);
or U2557 (N_2557,N_1756,N_1436);
nand U2558 (N_2558,N_1523,N_1857);
and U2559 (N_2559,N_1611,N_1711);
and U2560 (N_2560,N_1378,N_1272);
nor U2561 (N_2561,N_1499,N_1512);
or U2562 (N_2562,N_1308,N_1686);
or U2563 (N_2563,N_1740,N_1845);
nand U2564 (N_2564,N_1902,N_1747);
and U2565 (N_2565,N_1093,N_1391);
or U2566 (N_2566,N_1900,N_1943);
nor U2567 (N_2567,N_1419,N_1630);
nor U2568 (N_2568,N_1875,N_1275);
nand U2569 (N_2569,N_1780,N_1762);
or U2570 (N_2570,N_1729,N_1348);
nand U2571 (N_2571,N_1730,N_1657);
or U2572 (N_2572,N_1014,N_1482);
and U2573 (N_2573,N_1403,N_1556);
or U2574 (N_2574,N_1190,N_1305);
and U2575 (N_2575,N_1008,N_1464);
nand U2576 (N_2576,N_1811,N_1194);
nor U2577 (N_2577,N_1344,N_1223);
nor U2578 (N_2578,N_1523,N_1713);
and U2579 (N_2579,N_1659,N_1090);
or U2580 (N_2580,N_1346,N_1228);
nand U2581 (N_2581,N_1457,N_1251);
nand U2582 (N_2582,N_1828,N_1069);
xor U2583 (N_2583,N_1582,N_1681);
or U2584 (N_2584,N_1942,N_1683);
nand U2585 (N_2585,N_1429,N_1895);
and U2586 (N_2586,N_1666,N_1452);
nand U2587 (N_2587,N_1586,N_1621);
or U2588 (N_2588,N_1456,N_1034);
and U2589 (N_2589,N_1908,N_1599);
nand U2590 (N_2590,N_1301,N_1140);
or U2591 (N_2591,N_1603,N_1047);
or U2592 (N_2592,N_1357,N_1586);
nor U2593 (N_2593,N_1101,N_1311);
and U2594 (N_2594,N_1856,N_1683);
or U2595 (N_2595,N_1605,N_1561);
or U2596 (N_2596,N_1165,N_1993);
nand U2597 (N_2597,N_1957,N_1707);
nor U2598 (N_2598,N_1247,N_1634);
nand U2599 (N_2599,N_1863,N_1932);
nand U2600 (N_2600,N_1669,N_1071);
nor U2601 (N_2601,N_1886,N_1595);
nand U2602 (N_2602,N_1209,N_1855);
xnor U2603 (N_2603,N_1896,N_1464);
nand U2604 (N_2604,N_1483,N_1654);
nand U2605 (N_2605,N_1670,N_1190);
nor U2606 (N_2606,N_1974,N_1105);
or U2607 (N_2607,N_1912,N_1334);
and U2608 (N_2608,N_1983,N_1840);
nand U2609 (N_2609,N_1825,N_1908);
nor U2610 (N_2610,N_1130,N_1758);
and U2611 (N_2611,N_1932,N_1426);
nand U2612 (N_2612,N_1138,N_1024);
or U2613 (N_2613,N_1632,N_1978);
xor U2614 (N_2614,N_1028,N_1950);
or U2615 (N_2615,N_1948,N_1514);
nor U2616 (N_2616,N_1508,N_1149);
nand U2617 (N_2617,N_1355,N_1152);
nand U2618 (N_2618,N_1340,N_1256);
or U2619 (N_2619,N_1088,N_1290);
and U2620 (N_2620,N_1659,N_1572);
and U2621 (N_2621,N_1821,N_1651);
nor U2622 (N_2622,N_1590,N_1266);
or U2623 (N_2623,N_1299,N_1581);
or U2624 (N_2624,N_1100,N_1135);
nor U2625 (N_2625,N_1889,N_1270);
or U2626 (N_2626,N_1586,N_1477);
nand U2627 (N_2627,N_1107,N_1405);
and U2628 (N_2628,N_1607,N_1078);
and U2629 (N_2629,N_1936,N_1821);
nor U2630 (N_2630,N_1531,N_1603);
nand U2631 (N_2631,N_1425,N_1229);
and U2632 (N_2632,N_1515,N_1211);
or U2633 (N_2633,N_1002,N_1472);
nand U2634 (N_2634,N_1522,N_1372);
or U2635 (N_2635,N_1179,N_1753);
and U2636 (N_2636,N_1985,N_1703);
nor U2637 (N_2637,N_1120,N_1221);
nor U2638 (N_2638,N_1795,N_1323);
and U2639 (N_2639,N_1694,N_1130);
nand U2640 (N_2640,N_1775,N_1143);
and U2641 (N_2641,N_1159,N_1239);
and U2642 (N_2642,N_1682,N_1902);
or U2643 (N_2643,N_1901,N_1933);
nor U2644 (N_2644,N_1051,N_1544);
and U2645 (N_2645,N_1249,N_1850);
or U2646 (N_2646,N_1175,N_1702);
and U2647 (N_2647,N_1652,N_1826);
or U2648 (N_2648,N_1116,N_1517);
nand U2649 (N_2649,N_1762,N_1814);
nor U2650 (N_2650,N_1507,N_1360);
nand U2651 (N_2651,N_1078,N_1549);
nand U2652 (N_2652,N_1572,N_1412);
or U2653 (N_2653,N_1249,N_1252);
or U2654 (N_2654,N_1834,N_1180);
or U2655 (N_2655,N_1458,N_1294);
nand U2656 (N_2656,N_1106,N_1153);
nor U2657 (N_2657,N_1116,N_1061);
nor U2658 (N_2658,N_1480,N_1947);
or U2659 (N_2659,N_1609,N_1708);
nand U2660 (N_2660,N_1068,N_1064);
nand U2661 (N_2661,N_1701,N_1273);
or U2662 (N_2662,N_1103,N_1360);
nor U2663 (N_2663,N_1347,N_1216);
and U2664 (N_2664,N_1868,N_1719);
and U2665 (N_2665,N_1209,N_1003);
nand U2666 (N_2666,N_1279,N_1032);
nand U2667 (N_2667,N_1941,N_1672);
nor U2668 (N_2668,N_1227,N_1437);
or U2669 (N_2669,N_1645,N_1909);
nor U2670 (N_2670,N_1277,N_1335);
nand U2671 (N_2671,N_1164,N_1912);
or U2672 (N_2672,N_1334,N_1276);
nand U2673 (N_2673,N_1307,N_1420);
or U2674 (N_2674,N_1385,N_1630);
or U2675 (N_2675,N_1533,N_1505);
nand U2676 (N_2676,N_1902,N_1272);
nor U2677 (N_2677,N_1677,N_1133);
and U2678 (N_2678,N_1763,N_1548);
or U2679 (N_2679,N_1745,N_1057);
nor U2680 (N_2680,N_1159,N_1743);
and U2681 (N_2681,N_1553,N_1618);
and U2682 (N_2682,N_1285,N_1688);
nand U2683 (N_2683,N_1380,N_1103);
nand U2684 (N_2684,N_1693,N_1419);
or U2685 (N_2685,N_1650,N_1921);
or U2686 (N_2686,N_1343,N_1856);
and U2687 (N_2687,N_1051,N_1945);
nand U2688 (N_2688,N_1198,N_1436);
and U2689 (N_2689,N_1928,N_1705);
nor U2690 (N_2690,N_1844,N_1570);
or U2691 (N_2691,N_1507,N_1891);
nor U2692 (N_2692,N_1146,N_1419);
nor U2693 (N_2693,N_1922,N_1366);
nand U2694 (N_2694,N_1470,N_1066);
nand U2695 (N_2695,N_1672,N_1805);
or U2696 (N_2696,N_1161,N_1188);
nor U2697 (N_2697,N_1021,N_1133);
nor U2698 (N_2698,N_1177,N_1692);
nand U2699 (N_2699,N_1748,N_1109);
and U2700 (N_2700,N_1722,N_1252);
nand U2701 (N_2701,N_1951,N_1695);
or U2702 (N_2702,N_1087,N_1600);
or U2703 (N_2703,N_1058,N_1272);
or U2704 (N_2704,N_1201,N_1909);
and U2705 (N_2705,N_1710,N_1553);
nor U2706 (N_2706,N_1718,N_1209);
or U2707 (N_2707,N_1872,N_1374);
nor U2708 (N_2708,N_1218,N_1462);
and U2709 (N_2709,N_1101,N_1061);
and U2710 (N_2710,N_1025,N_1153);
or U2711 (N_2711,N_1531,N_1244);
or U2712 (N_2712,N_1141,N_1512);
or U2713 (N_2713,N_1584,N_1822);
nand U2714 (N_2714,N_1623,N_1283);
nand U2715 (N_2715,N_1033,N_1573);
nor U2716 (N_2716,N_1298,N_1710);
xor U2717 (N_2717,N_1728,N_1760);
or U2718 (N_2718,N_1527,N_1307);
and U2719 (N_2719,N_1134,N_1207);
and U2720 (N_2720,N_1539,N_1445);
nand U2721 (N_2721,N_1857,N_1867);
nand U2722 (N_2722,N_1885,N_1776);
nand U2723 (N_2723,N_1832,N_1130);
or U2724 (N_2724,N_1049,N_1976);
nor U2725 (N_2725,N_1881,N_1369);
nor U2726 (N_2726,N_1873,N_1075);
and U2727 (N_2727,N_1825,N_1848);
and U2728 (N_2728,N_1561,N_1094);
xor U2729 (N_2729,N_1105,N_1551);
nor U2730 (N_2730,N_1191,N_1685);
or U2731 (N_2731,N_1816,N_1735);
nand U2732 (N_2732,N_1120,N_1735);
nand U2733 (N_2733,N_1570,N_1750);
nor U2734 (N_2734,N_1590,N_1173);
or U2735 (N_2735,N_1528,N_1818);
and U2736 (N_2736,N_1940,N_1999);
nor U2737 (N_2737,N_1194,N_1673);
nor U2738 (N_2738,N_1489,N_1345);
or U2739 (N_2739,N_1145,N_1105);
nand U2740 (N_2740,N_1057,N_1552);
or U2741 (N_2741,N_1290,N_1366);
and U2742 (N_2742,N_1511,N_1941);
and U2743 (N_2743,N_1092,N_1543);
nand U2744 (N_2744,N_1129,N_1346);
nor U2745 (N_2745,N_1675,N_1080);
nand U2746 (N_2746,N_1132,N_1811);
and U2747 (N_2747,N_1014,N_1976);
or U2748 (N_2748,N_1298,N_1165);
or U2749 (N_2749,N_1465,N_1587);
and U2750 (N_2750,N_1139,N_1120);
and U2751 (N_2751,N_1747,N_1512);
xnor U2752 (N_2752,N_1482,N_1447);
nor U2753 (N_2753,N_1622,N_1482);
nor U2754 (N_2754,N_1588,N_1803);
or U2755 (N_2755,N_1344,N_1954);
or U2756 (N_2756,N_1645,N_1898);
nand U2757 (N_2757,N_1647,N_1950);
xor U2758 (N_2758,N_1631,N_1909);
xor U2759 (N_2759,N_1129,N_1054);
or U2760 (N_2760,N_1860,N_1540);
nor U2761 (N_2761,N_1562,N_1722);
and U2762 (N_2762,N_1476,N_1362);
and U2763 (N_2763,N_1338,N_1215);
or U2764 (N_2764,N_1334,N_1875);
nand U2765 (N_2765,N_1145,N_1959);
nor U2766 (N_2766,N_1511,N_1142);
nor U2767 (N_2767,N_1146,N_1226);
or U2768 (N_2768,N_1962,N_1998);
nor U2769 (N_2769,N_1439,N_1312);
and U2770 (N_2770,N_1132,N_1111);
nand U2771 (N_2771,N_1746,N_1546);
nor U2772 (N_2772,N_1178,N_1103);
nand U2773 (N_2773,N_1593,N_1423);
or U2774 (N_2774,N_1306,N_1694);
or U2775 (N_2775,N_1901,N_1925);
nand U2776 (N_2776,N_1138,N_1838);
nand U2777 (N_2777,N_1550,N_1480);
nand U2778 (N_2778,N_1323,N_1297);
or U2779 (N_2779,N_1095,N_1857);
or U2780 (N_2780,N_1185,N_1162);
or U2781 (N_2781,N_1184,N_1520);
or U2782 (N_2782,N_1971,N_1539);
or U2783 (N_2783,N_1300,N_1447);
nand U2784 (N_2784,N_1687,N_1048);
and U2785 (N_2785,N_1369,N_1937);
nor U2786 (N_2786,N_1181,N_1498);
nor U2787 (N_2787,N_1261,N_1954);
nand U2788 (N_2788,N_1060,N_1716);
and U2789 (N_2789,N_1535,N_1012);
and U2790 (N_2790,N_1458,N_1137);
and U2791 (N_2791,N_1823,N_1561);
nand U2792 (N_2792,N_1724,N_1032);
and U2793 (N_2793,N_1923,N_1574);
nor U2794 (N_2794,N_1375,N_1600);
nand U2795 (N_2795,N_1212,N_1367);
and U2796 (N_2796,N_1139,N_1722);
and U2797 (N_2797,N_1670,N_1808);
and U2798 (N_2798,N_1641,N_1017);
nand U2799 (N_2799,N_1909,N_1899);
nor U2800 (N_2800,N_1761,N_1558);
nor U2801 (N_2801,N_1980,N_1191);
and U2802 (N_2802,N_1209,N_1396);
xor U2803 (N_2803,N_1655,N_1017);
and U2804 (N_2804,N_1730,N_1569);
nand U2805 (N_2805,N_1030,N_1672);
nor U2806 (N_2806,N_1033,N_1714);
or U2807 (N_2807,N_1857,N_1076);
or U2808 (N_2808,N_1973,N_1626);
and U2809 (N_2809,N_1311,N_1398);
or U2810 (N_2810,N_1690,N_1327);
nor U2811 (N_2811,N_1523,N_1612);
nand U2812 (N_2812,N_1359,N_1745);
nand U2813 (N_2813,N_1426,N_1835);
or U2814 (N_2814,N_1524,N_1822);
and U2815 (N_2815,N_1516,N_1251);
or U2816 (N_2816,N_1101,N_1565);
and U2817 (N_2817,N_1597,N_1782);
and U2818 (N_2818,N_1351,N_1940);
nand U2819 (N_2819,N_1696,N_1663);
xor U2820 (N_2820,N_1987,N_1318);
nor U2821 (N_2821,N_1231,N_1371);
nor U2822 (N_2822,N_1055,N_1725);
nand U2823 (N_2823,N_1192,N_1884);
nor U2824 (N_2824,N_1839,N_1596);
nand U2825 (N_2825,N_1133,N_1785);
and U2826 (N_2826,N_1178,N_1533);
nor U2827 (N_2827,N_1466,N_1868);
and U2828 (N_2828,N_1636,N_1389);
nand U2829 (N_2829,N_1484,N_1998);
and U2830 (N_2830,N_1651,N_1313);
nor U2831 (N_2831,N_1676,N_1957);
nand U2832 (N_2832,N_1864,N_1395);
or U2833 (N_2833,N_1706,N_1236);
nor U2834 (N_2834,N_1928,N_1825);
nor U2835 (N_2835,N_1040,N_1434);
nor U2836 (N_2836,N_1116,N_1249);
nand U2837 (N_2837,N_1044,N_1197);
nand U2838 (N_2838,N_1292,N_1591);
nor U2839 (N_2839,N_1990,N_1266);
or U2840 (N_2840,N_1964,N_1137);
and U2841 (N_2841,N_1689,N_1693);
or U2842 (N_2842,N_1820,N_1327);
or U2843 (N_2843,N_1311,N_1855);
nand U2844 (N_2844,N_1091,N_1607);
and U2845 (N_2845,N_1849,N_1002);
nand U2846 (N_2846,N_1084,N_1482);
xor U2847 (N_2847,N_1032,N_1460);
nor U2848 (N_2848,N_1525,N_1510);
nor U2849 (N_2849,N_1492,N_1827);
nand U2850 (N_2850,N_1523,N_1317);
nor U2851 (N_2851,N_1000,N_1174);
and U2852 (N_2852,N_1891,N_1594);
nand U2853 (N_2853,N_1806,N_1065);
nor U2854 (N_2854,N_1820,N_1211);
nor U2855 (N_2855,N_1541,N_1673);
and U2856 (N_2856,N_1952,N_1721);
or U2857 (N_2857,N_1529,N_1265);
nor U2858 (N_2858,N_1571,N_1283);
or U2859 (N_2859,N_1678,N_1526);
or U2860 (N_2860,N_1162,N_1587);
or U2861 (N_2861,N_1300,N_1705);
or U2862 (N_2862,N_1031,N_1667);
nor U2863 (N_2863,N_1625,N_1316);
or U2864 (N_2864,N_1635,N_1874);
and U2865 (N_2865,N_1936,N_1139);
nor U2866 (N_2866,N_1455,N_1709);
or U2867 (N_2867,N_1323,N_1527);
or U2868 (N_2868,N_1108,N_1592);
nand U2869 (N_2869,N_1499,N_1733);
and U2870 (N_2870,N_1567,N_1959);
and U2871 (N_2871,N_1395,N_1371);
nand U2872 (N_2872,N_1220,N_1688);
and U2873 (N_2873,N_1834,N_1697);
nor U2874 (N_2874,N_1669,N_1182);
nor U2875 (N_2875,N_1186,N_1139);
or U2876 (N_2876,N_1468,N_1249);
or U2877 (N_2877,N_1952,N_1608);
nor U2878 (N_2878,N_1257,N_1408);
nor U2879 (N_2879,N_1224,N_1593);
nand U2880 (N_2880,N_1762,N_1002);
and U2881 (N_2881,N_1586,N_1289);
and U2882 (N_2882,N_1060,N_1169);
or U2883 (N_2883,N_1339,N_1071);
nor U2884 (N_2884,N_1158,N_1968);
nor U2885 (N_2885,N_1239,N_1188);
and U2886 (N_2886,N_1030,N_1366);
and U2887 (N_2887,N_1788,N_1390);
and U2888 (N_2888,N_1833,N_1980);
nand U2889 (N_2889,N_1429,N_1629);
and U2890 (N_2890,N_1183,N_1208);
and U2891 (N_2891,N_1896,N_1943);
nor U2892 (N_2892,N_1932,N_1234);
nand U2893 (N_2893,N_1712,N_1852);
or U2894 (N_2894,N_1907,N_1153);
nor U2895 (N_2895,N_1591,N_1646);
or U2896 (N_2896,N_1427,N_1937);
nand U2897 (N_2897,N_1575,N_1339);
and U2898 (N_2898,N_1430,N_1010);
or U2899 (N_2899,N_1716,N_1437);
nand U2900 (N_2900,N_1751,N_1172);
nor U2901 (N_2901,N_1724,N_1435);
nand U2902 (N_2902,N_1169,N_1785);
or U2903 (N_2903,N_1040,N_1753);
nor U2904 (N_2904,N_1479,N_1818);
and U2905 (N_2905,N_1820,N_1418);
or U2906 (N_2906,N_1746,N_1736);
or U2907 (N_2907,N_1030,N_1862);
nor U2908 (N_2908,N_1813,N_1893);
and U2909 (N_2909,N_1240,N_1701);
nor U2910 (N_2910,N_1156,N_1534);
nand U2911 (N_2911,N_1037,N_1904);
and U2912 (N_2912,N_1794,N_1243);
and U2913 (N_2913,N_1586,N_1265);
nor U2914 (N_2914,N_1228,N_1642);
nand U2915 (N_2915,N_1921,N_1181);
nor U2916 (N_2916,N_1022,N_1493);
nor U2917 (N_2917,N_1128,N_1469);
xor U2918 (N_2918,N_1023,N_1240);
and U2919 (N_2919,N_1612,N_1110);
nor U2920 (N_2920,N_1978,N_1136);
or U2921 (N_2921,N_1283,N_1285);
nand U2922 (N_2922,N_1619,N_1250);
and U2923 (N_2923,N_1636,N_1670);
xnor U2924 (N_2924,N_1158,N_1226);
nand U2925 (N_2925,N_1445,N_1458);
nor U2926 (N_2926,N_1306,N_1337);
nor U2927 (N_2927,N_1339,N_1162);
nand U2928 (N_2928,N_1642,N_1754);
nand U2929 (N_2929,N_1309,N_1542);
nand U2930 (N_2930,N_1194,N_1785);
nor U2931 (N_2931,N_1673,N_1932);
xor U2932 (N_2932,N_1686,N_1470);
and U2933 (N_2933,N_1316,N_1497);
nor U2934 (N_2934,N_1294,N_1651);
or U2935 (N_2935,N_1311,N_1288);
and U2936 (N_2936,N_1560,N_1641);
or U2937 (N_2937,N_1616,N_1518);
nand U2938 (N_2938,N_1083,N_1016);
nand U2939 (N_2939,N_1386,N_1727);
or U2940 (N_2940,N_1767,N_1536);
nor U2941 (N_2941,N_1734,N_1188);
nand U2942 (N_2942,N_1320,N_1692);
or U2943 (N_2943,N_1475,N_1981);
nor U2944 (N_2944,N_1059,N_1280);
nor U2945 (N_2945,N_1844,N_1816);
nor U2946 (N_2946,N_1076,N_1303);
and U2947 (N_2947,N_1672,N_1059);
and U2948 (N_2948,N_1704,N_1279);
or U2949 (N_2949,N_1163,N_1884);
nor U2950 (N_2950,N_1082,N_1260);
nand U2951 (N_2951,N_1019,N_1499);
and U2952 (N_2952,N_1310,N_1296);
or U2953 (N_2953,N_1686,N_1968);
and U2954 (N_2954,N_1965,N_1748);
or U2955 (N_2955,N_1803,N_1677);
nor U2956 (N_2956,N_1960,N_1106);
nor U2957 (N_2957,N_1115,N_1164);
nor U2958 (N_2958,N_1785,N_1460);
nand U2959 (N_2959,N_1970,N_1589);
nand U2960 (N_2960,N_1271,N_1096);
nand U2961 (N_2961,N_1461,N_1807);
nor U2962 (N_2962,N_1685,N_1341);
nand U2963 (N_2963,N_1143,N_1310);
nand U2964 (N_2964,N_1486,N_1162);
nor U2965 (N_2965,N_1658,N_1541);
nor U2966 (N_2966,N_1128,N_1702);
nand U2967 (N_2967,N_1957,N_1948);
or U2968 (N_2968,N_1391,N_1682);
and U2969 (N_2969,N_1647,N_1151);
nand U2970 (N_2970,N_1253,N_1633);
or U2971 (N_2971,N_1822,N_1441);
and U2972 (N_2972,N_1613,N_1549);
nand U2973 (N_2973,N_1912,N_1855);
nor U2974 (N_2974,N_1301,N_1835);
nand U2975 (N_2975,N_1132,N_1922);
and U2976 (N_2976,N_1481,N_1437);
and U2977 (N_2977,N_1845,N_1860);
nand U2978 (N_2978,N_1897,N_1247);
or U2979 (N_2979,N_1247,N_1733);
and U2980 (N_2980,N_1745,N_1720);
nand U2981 (N_2981,N_1751,N_1426);
nand U2982 (N_2982,N_1149,N_1066);
and U2983 (N_2983,N_1705,N_1233);
or U2984 (N_2984,N_1817,N_1279);
xnor U2985 (N_2985,N_1708,N_1259);
nor U2986 (N_2986,N_1057,N_1115);
nand U2987 (N_2987,N_1282,N_1033);
and U2988 (N_2988,N_1981,N_1694);
or U2989 (N_2989,N_1195,N_1208);
nand U2990 (N_2990,N_1659,N_1041);
and U2991 (N_2991,N_1342,N_1849);
nor U2992 (N_2992,N_1762,N_1470);
or U2993 (N_2993,N_1104,N_1604);
nor U2994 (N_2994,N_1178,N_1613);
and U2995 (N_2995,N_1690,N_1178);
and U2996 (N_2996,N_1973,N_1676);
nand U2997 (N_2997,N_1616,N_1085);
or U2998 (N_2998,N_1383,N_1378);
xnor U2999 (N_2999,N_1317,N_1367);
nor U3000 (N_3000,N_2402,N_2956);
nand U3001 (N_3001,N_2578,N_2069);
and U3002 (N_3002,N_2879,N_2000);
nand U3003 (N_3003,N_2110,N_2464);
nand U3004 (N_3004,N_2650,N_2266);
or U3005 (N_3005,N_2176,N_2157);
nand U3006 (N_3006,N_2033,N_2940);
or U3007 (N_3007,N_2821,N_2762);
xor U3008 (N_3008,N_2324,N_2703);
or U3009 (N_3009,N_2507,N_2630);
and U3010 (N_3010,N_2187,N_2674);
or U3011 (N_3011,N_2895,N_2197);
or U3012 (N_3012,N_2383,N_2700);
or U3013 (N_3013,N_2095,N_2531);
nand U3014 (N_3014,N_2035,N_2226);
nand U3015 (N_3015,N_2947,N_2004);
and U3016 (N_3016,N_2482,N_2448);
xor U3017 (N_3017,N_2679,N_2795);
nand U3018 (N_3018,N_2787,N_2306);
xnor U3019 (N_3019,N_2686,N_2583);
or U3020 (N_3020,N_2294,N_2493);
nor U3021 (N_3021,N_2455,N_2677);
xnor U3022 (N_3022,N_2903,N_2367);
and U3023 (N_3023,N_2883,N_2437);
nor U3024 (N_3024,N_2620,N_2627);
and U3025 (N_3025,N_2436,N_2721);
and U3026 (N_3026,N_2692,N_2673);
nand U3027 (N_3027,N_2162,N_2124);
nand U3028 (N_3028,N_2459,N_2327);
and U3029 (N_3029,N_2657,N_2639);
nor U3030 (N_3030,N_2667,N_2793);
or U3031 (N_3031,N_2812,N_2076);
and U3032 (N_3032,N_2648,N_2575);
or U3033 (N_3033,N_2789,N_2325);
nand U3034 (N_3034,N_2732,N_2345);
nor U3035 (N_3035,N_2937,N_2952);
nand U3036 (N_3036,N_2872,N_2736);
nand U3037 (N_3037,N_2598,N_2855);
nand U3038 (N_3038,N_2709,N_2591);
nand U3039 (N_3039,N_2473,N_2468);
and U3040 (N_3040,N_2103,N_2751);
and U3041 (N_3041,N_2061,N_2340);
or U3042 (N_3042,N_2082,N_2715);
nor U3043 (N_3043,N_2057,N_2809);
nor U3044 (N_3044,N_2240,N_2518);
and U3045 (N_3045,N_2605,N_2801);
and U3046 (N_3046,N_2961,N_2869);
nand U3047 (N_3047,N_2857,N_2764);
nor U3048 (N_3048,N_2411,N_2900);
nand U3049 (N_3049,N_2746,N_2156);
nand U3050 (N_3050,N_2585,N_2218);
and U3051 (N_3051,N_2376,N_2782);
and U3052 (N_3052,N_2768,N_2151);
and U3053 (N_3053,N_2091,N_2971);
or U3054 (N_3054,N_2353,N_2177);
or U3055 (N_3055,N_2001,N_2817);
and U3056 (N_3056,N_2009,N_2860);
nand U3057 (N_3057,N_2036,N_2923);
nand U3058 (N_3058,N_2342,N_2118);
or U3059 (N_3059,N_2698,N_2668);
or U3060 (N_3060,N_2790,N_2127);
nor U3061 (N_3061,N_2239,N_2007);
nand U3062 (N_3062,N_2344,N_2569);
nand U3063 (N_3063,N_2757,N_2930);
nor U3064 (N_3064,N_2395,N_2910);
or U3065 (N_3065,N_2726,N_2731);
nand U3066 (N_3066,N_2904,N_2121);
or U3067 (N_3067,N_2547,N_2488);
or U3068 (N_3068,N_2143,N_2804);
xnor U3069 (N_3069,N_2180,N_2435);
nand U3070 (N_3070,N_2363,N_2564);
nand U3071 (N_3071,N_2577,N_2765);
or U3072 (N_3072,N_2944,N_2894);
nor U3073 (N_3073,N_2548,N_2481);
nand U3074 (N_3074,N_2638,N_2109);
xor U3075 (N_3075,N_2675,N_2823);
nand U3076 (N_3076,N_2561,N_2465);
and U3077 (N_3077,N_2893,N_2797);
nand U3078 (N_3078,N_2926,N_2038);
or U3079 (N_3079,N_2070,N_2916);
nor U3080 (N_3080,N_2633,N_2168);
nor U3081 (N_3081,N_2539,N_2415);
or U3082 (N_3082,N_2773,N_2412);
or U3083 (N_3083,N_2943,N_2502);
and U3084 (N_3084,N_2398,N_2298);
nand U3085 (N_3085,N_2771,N_2310);
and U3086 (N_3086,N_2311,N_2553);
and U3087 (N_3087,N_2031,N_2166);
nand U3088 (N_3088,N_2358,N_2545);
or U3089 (N_3089,N_2831,N_2207);
xnor U3090 (N_3090,N_2421,N_2497);
nand U3091 (N_3091,N_2409,N_2687);
nor U3092 (N_3092,N_2217,N_2615);
or U3093 (N_3093,N_2037,N_2593);
or U3094 (N_3094,N_2949,N_2958);
nor U3095 (N_3095,N_2735,N_2044);
nand U3096 (N_3096,N_2443,N_2614);
nor U3097 (N_3097,N_2484,N_2800);
nand U3098 (N_3098,N_2612,N_2466);
nand U3099 (N_3099,N_2631,N_2955);
nor U3100 (N_3100,N_2719,N_2695);
and U3101 (N_3101,N_2020,N_2053);
nor U3102 (N_3102,N_2802,N_2529);
and U3103 (N_3103,N_2242,N_2186);
nor U3104 (N_3104,N_2030,N_2932);
and U3105 (N_3105,N_2541,N_2505);
and U3106 (N_3106,N_2832,N_2661);
and U3107 (N_3107,N_2935,N_2866);
and U3108 (N_3108,N_2595,N_2431);
and U3109 (N_3109,N_2097,N_2305);
or U3110 (N_3110,N_2806,N_2604);
or U3111 (N_3111,N_2780,N_2382);
nor U3112 (N_3112,N_2265,N_2978);
or U3113 (N_3113,N_2406,N_2196);
or U3114 (N_3114,N_2445,N_2556);
and U3115 (N_3115,N_2369,N_2193);
or U3116 (N_3116,N_2563,N_2424);
xnor U3117 (N_3117,N_2141,N_2597);
nor U3118 (N_3118,N_2254,N_2767);
or U3119 (N_3119,N_2694,N_2050);
or U3120 (N_3120,N_2144,N_2273);
and U3121 (N_3121,N_2815,N_2471);
and U3122 (N_3122,N_2241,N_2205);
and U3123 (N_3123,N_2316,N_2995);
or U3124 (N_3124,N_2028,N_2898);
nor U3125 (N_3125,N_2368,N_2308);
nand U3126 (N_3126,N_2418,N_2389);
or U3127 (N_3127,N_2642,N_2984);
or U3128 (N_3128,N_2624,N_2610);
and U3129 (N_3129,N_2979,N_2927);
nand U3130 (N_3130,N_2938,N_2770);
and U3131 (N_3131,N_2999,N_2514);
and U3132 (N_3132,N_2986,N_2691);
and U3133 (N_3133,N_2199,N_2158);
or U3134 (N_3134,N_2364,N_2613);
or U3135 (N_3135,N_2512,N_2813);
nor U3136 (N_3136,N_2798,N_2702);
and U3137 (N_3137,N_2211,N_2003);
nor U3138 (N_3138,N_2974,N_2783);
and U3139 (N_3139,N_2326,N_2527);
and U3140 (N_3140,N_2587,N_2796);
nor U3141 (N_3141,N_2623,N_2524);
nor U3142 (N_3142,N_2863,N_2704);
xor U3143 (N_3143,N_2077,N_2078);
nor U3144 (N_3144,N_2617,N_2963);
nand U3145 (N_3145,N_2915,N_2272);
nor U3146 (N_3146,N_2351,N_2046);
nand U3147 (N_3147,N_2234,N_2034);
and U3148 (N_3148,N_2745,N_2244);
xnor U3149 (N_3149,N_2808,N_2608);
and U3150 (N_3150,N_2526,N_2022);
and U3151 (N_3151,N_2554,N_2948);
nand U3152 (N_3152,N_2059,N_2132);
nor U3153 (N_3153,N_2432,N_2063);
and U3154 (N_3154,N_2341,N_2741);
nor U3155 (N_3155,N_2339,N_2139);
nand U3156 (N_3156,N_2092,N_2820);
xor U3157 (N_3157,N_2877,N_2589);
or U3158 (N_3158,N_2286,N_2519);
nand U3159 (N_3159,N_2774,N_2438);
xnor U3160 (N_3160,N_2334,N_2075);
xor U3161 (N_3161,N_2551,N_2985);
or U3162 (N_3162,N_2475,N_2149);
nor U3163 (N_3163,N_2029,N_2346);
or U3164 (N_3164,N_2159,N_2772);
nand U3165 (N_3165,N_2085,N_2622);
nand U3166 (N_3166,N_2784,N_2290);
or U3167 (N_3167,N_2896,N_2665);
or U3168 (N_3168,N_2912,N_2045);
xor U3169 (N_3169,N_2039,N_2452);
xor U3170 (N_3170,N_2106,N_2881);
or U3171 (N_3171,N_2429,N_2015);
nand U3172 (N_3172,N_2565,N_2439);
nand U3173 (N_3173,N_2534,N_2901);
or U3174 (N_3174,N_2213,N_2403);
and U3175 (N_3175,N_2084,N_2338);
nor U3176 (N_3176,N_2536,N_2906);
or U3177 (N_3177,N_2047,N_2739);
nand U3178 (N_3178,N_2396,N_2490);
nand U3179 (N_3179,N_2041,N_2018);
xor U3180 (N_3180,N_2954,N_2333);
nand U3181 (N_3181,N_2716,N_2275);
and U3182 (N_3182,N_2192,N_2147);
nor U3183 (N_3183,N_2641,N_2449);
and U3184 (N_3184,N_2861,N_2822);
and U3185 (N_3185,N_2463,N_2755);
and U3186 (N_3186,N_2011,N_2469);
nand U3187 (N_3187,N_2130,N_2479);
or U3188 (N_3188,N_2251,N_2165);
or U3189 (N_3189,N_2073,N_2387);
or U3190 (N_3190,N_2191,N_2837);
and U3191 (N_3191,N_2580,N_2330);
and U3192 (N_3192,N_2530,N_2865);
nand U3193 (N_3193,N_2884,N_2384);
nand U3194 (N_3194,N_2150,N_2889);
and U3195 (N_3195,N_2705,N_2182);
and U3196 (N_3196,N_2697,N_2173);
and U3197 (N_3197,N_2523,N_2319);
nor U3198 (N_3198,N_2289,N_2775);
xnor U3199 (N_3199,N_2343,N_2742);
and U3200 (N_3200,N_2131,N_2042);
nor U3201 (N_3201,N_2946,N_2905);
nand U3202 (N_3202,N_2748,N_2891);
or U3203 (N_3203,N_2397,N_2281);
or U3204 (N_3204,N_2611,N_2981);
nor U3205 (N_3205,N_2992,N_2257);
and U3206 (N_3206,N_2828,N_2747);
and U3207 (N_3207,N_2404,N_2458);
nor U3208 (N_3208,N_2055,N_2743);
nor U3209 (N_3209,N_2887,N_2522);
nor U3210 (N_3210,N_2581,N_2181);
nand U3211 (N_3211,N_2645,N_2964);
and U3212 (N_3212,N_2495,N_2811);
or U3213 (N_3213,N_2803,N_2474);
or U3214 (N_3214,N_2164,N_2880);
and U3215 (N_3215,N_2799,N_2440);
and U3216 (N_3216,N_2867,N_2267);
or U3217 (N_3217,N_2349,N_2447);
nor U3218 (N_3218,N_2087,N_2560);
and U3219 (N_3219,N_2568,N_2072);
nor U3220 (N_3220,N_2284,N_2834);
and U3221 (N_3221,N_2013,N_2924);
nor U3222 (N_3222,N_2997,N_2049);
xnor U3223 (N_3223,N_2461,N_2043);
nand U3224 (N_3224,N_2202,N_2122);
nand U3225 (N_3225,N_2525,N_2080);
and U3226 (N_3226,N_2385,N_2026);
nor U3227 (N_3227,N_2678,N_2725);
nand U3228 (N_3228,N_2271,N_2951);
nor U3229 (N_3229,N_2320,N_2566);
nand U3230 (N_3230,N_2111,N_2573);
and U3231 (N_3231,N_2658,N_2021);
nand U3232 (N_3232,N_2256,N_2322);
nand U3233 (N_3233,N_2666,N_2391);
xor U3234 (N_3234,N_2752,N_2816);
nand U3235 (N_3235,N_2220,N_2183);
or U3236 (N_3236,N_2838,N_2652);
and U3237 (N_3237,N_2285,N_2683);
xnor U3238 (N_3238,N_2847,N_2052);
or U3239 (N_3239,N_2138,N_2939);
or U3240 (N_3240,N_2989,N_2331);
nand U3241 (N_3241,N_2094,N_2224);
nand U3242 (N_3242,N_2017,N_2048);
nor U3243 (N_3243,N_2304,N_2172);
or U3244 (N_3244,N_2504,N_2909);
or U3245 (N_3245,N_2067,N_2014);
nor U3246 (N_3246,N_2921,N_2761);
and U3247 (N_3247,N_2386,N_2462);
and U3248 (N_3248,N_2178,N_2380);
nand U3249 (N_3249,N_2225,N_2203);
nor U3250 (N_3250,N_2329,N_2791);
or U3251 (N_3251,N_2212,N_2637);
nand U3252 (N_3252,N_2843,N_2788);
nand U3253 (N_3253,N_2407,N_2381);
or U3254 (N_3254,N_2291,N_2301);
nand U3255 (N_3255,N_2712,N_2002);
and U3256 (N_3256,N_2934,N_2546);
and U3257 (N_3257,N_2537,N_2390);
or U3258 (N_3258,N_2019,N_2646);
nor U3259 (N_3259,N_2786,N_2315);
or U3260 (N_3260,N_2517,N_2129);
nand U3261 (N_3261,N_2988,N_2140);
or U3262 (N_3262,N_2701,N_2259);
nand U3263 (N_3263,N_2231,N_2508);
nor U3264 (N_3264,N_2859,N_2662);
and U3265 (N_3265,N_2270,N_2635);
nor U3266 (N_3266,N_2312,N_2054);
nand U3267 (N_3267,N_2235,N_2025);
or U3268 (N_3268,N_2426,N_2253);
and U3269 (N_3269,N_2763,N_2478);
nand U3270 (N_3270,N_2247,N_2420);
xor U3271 (N_3271,N_2965,N_2886);
and U3272 (N_3272,N_2416,N_2260);
and U3273 (N_3273,N_2562,N_2393);
nor U3274 (N_3274,N_2169,N_2684);
nor U3275 (N_3275,N_2664,N_2875);
and U3276 (N_3276,N_2681,N_2920);
and U3277 (N_3277,N_2125,N_2606);
and U3278 (N_3278,N_2826,N_2829);
xnor U3279 (N_3279,N_2317,N_2819);
nor U3280 (N_3280,N_2016,N_2676);
or U3281 (N_3281,N_2972,N_2010);
and U3282 (N_3282,N_2467,N_2264);
nor U3283 (N_3283,N_2074,N_2706);
or U3284 (N_3284,N_2313,N_2137);
nand U3285 (N_3285,N_2457,N_2730);
nand U3286 (N_3286,N_2874,N_2051);
nor U3287 (N_3287,N_2347,N_2987);
nand U3288 (N_3288,N_2274,N_2753);
nor U3289 (N_3289,N_2135,N_2472);
and U3290 (N_3290,N_2119,N_2660);
xnor U3291 (N_3291,N_2370,N_2890);
and U3292 (N_3292,N_2012,N_2071);
nand U3293 (N_3293,N_2088,N_2555);
and U3294 (N_3294,N_2827,N_2852);
nor U3295 (N_3295,N_2328,N_2104);
or U3296 (N_3296,N_2552,N_2167);
and U3297 (N_3297,N_2064,N_2348);
or U3298 (N_3298,N_2410,N_2496);
and U3299 (N_3299,N_2332,N_2194);
nand U3300 (N_3300,N_2366,N_2629);
and U3301 (N_3301,N_2509,N_2671);
or U3302 (N_3302,N_2008,N_2922);
and U3303 (N_3303,N_2814,N_2230);
xor U3304 (N_3304,N_2388,N_2499);
or U3305 (N_3305,N_2897,N_2856);
nor U3306 (N_3306,N_2618,N_2559);
nand U3307 (N_3307,N_2371,N_2734);
nand U3308 (N_3308,N_2221,N_2841);
or U3309 (N_3309,N_2277,N_2441);
nand U3310 (N_3310,N_2532,N_2163);
nand U3311 (N_3311,N_2250,N_2544);
or U3312 (N_3312,N_2713,N_2925);
xor U3313 (N_3313,N_2685,N_2302);
and U3314 (N_3314,N_2006,N_2836);
or U3315 (N_3315,N_2998,N_2533);
or U3316 (N_3316,N_2628,N_2873);
or U3317 (N_3317,N_2114,N_2200);
xnor U3318 (N_3318,N_2210,N_2400);
and U3319 (N_3319,N_2198,N_2179);
and U3320 (N_3320,N_2093,N_2557);
and U3321 (N_3321,N_2848,N_2871);
nand U3322 (N_3322,N_2146,N_2835);
or U3323 (N_3323,N_2056,N_2243);
nor U3324 (N_3324,N_2969,N_2807);
nand U3325 (N_3325,N_2487,N_2280);
or U3326 (N_3326,N_2433,N_2669);
nand U3327 (N_3327,N_2749,N_2268);
nand U3328 (N_3328,N_2219,N_2249);
nand U3329 (N_3329,N_2255,N_2292);
nor U3330 (N_3330,N_2405,N_2659);
nand U3331 (N_3331,N_2195,N_2204);
xnor U3332 (N_3332,N_2511,N_2818);
nor U3333 (N_3333,N_2350,N_2501);
nor U3334 (N_3334,N_2689,N_2456);
nand U3335 (N_3335,N_2851,N_2711);
nor U3336 (N_3336,N_2663,N_2263);
or U3337 (N_3337,N_2878,N_2876);
or U3338 (N_3338,N_2483,N_2083);
nor U3339 (N_3339,N_2160,N_2967);
and U3340 (N_3340,N_2602,N_2616);
and U3341 (N_3341,N_2378,N_2261);
nand U3342 (N_3342,N_2699,N_2128);
nor U3343 (N_3343,N_2754,N_2336);
nand U3344 (N_3344,N_2579,N_2805);
or U3345 (N_3345,N_2117,N_2973);
or U3346 (N_3346,N_2521,N_2991);
or U3347 (N_3347,N_2005,N_2399);
or U3348 (N_3348,N_2237,N_2278);
and U3349 (N_3349,N_2550,N_2116);
and U3350 (N_3350,N_2592,N_2223);
and U3351 (N_3351,N_2510,N_2928);
nand U3352 (N_3352,N_2759,N_2607);
or U3353 (N_3353,N_2171,N_2892);
and U3354 (N_3354,N_2824,N_2888);
nor U3355 (N_3355,N_2941,N_2643);
or U3356 (N_3356,N_2833,N_2931);
and U3357 (N_3357,N_2089,N_2756);
nor U3358 (N_3358,N_2372,N_2201);
nor U3359 (N_3359,N_2722,N_2572);
xnor U3360 (N_3360,N_2649,N_2810);
nand U3361 (N_3361,N_2586,N_2090);
and U3362 (N_3362,N_2480,N_2287);
nor U3363 (N_3363,N_2238,N_2335);
or U3364 (N_3364,N_2609,N_2105);
nor U3365 (N_3365,N_2626,N_2318);
and U3366 (N_3366,N_2228,N_2506);
nand U3367 (N_3367,N_2477,N_2027);
or U3368 (N_3368,N_2723,N_2760);
nor U3369 (N_3369,N_2738,N_2968);
nand U3370 (N_3370,N_2354,N_2724);
nand U3371 (N_3371,N_2101,N_2858);
nand U3372 (N_3372,N_2236,N_2990);
nand U3373 (N_3373,N_2902,N_2491);
nand U3374 (N_3374,N_2428,N_2108);
or U3375 (N_3375,N_2942,N_2214);
nand U3376 (N_3376,N_2936,N_2269);
and U3377 (N_3377,N_2222,N_2516);
or U3378 (N_3378,N_2542,N_2654);
nor U3379 (N_3379,N_2245,N_2794);
nor U3380 (N_3380,N_2423,N_2885);
and U3381 (N_3381,N_2161,N_2543);
and U3382 (N_3382,N_2392,N_2123);
and U3383 (N_3383,N_2917,N_2778);
or U3384 (N_3384,N_2779,N_2549);
nand U3385 (N_3385,N_2977,N_2414);
or U3386 (N_3386,N_2766,N_2913);
and U3387 (N_3387,N_2846,N_2081);
and U3388 (N_3388,N_2582,N_2227);
or U3389 (N_3389,N_2229,N_2188);
nand U3390 (N_3390,N_2209,N_2494);
or U3391 (N_3391,N_2476,N_2850);
nand U3392 (N_3392,N_2682,N_2337);
nor U3393 (N_3393,N_2574,N_2634);
nor U3394 (N_3394,N_2184,N_2950);
nor U3395 (N_3395,N_2744,N_2434);
or U3396 (N_3396,N_2361,N_2148);
nand U3397 (N_3397,N_2296,N_2215);
nor U3398 (N_3398,N_2717,N_2590);
and U3399 (N_3399,N_2688,N_2599);
xor U3400 (N_3400,N_2145,N_2933);
and U3401 (N_3401,N_2058,N_2401);
nand U3402 (N_3402,N_2040,N_2769);
xnor U3403 (N_3403,N_2113,N_2707);
nor U3404 (N_3404,N_2945,N_2870);
or U3405 (N_3405,N_2714,N_2185);
and U3406 (N_3406,N_2750,N_2601);
nand U3407 (N_3407,N_2588,N_2098);
and U3408 (N_3408,N_2153,N_2538);
nand U3409 (N_3409,N_2099,N_2307);
and U3410 (N_3410,N_2596,N_2252);
nor U3411 (N_3411,N_2379,N_2727);
and U3412 (N_3412,N_2740,N_2190);
or U3413 (N_3413,N_2068,N_2728);
and U3414 (N_3414,N_2503,N_2982);
or U3415 (N_3415,N_2216,N_2983);
nor U3416 (N_3416,N_2232,N_2849);
and U3417 (N_3417,N_2102,N_2929);
and U3418 (N_3418,N_2446,N_2840);
or U3419 (N_3419,N_2993,N_2647);
or U3420 (N_3420,N_2844,N_2737);
nand U3421 (N_3421,N_2115,N_2417);
xnor U3422 (N_3422,N_2792,N_2134);
nand U3423 (N_3423,N_2980,N_2460);
nor U3424 (N_3424,N_2422,N_2644);
and U3425 (N_3425,N_2258,N_2086);
and U3426 (N_3426,N_2696,N_2206);
or U3427 (N_3427,N_2451,N_2853);
nand U3428 (N_3428,N_2670,N_2603);
nor U3429 (N_3429,N_2758,N_2377);
nor U3430 (N_3430,N_2133,N_2842);
and U3431 (N_3431,N_2619,N_2854);
nand U3432 (N_3432,N_2066,N_2155);
or U3433 (N_3433,N_2500,N_2425);
xnor U3434 (N_3434,N_2233,N_2962);
nor U3435 (N_3435,N_2830,N_2919);
or U3436 (N_3436,N_2540,N_2845);
nand U3437 (N_3437,N_2175,N_2096);
or U3438 (N_3438,N_2314,N_2024);
and U3439 (N_3439,N_2571,N_2374);
nand U3440 (N_3440,N_2899,N_2444);
and U3441 (N_3441,N_2365,N_2720);
or U3442 (N_3442,N_2970,N_2293);
or U3443 (N_3443,N_2170,N_2279);
nor U3444 (N_3444,N_2126,N_2283);
and U3445 (N_3445,N_2454,N_2136);
and U3446 (N_3446,N_2032,N_2394);
nand U3447 (N_3447,N_2489,N_2966);
or U3448 (N_3448,N_2975,N_2413);
xor U3449 (N_3449,N_2918,N_2154);
nand U3450 (N_3450,N_2282,N_2453);
or U3451 (N_3451,N_2655,N_2570);
nand U3452 (N_3452,N_2733,N_2375);
and U3453 (N_3453,N_2653,N_2656);
nor U3454 (N_3454,N_2486,N_2959);
and U3455 (N_3455,N_2680,N_2632);
nor U3456 (N_3456,N_2864,N_2485);
or U3457 (N_3457,N_2100,N_2300);
and U3458 (N_3458,N_2060,N_2708);
nor U3459 (N_3459,N_2208,N_2112);
or U3460 (N_3460,N_2957,N_2174);
nor U3461 (N_3461,N_2189,N_2868);
nand U3462 (N_3462,N_2352,N_2594);
and U3463 (N_3463,N_2693,N_2528);
nor U3464 (N_3464,N_2299,N_2960);
and U3465 (N_3465,N_2356,N_2882);
and U3466 (N_3466,N_2419,N_2994);
and U3467 (N_3467,N_2142,N_2839);
nor U3468 (N_3468,N_2576,N_2584);
xnor U3469 (N_3469,N_2430,N_2718);
nor U3470 (N_3470,N_2023,N_2636);
and U3471 (N_3471,N_2427,N_2408);
nor U3472 (N_3472,N_2470,N_2907);
nor U3473 (N_3473,N_2079,N_2498);
or U3474 (N_3474,N_2120,N_2785);
nand U3475 (N_3475,N_2908,N_2107);
nor U3476 (N_3476,N_2621,N_2323);
and U3477 (N_3477,N_2911,N_2651);
nand U3478 (N_3478,N_2262,N_2862);
nand U3479 (N_3479,N_2062,N_2355);
xor U3480 (N_3480,N_2492,N_2357);
nand U3481 (N_3481,N_2450,N_2672);
nor U3482 (N_3482,N_2690,N_2953);
nor U3483 (N_3483,N_2362,N_2567);
nand U3484 (N_3484,N_2625,N_2513);
or U3485 (N_3485,N_2295,N_2373);
nor U3486 (N_3486,N_2288,N_2776);
nor U3487 (N_3487,N_2825,N_2777);
nor U3488 (N_3488,N_2710,N_2360);
nor U3489 (N_3489,N_2303,N_2515);
nand U3490 (N_3490,N_2520,N_2276);
nor U3491 (N_3491,N_2558,N_2996);
nor U3492 (N_3492,N_2640,N_2914);
and U3493 (N_3493,N_2297,N_2248);
nand U3494 (N_3494,N_2976,N_2309);
or U3495 (N_3495,N_2152,N_2246);
or U3496 (N_3496,N_2600,N_2442);
or U3497 (N_3497,N_2729,N_2535);
nand U3498 (N_3498,N_2359,N_2065);
and U3499 (N_3499,N_2321,N_2781);
or U3500 (N_3500,N_2911,N_2950);
and U3501 (N_3501,N_2865,N_2887);
nor U3502 (N_3502,N_2252,N_2557);
and U3503 (N_3503,N_2858,N_2573);
and U3504 (N_3504,N_2206,N_2414);
and U3505 (N_3505,N_2427,N_2009);
nor U3506 (N_3506,N_2699,N_2280);
and U3507 (N_3507,N_2958,N_2034);
nand U3508 (N_3508,N_2685,N_2153);
or U3509 (N_3509,N_2642,N_2480);
nand U3510 (N_3510,N_2072,N_2320);
nor U3511 (N_3511,N_2244,N_2128);
xnor U3512 (N_3512,N_2349,N_2354);
or U3513 (N_3513,N_2690,N_2995);
nand U3514 (N_3514,N_2674,N_2596);
and U3515 (N_3515,N_2314,N_2216);
nor U3516 (N_3516,N_2618,N_2998);
and U3517 (N_3517,N_2167,N_2603);
or U3518 (N_3518,N_2437,N_2516);
nor U3519 (N_3519,N_2263,N_2875);
nand U3520 (N_3520,N_2613,N_2157);
and U3521 (N_3521,N_2756,N_2151);
and U3522 (N_3522,N_2646,N_2649);
and U3523 (N_3523,N_2350,N_2970);
nand U3524 (N_3524,N_2876,N_2563);
or U3525 (N_3525,N_2682,N_2608);
nor U3526 (N_3526,N_2797,N_2325);
nand U3527 (N_3527,N_2747,N_2409);
nor U3528 (N_3528,N_2351,N_2056);
or U3529 (N_3529,N_2768,N_2840);
nor U3530 (N_3530,N_2404,N_2936);
or U3531 (N_3531,N_2437,N_2434);
and U3532 (N_3532,N_2487,N_2536);
nand U3533 (N_3533,N_2337,N_2877);
nor U3534 (N_3534,N_2329,N_2834);
nor U3535 (N_3535,N_2688,N_2068);
and U3536 (N_3536,N_2219,N_2372);
or U3537 (N_3537,N_2626,N_2693);
and U3538 (N_3538,N_2037,N_2898);
nor U3539 (N_3539,N_2964,N_2492);
and U3540 (N_3540,N_2486,N_2466);
and U3541 (N_3541,N_2801,N_2538);
and U3542 (N_3542,N_2900,N_2808);
and U3543 (N_3543,N_2365,N_2197);
nor U3544 (N_3544,N_2932,N_2085);
or U3545 (N_3545,N_2197,N_2087);
and U3546 (N_3546,N_2866,N_2798);
nor U3547 (N_3547,N_2291,N_2953);
or U3548 (N_3548,N_2391,N_2687);
or U3549 (N_3549,N_2436,N_2168);
nand U3550 (N_3550,N_2974,N_2180);
nand U3551 (N_3551,N_2150,N_2922);
nand U3552 (N_3552,N_2364,N_2197);
nor U3553 (N_3553,N_2702,N_2741);
nor U3554 (N_3554,N_2964,N_2626);
and U3555 (N_3555,N_2036,N_2575);
nand U3556 (N_3556,N_2651,N_2404);
and U3557 (N_3557,N_2839,N_2353);
nor U3558 (N_3558,N_2866,N_2478);
and U3559 (N_3559,N_2854,N_2200);
nand U3560 (N_3560,N_2361,N_2067);
and U3561 (N_3561,N_2296,N_2627);
and U3562 (N_3562,N_2849,N_2838);
nor U3563 (N_3563,N_2696,N_2945);
and U3564 (N_3564,N_2883,N_2783);
and U3565 (N_3565,N_2043,N_2481);
or U3566 (N_3566,N_2597,N_2109);
nor U3567 (N_3567,N_2106,N_2260);
nand U3568 (N_3568,N_2118,N_2417);
nand U3569 (N_3569,N_2650,N_2822);
or U3570 (N_3570,N_2707,N_2761);
and U3571 (N_3571,N_2440,N_2549);
nand U3572 (N_3572,N_2652,N_2038);
or U3573 (N_3573,N_2996,N_2109);
or U3574 (N_3574,N_2736,N_2399);
and U3575 (N_3575,N_2417,N_2501);
nor U3576 (N_3576,N_2620,N_2344);
nor U3577 (N_3577,N_2226,N_2639);
xor U3578 (N_3578,N_2358,N_2649);
nand U3579 (N_3579,N_2835,N_2107);
nor U3580 (N_3580,N_2353,N_2739);
or U3581 (N_3581,N_2558,N_2382);
nand U3582 (N_3582,N_2674,N_2890);
and U3583 (N_3583,N_2406,N_2454);
or U3584 (N_3584,N_2126,N_2003);
nor U3585 (N_3585,N_2811,N_2263);
nand U3586 (N_3586,N_2264,N_2600);
and U3587 (N_3587,N_2153,N_2329);
xnor U3588 (N_3588,N_2681,N_2869);
or U3589 (N_3589,N_2627,N_2097);
nand U3590 (N_3590,N_2659,N_2440);
nand U3591 (N_3591,N_2726,N_2851);
nor U3592 (N_3592,N_2513,N_2856);
xnor U3593 (N_3593,N_2446,N_2477);
nand U3594 (N_3594,N_2465,N_2642);
nand U3595 (N_3595,N_2758,N_2699);
and U3596 (N_3596,N_2029,N_2815);
nand U3597 (N_3597,N_2771,N_2465);
or U3598 (N_3598,N_2044,N_2233);
and U3599 (N_3599,N_2770,N_2337);
nand U3600 (N_3600,N_2115,N_2327);
or U3601 (N_3601,N_2221,N_2366);
nor U3602 (N_3602,N_2029,N_2926);
nand U3603 (N_3603,N_2090,N_2374);
nor U3604 (N_3604,N_2976,N_2671);
nand U3605 (N_3605,N_2658,N_2646);
or U3606 (N_3606,N_2546,N_2007);
and U3607 (N_3607,N_2982,N_2498);
and U3608 (N_3608,N_2817,N_2674);
and U3609 (N_3609,N_2658,N_2243);
nor U3610 (N_3610,N_2632,N_2549);
or U3611 (N_3611,N_2689,N_2003);
nor U3612 (N_3612,N_2996,N_2635);
nand U3613 (N_3613,N_2577,N_2920);
and U3614 (N_3614,N_2162,N_2138);
nor U3615 (N_3615,N_2595,N_2504);
nor U3616 (N_3616,N_2031,N_2378);
nor U3617 (N_3617,N_2087,N_2001);
nor U3618 (N_3618,N_2309,N_2115);
nand U3619 (N_3619,N_2787,N_2101);
nand U3620 (N_3620,N_2166,N_2217);
nand U3621 (N_3621,N_2933,N_2299);
and U3622 (N_3622,N_2396,N_2446);
nand U3623 (N_3623,N_2528,N_2996);
and U3624 (N_3624,N_2149,N_2659);
and U3625 (N_3625,N_2095,N_2791);
nand U3626 (N_3626,N_2213,N_2965);
nand U3627 (N_3627,N_2298,N_2283);
nand U3628 (N_3628,N_2376,N_2488);
and U3629 (N_3629,N_2761,N_2506);
nand U3630 (N_3630,N_2369,N_2367);
nand U3631 (N_3631,N_2917,N_2745);
and U3632 (N_3632,N_2509,N_2163);
nand U3633 (N_3633,N_2360,N_2361);
nand U3634 (N_3634,N_2412,N_2879);
nand U3635 (N_3635,N_2471,N_2375);
and U3636 (N_3636,N_2322,N_2339);
or U3637 (N_3637,N_2787,N_2703);
or U3638 (N_3638,N_2089,N_2145);
nor U3639 (N_3639,N_2211,N_2529);
or U3640 (N_3640,N_2148,N_2193);
or U3641 (N_3641,N_2278,N_2573);
nor U3642 (N_3642,N_2668,N_2982);
nand U3643 (N_3643,N_2705,N_2396);
nor U3644 (N_3644,N_2897,N_2265);
or U3645 (N_3645,N_2909,N_2225);
nand U3646 (N_3646,N_2115,N_2268);
nand U3647 (N_3647,N_2846,N_2578);
nor U3648 (N_3648,N_2424,N_2922);
and U3649 (N_3649,N_2405,N_2892);
or U3650 (N_3650,N_2269,N_2102);
or U3651 (N_3651,N_2369,N_2516);
nor U3652 (N_3652,N_2600,N_2851);
nor U3653 (N_3653,N_2495,N_2742);
and U3654 (N_3654,N_2147,N_2472);
xor U3655 (N_3655,N_2893,N_2661);
or U3656 (N_3656,N_2839,N_2918);
nand U3657 (N_3657,N_2209,N_2656);
and U3658 (N_3658,N_2076,N_2199);
nand U3659 (N_3659,N_2392,N_2473);
and U3660 (N_3660,N_2353,N_2926);
nor U3661 (N_3661,N_2181,N_2478);
nand U3662 (N_3662,N_2295,N_2440);
and U3663 (N_3663,N_2088,N_2572);
or U3664 (N_3664,N_2806,N_2627);
nand U3665 (N_3665,N_2906,N_2792);
nor U3666 (N_3666,N_2669,N_2351);
or U3667 (N_3667,N_2734,N_2254);
and U3668 (N_3668,N_2670,N_2320);
or U3669 (N_3669,N_2260,N_2250);
and U3670 (N_3670,N_2382,N_2069);
nand U3671 (N_3671,N_2814,N_2181);
xor U3672 (N_3672,N_2076,N_2816);
nor U3673 (N_3673,N_2054,N_2727);
and U3674 (N_3674,N_2195,N_2754);
nor U3675 (N_3675,N_2844,N_2120);
nor U3676 (N_3676,N_2182,N_2628);
and U3677 (N_3677,N_2954,N_2776);
xor U3678 (N_3678,N_2229,N_2496);
nor U3679 (N_3679,N_2711,N_2941);
and U3680 (N_3680,N_2121,N_2243);
or U3681 (N_3681,N_2600,N_2270);
nor U3682 (N_3682,N_2420,N_2218);
and U3683 (N_3683,N_2503,N_2364);
nor U3684 (N_3684,N_2351,N_2353);
or U3685 (N_3685,N_2106,N_2497);
nor U3686 (N_3686,N_2091,N_2176);
or U3687 (N_3687,N_2171,N_2963);
nand U3688 (N_3688,N_2625,N_2300);
and U3689 (N_3689,N_2461,N_2276);
nor U3690 (N_3690,N_2028,N_2430);
nand U3691 (N_3691,N_2459,N_2958);
and U3692 (N_3692,N_2346,N_2588);
or U3693 (N_3693,N_2275,N_2352);
nand U3694 (N_3694,N_2705,N_2181);
nor U3695 (N_3695,N_2300,N_2744);
or U3696 (N_3696,N_2888,N_2996);
or U3697 (N_3697,N_2404,N_2487);
and U3698 (N_3698,N_2880,N_2637);
xor U3699 (N_3699,N_2786,N_2848);
and U3700 (N_3700,N_2042,N_2236);
nor U3701 (N_3701,N_2529,N_2940);
and U3702 (N_3702,N_2116,N_2201);
and U3703 (N_3703,N_2598,N_2790);
or U3704 (N_3704,N_2415,N_2156);
nor U3705 (N_3705,N_2823,N_2661);
or U3706 (N_3706,N_2911,N_2901);
or U3707 (N_3707,N_2207,N_2936);
or U3708 (N_3708,N_2752,N_2459);
nand U3709 (N_3709,N_2200,N_2495);
nand U3710 (N_3710,N_2161,N_2561);
nand U3711 (N_3711,N_2943,N_2118);
nand U3712 (N_3712,N_2774,N_2586);
nand U3713 (N_3713,N_2085,N_2524);
and U3714 (N_3714,N_2710,N_2324);
xnor U3715 (N_3715,N_2579,N_2893);
nor U3716 (N_3716,N_2576,N_2725);
nor U3717 (N_3717,N_2168,N_2429);
nor U3718 (N_3718,N_2531,N_2721);
and U3719 (N_3719,N_2062,N_2662);
nand U3720 (N_3720,N_2698,N_2238);
or U3721 (N_3721,N_2000,N_2358);
nor U3722 (N_3722,N_2248,N_2018);
nor U3723 (N_3723,N_2003,N_2488);
nor U3724 (N_3724,N_2903,N_2451);
nand U3725 (N_3725,N_2256,N_2706);
xnor U3726 (N_3726,N_2955,N_2303);
nor U3727 (N_3727,N_2386,N_2774);
nand U3728 (N_3728,N_2377,N_2493);
and U3729 (N_3729,N_2605,N_2276);
nor U3730 (N_3730,N_2010,N_2611);
or U3731 (N_3731,N_2085,N_2936);
or U3732 (N_3732,N_2364,N_2369);
nor U3733 (N_3733,N_2988,N_2297);
and U3734 (N_3734,N_2451,N_2604);
nor U3735 (N_3735,N_2642,N_2054);
nand U3736 (N_3736,N_2972,N_2845);
nor U3737 (N_3737,N_2816,N_2421);
nor U3738 (N_3738,N_2652,N_2897);
and U3739 (N_3739,N_2462,N_2821);
xor U3740 (N_3740,N_2336,N_2418);
xor U3741 (N_3741,N_2239,N_2456);
and U3742 (N_3742,N_2176,N_2006);
or U3743 (N_3743,N_2147,N_2874);
and U3744 (N_3744,N_2454,N_2042);
nor U3745 (N_3745,N_2820,N_2395);
nand U3746 (N_3746,N_2507,N_2198);
nand U3747 (N_3747,N_2666,N_2542);
nand U3748 (N_3748,N_2907,N_2536);
and U3749 (N_3749,N_2935,N_2430);
and U3750 (N_3750,N_2887,N_2975);
or U3751 (N_3751,N_2407,N_2889);
or U3752 (N_3752,N_2663,N_2709);
nor U3753 (N_3753,N_2155,N_2138);
nor U3754 (N_3754,N_2340,N_2283);
and U3755 (N_3755,N_2071,N_2304);
xnor U3756 (N_3756,N_2826,N_2239);
and U3757 (N_3757,N_2207,N_2523);
nor U3758 (N_3758,N_2959,N_2756);
nor U3759 (N_3759,N_2128,N_2014);
nor U3760 (N_3760,N_2989,N_2878);
and U3761 (N_3761,N_2144,N_2593);
and U3762 (N_3762,N_2554,N_2222);
nor U3763 (N_3763,N_2568,N_2015);
nand U3764 (N_3764,N_2716,N_2277);
and U3765 (N_3765,N_2074,N_2697);
or U3766 (N_3766,N_2947,N_2667);
and U3767 (N_3767,N_2374,N_2238);
and U3768 (N_3768,N_2964,N_2671);
or U3769 (N_3769,N_2319,N_2746);
xnor U3770 (N_3770,N_2691,N_2348);
nor U3771 (N_3771,N_2196,N_2503);
or U3772 (N_3772,N_2601,N_2248);
or U3773 (N_3773,N_2186,N_2416);
or U3774 (N_3774,N_2960,N_2526);
nor U3775 (N_3775,N_2808,N_2433);
nand U3776 (N_3776,N_2913,N_2268);
nor U3777 (N_3777,N_2681,N_2452);
or U3778 (N_3778,N_2317,N_2098);
and U3779 (N_3779,N_2488,N_2982);
or U3780 (N_3780,N_2245,N_2317);
nor U3781 (N_3781,N_2678,N_2190);
nor U3782 (N_3782,N_2997,N_2540);
nor U3783 (N_3783,N_2781,N_2735);
nor U3784 (N_3784,N_2350,N_2960);
and U3785 (N_3785,N_2943,N_2985);
and U3786 (N_3786,N_2362,N_2080);
and U3787 (N_3787,N_2096,N_2214);
or U3788 (N_3788,N_2582,N_2922);
nand U3789 (N_3789,N_2220,N_2047);
nand U3790 (N_3790,N_2047,N_2957);
and U3791 (N_3791,N_2014,N_2764);
or U3792 (N_3792,N_2832,N_2527);
nand U3793 (N_3793,N_2664,N_2997);
nor U3794 (N_3794,N_2073,N_2773);
nand U3795 (N_3795,N_2087,N_2684);
and U3796 (N_3796,N_2772,N_2712);
or U3797 (N_3797,N_2343,N_2619);
or U3798 (N_3798,N_2249,N_2230);
or U3799 (N_3799,N_2896,N_2501);
nor U3800 (N_3800,N_2813,N_2595);
nand U3801 (N_3801,N_2511,N_2961);
nand U3802 (N_3802,N_2335,N_2629);
and U3803 (N_3803,N_2616,N_2781);
nand U3804 (N_3804,N_2922,N_2777);
or U3805 (N_3805,N_2197,N_2697);
nor U3806 (N_3806,N_2082,N_2081);
nor U3807 (N_3807,N_2989,N_2285);
nor U3808 (N_3808,N_2598,N_2049);
nor U3809 (N_3809,N_2011,N_2821);
xor U3810 (N_3810,N_2453,N_2194);
nor U3811 (N_3811,N_2489,N_2601);
and U3812 (N_3812,N_2631,N_2799);
nor U3813 (N_3813,N_2501,N_2720);
nand U3814 (N_3814,N_2700,N_2006);
nand U3815 (N_3815,N_2023,N_2711);
nor U3816 (N_3816,N_2858,N_2983);
nor U3817 (N_3817,N_2915,N_2661);
nor U3818 (N_3818,N_2470,N_2306);
and U3819 (N_3819,N_2773,N_2996);
nand U3820 (N_3820,N_2859,N_2314);
or U3821 (N_3821,N_2248,N_2387);
or U3822 (N_3822,N_2457,N_2948);
nand U3823 (N_3823,N_2901,N_2360);
or U3824 (N_3824,N_2430,N_2486);
or U3825 (N_3825,N_2130,N_2294);
nor U3826 (N_3826,N_2646,N_2578);
xor U3827 (N_3827,N_2820,N_2258);
or U3828 (N_3828,N_2084,N_2557);
and U3829 (N_3829,N_2407,N_2835);
and U3830 (N_3830,N_2471,N_2611);
nand U3831 (N_3831,N_2230,N_2161);
and U3832 (N_3832,N_2185,N_2374);
nor U3833 (N_3833,N_2091,N_2494);
nand U3834 (N_3834,N_2777,N_2838);
nand U3835 (N_3835,N_2481,N_2726);
and U3836 (N_3836,N_2165,N_2292);
or U3837 (N_3837,N_2423,N_2891);
or U3838 (N_3838,N_2221,N_2032);
and U3839 (N_3839,N_2667,N_2010);
nand U3840 (N_3840,N_2405,N_2956);
nand U3841 (N_3841,N_2578,N_2494);
nand U3842 (N_3842,N_2150,N_2079);
and U3843 (N_3843,N_2656,N_2411);
nand U3844 (N_3844,N_2545,N_2603);
nand U3845 (N_3845,N_2102,N_2736);
or U3846 (N_3846,N_2838,N_2546);
and U3847 (N_3847,N_2018,N_2873);
and U3848 (N_3848,N_2574,N_2977);
nand U3849 (N_3849,N_2800,N_2033);
and U3850 (N_3850,N_2246,N_2425);
and U3851 (N_3851,N_2166,N_2968);
and U3852 (N_3852,N_2428,N_2710);
and U3853 (N_3853,N_2651,N_2395);
or U3854 (N_3854,N_2916,N_2928);
nand U3855 (N_3855,N_2396,N_2948);
or U3856 (N_3856,N_2156,N_2501);
or U3857 (N_3857,N_2765,N_2214);
and U3858 (N_3858,N_2240,N_2923);
and U3859 (N_3859,N_2561,N_2788);
or U3860 (N_3860,N_2219,N_2417);
and U3861 (N_3861,N_2038,N_2186);
or U3862 (N_3862,N_2150,N_2284);
nand U3863 (N_3863,N_2219,N_2089);
or U3864 (N_3864,N_2431,N_2990);
or U3865 (N_3865,N_2434,N_2363);
nand U3866 (N_3866,N_2658,N_2898);
or U3867 (N_3867,N_2613,N_2988);
nand U3868 (N_3868,N_2489,N_2968);
or U3869 (N_3869,N_2669,N_2151);
nand U3870 (N_3870,N_2049,N_2609);
and U3871 (N_3871,N_2173,N_2731);
nand U3872 (N_3872,N_2054,N_2706);
or U3873 (N_3873,N_2085,N_2844);
nor U3874 (N_3874,N_2495,N_2906);
and U3875 (N_3875,N_2605,N_2546);
nand U3876 (N_3876,N_2703,N_2598);
or U3877 (N_3877,N_2257,N_2737);
nand U3878 (N_3878,N_2149,N_2539);
or U3879 (N_3879,N_2892,N_2668);
and U3880 (N_3880,N_2118,N_2401);
and U3881 (N_3881,N_2834,N_2266);
nor U3882 (N_3882,N_2337,N_2863);
nand U3883 (N_3883,N_2095,N_2727);
and U3884 (N_3884,N_2376,N_2838);
or U3885 (N_3885,N_2236,N_2484);
and U3886 (N_3886,N_2809,N_2662);
or U3887 (N_3887,N_2093,N_2122);
or U3888 (N_3888,N_2573,N_2658);
xor U3889 (N_3889,N_2679,N_2758);
nand U3890 (N_3890,N_2001,N_2212);
nor U3891 (N_3891,N_2979,N_2961);
and U3892 (N_3892,N_2472,N_2413);
nand U3893 (N_3893,N_2483,N_2063);
or U3894 (N_3894,N_2097,N_2205);
nor U3895 (N_3895,N_2246,N_2987);
or U3896 (N_3896,N_2974,N_2426);
and U3897 (N_3897,N_2254,N_2104);
or U3898 (N_3898,N_2793,N_2807);
or U3899 (N_3899,N_2853,N_2519);
nand U3900 (N_3900,N_2728,N_2229);
nor U3901 (N_3901,N_2356,N_2703);
and U3902 (N_3902,N_2198,N_2537);
nand U3903 (N_3903,N_2973,N_2214);
nand U3904 (N_3904,N_2355,N_2615);
nor U3905 (N_3905,N_2686,N_2956);
nand U3906 (N_3906,N_2152,N_2129);
or U3907 (N_3907,N_2313,N_2686);
and U3908 (N_3908,N_2381,N_2198);
and U3909 (N_3909,N_2318,N_2069);
or U3910 (N_3910,N_2243,N_2879);
and U3911 (N_3911,N_2020,N_2492);
nor U3912 (N_3912,N_2014,N_2040);
nand U3913 (N_3913,N_2021,N_2137);
nor U3914 (N_3914,N_2097,N_2838);
nor U3915 (N_3915,N_2521,N_2262);
nand U3916 (N_3916,N_2361,N_2877);
nand U3917 (N_3917,N_2067,N_2820);
nor U3918 (N_3918,N_2013,N_2463);
nor U3919 (N_3919,N_2543,N_2961);
and U3920 (N_3920,N_2203,N_2533);
nand U3921 (N_3921,N_2191,N_2629);
nand U3922 (N_3922,N_2712,N_2880);
and U3923 (N_3923,N_2382,N_2712);
or U3924 (N_3924,N_2562,N_2298);
or U3925 (N_3925,N_2636,N_2497);
nand U3926 (N_3926,N_2209,N_2065);
or U3927 (N_3927,N_2490,N_2975);
nor U3928 (N_3928,N_2207,N_2021);
nor U3929 (N_3929,N_2361,N_2347);
nor U3930 (N_3930,N_2589,N_2024);
nand U3931 (N_3931,N_2567,N_2368);
and U3932 (N_3932,N_2145,N_2126);
and U3933 (N_3933,N_2482,N_2052);
and U3934 (N_3934,N_2463,N_2476);
or U3935 (N_3935,N_2459,N_2082);
or U3936 (N_3936,N_2525,N_2031);
and U3937 (N_3937,N_2645,N_2789);
nand U3938 (N_3938,N_2794,N_2380);
nand U3939 (N_3939,N_2590,N_2322);
or U3940 (N_3940,N_2995,N_2666);
and U3941 (N_3941,N_2828,N_2195);
nor U3942 (N_3942,N_2630,N_2838);
nor U3943 (N_3943,N_2143,N_2327);
nor U3944 (N_3944,N_2163,N_2220);
and U3945 (N_3945,N_2456,N_2748);
nand U3946 (N_3946,N_2628,N_2214);
nor U3947 (N_3947,N_2285,N_2200);
nor U3948 (N_3948,N_2103,N_2843);
nand U3949 (N_3949,N_2507,N_2825);
or U3950 (N_3950,N_2006,N_2883);
nand U3951 (N_3951,N_2843,N_2347);
nand U3952 (N_3952,N_2092,N_2209);
nand U3953 (N_3953,N_2171,N_2897);
and U3954 (N_3954,N_2265,N_2111);
nor U3955 (N_3955,N_2991,N_2894);
or U3956 (N_3956,N_2375,N_2549);
nand U3957 (N_3957,N_2842,N_2660);
nand U3958 (N_3958,N_2353,N_2180);
nand U3959 (N_3959,N_2943,N_2408);
and U3960 (N_3960,N_2173,N_2667);
nor U3961 (N_3961,N_2415,N_2089);
nor U3962 (N_3962,N_2890,N_2019);
nor U3963 (N_3963,N_2560,N_2311);
and U3964 (N_3964,N_2060,N_2640);
nor U3965 (N_3965,N_2007,N_2190);
or U3966 (N_3966,N_2240,N_2560);
nand U3967 (N_3967,N_2056,N_2022);
and U3968 (N_3968,N_2596,N_2985);
nand U3969 (N_3969,N_2591,N_2439);
nand U3970 (N_3970,N_2245,N_2374);
or U3971 (N_3971,N_2030,N_2311);
nand U3972 (N_3972,N_2856,N_2862);
and U3973 (N_3973,N_2237,N_2616);
nor U3974 (N_3974,N_2073,N_2647);
or U3975 (N_3975,N_2649,N_2217);
nand U3976 (N_3976,N_2681,N_2050);
or U3977 (N_3977,N_2175,N_2162);
xnor U3978 (N_3978,N_2670,N_2464);
and U3979 (N_3979,N_2251,N_2641);
and U3980 (N_3980,N_2517,N_2099);
xnor U3981 (N_3981,N_2860,N_2837);
nor U3982 (N_3982,N_2677,N_2791);
and U3983 (N_3983,N_2716,N_2403);
nor U3984 (N_3984,N_2105,N_2530);
and U3985 (N_3985,N_2550,N_2621);
nand U3986 (N_3986,N_2223,N_2306);
nor U3987 (N_3987,N_2707,N_2759);
and U3988 (N_3988,N_2319,N_2889);
or U3989 (N_3989,N_2730,N_2665);
and U3990 (N_3990,N_2283,N_2228);
nor U3991 (N_3991,N_2070,N_2692);
and U3992 (N_3992,N_2368,N_2050);
nand U3993 (N_3993,N_2691,N_2526);
or U3994 (N_3994,N_2166,N_2454);
nor U3995 (N_3995,N_2537,N_2164);
and U3996 (N_3996,N_2188,N_2241);
and U3997 (N_3997,N_2933,N_2128);
nor U3998 (N_3998,N_2241,N_2409);
nand U3999 (N_3999,N_2665,N_2237);
nand U4000 (N_4000,N_3969,N_3475);
nor U4001 (N_4001,N_3585,N_3326);
or U4002 (N_4002,N_3520,N_3164);
nand U4003 (N_4003,N_3329,N_3421);
nand U4004 (N_4004,N_3111,N_3627);
or U4005 (N_4005,N_3407,N_3169);
or U4006 (N_4006,N_3967,N_3268);
or U4007 (N_4007,N_3492,N_3124);
xor U4008 (N_4008,N_3256,N_3479);
nand U4009 (N_4009,N_3104,N_3952);
nor U4010 (N_4010,N_3081,N_3241);
or U4011 (N_4011,N_3198,N_3537);
nor U4012 (N_4012,N_3675,N_3197);
nor U4013 (N_4013,N_3316,N_3708);
xnor U4014 (N_4014,N_3784,N_3626);
and U4015 (N_4015,N_3714,N_3925);
and U4016 (N_4016,N_3077,N_3348);
and U4017 (N_4017,N_3338,N_3002);
nor U4018 (N_4018,N_3828,N_3785);
nor U4019 (N_4019,N_3181,N_3919);
or U4020 (N_4020,N_3279,N_3194);
or U4021 (N_4021,N_3861,N_3078);
and U4022 (N_4022,N_3090,N_3727);
or U4023 (N_4023,N_3245,N_3551);
nor U4024 (N_4024,N_3362,N_3143);
nand U4025 (N_4025,N_3762,N_3936);
nor U4026 (N_4026,N_3183,N_3100);
or U4027 (N_4027,N_3232,N_3276);
nor U4028 (N_4028,N_3655,N_3607);
nand U4029 (N_4029,N_3014,N_3695);
nor U4030 (N_4030,N_3435,N_3021);
nand U4031 (N_4031,N_3017,N_3712);
nand U4032 (N_4032,N_3039,N_3775);
and U4033 (N_4033,N_3909,N_3369);
or U4034 (N_4034,N_3820,N_3176);
or U4035 (N_4035,N_3765,N_3796);
nor U4036 (N_4036,N_3223,N_3290);
and U4037 (N_4037,N_3965,N_3233);
nor U4038 (N_4038,N_3532,N_3360);
nand U4039 (N_4039,N_3342,N_3953);
and U4040 (N_4040,N_3476,N_3167);
nand U4041 (N_4041,N_3343,N_3050);
nor U4042 (N_4042,N_3672,N_3184);
or U4043 (N_4043,N_3071,N_3844);
nor U4044 (N_4044,N_3696,N_3751);
or U4045 (N_4045,N_3347,N_3452);
nor U4046 (N_4046,N_3913,N_3653);
nand U4047 (N_4047,N_3313,N_3154);
nand U4048 (N_4048,N_3906,N_3069);
nor U4049 (N_4049,N_3892,N_3526);
and U4050 (N_4050,N_3036,N_3642);
and U4051 (N_4051,N_3063,N_3240);
or U4052 (N_4052,N_3948,N_3266);
nand U4053 (N_4053,N_3257,N_3331);
nand U4054 (N_4054,N_3987,N_3150);
and U4055 (N_4055,N_3140,N_3383);
nand U4056 (N_4056,N_3813,N_3157);
nand U4057 (N_4057,N_3064,N_3651);
or U4058 (N_4058,N_3344,N_3898);
nand U4059 (N_4059,N_3885,N_3778);
xor U4060 (N_4060,N_3067,N_3195);
nand U4061 (N_4061,N_3450,N_3959);
and U4062 (N_4062,N_3059,N_3246);
nand U4063 (N_4063,N_3022,N_3776);
nor U4064 (N_4064,N_3399,N_3750);
nor U4065 (N_4065,N_3589,N_3384);
and U4066 (N_4066,N_3699,N_3193);
or U4067 (N_4067,N_3519,N_3262);
nand U4068 (N_4068,N_3267,N_3875);
nand U4069 (N_4069,N_3380,N_3853);
and U4070 (N_4070,N_3337,N_3464);
and U4071 (N_4071,N_3949,N_3920);
and U4072 (N_4072,N_3872,N_3914);
or U4073 (N_4073,N_3471,N_3812);
nand U4074 (N_4074,N_3504,N_3503);
and U4075 (N_4075,N_3336,N_3349);
and U4076 (N_4076,N_3971,N_3145);
and U4077 (N_4077,N_3803,N_3698);
and U4078 (N_4078,N_3926,N_3204);
nand U4079 (N_4079,N_3320,N_3954);
nand U4080 (N_4080,N_3544,N_3229);
nor U4081 (N_4081,N_3173,N_3260);
and U4082 (N_4082,N_3402,N_3951);
and U4083 (N_4083,N_3355,N_3255);
and U4084 (N_4084,N_3187,N_3249);
or U4085 (N_4085,N_3190,N_3389);
or U4086 (N_4086,N_3112,N_3568);
and U4087 (N_4087,N_3740,N_3060);
nor U4088 (N_4088,N_3427,N_3049);
and U4089 (N_4089,N_3016,N_3999);
and U4090 (N_4090,N_3066,N_3702);
and U4091 (N_4091,N_3045,N_3841);
or U4092 (N_4092,N_3613,N_3174);
and U4093 (N_4093,N_3908,N_3935);
xor U4094 (N_4094,N_3263,N_3426);
nor U4095 (N_4095,N_3089,N_3917);
or U4096 (N_4096,N_3725,N_3911);
nor U4097 (N_4097,N_3284,N_3491);
nand U4098 (N_4098,N_3324,N_3700);
and U4099 (N_4099,N_3634,N_3274);
nor U4100 (N_4100,N_3603,N_3583);
or U4101 (N_4101,N_3390,N_3761);
xor U4102 (N_4102,N_3010,N_3024);
nor U4103 (N_4103,N_3946,N_3582);
nand U4104 (N_4104,N_3618,N_3110);
or U4105 (N_4105,N_3494,N_3735);
and U4106 (N_4106,N_3298,N_3625);
and U4107 (N_4107,N_3209,N_3561);
nand U4108 (N_4108,N_3545,N_3990);
and U4109 (N_4109,N_3644,N_3539);
nor U4110 (N_4110,N_3300,N_3612);
and U4111 (N_4111,N_3810,N_3213);
and U4112 (N_4112,N_3029,N_3599);
nand U4113 (N_4113,N_3217,N_3447);
nor U4114 (N_4114,N_3912,N_3535);
nand U4115 (N_4115,N_3522,N_3474);
nand U4116 (N_4116,N_3448,N_3608);
or U4117 (N_4117,N_3837,N_3147);
and U4118 (N_4118,N_3887,N_3648);
and U4119 (N_4119,N_3604,N_3117);
and U4120 (N_4120,N_3947,N_3499);
nor U4121 (N_4121,N_3053,N_3681);
or U4122 (N_4122,N_3477,N_3172);
nand U4123 (N_4123,N_3554,N_3871);
nor U4124 (N_4124,N_3941,N_3731);
or U4125 (N_4125,N_3856,N_3107);
or U4126 (N_4126,N_3034,N_3557);
nor U4127 (N_4127,N_3040,N_3170);
and U4128 (N_4128,N_3786,N_3849);
nor U4129 (N_4129,N_3905,N_3596);
and U4130 (N_4130,N_3701,N_3317);
nor U4131 (N_4131,N_3955,N_3041);
or U4132 (N_4132,N_3141,N_3674);
and U4133 (N_4133,N_3543,N_3753);
nand U4134 (N_4134,N_3839,N_3237);
or U4135 (N_4135,N_3883,N_3026);
nand U4136 (N_4136,N_3662,N_3381);
and U4137 (N_4137,N_3822,N_3834);
nand U4138 (N_4138,N_3502,N_3253);
or U4139 (N_4139,N_3549,N_3079);
or U4140 (N_4140,N_3845,N_3496);
and U4141 (N_4141,N_3848,N_3556);
nor U4142 (N_4142,N_3484,N_3802);
nand U4143 (N_4143,N_3322,N_3231);
nor U4144 (N_4144,N_3043,N_3523);
nand U4145 (N_4145,N_3118,N_3835);
nor U4146 (N_4146,N_3904,N_3061);
nand U4147 (N_4147,N_3414,N_3606);
nand U4148 (N_4148,N_3437,N_3244);
and U4149 (N_4149,N_3033,N_3619);
and U4150 (N_4150,N_3028,N_3308);
nand U4151 (N_4151,N_3108,N_3005);
nor U4152 (N_4152,N_3921,N_3306);
nor U4153 (N_4153,N_3594,N_3646);
nor U4154 (N_4154,N_3472,N_3062);
nand U4155 (N_4155,N_3149,N_3956);
or U4156 (N_4156,N_3873,N_3424);
or U4157 (N_4157,N_3972,N_3465);
nand U4158 (N_4158,N_3610,N_3046);
or U4159 (N_4159,N_3756,N_3558);
xnor U4160 (N_4160,N_3483,N_3962);
or U4161 (N_4161,N_3098,N_3983);
or U4162 (N_4162,N_3616,N_3763);
or U4163 (N_4163,N_3964,N_3710);
nand U4164 (N_4164,N_3467,N_3457);
or U4165 (N_4165,N_3481,N_3534);
nor U4166 (N_4166,N_3927,N_3746);
and U4167 (N_4167,N_3995,N_3893);
or U4168 (N_4168,N_3304,N_3752);
nand U4169 (N_4169,N_3311,N_3418);
or U4170 (N_4170,N_3718,N_3628);
nor U4171 (N_4171,N_3413,N_3321);
and U4172 (N_4172,N_3876,N_3470);
nand U4173 (N_4173,N_3547,N_3131);
and U4174 (N_4174,N_3023,N_3823);
and U4175 (N_4175,N_3092,N_3747);
or U4176 (N_4176,N_3272,N_3333);
or U4177 (N_4177,N_3278,N_3048);
nor U4178 (N_4178,N_3720,N_3387);
or U4179 (N_4179,N_3236,N_3847);
and U4180 (N_4180,N_3136,N_3259);
nand U4181 (N_4181,N_3722,N_3570);
nand U4182 (N_4182,N_3189,N_3728);
nand U4183 (N_4183,N_3388,N_3215);
nor U4184 (N_4184,N_3391,N_3573);
or U4185 (N_4185,N_3461,N_3637);
nand U4186 (N_4186,N_3766,N_3989);
nor U4187 (N_4187,N_3578,N_3431);
nor U4188 (N_4188,N_3992,N_3374);
and U4189 (N_4189,N_3264,N_3788);
nand U4190 (N_4190,N_3487,N_3711);
and U4191 (N_4191,N_3564,N_3030);
nand U4192 (N_4192,N_3423,N_3091);
nand U4193 (N_4193,N_3428,N_3678);
nand U4194 (N_4194,N_3975,N_3748);
or U4195 (N_4195,N_3175,N_3218);
or U4196 (N_4196,N_3439,N_3351);
or U4197 (N_4197,N_3797,N_3515);
and U4198 (N_4198,N_3000,N_3622);
nand U4199 (N_4199,N_3006,N_3196);
or U4200 (N_4200,N_3665,N_3130);
nand U4201 (N_4201,N_3212,N_3799);
or U4202 (N_4202,N_3162,N_3758);
and U4203 (N_4203,N_3417,N_3330);
and U4204 (N_4204,N_3996,N_3840);
or U4205 (N_4205,N_3047,N_3392);
or U4206 (N_4206,N_3986,N_3295);
and U4207 (N_4207,N_3770,N_3393);
and U4208 (N_4208,N_3726,N_3134);
xnor U4209 (N_4209,N_3035,N_3357);
nand U4210 (N_4210,N_3419,N_3716);
nand U4211 (N_4211,N_3531,N_3787);
and U4212 (N_4212,N_3782,N_3930);
nand U4213 (N_4213,N_3307,N_3806);
nand U4214 (N_4214,N_3303,N_3654);
and U4215 (N_4215,N_3121,N_3151);
and U4216 (N_4216,N_3283,N_3888);
or U4217 (N_4217,N_3294,N_3230);
nand U4218 (N_4218,N_3025,N_3924);
or U4219 (N_4219,N_3656,N_3445);
nor U4220 (N_4220,N_3692,N_3238);
and U4221 (N_4221,N_3186,N_3404);
or U4222 (N_4222,N_3314,N_3895);
or U4223 (N_4223,N_3354,N_3824);
nand U4224 (N_4224,N_3182,N_3635);
or U4225 (N_4225,N_3070,N_3301);
nand U4226 (N_4226,N_3395,N_3243);
and U4227 (N_4227,N_3540,N_3125);
or U4228 (N_4228,N_3833,N_3291);
or U4229 (N_4229,N_3667,N_3438);
xor U4230 (N_4230,N_3693,N_3529);
nor U4231 (N_4231,N_3441,N_3994);
xor U4232 (N_4232,N_3054,N_3730);
nand U4233 (N_4233,N_3817,N_3055);
nand U4234 (N_4234,N_3297,N_3944);
nor U4235 (N_4235,N_3180,N_3816);
and U4236 (N_4236,N_3429,N_3772);
nand U4237 (N_4237,N_3058,N_3072);
or U4238 (N_4238,N_3633,N_3846);
nand U4239 (N_4239,N_3581,N_3500);
nand U4240 (N_4240,N_3292,N_3370);
and U4241 (N_4241,N_3097,N_3736);
nand U4242 (N_4242,N_3270,N_3334);
or U4243 (N_4243,N_3252,N_3783);
nor U4244 (N_4244,N_3598,N_3794);
xnor U4245 (N_4245,N_3790,N_3767);
nor U4246 (N_4246,N_3269,N_3550);
nor U4247 (N_4247,N_3261,N_3670);
or U4248 (N_4248,N_3299,N_3444);
nor U4249 (N_4249,N_3838,N_3528);
nand U4250 (N_4250,N_3814,N_3852);
and U4251 (N_4251,N_3210,N_3660);
or U4252 (N_4252,N_3863,N_3155);
or U4253 (N_4253,N_3168,N_3825);
or U4254 (N_4254,N_3850,N_3469);
nand U4255 (N_4255,N_3979,N_3411);
and U4256 (N_4256,N_3473,N_3680);
nor U4257 (N_4257,N_3051,N_3771);
nor U4258 (N_4258,N_3376,N_3900);
nor U4259 (N_4259,N_3577,N_3982);
nand U4260 (N_4260,N_3829,N_3928);
nor U4261 (N_4261,N_3234,N_3862);
nor U4262 (N_4262,N_3013,N_3569);
and U4263 (N_4263,N_3842,N_3011);
and U4264 (N_4264,N_3372,N_3691);
nor U4265 (N_4265,N_3791,N_3511);
nand U4266 (N_4266,N_3860,N_3517);
nor U4267 (N_4267,N_3724,N_3009);
nor U4268 (N_4268,N_3759,N_3804);
and U4269 (N_4269,N_3076,N_3382);
nor U4270 (N_4270,N_3356,N_3485);
nand U4271 (N_4271,N_3859,N_3942);
and U4272 (N_4272,N_3571,N_3227);
nor U4273 (N_4273,N_3225,N_3074);
nor U4274 (N_4274,N_3205,N_3686);
and U4275 (N_4275,N_3430,N_3880);
and U4276 (N_4276,N_3514,N_3922);
nor U4277 (N_4277,N_3536,N_3934);
nand U4278 (N_4278,N_3340,N_3505);
or U4279 (N_4279,N_3669,N_3588);
and U4280 (N_4280,N_3466,N_3918);
nand U4281 (N_4281,N_3801,N_3741);
or U4282 (N_4282,N_3903,N_3282);
nor U4283 (N_4283,N_3562,N_3401);
nand U4284 (N_4284,N_3617,N_3211);
nand U4285 (N_4285,N_3510,N_3226);
or U4286 (N_4286,N_3386,N_3508);
nor U4287 (N_4287,N_3805,N_3705);
or U4288 (N_4288,N_3614,N_3251);
nor U4289 (N_4289,N_3866,N_3339);
nand U4290 (N_4290,N_3273,N_3530);
or U4291 (N_4291,N_3978,N_3191);
nor U4292 (N_4292,N_3115,N_3289);
nor U4293 (N_4293,N_3285,N_3957);
and U4294 (N_4294,N_3738,N_3658);
nor U4295 (N_4295,N_3102,N_3734);
or U4296 (N_4296,N_3595,N_3302);
nor U4297 (N_4297,N_3683,N_3609);
nand U4298 (N_4298,N_3552,N_3179);
nor U4299 (N_4299,N_3052,N_3615);
or U4300 (N_4300,N_3235,N_3146);
or U4301 (N_4301,N_3984,N_3966);
nand U4302 (N_4302,N_3206,N_3456);
nand U4303 (N_4303,N_3901,N_3083);
nor U4304 (N_4304,N_3968,N_3960);
and U4305 (N_4305,N_3281,N_3165);
nand U4306 (N_4306,N_3855,N_3732);
nor U4307 (N_4307,N_3524,N_3621);
and U4308 (N_4308,N_3629,N_3498);
nor U4309 (N_4309,N_3495,N_3690);
or U4310 (N_4310,N_3403,N_3084);
and U4311 (N_4311,N_3420,N_3601);
nand U4312 (N_4312,N_3915,N_3371);
nor U4313 (N_4313,N_3673,N_3363);
nand U4314 (N_4314,N_3963,N_3798);
nand U4315 (N_4315,N_3793,N_3160);
or U4316 (N_4316,N_3630,N_3129);
nand U4317 (N_4317,N_3684,N_3795);
or U4318 (N_4318,N_3103,N_3042);
and U4319 (N_4319,N_3073,N_3202);
and U4320 (N_4320,N_3398,N_3085);
nor U4321 (N_4321,N_3507,N_3819);
and U4322 (N_4322,N_3088,N_3138);
nor U4323 (N_4323,N_3409,N_3755);
or U4324 (N_4324,N_3961,N_3001);
nor U4325 (N_4325,N_3497,N_3997);
nand U4326 (N_4326,N_3120,N_3639);
and U4327 (N_4327,N_3004,N_3600);
or U4328 (N_4328,N_3153,N_3114);
or U4329 (N_4329,N_3749,N_3265);
nand U4330 (N_4330,N_3199,N_3867);
and U4331 (N_4331,N_3137,N_3542);
and U4332 (N_4332,N_3881,N_3436);
xor U4333 (N_4333,N_3319,N_3572);
or U4334 (N_4334,N_3886,N_3679);
nand U4335 (N_4335,N_3239,N_3038);
nand U4336 (N_4336,N_3706,N_3159);
nor U4337 (N_4337,N_3509,N_3800);
and U4338 (N_4338,N_3988,N_3870);
and U4339 (N_4339,N_3415,N_3099);
or U4340 (N_4340,N_3087,N_3991);
xor U4341 (N_4341,N_3119,N_3777);
nor U4342 (N_4342,N_3451,N_3977);
nor U4343 (N_4343,N_3943,N_3144);
nand U4344 (N_4344,N_3019,N_3275);
and U4345 (N_4345,N_3742,N_3139);
nor U4346 (N_4346,N_3620,N_3332);
and U4347 (N_4347,N_3093,N_3869);
and U4348 (N_4348,N_3425,N_3937);
nor U4349 (N_4349,N_3353,N_3478);
and U4350 (N_4350,N_3567,N_3713);
or U4351 (N_4351,N_3228,N_3768);
nor U4352 (N_4352,N_3432,N_3764);
nor U4353 (N_4353,N_3688,N_3897);
or U4354 (N_4354,N_3541,N_3020);
or U4355 (N_4355,N_3843,N_3327);
or U4356 (N_4356,N_3135,N_3910);
and U4357 (N_4357,N_3396,N_3579);
or U4358 (N_4358,N_3003,N_3152);
nor U4359 (N_4359,N_3488,N_3874);
nand U4360 (N_4360,N_3586,N_3640);
nand U4361 (N_4361,N_3220,N_3224);
nand U4362 (N_4362,N_3821,N_3645);
nand U4363 (N_4363,N_3203,N_3976);
or U4364 (N_4364,N_3780,N_3974);
nor U4365 (N_4365,N_3636,N_3546);
and U4366 (N_4366,N_3493,N_3889);
and U4367 (N_4367,N_3123,N_3468);
or U4368 (N_4368,N_3288,N_3809);
or U4369 (N_4369,N_3221,N_3406);
or U4370 (N_4370,N_3884,N_3280);
and U4371 (N_4371,N_3486,N_3095);
xor U4372 (N_4372,N_3335,N_3566);
nand U4373 (N_4373,N_3985,N_3664);
nor U4374 (N_4374,N_3106,N_3744);
and U4375 (N_4375,N_3075,N_3012);
nand U4376 (N_4376,N_3373,N_3364);
nor U4377 (N_4377,N_3214,N_3027);
xor U4378 (N_4378,N_3757,N_3185);
nor U4379 (N_4379,N_3293,N_3538);
nand U4380 (N_4380,N_3970,N_3201);
nor U4381 (N_4381,N_3826,N_3932);
and U4382 (N_4382,N_3894,N_3341);
nor U4383 (N_4383,N_3703,N_3512);
or U4384 (N_4384,N_3584,N_3148);
or U4385 (N_4385,N_3981,N_3891);
nand U4386 (N_4386,N_3171,N_3080);
and U4387 (N_4387,N_3980,N_3623);
and U4388 (N_4388,N_3328,N_3877);
nor U4389 (N_4389,N_3950,N_3296);
or U4390 (N_4390,N_3807,N_3657);
and U4391 (N_4391,N_3574,N_3774);
nand U4392 (N_4392,N_3717,N_3394);
and U4393 (N_4393,N_3666,N_3525);
nor U4394 (N_4394,N_3808,N_3831);
or U4395 (N_4395,N_3548,N_3832);
or U4396 (N_4396,N_3754,N_3325);
nor U4397 (N_4397,N_3346,N_3133);
or U4398 (N_4398,N_3455,N_3200);
nand U4399 (N_4399,N_3521,N_3709);
nand U4400 (N_4400,N_3707,N_3132);
xnor U4401 (N_4401,N_3410,N_3094);
nor U4402 (N_4402,N_3443,N_3527);
and U4403 (N_4403,N_3449,N_3878);
nor U4404 (N_4404,N_3685,N_3811);
or U4405 (N_4405,N_3359,N_3661);
xnor U4406 (N_4406,N_3652,N_3769);
and U4407 (N_4407,N_3161,N_3649);
or U4408 (N_4408,N_3587,N_3638);
or U4409 (N_4409,N_3434,N_3408);
and U4410 (N_4410,N_3739,N_3659);
and U4411 (N_4411,N_3454,N_3057);
and U4412 (N_4412,N_3453,N_3518);
nand U4413 (N_4413,N_3086,N_3597);
nand U4414 (N_4414,N_3254,N_3694);
nor U4415 (N_4415,N_3459,N_3361);
nor U4416 (N_4416,N_3007,N_3575);
and U4417 (N_4417,N_3676,N_3277);
nor U4418 (N_4418,N_3126,N_3533);
and U4419 (N_4419,N_3858,N_3385);
nor U4420 (N_4420,N_3643,N_3258);
and U4421 (N_4421,N_3938,N_3591);
or U4422 (N_4422,N_3632,N_3851);
or U4423 (N_4423,N_3056,N_3737);
and U4424 (N_4424,N_3032,N_3400);
and U4425 (N_4425,N_3250,N_3365);
or U4426 (N_4426,N_3216,N_3318);
nand U4427 (N_4427,N_3462,N_3611);
nand U4428 (N_4428,N_3939,N_3560);
or U4429 (N_4429,N_3940,N_3433);
nor U4430 (N_4430,N_3677,N_3113);
nor U4431 (N_4431,N_3082,N_3463);
xor U4432 (N_4432,N_3689,N_3177);
or U4433 (N_4433,N_3933,N_3156);
and U4434 (N_4434,N_3178,N_3352);
nand U4435 (N_4435,N_3367,N_3312);
nand U4436 (N_4436,N_3719,N_3580);
or U4437 (N_4437,N_3015,N_3945);
nor U4438 (N_4438,N_3815,N_3907);
nand U4439 (N_4439,N_3854,N_3864);
or U4440 (N_4440,N_3366,N_3163);
and U4441 (N_4441,N_3008,N_3489);
nand U4442 (N_4442,N_3553,N_3687);
nor U4443 (N_4443,N_3368,N_3127);
nand U4444 (N_4444,N_3682,N_3882);
and U4445 (N_4445,N_3779,N_3789);
and U4446 (N_4446,N_3416,N_3641);
or U4447 (N_4447,N_3460,N_3650);
nand U4448 (N_4448,N_3375,N_3101);
and U4449 (N_4449,N_3902,N_3222);
and U4450 (N_4450,N_3890,N_3379);
xnor U4451 (N_4451,N_3310,N_3248);
or U4452 (N_4452,N_3105,N_3733);
or U4453 (N_4453,N_3490,N_3315);
or U4454 (N_4454,N_3745,N_3973);
or U4455 (N_4455,N_3242,N_3482);
or U4456 (N_4456,N_3458,N_3576);
or U4457 (N_4457,N_3422,N_3096);
or U4458 (N_4458,N_3513,N_3593);
or U4459 (N_4459,N_3836,N_3697);
or U4460 (N_4460,N_3286,N_3590);
and U4461 (N_4461,N_3309,N_3192);
nand U4462 (N_4462,N_3818,N_3208);
or U4463 (N_4463,N_3555,N_3830);
or U4464 (N_4464,N_3068,N_3345);
nand U4465 (N_4465,N_3715,N_3446);
and U4466 (N_4466,N_3122,N_3506);
nor U4467 (N_4467,N_3031,N_3857);
nor U4468 (N_4468,N_3668,N_3405);
and U4469 (N_4469,N_3868,N_3247);
nand U4470 (N_4470,N_3188,N_3792);
or U4471 (N_4471,N_3602,N_3350);
or U4472 (N_4472,N_3440,N_3412);
and U4473 (N_4473,N_3647,N_3704);
nand U4474 (N_4474,N_3563,N_3305);
nor U4475 (N_4475,N_3219,N_3671);
or U4476 (N_4476,N_3378,N_3879);
nand U4477 (N_4477,N_3018,N_3565);
nand U4478 (N_4478,N_3899,N_3109);
nor U4479 (N_4479,N_3743,N_3480);
or U4480 (N_4480,N_3592,N_3896);
and U4481 (N_4481,N_3929,N_3993);
and U4482 (N_4482,N_3397,N_3916);
and U4483 (N_4483,N_3721,N_3166);
nor U4484 (N_4484,N_3037,N_3781);
and U4485 (N_4485,N_3271,N_3958);
nor U4486 (N_4486,N_3158,N_3729);
nor U4487 (N_4487,N_3760,N_3516);
or U4488 (N_4488,N_3358,N_3663);
or U4489 (N_4489,N_3501,N_3723);
nand U4490 (N_4490,N_3605,N_3207);
nor U4491 (N_4491,N_3559,N_3044);
nand U4492 (N_4492,N_3827,N_3624);
and U4493 (N_4493,N_3065,N_3931);
nand U4494 (N_4494,N_3865,N_3923);
nand U4495 (N_4495,N_3116,N_3377);
and U4496 (N_4496,N_3287,N_3631);
and U4497 (N_4497,N_3442,N_3142);
and U4498 (N_4498,N_3998,N_3773);
or U4499 (N_4499,N_3128,N_3323);
and U4500 (N_4500,N_3790,N_3282);
or U4501 (N_4501,N_3118,N_3096);
nand U4502 (N_4502,N_3106,N_3808);
nand U4503 (N_4503,N_3358,N_3907);
nor U4504 (N_4504,N_3231,N_3510);
or U4505 (N_4505,N_3151,N_3314);
nor U4506 (N_4506,N_3861,N_3881);
or U4507 (N_4507,N_3717,N_3932);
nand U4508 (N_4508,N_3066,N_3747);
nand U4509 (N_4509,N_3529,N_3048);
and U4510 (N_4510,N_3676,N_3864);
nand U4511 (N_4511,N_3468,N_3578);
and U4512 (N_4512,N_3827,N_3944);
nand U4513 (N_4513,N_3003,N_3783);
nor U4514 (N_4514,N_3233,N_3331);
xor U4515 (N_4515,N_3782,N_3348);
or U4516 (N_4516,N_3134,N_3402);
or U4517 (N_4517,N_3671,N_3263);
nand U4518 (N_4518,N_3710,N_3856);
nand U4519 (N_4519,N_3997,N_3555);
and U4520 (N_4520,N_3027,N_3015);
nand U4521 (N_4521,N_3463,N_3294);
nand U4522 (N_4522,N_3039,N_3341);
nor U4523 (N_4523,N_3043,N_3212);
or U4524 (N_4524,N_3356,N_3672);
nand U4525 (N_4525,N_3154,N_3495);
and U4526 (N_4526,N_3510,N_3013);
nand U4527 (N_4527,N_3659,N_3602);
and U4528 (N_4528,N_3451,N_3580);
nor U4529 (N_4529,N_3598,N_3209);
nand U4530 (N_4530,N_3458,N_3404);
or U4531 (N_4531,N_3012,N_3852);
xor U4532 (N_4532,N_3308,N_3736);
or U4533 (N_4533,N_3719,N_3126);
nor U4534 (N_4534,N_3198,N_3113);
nand U4535 (N_4535,N_3466,N_3070);
and U4536 (N_4536,N_3302,N_3482);
nor U4537 (N_4537,N_3825,N_3627);
nand U4538 (N_4538,N_3757,N_3134);
or U4539 (N_4539,N_3271,N_3371);
nand U4540 (N_4540,N_3589,N_3172);
nand U4541 (N_4541,N_3834,N_3171);
and U4542 (N_4542,N_3406,N_3724);
nand U4543 (N_4543,N_3128,N_3852);
and U4544 (N_4544,N_3049,N_3234);
or U4545 (N_4545,N_3628,N_3382);
or U4546 (N_4546,N_3553,N_3110);
or U4547 (N_4547,N_3551,N_3604);
nand U4548 (N_4548,N_3663,N_3185);
or U4549 (N_4549,N_3525,N_3095);
nor U4550 (N_4550,N_3819,N_3001);
or U4551 (N_4551,N_3010,N_3898);
nand U4552 (N_4552,N_3056,N_3011);
xnor U4553 (N_4553,N_3188,N_3026);
and U4554 (N_4554,N_3883,N_3201);
or U4555 (N_4555,N_3057,N_3242);
nand U4556 (N_4556,N_3889,N_3751);
nor U4557 (N_4557,N_3025,N_3390);
nand U4558 (N_4558,N_3353,N_3202);
or U4559 (N_4559,N_3065,N_3739);
nand U4560 (N_4560,N_3953,N_3192);
and U4561 (N_4561,N_3286,N_3652);
or U4562 (N_4562,N_3002,N_3652);
nor U4563 (N_4563,N_3581,N_3389);
or U4564 (N_4564,N_3210,N_3516);
nand U4565 (N_4565,N_3146,N_3191);
nor U4566 (N_4566,N_3256,N_3843);
and U4567 (N_4567,N_3732,N_3457);
nor U4568 (N_4568,N_3330,N_3026);
or U4569 (N_4569,N_3038,N_3747);
or U4570 (N_4570,N_3759,N_3983);
nor U4571 (N_4571,N_3597,N_3556);
nand U4572 (N_4572,N_3303,N_3806);
nor U4573 (N_4573,N_3381,N_3377);
or U4574 (N_4574,N_3924,N_3201);
nor U4575 (N_4575,N_3341,N_3888);
nor U4576 (N_4576,N_3027,N_3682);
and U4577 (N_4577,N_3314,N_3441);
nand U4578 (N_4578,N_3949,N_3314);
nor U4579 (N_4579,N_3641,N_3551);
and U4580 (N_4580,N_3785,N_3351);
or U4581 (N_4581,N_3977,N_3461);
or U4582 (N_4582,N_3853,N_3740);
or U4583 (N_4583,N_3708,N_3180);
nor U4584 (N_4584,N_3058,N_3389);
nand U4585 (N_4585,N_3688,N_3411);
or U4586 (N_4586,N_3973,N_3318);
nand U4587 (N_4587,N_3347,N_3958);
or U4588 (N_4588,N_3759,N_3891);
or U4589 (N_4589,N_3359,N_3418);
and U4590 (N_4590,N_3660,N_3026);
nand U4591 (N_4591,N_3044,N_3414);
and U4592 (N_4592,N_3296,N_3323);
and U4593 (N_4593,N_3264,N_3450);
or U4594 (N_4594,N_3617,N_3865);
and U4595 (N_4595,N_3083,N_3240);
and U4596 (N_4596,N_3059,N_3680);
and U4597 (N_4597,N_3948,N_3822);
nor U4598 (N_4598,N_3910,N_3678);
nand U4599 (N_4599,N_3169,N_3145);
or U4600 (N_4600,N_3225,N_3197);
nor U4601 (N_4601,N_3081,N_3918);
and U4602 (N_4602,N_3082,N_3290);
or U4603 (N_4603,N_3589,N_3908);
nor U4604 (N_4604,N_3920,N_3406);
nor U4605 (N_4605,N_3184,N_3142);
and U4606 (N_4606,N_3880,N_3868);
or U4607 (N_4607,N_3439,N_3795);
nor U4608 (N_4608,N_3657,N_3044);
and U4609 (N_4609,N_3049,N_3184);
and U4610 (N_4610,N_3997,N_3556);
nand U4611 (N_4611,N_3189,N_3590);
or U4612 (N_4612,N_3693,N_3813);
and U4613 (N_4613,N_3049,N_3388);
or U4614 (N_4614,N_3228,N_3630);
or U4615 (N_4615,N_3419,N_3591);
and U4616 (N_4616,N_3009,N_3468);
or U4617 (N_4617,N_3261,N_3780);
xor U4618 (N_4618,N_3502,N_3272);
xnor U4619 (N_4619,N_3642,N_3102);
and U4620 (N_4620,N_3276,N_3038);
nand U4621 (N_4621,N_3504,N_3877);
or U4622 (N_4622,N_3508,N_3616);
or U4623 (N_4623,N_3063,N_3805);
or U4624 (N_4624,N_3450,N_3980);
and U4625 (N_4625,N_3421,N_3416);
nor U4626 (N_4626,N_3880,N_3122);
or U4627 (N_4627,N_3127,N_3819);
and U4628 (N_4628,N_3902,N_3101);
or U4629 (N_4629,N_3508,N_3163);
nor U4630 (N_4630,N_3975,N_3321);
and U4631 (N_4631,N_3129,N_3308);
xor U4632 (N_4632,N_3724,N_3717);
nor U4633 (N_4633,N_3076,N_3703);
and U4634 (N_4634,N_3683,N_3527);
nand U4635 (N_4635,N_3071,N_3744);
nand U4636 (N_4636,N_3523,N_3935);
nor U4637 (N_4637,N_3466,N_3290);
nand U4638 (N_4638,N_3363,N_3520);
or U4639 (N_4639,N_3925,N_3296);
nor U4640 (N_4640,N_3520,N_3591);
and U4641 (N_4641,N_3238,N_3671);
nand U4642 (N_4642,N_3699,N_3823);
nor U4643 (N_4643,N_3366,N_3674);
and U4644 (N_4644,N_3483,N_3845);
or U4645 (N_4645,N_3957,N_3438);
xor U4646 (N_4646,N_3531,N_3369);
and U4647 (N_4647,N_3895,N_3420);
nor U4648 (N_4648,N_3564,N_3169);
nand U4649 (N_4649,N_3239,N_3527);
nand U4650 (N_4650,N_3024,N_3774);
or U4651 (N_4651,N_3470,N_3583);
nand U4652 (N_4652,N_3506,N_3462);
or U4653 (N_4653,N_3176,N_3603);
xor U4654 (N_4654,N_3487,N_3675);
nor U4655 (N_4655,N_3487,N_3592);
nor U4656 (N_4656,N_3169,N_3245);
nand U4657 (N_4657,N_3704,N_3557);
nor U4658 (N_4658,N_3194,N_3484);
nor U4659 (N_4659,N_3645,N_3029);
and U4660 (N_4660,N_3636,N_3660);
and U4661 (N_4661,N_3743,N_3894);
nor U4662 (N_4662,N_3237,N_3000);
or U4663 (N_4663,N_3944,N_3035);
and U4664 (N_4664,N_3344,N_3407);
or U4665 (N_4665,N_3149,N_3353);
nand U4666 (N_4666,N_3821,N_3473);
nor U4667 (N_4667,N_3749,N_3048);
or U4668 (N_4668,N_3763,N_3916);
or U4669 (N_4669,N_3698,N_3144);
nor U4670 (N_4670,N_3077,N_3177);
nor U4671 (N_4671,N_3151,N_3719);
or U4672 (N_4672,N_3036,N_3536);
nor U4673 (N_4673,N_3550,N_3979);
nor U4674 (N_4674,N_3799,N_3253);
nor U4675 (N_4675,N_3653,N_3562);
or U4676 (N_4676,N_3601,N_3388);
or U4677 (N_4677,N_3300,N_3248);
and U4678 (N_4678,N_3679,N_3307);
nand U4679 (N_4679,N_3812,N_3185);
nor U4680 (N_4680,N_3013,N_3462);
nand U4681 (N_4681,N_3476,N_3906);
and U4682 (N_4682,N_3429,N_3833);
and U4683 (N_4683,N_3857,N_3674);
and U4684 (N_4684,N_3861,N_3718);
nand U4685 (N_4685,N_3408,N_3748);
and U4686 (N_4686,N_3974,N_3016);
nor U4687 (N_4687,N_3515,N_3606);
or U4688 (N_4688,N_3807,N_3254);
nor U4689 (N_4689,N_3262,N_3787);
or U4690 (N_4690,N_3072,N_3866);
or U4691 (N_4691,N_3197,N_3718);
nand U4692 (N_4692,N_3503,N_3596);
nor U4693 (N_4693,N_3210,N_3267);
or U4694 (N_4694,N_3289,N_3863);
and U4695 (N_4695,N_3807,N_3582);
or U4696 (N_4696,N_3601,N_3245);
or U4697 (N_4697,N_3055,N_3426);
or U4698 (N_4698,N_3410,N_3559);
or U4699 (N_4699,N_3536,N_3902);
or U4700 (N_4700,N_3106,N_3533);
and U4701 (N_4701,N_3861,N_3838);
nand U4702 (N_4702,N_3214,N_3476);
and U4703 (N_4703,N_3940,N_3989);
nor U4704 (N_4704,N_3567,N_3523);
and U4705 (N_4705,N_3297,N_3783);
nor U4706 (N_4706,N_3252,N_3962);
and U4707 (N_4707,N_3048,N_3748);
nand U4708 (N_4708,N_3771,N_3117);
nand U4709 (N_4709,N_3692,N_3784);
nor U4710 (N_4710,N_3082,N_3788);
or U4711 (N_4711,N_3990,N_3440);
or U4712 (N_4712,N_3179,N_3623);
nand U4713 (N_4713,N_3571,N_3367);
or U4714 (N_4714,N_3066,N_3262);
nor U4715 (N_4715,N_3407,N_3443);
nand U4716 (N_4716,N_3468,N_3652);
and U4717 (N_4717,N_3323,N_3848);
nor U4718 (N_4718,N_3793,N_3576);
and U4719 (N_4719,N_3475,N_3311);
or U4720 (N_4720,N_3287,N_3139);
or U4721 (N_4721,N_3353,N_3597);
nand U4722 (N_4722,N_3202,N_3080);
and U4723 (N_4723,N_3457,N_3112);
nor U4724 (N_4724,N_3686,N_3549);
nand U4725 (N_4725,N_3914,N_3300);
nand U4726 (N_4726,N_3240,N_3625);
and U4727 (N_4727,N_3186,N_3804);
xnor U4728 (N_4728,N_3556,N_3479);
nand U4729 (N_4729,N_3261,N_3652);
or U4730 (N_4730,N_3926,N_3121);
or U4731 (N_4731,N_3004,N_3499);
nand U4732 (N_4732,N_3354,N_3098);
xor U4733 (N_4733,N_3032,N_3824);
or U4734 (N_4734,N_3727,N_3849);
or U4735 (N_4735,N_3558,N_3936);
nand U4736 (N_4736,N_3934,N_3101);
nand U4737 (N_4737,N_3684,N_3045);
or U4738 (N_4738,N_3154,N_3815);
xor U4739 (N_4739,N_3558,N_3577);
nand U4740 (N_4740,N_3989,N_3024);
nor U4741 (N_4741,N_3561,N_3666);
xor U4742 (N_4742,N_3815,N_3587);
or U4743 (N_4743,N_3236,N_3790);
nand U4744 (N_4744,N_3534,N_3199);
or U4745 (N_4745,N_3055,N_3634);
or U4746 (N_4746,N_3027,N_3065);
or U4747 (N_4747,N_3303,N_3691);
or U4748 (N_4748,N_3722,N_3138);
nor U4749 (N_4749,N_3290,N_3213);
and U4750 (N_4750,N_3623,N_3868);
or U4751 (N_4751,N_3160,N_3542);
or U4752 (N_4752,N_3001,N_3969);
and U4753 (N_4753,N_3636,N_3142);
and U4754 (N_4754,N_3528,N_3590);
or U4755 (N_4755,N_3387,N_3441);
or U4756 (N_4756,N_3373,N_3629);
or U4757 (N_4757,N_3779,N_3705);
nand U4758 (N_4758,N_3940,N_3786);
and U4759 (N_4759,N_3945,N_3252);
nor U4760 (N_4760,N_3624,N_3473);
or U4761 (N_4761,N_3734,N_3111);
and U4762 (N_4762,N_3064,N_3667);
and U4763 (N_4763,N_3696,N_3425);
nand U4764 (N_4764,N_3869,N_3828);
and U4765 (N_4765,N_3809,N_3931);
nand U4766 (N_4766,N_3029,N_3373);
and U4767 (N_4767,N_3739,N_3859);
or U4768 (N_4768,N_3303,N_3416);
nor U4769 (N_4769,N_3441,N_3000);
or U4770 (N_4770,N_3611,N_3468);
or U4771 (N_4771,N_3318,N_3102);
or U4772 (N_4772,N_3814,N_3359);
nor U4773 (N_4773,N_3754,N_3860);
nand U4774 (N_4774,N_3811,N_3703);
nor U4775 (N_4775,N_3642,N_3549);
and U4776 (N_4776,N_3722,N_3483);
nand U4777 (N_4777,N_3016,N_3416);
or U4778 (N_4778,N_3468,N_3308);
nor U4779 (N_4779,N_3101,N_3653);
and U4780 (N_4780,N_3003,N_3736);
nor U4781 (N_4781,N_3968,N_3207);
and U4782 (N_4782,N_3860,N_3034);
nor U4783 (N_4783,N_3686,N_3695);
or U4784 (N_4784,N_3674,N_3689);
nor U4785 (N_4785,N_3340,N_3983);
or U4786 (N_4786,N_3231,N_3475);
or U4787 (N_4787,N_3853,N_3084);
nand U4788 (N_4788,N_3930,N_3937);
and U4789 (N_4789,N_3148,N_3746);
nand U4790 (N_4790,N_3760,N_3650);
or U4791 (N_4791,N_3816,N_3723);
and U4792 (N_4792,N_3926,N_3125);
or U4793 (N_4793,N_3170,N_3556);
nand U4794 (N_4794,N_3946,N_3988);
nand U4795 (N_4795,N_3280,N_3253);
and U4796 (N_4796,N_3450,N_3034);
nor U4797 (N_4797,N_3873,N_3097);
and U4798 (N_4798,N_3968,N_3246);
nor U4799 (N_4799,N_3988,N_3357);
nand U4800 (N_4800,N_3449,N_3394);
nor U4801 (N_4801,N_3254,N_3913);
or U4802 (N_4802,N_3511,N_3198);
or U4803 (N_4803,N_3692,N_3979);
nand U4804 (N_4804,N_3862,N_3965);
nand U4805 (N_4805,N_3009,N_3197);
and U4806 (N_4806,N_3159,N_3968);
or U4807 (N_4807,N_3308,N_3431);
nand U4808 (N_4808,N_3049,N_3753);
nor U4809 (N_4809,N_3507,N_3410);
xor U4810 (N_4810,N_3045,N_3018);
or U4811 (N_4811,N_3581,N_3366);
nand U4812 (N_4812,N_3793,N_3162);
and U4813 (N_4813,N_3481,N_3611);
or U4814 (N_4814,N_3013,N_3220);
or U4815 (N_4815,N_3497,N_3479);
nor U4816 (N_4816,N_3842,N_3163);
and U4817 (N_4817,N_3249,N_3506);
nor U4818 (N_4818,N_3203,N_3957);
and U4819 (N_4819,N_3038,N_3158);
or U4820 (N_4820,N_3140,N_3520);
or U4821 (N_4821,N_3709,N_3415);
nand U4822 (N_4822,N_3561,N_3825);
nand U4823 (N_4823,N_3167,N_3347);
or U4824 (N_4824,N_3197,N_3443);
nand U4825 (N_4825,N_3736,N_3486);
nor U4826 (N_4826,N_3955,N_3055);
nor U4827 (N_4827,N_3567,N_3240);
nor U4828 (N_4828,N_3823,N_3483);
and U4829 (N_4829,N_3173,N_3900);
and U4830 (N_4830,N_3472,N_3007);
or U4831 (N_4831,N_3852,N_3190);
or U4832 (N_4832,N_3683,N_3250);
nor U4833 (N_4833,N_3101,N_3077);
and U4834 (N_4834,N_3178,N_3904);
nand U4835 (N_4835,N_3302,N_3467);
and U4836 (N_4836,N_3844,N_3611);
or U4837 (N_4837,N_3381,N_3342);
nand U4838 (N_4838,N_3036,N_3935);
or U4839 (N_4839,N_3296,N_3743);
or U4840 (N_4840,N_3237,N_3534);
or U4841 (N_4841,N_3510,N_3366);
nor U4842 (N_4842,N_3816,N_3283);
nor U4843 (N_4843,N_3480,N_3516);
nor U4844 (N_4844,N_3354,N_3341);
nor U4845 (N_4845,N_3446,N_3395);
and U4846 (N_4846,N_3272,N_3804);
nand U4847 (N_4847,N_3731,N_3664);
nand U4848 (N_4848,N_3829,N_3206);
and U4849 (N_4849,N_3444,N_3784);
or U4850 (N_4850,N_3625,N_3130);
and U4851 (N_4851,N_3221,N_3795);
nand U4852 (N_4852,N_3219,N_3474);
nand U4853 (N_4853,N_3811,N_3637);
nand U4854 (N_4854,N_3836,N_3815);
nand U4855 (N_4855,N_3989,N_3529);
and U4856 (N_4856,N_3881,N_3214);
nor U4857 (N_4857,N_3471,N_3624);
and U4858 (N_4858,N_3820,N_3371);
nand U4859 (N_4859,N_3606,N_3939);
and U4860 (N_4860,N_3001,N_3772);
and U4861 (N_4861,N_3462,N_3467);
nor U4862 (N_4862,N_3628,N_3527);
nor U4863 (N_4863,N_3246,N_3392);
nor U4864 (N_4864,N_3464,N_3253);
nor U4865 (N_4865,N_3607,N_3307);
nor U4866 (N_4866,N_3705,N_3952);
or U4867 (N_4867,N_3306,N_3039);
and U4868 (N_4868,N_3730,N_3704);
nor U4869 (N_4869,N_3657,N_3411);
nor U4870 (N_4870,N_3957,N_3982);
nor U4871 (N_4871,N_3906,N_3931);
nor U4872 (N_4872,N_3158,N_3401);
nand U4873 (N_4873,N_3713,N_3944);
and U4874 (N_4874,N_3958,N_3224);
nor U4875 (N_4875,N_3109,N_3608);
nand U4876 (N_4876,N_3557,N_3707);
nor U4877 (N_4877,N_3853,N_3662);
or U4878 (N_4878,N_3010,N_3401);
nor U4879 (N_4879,N_3091,N_3680);
and U4880 (N_4880,N_3005,N_3531);
or U4881 (N_4881,N_3596,N_3809);
or U4882 (N_4882,N_3815,N_3118);
and U4883 (N_4883,N_3206,N_3543);
nor U4884 (N_4884,N_3049,N_3132);
nor U4885 (N_4885,N_3951,N_3881);
nor U4886 (N_4886,N_3921,N_3338);
nand U4887 (N_4887,N_3595,N_3166);
nand U4888 (N_4888,N_3218,N_3447);
and U4889 (N_4889,N_3042,N_3961);
and U4890 (N_4890,N_3182,N_3020);
and U4891 (N_4891,N_3747,N_3478);
nand U4892 (N_4892,N_3220,N_3555);
and U4893 (N_4893,N_3868,N_3704);
and U4894 (N_4894,N_3716,N_3833);
or U4895 (N_4895,N_3718,N_3329);
xnor U4896 (N_4896,N_3251,N_3637);
nor U4897 (N_4897,N_3295,N_3267);
nor U4898 (N_4898,N_3096,N_3002);
nor U4899 (N_4899,N_3862,N_3052);
or U4900 (N_4900,N_3576,N_3688);
and U4901 (N_4901,N_3490,N_3065);
or U4902 (N_4902,N_3801,N_3469);
nor U4903 (N_4903,N_3930,N_3470);
and U4904 (N_4904,N_3736,N_3176);
and U4905 (N_4905,N_3766,N_3213);
nand U4906 (N_4906,N_3218,N_3144);
nor U4907 (N_4907,N_3544,N_3431);
nor U4908 (N_4908,N_3890,N_3025);
nand U4909 (N_4909,N_3505,N_3352);
nand U4910 (N_4910,N_3438,N_3206);
or U4911 (N_4911,N_3088,N_3441);
nor U4912 (N_4912,N_3792,N_3091);
nor U4913 (N_4913,N_3648,N_3252);
and U4914 (N_4914,N_3366,N_3814);
nor U4915 (N_4915,N_3204,N_3928);
and U4916 (N_4916,N_3053,N_3601);
nor U4917 (N_4917,N_3509,N_3188);
and U4918 (N_4918,N_3980,N_3711);
and U4919 (N_4919,N_3297,N_3972);
nor U4920 (N_4920,N_3844,N_3636);
and U4921 (N_4921,N_3322,N_3821);
xor U4922 (N_4922,N_3675,N_3188);
and U4923 (N_4923,N_3526,N_3252);
nand U4924 (N_4924,N_3253,N_3756);
nand U4925 (N_4925,N_3596,N_3923);
nor U4926 (N_4926,N_3220,N_3577);
or U4927 (N_4927,N_3257,N_3237);
or U4928 (N_4928,N_3583,N_3486);
nor U4929 (N_4929,N_3080,N_3411);
nand U4930 (N_4930,N_3148,N_3603);
xor U4931 (N_4931,N_3362,N_3203);
xor U4932 (N_4932,N_3072,N_3863);
nor U4933 (N_4933,N_3032,N_3911);
nor U4934 (N_4934,N_3292,N_3060);
and U4935 (N_4935,N_3983,N_3317);
or U4936 (N_4936,N_3485,N_3951);
or U4937 (N_4937,N_3599,N_3806);
nor U4938 (N_4938,N_3574,N_3311);
or U4939 (N_4939,N_3882,N_3200);
and U4940 (N_4940,N_3557,N_3661);
or U4941 (N_4941,N_3439,N_3203);
nor U4942 (N_4942,N_3002,N_3014);
nor U4943 (N_4943,N_3619,N_3001);
and U4944 (N_4944,N_3704,N_3498);
nor U4945 (N_4945,N_3630,N_3303);
nand U4946 (N_4946,N_3196,N_3150);
and U4947 (N_4947,N_3967,N_3508);
or U4948 (N_4948,N_3645,N_3782);
or U4949 (N_4949,N_3353,N_3853);
or U4950 (N_4950,N_3095,N_3539);
nor U4951 (N_4951,N_3226,N_3784);
and U4952 (N_4952,N_3635,N_3645);
nand U4953 (N_4953,N_3661,N_3524);
or U4954 (N_4954,N_3099,N_3307);
nor U4955 (N_4955,N_3594,N_3997);
nand U4956 (N_4956,N_3129,N_3344);
nor U4957 (N_4957,N_3488,N_3959);
nand U4958 (N_4958,N_3724,N_3488);
and U4959 (N_4959,N_3802,N_3216);
or U4960 (N_4960,N_3098,N_3805);
or U4961 (N_4961,N_3899,N_3909);
nand U4962 (N_4962,N_3951,N_3283);
and U4963 (N_4963,N_3903,N_3298);
and U4964 (N_4964,N_3472,N_3217);
xor U4965 (N_4965,N_3543,N_3892);
nand U4966 (N_4966,N_3382,N_3372);
nand U4967 (N_4967,N_3143,N_3873);
nand U4968 (N_4968,N_3766,N_3715);
or U4969 (N_4969,N_3674,N_3826);
and U4970 (N_4970,N_3709,N_3956);
nand U4971 (N_4971,N_3168,N_3622);
nand U4972 (N_4972,N_3982,N_3215);
nor U4973 (N_4973,N_3949,N_3368);
nor U4974 (N_4974,N_3694,N_3942);
nor U4975 (N_4975,N_3153,N_3781);
or U4976 (N_4976,N_3086,N_3644);
nor U4977 (N_4977,N_3460,N_3974);
and U4978 (N_4978,N_3661,N_3871);
and U4979 (N_4979,N_3301,N_3017);
nand U4980 (N_4980,N_3725,N_3669);
or U4981 (N_4981,N_3819,N_3008);
nor U4982 (N_4982,N_3312,N_3013);
nor U4983 (N_4983,N_3057,N_3100);
nor U4984 (N_4984,N_3082,N_3038);
nor U4985 (N_4985,N_3078,N_3580);
nand U4986 (N_4986,N_3436,N_3559);
nor U4987 (N_4987,N_3054,N_3102);
nand U4988 (N_4988,N_3518,N_3484);
nor U4989 (N_4989,N_3160,N_3189);
nand U4990 (N_4990,N_3635,N_3312);
nor U4991 (N_4991,N_3069,N_3070);
and U4992 (N_4992,N_3379,N_3778);
or U4993 (N_4993,N_3293,N_3869);
or U4994 (N_4994,N_3424,N_3196);
nand U4995 (N_4995,N_3252,N_3927);
or U4996 (N_4996,N_3356,N_3230);
nor U4997 (N_4997,N_3759,N_3778);
or U4998 (N_4998,N_3110,N_3276);
and U4999 (N_4999,N_3575,N_3083);
nand U5000 (N_5000,N_4431,N_4030);
nand U5001 (N_5001,N_4757,N_4455);
nor U5002 (N_5002,N_4732,N_4653);
nor U5003 (N_5003,N_4530,N_4673);
nand U5004 (N_5004,N_4614,N_4780);
and U5005 (N_5005,N_4647,N_4630);
or U5006 (N_5006,N_4882,N_4237);
nand U5007 (N_5007,N_4177,N_4608);
and U5008 (N_5008,N_4395,N_4662);
xnor U5009 (N_5009,N_4928,N_4364);
nand U5010 (N_5010,N_4875,N_4546);
nor U5011 (N_5011,N_4547,N_4168);
nand U5012 (N_5012,N_4899,N_4008);
xor U5013 (N_5013,N_4373,N_4461);
nor U5014 (N_5014,N_4013,N_4678);
nor U5015 (N_5015,N_4725,N_4394);
or U5016 (N_5016,N_4404,N_4854);
and U5017 (N_5017,N_4606,N_4306);
nand U5018 (N_5018,N_4345,N_4528);
nand U5019 (N_5019,N_4629,N_4110);
nand U5020 (N_5020,N_4090,N_4343);
nor U5021 (N_5021,N_4269,N_4485);
and U5022 (N_5022,N_4275,N_4317);
and U5023 (N_5023,N_4487,N_4517);
and U5024 (N_5024,N_4223,N_4851);
nor U5025 (N_5025,N_4721,N_4765);
or U5026 (N_5026,N_4934,N_4557);
or U5027 (N_5027,N_4065,N_4739);
nor U5028 (N_5028,N_4255,N_4468);
nand U5029 (N_5029,N_4612,N_4883);
and U5030 (N_5030,N_4108,N_4143);
or U5031 (N_5031,N_4621,N_4607);
nor U5032 (N_5032,N_4704,N_4002);
nor U5033 (N_5033,N_4555,N_4178);
or U5034 (N_5034,N_4565,N_4610);
and U5035 (N_5035,N_4985,N_4412);
and U5036 (N_5036,N_4651,N_4241);
or U5037 (N_5037,N_4171,N_4714);
or U5038 (N_5038,N_4135,N_4533);
nand U5039 (N_5039,N_4675,N_4181);
or U5040 (N_5040,N_4832,N_4426);
xnor U5041 (N_5041,N_4545,N_4801);
and U5042 (N_5042,N_4045,N_4901);
nand U5043 (N_5043,N_4907,N_4756);
nor U5044 (N_5044,N_4666,N_4250);
and U5045 (N_5045,N_4462,N_4881);
or U5046 (N_5046,N_4146,N_4294);
and U5047 (N_5047,N_4843,N_4860);
nand U5048 (N_5048,N_4151,N_4897);
nor U5049 (N_5049,N_4198,N_4200);
and U5050 (N_5050,N_4482,N_4128);
nand U5051 (N_5051,N_4686,N_4878);
and U5052 (N_5052,N_4753,N_4945);
or U5053 (N_5053,N_4480,N_4025);
or U5054 (N_5054,N_4094,N_4968);
or U5055 (N_5055,N_4710,N_4292);
nand U5056 (N_5056,N_4604,N_4184);
nand U5057 (N_5057,N_4259,N_4773);
or U5058 (N_5058,N_4498,N_4060);
nor U5059 (N_5059,N_4116,N_4609);
and U5060 (N_5060,N_4516,N_4646);
and U5061 (N_5061,N_4434,N_4764);
nand U5062 (N_5062,N_4706,N_4232);
and U5063 (N_5063,N_4965,N_4526);
nand U5064 (N_5064,N_4082,N_4733);
and U5065 (N_5065,N_4271,N_4386);
nand U5066 (N_5066,N_4549,N_4332);
or U5067 (N_5067,N_4109,N_4367);
nor U5068 (N_5068,N_4137,N_4817);
nor U5069 (N_5069,N_4311,N_4974);
nand U5070 (N_5070,N_4486,N_4695);
nor U5071 (N_5071,N_4173,N_4515);
or U5072 (N_5072,N_4510,N_4284);
and U5073 (N_5073,N_4446,N_4833);
xnor U5074 (N_5074,N_4677,N_4210);
nand U5075 (N_5075,N_4585,N_4684);
or U5076 (N_5076,N_4236,N_4124);
nand U5077 (N_5077,N_4266,N_4014);
or U5078 (N_5078,N_4153,N_4514);
nor U5079 (N_5079,N_4349,N_4903);
and U5080 (N_5080,N_4382,N_4463);
nor U5081 (N_5081,N_4212,N_4297);
nor U5082 (N_5082,N_4844,N_4144);
nor U5083 (N_5083,N_4596,N_4460);
nand U5084 (N_5084,N_4478,N_4865);
nor U5085 (N_5085,N_4339,N_4942);
or U5086 (N_5086,N_4273,N_4385);
nand U5087 (N_5087,N_4272,N_4905);
or U5088 (N_5088,N_4326,N_4933);
or U5089 (N_5089,N_4348,N_4454);
or U5090 (N_5090,N_4493,N_4683);
xor U5091 (N_5091,N_4741,N_4053);
or U5092 (N_5092,N_4472,N_4372);
and U5093 (N_5093,N_4464,N_4083);
and U5094 (N_5094,N_4518,N_4619);
and U5095 (N_5095,N_4685,N_4257);
and U5096 (N_5096,N_4499,N_4477);
nand U5097 (N_5097,N_4894,N_4960);
or U5098 (N_5098,N_4481,N_4603);
nand U5099 (N_5099,N_4620,N_4365);
or U5100 (N_5100,N_4233,N_4270);
nand U5101 (N_5101,N_4010,N_4113);
or U5102 (N_5102,N_4605,N_4694);
and U5103 (N_5103,N_4229,N_4329);
nand U5104 (N_5104,N_4381,N_4017);
nand U5105 (N_5105,N_4952,N_4401);
nor U5106 (N_5106,N_4709,N_4738);
nor U5107 (N_5107,N_4003,N_4202);
or U5108 (N_5108,N_4012,N_4786);
or U5109 (N_5109,N_4838,N_4656);
nor U5110 (N_5110,N_4587,N_4736);
and U5111 (N_5111,N_4087,N_4595);
and U5112 (N_5112,N_4230,N_4433);
nand U5113 (N_5113,N_4783,N_4321);
and U5114 (N_5114,N_4577,N_4015);
nor U5115 (N_5115,N_4772,N_4203);
nand U5116 (N_5116,N_4961,N_4523);
and U5117 (N_5117,N_4479,N_4268);
and U5118 (N_5118,N_4635,N_4357);
nor U5119 (N_5119,N_4570,N_4866);
or U5120 (N_5120,N_4802,N_4323);
and U5121 (N_5121,N_4745,N_4403);
or U5122 (N_5122,N_4936,N_4906);
and U5123 (N_5123,N_4874,N_4123);
and U5124 (N_5124,N_4645,N_4283);
or U5125 (N_5125,N_4593,N_4615);
or U5126 (N_5126,N_4640,N_4876);
nand U5127 (N_5127,N_4328,N_4501);
and U5128 (N_5128,N_4421,N_4525);
xnor U5129 (N_5129,N_4409,N_4084);
nand U5130 (N_5130,N_4537,N_4247);
and U5131 (N_5131,N_4397,N_4959);
nor U5132 (N_5132,N_4892,N_4042);
xnor U5133 (N_5133,N_4160,N_4072);
or U5134 (N_5134,N_4338,N_4139);
or U5135 (N_5135,N_4320,N_4650);
nor U5136 (N_5136,N_4682,N_4588);
nor U5137 (N_5137,N_4127,N_4639);
and U5138 (N_5138,N_4162,N_4425);
or U5139 (N_5139,N_4375,N_4575);
nor U5140 (N_5140,N_4719,N_4943);
nand U5141 (N_5141,N_4506,N_4224);
nand U5142 (N_5142,N_4914,N_4490);
nor U5143 (N_5143,N_4318,N_4567);
or U5144 (N_5144,N_4359,N_4192);
nor U5145 (N_5145,N_4550,N_4638);
nand U5146 (N_5146,N_4862,N_4841);
xor U5147 (N_5147,N_4969,N_4778);
or U5148 (N_5148,N_4211,N_4950);
and U5149 (N_5149,N_4183,N_4659);
nand U5150 (N_5150,N_4774,N_4669);
nand U5151 (N_5151,N_4599,N_4561);
or U5152 (N_5152,N_4344,N_4652);
or U5153 (N_5153,N_4879,N_4019);
nor U5154 (N_5154,N_4024,N_4873);
nor U5155 (N_5155,N_4554,N_4055);
nand U5156 (N_5156,N_4234,N_4855);
and U5157 (N_5157,N_4798,N_4193);
or U5158 (N_5158,N_4444,N_4658);
nand U5159 (N_5159,N_4849,N_4459);
nor U5160 (N_5160,N_4448,N_4702);
nand U5161 (N_5161,N_4484,N_4697);
or U5162 (N_5162,N_4190,N_4799);
nor U5163 (N_5163,N_4712,N_4327);
nand U5164 (N_5164,N_4935,N_4842);
and U5165 (N_5165,N_4069,N_4107);
or U5166 (N_5166,N_4360,N_4004);
and U5167 (N_5167,N_4782,N_4520);
and U5168 (N_5168,N_4809,N_4141);
nand U5169 (N_5169,N_4443,N_4219);
and U5170 (N_5170,N_4885,N_4668);
nand U5171 (N_5171,N_4287,N_4663);
nand U5172 (N_5172,N_4281,N_4611);
nand U5173 (N_5173,N_4976,N_4680);
nand U5174 (N_5174,N_4857,N_4041);
or U5175 (N_5175,N_4191,N_4558);
and U5176 (N_5176,N_4660,N_4301);
nor U5177 (N_5177,N_4351,N_4752);
and U5178 (N_5178,N_4172,N_4073);
nor U5179 (N_5179,N_4166,N_4341);
nand U5180 (N_5180,N_4251,N_4924);
nand U5181 (N_5181,N_4589,N_4355);
and U5182 (N_5182,N_4507,N_4147);
nand U5183 (N_5183,N_4369,N_4331);
or U5184 (N_5184,N_4616,N_4504);
nor U5185 (N_5185,N_4717,N_4118);
nor U5186 (N_5186,N_4429,N_4185);
nor U5187 (N_5187,N_4804,N_4826);
nor U5188 (N_5188,N_4910,N_4541);
and U5189 (N_5189,N_4734,N_4204);
nand U5190 (N_5190,N_4856,N_4416);
and U5191 (N_5191,N_4913,N_4001);
xnor U5192 (N_5192,N_4845,N_4743);
nand U5193 (N_5193,N_4784,N_4793);
xor U5194 (N_5194,N_4674,N_4823);
or U5195 (N_5195,N_4532,N_4641);
nand U5196 (N_5196,N_4740,N_4762);
nor U5197 (N_5197,N_4228,N_4643);
or U5198 (N_5198,N_4114,N_4260);
and U5199 (N_5199,N_4637,N_4703);
xnor U5200 (N_5200,N_4342,N_4475);
or U5201 (N_5201,N_4417,N_4347);
nand U5202 (N_5202,N_4097,N_4303);
nand U5203 (N_5203,N_4729,N_4491);
nand U5204 (N_5204,N_4337,N_4869);
nand U5205 (N_5205,N_4904,N_4106);
and U5206 (N_5206,N_4028,N_4440);
nor U5207 (N_5207,N_4718,N_4676);
nand U5208 (N_5208,N_4927,N_4921);
or U5209 (N_5209,N_4699,N_4981);
and U5210 (N_5210,N_4781,N_4432);
nor U5211 (N_5211,N_4285,N_4340);
nand U5212 (N_5212,N_4992,N_4815);
nand U5213 (N_5213,N_4835,N_4973);
or U5214 (N_5214,N_4150,N_4154);
nor U5215 (N_5215,N_4189,N_4134);
nand U5216 (N_5216,N_4098,N_4451);
or U5217 (N_5217,N_4747,N_4280);
nor U5218 (N_5218,N_4672,N_4582);
and U5219 (N_5219,N_4552,N_4789);
nand U5220 (N_5220,N_4648,N_4966);
and U5221 (N_5221,N_4111,N_4947);
nor U5222 (N_5222,N_4671,N_4562);
and U5223 (N_5223,N_4982,N_4583);
or U5224 (N_5224,N_4182,N_4993);
or U5225 (N_5225,N_4670,N_4092);
xor U5226 (N_5226,N_4768,N_4626);
or U5227 (N_5227,N_4384,N_4129);
nand U5228 (N_5228,N_4602,N_4170);
nand U5229 (N_5229,N_4958,N_4744);
or U5230 (N_5230,N_4075,N_4578);
or U5231 (N_5231,N_4009,N_4370);
and U5232 (N_5232,N_4047,N_4792);
nand U5233 (N_5233,N_4022,N_4214);
nand U5234 (N_5234,N_4911,N_4220);
or U5235 (N_5235,N_4324,N_4388);
nand U5236 (N_5236,N_4046,N_4057);
and U5237 (N_5237,N_4536,N_4690);
nand U5238 (N_5238,N_4086,N_4419);
xnor U5239 (N_5239,N_4374,N_4556);
or U5240 (N_5240,N_4963,N_4180);
xor U5241 (N_5241,N_4186,N_4390);
or U5242 (N_5242,N_4877,N_4754);
and U5243 (N_5243,N_4760,N_4748);
nand U5244 (N_5244,N_4531,N_4298);
or U5245 (N_5245,N_4038,N_4422);
or U5246 (N_5246,N_4112,N_4824);
or U5247 (N_5247,N_4511,N_4896);
and U5248 (N_5248,N_4165,N_4867);
nand U5249 (N_5249,N_4465,N_4244);
xor U5250 (N_5250,N_4957,N_4050);
and U5251 (N_5251,N_4070,N_4566);
or U5252 (N_5252,N_4688,N_4474);
and U5253 (N_5253,N_4521,N_4415);
and U5254 (N_5254,N_4119,N_4850);
or U5255 (N_5255,N_4277,N_4316);
nand U5256 (N_5256,N_4095,N_4405);
nand U5257 (N_5257,N_4054,N_4380);
or U5258 (N_5258,N_4926,N_4972);
or U5259 (N_5259,N_4353,N_4218);
and U5260 (N_5260,N_4121,N_4722);
nand U5261 (N_5261,N_4217,N_4435);
or U5262 (N_5262,N_4356,N_4076);
nor U5263 (N_5263,N_4655,N_4563);
nand U5264 (N_5264,N_4148,N_4746);
nor U5265 (N_5265,N_4573,N_4564);
and U5266 (N_5266,N_4949,N_4667);
xor U5267 (N_5267,N_4392,N_4158);
or U5268 (N_5268,N_4983,N_4505);
nand U5269 (N_5269,N_4978,N_4399);
and U5270 (N_5270,N_4133,N_4400);
nor U5271 (N_5271,N_4037,N_4430);
nand U5272 (N_5272,N_4975,N_4693);
nand U5273 (N_5273,N_4551,N_4163);
or U5274 (N_5274,N_4758,N_4115);
nor U5275 (N_5275,N_4543,N_4997);
nor U5276 (N_5276,N_4040,N_4713);
or U5277 (N_5277,N_4995,N_4542);
nand U5278 (N_5278,N_4209,N_4253);
nor U5279 (N_5279,N_4059,N_4264);
nor U5280 (N_5280,N_4948,N_4836);
nand U5281 (N_5281,N_4293,N_4822);
or U5282 (N_5282,N_4377,N_4290);
nand U5283 (N_5283,N_4735,N_4770);
nand U5284 (N_5284,N_4502,N_4918);
nand U5285 (N_5285,N_4174,N_4007);
or U5286 (N_5286,N_4512,N_4777);
nand U5287 (N_5287,N_4081,N_4061);
or U5288 (N_5288,N_4807,N_4383);
and U5289 (N_5289,N_4813,N_4938);
nand U5290 (N_5290,N_4393,N_4408);
nand U5291 (N_5291,N_4503,N_4276);
nand U5292 (N_5292,N_4424,N_4391);
nor U5293 (N_5293,N_4571,N_4586);
nor U5294 (N_5294,N_4201,N_4681);
nand U5295 (N_5295,N_4977,N_4362);
nand U5296 (N_5296,N_4452,N_4853);
or U5297 (N_5297,N_4954,N_4445);
nand U5298 (N_5298,N_4785,N_4755);
or U5299 (N_5299,N_4221,N_4691);
or U5300 (N_5300,N_4021,N_4314);
or U5301 (N_5301,N_4767,N_4175);
or U5302 (N_5302,N_4908,N_4791);
nor U5303 (N_5303,N_4363,N_4979);
and U5304 (N_5304,N_4058,N_4909);
nor U5305 (N_5305,N_4636,N_4023);
nor U5306 (N_5306,N_4299,N_4569);
nand U5307 (N_5307,N_4529,N_4991);
nand U5308 (N_5308,N_4946,N_4354);
or U5309 (N_5309,N_4900,N_4750);
nand U5310 (N_5310,N_4806,N_4295);
nor U5311 (N_5311,N_4000,N_4967);
or U5312 (N_5312,N_4937,N_4225);
nor U5313 (N_5313,N_4999,N_4387);
or U5314 (N_5314,N_4705,N_4846);
nor U5315 (N_5315,N_4581,N_4282);
and U5316 (N_5316,N_4970,N_4818);
nor U5317 (N_5317,N_4368,N_4441);
and U5318 (N_5318,N_4248,N_4628);
or U5319 (N_5319,N_4613,N_4700);
nand U5320 (N_5320,N_4207,N_4898);
nand U5321 (N_5321,N_4893,N_4044);
nor U5322 (N_5322,N_4313,N_4427);
nor U5323 (N_5323,N_4821,N_4043);
nor U5324 (N_5324,N_4438,N_4941);
and U5325 (N_5325,N_4779,N_4559);
nor U5326 (N_5326,N_4026,N_4687);
and U5327 (N_5327,N_4984,N_4771);
nor U5328 (N_5328,N_4590,N_4895);
and U5329 (N_5329,N_4707,N_4737);
and U5330 (N_5330,N_4447,N_4986);
nor U5331 (N_5331,N_4795,N_4820);
or U5332 (N_5332,N_4888,N_4912);
and U5333 (N_5333,N_4955,N_4265);
nand U5334 (N_5334,N_4291,N_4534);
nor U5335 (N_5335,N_4953,N_4125);
or U5336 (N_5336,N_4246,N_4398);
nor U5337 (N_5337,N_4592,N_4489);
or U5338 (N_5338,N_4018,N_4483);
and U5339 (N_5339,N_4199,N_4539);
or U5340 (N_5340,N_4964,N_4187);
or U5341 (N_5341,N_4256,N_4796);
or U5342 (N_5342,N_4711,N_4940);
or U5343 (N_5343,N_4423,N_4215);
nor U5344 (N_5344,N_4810,N_4205);
or U5345 (N_5345,N_4708,N_4074);
or U5346 (N_5346,N_4932,N_4724);
and U5347 (N_5347,N_4916,N_4197);
nor U5348 (N_5348,N_4889,N_4548);
nand U5349 (N_5349,N_4829,N_4469);
or U5350 (N_5350,N_4723,N_4300);
nand U5351 (N_5351,N_4195,N_4439);
and U5352 (N_5352,N_4890,N_4880);
and U5353 (N_5353,N_4105,N_4120);
or U5354 (N_5354,N_4597,N_4864);
nand U5355 (N_5355,N_4138,N_4998);
and U5356 (N_5356,N_4376,N_4450);
nand U5357 (N_5357,N_4830,N_4305);
and U5358 (N_5358,N_4034,N_4692);
and U5359 (N_5359,N_4406,N_4176);
and U5360 (N_5360,N_4508,N_4990);
nor U5361 (N_5361,N_4267,N_4679);
nand U5362 (N_5362,N_4980,N_4863);
and U5363 (N_5363,N_4242,N_4726);
nor U5364 (N_5364,N_4302,N_4576);
or U5365 (N_5365,N_4100,N_4664);
nor U5366 (N_5366,N_4103,N_4776);
or U5367 (N_5367,N_4797,N_4891);
and U5368 (N_5368,N_4872,N_4458);
nand U5369 (N_5369,N_4319,N_4261);
nand U5370 (N_5370,N_4831,N_4827);
or U5371 (N_5371,N_4334,N_4254);
nand U5372 (N_5372,N_4467,N_4414);
nand U5373 (N_5373,N_4179,N_4852);
or U5374 (N_5374,N_4033,N_4145);
and U5375 (N_5375,N_4715,N_4473);
and U5376 (N_5376,N_4307,N_4816);
nor U5377 (N_5377,N_4618,N_4847);
and U5378 (N_5378,N_4031,N_4011);
nand U5379 (N_5379,N_4728,N_4622);
or U5380 (N_5380,N_4308,N_4407);
or U5381 (N_5381,N_4325,N_4632);
nand U5382 (N_5382,N_4239,N_4068);
or U5383 (N_5383,N_4152,N_4915);
and U5384 (N_5384,N_4601,N_4625);
nand U5385 (N_5385,N_4837,N_4336);
nand U5386 (N_5386,N_4213,N_4720);
and U5387 (N_5387,N_4208,N_4617);
nor U5388 (N_5388,N_4096,N_4036);
nand U5389 (N_5389,N_4811,N_4665);
and U5390 (N_5390,N_4091,N_4996);
nor U5391 (N_5391,N_4598,N_4513);
nand U5392 (N_5392,N_4066,N_4759);
nand U5393 (N_5393,N_4496,N_4930);
nand U5394 (N_5394,N_4457,N_4654);
and U5395 (N_5395,N_4006,N_4868);
and U5396 (N_5396,N_4931,N_4840);
nand U5397 (N_5397,N_4278,N_4500);
nand U5398 (N_5398,N_4730,N_4051);
nor U5399 (N_5399,N_4456,N_4196);
or U5400 (N_5400,N_4088,N_4159);
nor U5401 (N_5401,N_4535,N_4634);
nand U5402 (N_5402,N_4584,N_4572);
or U5403 (N_5403,N_4453,N_4032);
nand U5404 (N_5404,N_4627,N_4102);
nor U5405 (N_5405,N_4470,N_4766);
or U5406 (N_5406,N_4449,N_4494);
and U5407 (N_5407,N_4527,N_4413);
or U5408 (N_5408,N_4971,N_4005);
or U5409 (N_5409,N_4312,N_4929);
and U5410 (N_5410,N_4812,N_4288);
and U5411 (N_5411,N_4805,N_4887);
nand U5412 (N_5412,N_4379,N_4631);
nor U5413 (N_5413,N_4131,N_4560);
and U5414 (N_5414,N_4243,N_4828);
nor U5415 (N_5415,N_4731,N_4870);
nor U5416 (N_5416,N_4962,N_4063);
or U5417 (N_5417,N_4167,N_4330);
and U5418 (N_5418,N_4117,N_4689);
or U5419 (N_5419,N_4579,N_4803);
and U5420 (N_5420,N_4289,N_4194);
nor U5421 (N_5421,N_4442,N_4989);
nand U5422 (N_5422,N_4262,N_4350);
or U5423 (N_5423,N_4089,N_4495);
or U5424 (N_5424,N_4819,N_4951);
nor U5425 (N_5425,N_4052,N_4574);
and U5426 (N_5426,N_4859,N_4788);
xnor U5427 (N_5427,N_4304,N_4839);
nor U5428 (N_5428,N_4140,N_4988);
nor U5429 (N_5429,N_4226,N_4808);
nand U5430 (N_5430,N_4077,N_4418);
xnor U5431 (N_5431,N_4240,N_4080);
nor U5432 (N_5432,N_4263,N_4919);
and U5433 (N_5433,N_4871,N_4039);
and U5434 (N_5434,N_4402,N_4378);
or U5435 (N_5435,N_4222,N_4389);
nor U5436 (N_5436,N_4944,N_4519);
and U5437 (N_5437,N_4509,N_4716);
nor U5438 (N_5438,N_4696,N_4396);
and U5439 (N_5439,N_4161,N_4067);
or U5440 (N_5440,N_4064,N_4591);
or U5441 (N_5441,N_4371,N_4727);
nor U5442 (N_5442,N_4049,N_4020);
nand U5443 (N_5443,N_4939,N_4538);
or U5444 (N_5444,N_4157,N_4471);
or U5445 (N_5445,N_4296,N_4027);
nand U5446 (N_5446,N_4858,N_4258);
or U5447 (N_5447,N_4235,N_4155);
nor U5448 (N_5448,N_4136,N_4661);
or U5449 (N_5449,N_4920,N_4787);
or U5450 (N_5450,N_4994,N_4834);
or U5451 (N_5451,N_4644,N_4206);
or U5452 (N_5452,N_4794,N_4436);
or U5453 (N_5453,N_4315,N_4016);
and U5454 (N_5454,N_4035,N_4761);
nor U5455 (N_5455,N_4902,N_4923);
and U5456 (N_5456,N_4524,N_4361);
xnor U5457 (N_5457,N_4286,N_4568);
nor U5458 (N_5458,N_4848,N_4104);
and U5459 (N_5459,N_4825,N_4101);
nor U5460 (N_5460,N_4763,N_4245);
and U5461 (N_5461,N_4358,N_4540);
nand U5462 (N_5462,N_4886,N_4149);
and U5463 (N_5463,N_4814,N_4085);
nand U5464 (N_5464,N_4279,N_4956);
nand U5465 (N_5465,N_4231,N_4188);
nand U5466 (N_5466,N_4309,N_4062);
nand U5467 (N_5467,N_4698,N_4861);
and U5468 (N_5468,N_4366,N_4164);
nand U5469 (N_5469,N_4420,N_4078);
or U5470 (N_5470,N_4249,N_4156);
or U5471 (N_5471,N_4642,N_4428);
and U5472 (N_5472,N_4142,N_4917);
nor U5473 (N_5473,N_4775,N_4079);
nor U5474 (N_5474,N_4333,N_4335);
nand U5475 (N_5475,N_4227,N_4126);
and U5476 (N_5476,N_4800,N_4093);
nand U5477 (N_5477,N_4048,N_4925);
nor U5478 (N_5478,N_4544,N_4553);
nand U5479 (N_5479,N_4122,N_4657);
or U5480 (N_5480,N_4488,N_4623);
or U5481 (N_5481,N_4411,N_4749);
and U5482 (N_5482,N_4099,N_4132);
or U5483 (N_5483,N_4633,N_4169);
nand U5484 (N_5484,N_4594,N_4624);
xor U5485 (N_5485,N_4580,N_4522);
nand U5486 (N_5486,N_4274,N_4790);
and U5487 (N_5487,N_4029,N_4310);
or U5488 (N_5488,N_4769,N_4056);
nand U5489 (N_5489,N_4352,N_4130);
nor U5490 (N_5490,N_4410,N_4884);
or U5491 (N_5491,N_4497,N_4701);
and U5492 (N_5492,N_4466,N_4476);
or U5493 (N_5493,N_4346,N_4492);
and U5494 (N_5494,N_4742,N_4252);
and U5495 (N_5495,N_4987,N_4071);
nor U5496 (N_5496,N_4322,N_4751);
nor U5497 (N_5497,N_4922,N_4437);
nand U5498 (N_5498,N_4649,N_4216);
nand U5499 (N_5499,N_4600,N_4238);
nand U5500 (N_5500,N_4743,N_4711);
nand U5501 (N_5501,N_4414,N_4888);
nand U5502 (N_5502,N_4214,N_4903);
and U5503 (N_5503,N_4698,N_4867);
or U5504 (N_5504,N_4345,N_4831);
and U5505 (N_5505,N_4597,N_4471);
and U5506 (N_5506,N_4725,N_4215);
nor U5507 (N_5507,N_4687,N_4615);
and U5508 (N_5508,N_4803,N_4205);
xor U5509 (N_5509,N_4469,N_4385);
and U5510 (N_5510,N_4229,N_4263);
or U5511 (N_5511,N_4812,N_4348);
nor U5512 (N_5512,N_4159,N_4552);
nand U5513 (N_5513,N_4330,N_4883);
nor U5514 (N_5514,N_4251,N_4527);
and U5515 (N_5515,N_4774,N_4970);
nor U5516 (N_5516,N_4661,N_4330);
nand U5517 (N_5517,N_4517,N_4636);
nor U5518 (N_5518,N_4440,N_4748);
nand U5519 (N_5519,N_4147,N_4142);
and U5520 (N_5520,N_4451,N_4966);
or U5521 (N_5521,N_4235,N_4167);
and U5522 (N_5522,N_4059,N_4540);
and U5523 (N_5523,N_4753,N_4147);
nor U5524 (N_5524,N_4551,N_4237);
nand U5525 (N_5525,N_4815,N_4164);
and U5526 (N_5526,N_4162,N_4025);
xnor U5527 (N_5527,N_4513,N_4129);
nand U5528 (N_5528,N_4038,N_4814);
nor U5529 (N_5529,N_4680,N_4090);
and U5530 (N_5530,N_4961,N_4512);
or U5531 (N_5531,N_4159,N_4825);
or U5532 (N_5532,N_4366,N_4872);
xnor U5533 (N_5533,N_4895,N_4629);
and U5534 (N_5534,N_4004,N_4140);
or U5535 (N_5535,N_4814,N_4884);
and U5536 (N_5536,N_4421,N_4123);
nand U5537 (N_5537,N_4242,N_4412);
or U5538 (N_5538,N_4967,N_4478);
and U5539 (N_5539,N_4742,N_4632);
nor U5540 (N_5540,N_4517,N_4254);
and U5541 (N_5541,N_4545,N_4739);
and U5542 (N_5542,N_4970,N_4768);
or U5543 (N_5543,N_4352,N_4659);
nand U5544 (N_5544,N_4453,N_4057);
nor U5545 (N_5545,N_4295,N_4254);
nand U5546 (N_5546,N_4406,N_4606);
or U5547 (N_5547,N_4944,N_4847);
and U5548 (N_5548,N_4903,N_4262);
nand U5549 (N_5549,N_4040,N_4747);
nor U5550 (N_5550,N_4396,N_4678);
nand U5551 (N_5551,N_4334,N_4155);
or U5552 (N_5552,N_4515,N_4367);
and U5553 (N_5553,N_4024,N_4681);
and U5554 (N_5554,N_4880,N_4859);
nand U5555 (N_5555,N_4191,N_4716);
or U5556 (N_5556,N_4318,N_4613);
nand U5557 (N_5557,N_4615,N_4276);
or U5558 (N_5558,N_4457,N_4193);
nor U5559 (N_5559,N_4334,N_4132);
or U5560 (N_5560,N_4339,N_4582);
nor U5561 (N_5561,N_4645,N_4618);
and U5562 (N_5562,N_4968,N_4789);
or U5563 (N_5563,N_4501,N_4494);
nor U5564 (N_5564,N_4677,N_4921);
xor U5565 (N_5565,N_4272,N_4089);
nor U5566 (N_5566,N_4788,N_4193);
nor U5567 (N_5567,N_4921,N_4615);
nand U5568 (N_5568,N_4134,N_4193);
nand U5569 (N_5569,N_4387,N_4959);
and U5570 (N_5570,N_4111,N_4168);
and U5571 (N_5571,N_4204,N_4554);
nand U5572 (N_5572,N_4991,N_4969);
and U5573 (N_5573,N_4461,N_4684);
nand U5574 (N_5574,N_4735,N_4612);
nor U5575 (N_5575,N_4022,N_4838);
nor U5576 (N_5576,N_4896,N_4244);
nor U5577 (N_5577,N_4575,N_4642);
or U5578 (N_5578,N_4302,N_4356);
nand U5579 (N_5579,N_4628,N_4524);
nor U5580 (N_5580,N_4714,N_4067);
and U5581 (N_5581,N_4921,N_4097);
nand U5582 (N_5582,N_4495,N_4621);
or U5583 (N_5583,N_4583,N_4934);
nand U5584 (N_5584,N_4699,N_4604);
and U5585 (N_5585,N_4868,N_4317);
xnor U5586 (N_5586,N_4992,N_4185);
nor U5587 (N_5587,N_4415,N_4170);
and U5588 (N_5588,N_4242,N_4992);
or U5589 (N_5589,N_4098,N_4129);
nand U5590 (N_5590,N_4117,N_4044);
xnor U5591 (N_5591,N_4213,N_4965);
nand U5592 (N_5592,N_4896,N_4766);
and U5593 (N_5593,N_4440,N_4508);
and U5594 (N_5594,N_4439,N_4899);
nand U5595 (N_5595,N_4736,N_4629);
and U5596 (N_5596,N_4885,N_4605);
or U5597 (N_5597,N_4310,N_4507);
or U5598 (N_5598,N_4681,N_4849);
and U5599 (N_5599,N_4174,N_4788);
or U5600 (N_5600,N_4227,N_4546);
or U5601 (N_5601,N_4943,N_4788);
and U5602 (N_5602,N_4587,N_4140);
or U5603 (N_5603,N_4374,N_4289);
or U5604 (N_5604,N_4422,N_4347);
nor U5605 (N_5605,N_4144,N_4289);
nor U5606 (N_5606,N_4564,N_4938);
nor U5607 (N_5607,N_4907,N_4191);
and U5608 (N_5608,N_4900,N_4557);
and U5609 (N_5609,N_4158,N_4932);
and U5610 (N_5610,N_4202,N_4574);
or U5611 (N_5611,N_4860,N_4990);
or U5612 (N_5612,N_4051,N_4824);
and U5613 (N_5613,N_4290,N_4968);
or U5614 (N_5614,N_4972,N_4598);
and U5615 (N_5615,N_4392,N_4202);
nor U5616 (N_5616,N_4508,N_4850);
and U5617 (N_5617,N_4335,N_4864);
or U5618 (N_5618,N_4875,N_4887);
and U5619 (N_5619,N_4527,N_4711);
or U5620 (N_5620,N_4366,N_4764);
and U5621 (N_5621,N_4381,N_4012);
nand U5622 (N_5622,N_4900,N_4957);
and U5623 (N_5623,N_4914,N_4883);
or U5624 (N_5624,N_4098,N_4902);
nor U5625 (N_5625,N_4747,N_4249);
or U5626 (N_5626,N_4366,N_4003);
and U5627 (N_5627,N_4145,N_4490);
and U5628 (N_5628,N_4068,N_4021);
nand U5629 (N_5629,N_4822,N_4215);
and U5630 (N_5630,N_4676,N_4034);
and U5631 (N_5631,N_4921,N_4064);
or U5632 (N_5632,N_4114,N_4419);
nand U5633 (N_5633,N_4099,N_4811);
and U5634 (N_5634,N_4348,N_4060);
and U5635 (N_5635,N_4960,N_4542);
and U5636 (N_5636,N_4232,N_4433);
or U5637 (N_5637,N_4352,N_4166);
nor U5638 (N_5638,N_4069,N_4449);
nand U5639 (N_5639,N_4884,N_4459);
nand U5640 (N_5640,N_4661,N_4799);
and U5641 (N_5641,N_4528,N_4914);
or U5642 (N_5642,N_4271,N_4922);
nand U5643 (N_5643,N_4800,N_4394);
nand U5644 (N_5644,N_4045,N_4263);
or U5645 (N_5645,N_4139,N_4571);
nor U5646 (N_5646,N_4043,N_4721);
nor U5647 (N_5647,N_4527,N_4162);
nand U5648 (N_5648,N_4441,N_4755);
nor U5649 (N_5649,N_4396,N_4574);
nand U5650 (N_5650,N_4174,N_4423);
nor U5651 (N_5651,N_4839,N_4845);
nand U5652 (N_5652,N_4470,N_4965);
nor U5653 (N_5653,N_4455,N_4642);
or U5654 (N_5654,N_4945,N_4254);
and U5655 (N_5655,N_4059,N_4675);
nand U5656 (N_5656,N_4843,N_4971);
or U5657 (N_5657,N_4591,N_4588);
and U5658 (N_5658,N_4930,N_4060);
and U5659 (N_5659,N_4789,N_4644);
and U5660 (N_5660,N_4908,N_4249);
xnor U5661 (N_5661,N_4615,N_4473);
and U5662 (N_5662,N_4952,N_4944);
nor U5663 (N_5663,N_4533,N_4978);
or U5664 (N_5664,N_4156,N_4435);
nand U5665 (N_5665,N_4963,N_4236);
nor U5666 (N_5666,N_4536,N_4635);
nor U5667 (N_5667,N_4023,N_4278);
nor U5668 (N_5668,N_4666,N_4494);
and U5669 (N_5669,N_4923,N_4681);
or U5670 (N_5670,N_4546,N_4830);
and U5671 (N_5671,N_4172,N_4103);
or U5672 (N_5672,N_4138,N_4792);
nor U5673 (N_5673,N_4493,N_4817);
nand U5674 (N_5674,N_4419,N_4905);
or U5675 (N_5675,N_4376,N_4577);
or U5676 (N_5676,N_4737,N_4381);
and U5677 (N_5677,N_4631,N_4853);
nand U5678 (N_5678,N_4367,N_4150);
or U5679 (N_5679,N_4131,N_4112);
or U5680 (N_5680,N_4350,N_4395);
or U5681 (N_5681,N_4753,N_4137);
nor U5682 (N_5682,N_4528,N_4102);
nand U5683 (N_5683,N_4389,N_4263);
nand U5684 (N_5684,N_4067,N_4735);
xnor U5685 (N_5685,N_4728,N_4992);
and U5686 (N_5686,N_4860,N_4070);
nand U5687 (N_5687,N_4258,N_4260);
or U5688 (N_5688,N_4286,N_4778);
xnor U5689 (N_5689,N_4743,N_4745);
or U5690 (N_5690,N_4140,N_4125);
and U5691 (N_5691,N_4567,N_4901);
nand U5692 (N_5692,N_4820,N_4390);
and U5693 (N_5693,N_4587,N_4906);
and U5694 (N_5694,N_4282,N_4763);
nand U5695 (N_5695,N_4028,N_4550);
nand U5696 (N_5696,N_4428,N_4827);
nand U5697 (N_5697,N_4052,N_4988);
nand U5698 (N_5698,N_4829,N_4247);
nor U5699 (N_5699,N_4902,N_4315);
nand U5700 (N_5700,N_4272,N_4742);
nand U5701 (N_5701,N_4155,N_4575);
nor U5702 (N_5702,N_4126,N_4611);
nand U5703 (N_5703,N_4373,N_4744);
nand U5704 (N_5704,N_4886,N_4466);
nor U5705 (N_5705,N_4264,N_4671);
nor U5706 (N_5706,N_4962,N_4437);
nor U5707 (N_5707,N_4132,N_4998);
nor U5708 (N_5708,N_4089,N_4461);
and U5709 (N_5709,N_4221,N_4209);
nand U5710 (N_5710,N_4722,N_4231);
and U5711 (N_5711,N_4205,N_4984);
nor U5712 (N_5712,N_4920,N_4922);
or U5713 (N_5713,N_4776,N_4829);
and U5714 (N_5714,N_4621,N_4892);
nand U5715 (N_5715,N_4551,N_4364);
nor U5716 (N_5716,N_4753,N_4183);
nor U5717 (N_5717,N_4989,N_4891);
nor U5718 (N_5718,N_4694,N_4851);
or U5719 (N_5719,N_4714,N_4338);
or U5720 (N_5720,N_4475,N_4909);
nand U5721 (N_5721,N_4851,N_4796);
nand U5722 (N_5722,N_4258,N_4229);
or U5723 (N_5723,N_4350,N_4017);
nor U5724 (N_5724,N_4782,N_4948);
and U5725 (N_5725,N_4780,N_4296);
nand U5726 (N_5726,N_4361,N_4882);
or U5727 (N_5727,N_4059,N_4688);
nor U5728 (N_5728,N_4012,N_4657);
nor U5729 (N_5729,N_4908,N_4414);
and U5730 (N_5730,N_4343,N_4266);
xor U5731 (N_5731,N_4180,N_4951);
nand U5732 (N_5732,N_4998,N_4628);
nor U5733 (N_5733,N_4849,N_4829);
nand U5734 (N_5734,N_4328,N_4538);
nor U5735 (N_5735,N_4613,N_4986);
nand U5736 (N_5736,N_4303,N_4685);
nor U5737 (N_5737,N_4470,N_4840);
and U5738 (N_5738,N_4634,N_4376);
nor U5739 (N_5739,N_4616,N_4120);
xnor U5740 (N_5740,N_4526,N_4937);
nor U5741 (N_5741,N_4408,N_4015);
nor U5742 (N_5742,N_4522,N_4395);
nor U5743 (N_5743,N_4598,N_4541);
nor U5744 (N_5744,N_4754,N_4177);
and U5745 (N_5745,N_4113,N_4791);
nor U5746 (N_5746,N_4533,N_4474);
or U5747 (N_5747,N_4273,N_4418);
nand U5748 (N_5748,N_4365,N_4718);
nand U5749 (N_5749,N_4071,N_4488);
or U5750 (N_5750,N_4999,N_4471);
nand U5751 (N_5751,N_4298,N_4488);
nor U5752 (N_5752,N_4630,N_4574);
nand U5753 (N_5753,N_4137,N_4500);
and U5754 (N_5754,N_4536,N_4005);
nor U5755 (N_5755,N_4658,N_4708);
nor U5756 (N_5756,N_4327,N_4580);
nand U5757 (N_5757,N_4668,N_4966);
nand U5758 (N_5758,N_4675,N_4888);
nand U5759 (N_5759,N_4010,N_4879);
or U5760 (N_5760,N_4580,N_4107);
or U5761 (N_5761,N_4017,N_4854);
nor U5762 (N_5762,N_4054,N_4396);
nor U5763 (N_5763,N_4176,N_4110);
nor U5764 (N_5764,N_4051,N_4461);
nor U5765 (N_5765,N_4381,N_4101);
xnor U5766 (N_5766,N_4788,N_4119);
nor U5767 (N_5767,N_4165,N_4876);
nor U5768 (N_5768,N_4300,N_4254);
and U5769 (N_5769,N_4429,N_4469);
nor U5770 (N_5770,N_4848,N_4164);
or U5771 (N_5771,N_4570,N_4901);
and U5772 (N_5772,N_4183,N_4389);
nand U5773 (N_5773,N_4826,N_4351);
or U5774 (N_5774,N_4163,N_4573);
nor U5775 (N_5775,N_4526,N_4878);
and U5776 (N_5776,N_4660,N_4053);
or U5777 (N_5777,N_4616,N_4737);
nand U5778 (N_5778,N_4218,N_4560);
and U5779 (N_5779,N_4397,N_4895);
nor U5780 (N_5780,N_4315,N_4548);
or U5781 (N_5781,N_4603,N_4495);
and U5782 (N_5782,N_4763,N_4935);
xor U5783 (N_5783,N_4695,N_4786);
and U5784 (N_5784,N_4952,N_4329);
nand U5785 (N_5785,N_4617,N_4527);
nand U5786 (N_5786,N_4152,N_4087);
nor U5787 (N_5787,N_4624,N_4195);
and U5788 (N_5788,N_4776,N_4505);
nor U5789 (N_5789,N_4648,N_4372);
or U5790 (N_5790,N_4581,N_4538);
or U5791 (N_5791,N_4625,N_4921);
nor U5792 (N_5792,N_4516,N_4778);
nor U5793 (N_5793,N_4404,N_4817);
nor U5794 (N_5794,N_4004,N_4288);
and U5795 (N_5795,N_4437,N_4304);
nor U5796 (N_5796,N_4581,N_4464);
and U5797 (N_5797,N_4646,N_4589);
or U5798 (N_5798,N_4524,N_4364);
or U5799 (N_5799,N_4898,N_4040);
or U5800 (N_5800,N_4980,N_4518);
or U5801 (N_5801,N_4725,N_4380);
and U5802 (N_5802,N_4268,N_4224);
nand U5803 (N_5803,N_4565,N_4200);
or U5804 (N_5804,N_4486,N_4220);
nand U5805 (N_5805,N_4088,N_4891);
nand U5806 (N_5806,N_4009,N_4526);
or U5807 (N_5807,N_4169,N_4058);
nand U5808 (N_5808,N_4774,N_4363);
and U5809 (N_5809,N_4403,N_4762);
and U5810 (N_5810,N_4945,N_4576);
and U5811 (N_5811,N_4043,N_4401);
xor U5812 (N_5812,N_4264,N_4617);
nand U5813 (N_5813,N_4487,N_4826);
nand U5814 (N_5814,N_4017,N_4265);
nand U5815 (N_5815,N_4257,N_4007);
nand U5816 (N_5816,N_4251,N_4140);
and U5817 (N_5817,N_4166,N_4780);
and U5818 (N_5818,N_4043,N_4238);
and U5819 (N_5819,N_4677,N_4605);
or U5820 (N_5820,N_4944,N_4210);
and U5821 (N_5821,N_4923,N_4012);
and U5822 (N_5822,N_4887,N_4483);
nor U5823 (N_5823,N_4641,N_4519);
nand U5824 (N_5824,N_4178,N_4493);
or U5825 (N_5825,N_4723,N_4608);
nor U5826 (N_5826,N_4332,N_4301);
and U5827 (N_5827,N_4203,N_4186);
nor U5828 (N_5828,N_4619,N_4083);
nand U5829 (N_5829,N_4634,N_4093);
nor U5830 (N_5830,N_4986,N_4344);
and U5831 (N_5831,N_4949,N_4488);
nand U5832 (N_5832,N_4042,N_4902);
nor U5833 (N_5833,N_4040,N_4078);
xor U5834 (N_5834,N_4945,N_4926);
nor U5835 (N_5835,N_4901,N_4773);
or U5836 (N_5836,N_4162,N_4121);
nor U5837 (N_5837,N_4150,N_4892);
and U5838 (N_5838,N_4155,N_4468);
nor U5839 (N_5839,N_4501,N_4566);
nand U5840 (N_5840,N_4210,N_4439);
and U5841 (N_5841,N_4201,N_4753);
nand U5842 (N_5842,N_4237,N_4619);
nand U5843 (N_5843,N_4291,N_4368);
or U5844 (N_5844,N_4980,N_4419);
nor U5845 (N_5845,N_4080,N_4670);
nor U5846 (N_5846,N_4283,N_4848);
or U5847 (N_5847,N_4641,N_4604);
nor U5848 (N_5848,N_4705,N_4382);
nor U5849 (N_5849,N_4794,N_4077);
nor U5850 (N_5850,N_4222,N_4650);
nor U5851 (N_5851,N_4820,N_4603);
and U5852 (N_5852,N_4199,N_4613);
nand U5853 (N_5853,N_4993,N_4961);
or U5854 (N_5854,N_4249,N_4186);
nand U5855 (N_5855,N_4226,N_4280);
nand U5856 (N_5856,N_4377,N_4175);
nand U5857 (N_5857,N_4217,N_4867);
nand U5858 (N_5858,N_4618,N_4990);
or U5859 (N_5859,N_4013,N_4859);
nor U5860 (N_5860,N_4638,N_4061);
and U5861 (N_5861,N_4036,N_4037);
and U5862 (N_5862,N_4257,N_4438);
or U5863 (N_5863,N_4281,N_4654);
nor U5864 (N_5864,N_4573,N_4462);
nor U5865 (N_5865,N_4518,N_4748);
and U5866 (N_5866,N_4418,N_4288);
or U5867 (N_5867,N_4855,N_4801);
nor U5868 (N_5868,N_4932,N_4878);
nand U5869 (N_5869,N_4616,N_4592);
or U5870 (N_5870,N_4550,N_4371);
and U5871 (N_5871,N_4496,N_4626);
or U5872 (N_5872,N_4192,N_4341);
or U5873 (N_5873,N_4883,N_4834);
and U5874 (N_5874,N_4699,N_4075);
nand U5875 (N_5875,N_4728,N_4253);
and U5876 (N_5876,N_4998,N_4263);
or U5877 (N_5877,N_4414,N_4804);
and U5878 (N_5878,N_4791,N_4181);
nor U5879 (N_5879,N_4048,N_4815);
and U5880 (N_5880,N_4560,N_4319);
nor U5881 (N_5881,N_4214,N_4739);
and U5882 (N_5882,N_4920,N_4697);
nor U5883 (N_5883,N_4713,N_4883);
nand U5884 (N_5884,N_4514,N_4677);
nor U5885 (N_5885,N_4082,N_4409);
or U5886 (N_5886,N_4092,N_4819);
or U5887 (N_5887,N_4282,N_4693);
nand U5888 (N_5888,N_4614,N_4251);
and U5889 (N_5889,N_4948,N_4800);
or U5890 (N_5890,N_4910,N_4778);
nor U5891 (N_5891,N_4130,N_4617);
or U5892 (N_5892,N_4897,N_4832);
xor U5893 (N_5893,N_4933,N_4534);
and U5894 (N_5894,N_4339,N_4115);
nor U5895 (N_5895,N_4817,N_4068);
nor U5896 (N_5896,N_4718,N_4650);
nand U5897 (N_5897,N_4262,N_4554);
nor U5898 (N_5898,N_4217,N_4624);
or U5899 (N_5899,N_4573,N_4453);
nor U5900 (N_5900,N_4388,N_4514);
nor U5901 (N_5901,N_4571,N_4212);
and U5902 (N_5902,N_4428,N_4188);
and U5903 (N_5903,N_4575,N_4491);
nor U5904 (N_5904,N_4290,N_4956);
or U5905 (N_5905,N_4895,N_4542);
and U5906 (N_5906,N_4976,N_4799);
nand U5907 (N_5907,N_4934,N_4538);
and U5908 (N_5908,N_4479,N_4164);
and U5909 (N_5909,N_4283,N_4275);
and U5910 (N_5910,N_4596,N_4031);
and U5911 (N_5911,N_4367,N_4135);
or U5912 (N_5912,N_4725,N_4560);
nor U5913 (N_5913,N_4794,N_4486);
and U5914 (N_5914,N_4808,N_4111);
nor U5915 (N_5915,N_4725,N_4907);
or U5916 (N_5916,N_4974,N_4833);
nand U5917 (N_5917,N_4375,N_4598);
nor U5918 (N_5918,N_4063,N_4139);
or U5919 (N_5919,N_4633,N_4036);
or U5920 (N_5920,N_4684,N_4168);
nor U5921 (N_5921,N_4990,N_4709);
nor U5922 (N_5922,N_4585,N_4594);
or U5923 (N_5923,N_4575,N_4453);
nor U5924 (N_5924,N_4068,N_4884);
or U5925 (N_5925,N_4158,N_4684);
or U5926 (N_5926,N_4919,N_4981);
and U5927 (N_5927,N_4869,N_4744);
and U5928 (N_5928,N_4370,N_4820);
and U5929 (N_5929,N_4353,N_4023);
or U5930 (N_5930,N_4789,N_4855);
nand U5931 (N_5931,N_4223,N_4665);
and U5932 (N_5932,N_4792,N_4915);
nor U5933 (N_5933,N_4855,N_4695);
and U5934 (N_5934,N_4935,N_4266);
nor U5935 (N_5935,N_4099,N_4496);
nand U5936 (N_5936,N_4877,N_4263);
or U5937 (N_5937,N_4699,N_4370);
nor U5938 (N_5938,N_4472,N_4040);
and U5939 (N_5939,N_4526,N_4933);
and U5940 (N_5940,N_4566,N_4004);
nor U5941 (N_5941,N_4255,N_4560);
or U5942 (N_5942,N_4231,N_4694);
nand U5943 (N_5943,N_4742,N_4730);
nand U5944 (N_5944,N_4952,N_4732);
nor U5945 (N_5945,N_4807,N_4951);
nand U5946 (N_5946,N_4090,N_4668);
nand U5947 (N_5947,N_4034,N_4070);
nor U5948 (N_5948,N_4024,N_4041);
and U5949 (N_5949,N_4547,N_4185);
or U5950 (N_5950,N_4608,N_4101);
nor U5951 (N_5951,N_4711,N_4285);
nor U5952 (N_5952,N_4579,N_4572);
nor U5953 (N_5953,N_4592,N_4487);
or U5954 (N_5954,N_4905,N_4833);
and U5955 (N_5955,N_4180,N_4497);
nor U5956 (N_5956,N_4627,N_4877);
or U5957 (N_5957,N_4506,N_4680);
or U5958 (N_5958,N_4260,N_4063);
nor U5959 (N_5959,N_4213,N_4643);
nor U5960 (N_5960,N_4294,N_4459);
or U5961 (N_5961,N_4825,N_4278);
and U5962 (N_5962,N_4212,N_4490);
nand U5963 (N_5963,N_4006,N_4875);
xnor U5964 (N_5964,N_4827,N_4077);
nor U5965 (N_5965,N_4555,N_4769);
nor U5966 (N_5966,N_4609,N_4219);
and U5967 (N_5967,N_4201,N_4092);
nand U5968 (N_5968,N_4944,N_4335);
nor U5969 (N_5969,N_4071,N_4327);
xor U5970 (N_5970,N_4239,N_4088);
nand U5971 (N_5971,N_4848,N_4423);
and U5972 (N_5972,N_4107,N_4667);
xor U5973 (N_5973,N_4660,N_4369);
nand U5974 (N_5974,N_4672,N_4079);
nor U5975 (N_5975,N_4385,N_4816);
and U5976 (N_5976,N_4026,N_4160);
nand U5977 (N_5977,N_4498,N_4282);
or U5978 (N_5978,N_4629,N_4893);
nand U5979 (N_5979,N_4145,N_4500);
nand U5980 (N_5980,N_4477,N_4459);
and U5981 (N_5981,N_4702,N_4344);
or U5982 (N_5982,N_4324,N_4442);
or U5983 (N_5983,N_4885,N_4340);
nand U5984 (N_5984,N_4011,N_4732);
and U5985 (N_5985,N_4426,N_4165);
nor U5986 (N_5986,N_4595,N_4476);
and U5987 (N_5987,N_4853,N_4172);
nor U5988 (N_5988,N_4816,N_4558);
nand U5989 (N_5989,N_4319,N_4546);
nor U5990 (N_5990,N_4961,N_4283);
and U5991 (N_5991,N_4981,N_4020);
nor U5992 (N_5992,N_4139,N_4532);
and U5993 (N_5993,N_4083,N_4419);
and U5994 (N_5994,N_4517,N_4135);
nor U5995 (N_5995,N_4247,N_4789);
nor U5996 (N_5996,N_4974,N_4076);
or U5997 (N_5997,N_4687,N_4818);
or U5998 (N_5998,N_4452,N_4617);
nor U5999 (N_5999,N_4102,N_4267);
nor U6000 (N_6000,N_5730,N_5246);
nor U6001 (N_6001,N_5256,N_5158);
nand U6002 (N_6002,N_5528,N_5919);
nor U6003 (N_6003,N_5415,N_5386);
and U6004 (N_6004,N_5804,N_5550);
nand U6005 (N_6005,N_5122,N_5400);
nor U6006 (N_6006,N_5947,N_5013);
or U6007 (N_6007,N_5966,N_5992);
nor U6008 (N_6008,N_5378,N_5064);
nand U6009 (N_6009,N_5327,N_5712);
nand U6010 (N_6010,N_5551,N_5505);
and U6011 (N_6011,N_5601,N_5424);
and U6012 (N_6012,N_5135,N_5693);
or U6013 (N_6013,N_5828,N_5362);
and U6014 (N_6014,N_5278,N_5187);
or U6015 (N_6015,N_5879,N_5057);
or U6016 (N_6016,N_5244,N_5124);
nor U6017 (N_6017,N_5322,N_5318);
or U6018 (N_6018,N_5680,N_5722);
nor U6019 (N_6019,N_5569,N_5502);
nor U6020 (N_6020,N_5731,N_5972);
and U6021 (N_6021,N_5269,N_5771);
nor U6022 (N_6022,N_5032,N_5222);
nand U6023 (N_6023,N_5952,N_5916);
nand U6024 (N_6024,N_5240,N_5797);
nor U6025 (N_6025,N_5118,N_5822);
or U6026 (N_6026,N_5204,N_5454);
or U6027 (N_6027,N_5364,N_5393);
nor U6028 (N_6028,N_5043,N_5787);
or U6029 (N_6029,N_5396,N_5446);
or U6030 (N_6030,N_5727,N_5990);
nand U6031 (N_6031,N_5979,N_5027);
and U6032 (N_6032,N_5908,N_5700);
and U6033 (N_6033,N_5156,N_5753);
or U6034 (N_6034,N_5084,N_5615);
and U6035 (N_6035,N_5482,N_5299);
nor U6036 (N_6036,N_5332,N_5785);
and U6037 (N_6037,N_5419,N_5366);
or U6038 (N_6038,N_5850,N_5655);
nor U6039 (N_6039,N_5997,N_5300);
nand U6040 (N_6040,N_5884,N_5987);
and U6041 (N_6041,N_5173,N_5874);
or U6042 (N_6042,N_5654,N_5137);
nor U6043 (N_6043,N_5637,N_5563);
or U6044 (N_6044,N_5737,N_5497);
nand U6045 (N_6045,N_5086,N_5986);
and U6046 (N_6046,N_5112,N_5520);
xnor U6047 (N_6047,N_5420,N_5455);
nand U6048 (N_6048,N_5592,N_5429);
or U6049 (N_6049,N_5447,N_5851);
and U6050 (N_6050,N_5511,N_5843);
nand U6051 (N_6051,N_5656,N_5763);
or U6052 (N_6052,N_5766,N_5684);
or U6053 (N_6053,N_5075,N_5252);
nor U6054 (N_6054,N_5599,N_5573);
or U6055 (N_6055,N_5167,N_5148);
and U6056 (N_6056,N_5006,N_5307);
nor U6057 (N_6057,N_5401,N_5208);
or U6058 (N_6058,N_5186,N_5630);
and U6059 (N_6059,N_5088,N_5217);
or U6060 (N_6060,N_5469,N_5690);
nand U6061 (N_6061,N_5260,N_5312);
nor U6062 (N_6062,N_5263,N_5005);
nand U6063 (N_6063,N_5163,N_5097);
nand U6064 (N_6064,N_5311,N_5930);
and U6065 (N_6065,N_5212,N_5036);
or U6066 (N_6066,N_5931,N_5848);
nand U6067 (N_6067,N_5477,N_5099);
nor U6068 (N_6068,N_5869,N_5872);
nand U6069 (N_6069,N_5669,N_5957);
or U6070 (N_6070,N_5658,N_5819);
and U6071 (N_6071,N_5767,N_5677);
nor U6072 (N_6072,N_5568,N_5255);
or U6073 (N_6073,N_5522,N_5954);
nand U6074 (N_6074,N_5570,N_5679);
or U6075 (N_6075,N_5127,N_5344);
or U6076 (N_6076,N_5800,N_5335);
xor U6077 (N_6077,N_5642,N_5540);
nor U6078 (N_6078,N_5302,N_5154);
or U6079 (N_6079,N_5219,N_5232);
nand U6080 (N_6080,N_5868,N_5065);
nor U6081 (N_6081,N_5385,N_5659);
or U6082 (N_6082,N_5471,N_5985);
or U6083 (N_6083,N_5503,N_5705);
nand U6084 (N_6084,N_5932,N_5309);
nor U6085 (N_6085,N_5545,N_5912);
nor U6086 (N_6086,N_5428,N_5634);
nand U6087 (N_6087,N_5604,N_5360);
and U6088 (N_6088,N_5710,N_5228);
or U6089 (N_6089,N_5350,N_5751);
nand U6090 (N_6090,N_5081,N_5685);
nand U6091 (N_6091,N_5392,N_5480);
or U6092 (N_6092,N_5431,N_5574);
and U6093 (N_6093,N_5319,N_5498);
or U6094 (N_6094,N_5144,N_5519);
nand U6095 (N_6095,N_5418,N_5698);
nor U6096 (N_6096,N_5936,N_5793);
xor U6097 (N_6097,N_5649,N_5547);
nor U6098 (N_6098,N_5702,N_5775);
or U6099 (N_6099,N_5190,N_5661);
and U6100 (N_6100,N_5092,N_5166);
nor U6101 (N_6101,N_5918,N_5830);
and U6102 (N_6102,N_5821,N_5998);
nor U6103 (N_6103,N_5399,N_5372);
and U6104 (N_6104,N_5609,N_5953);
xor U6105 (N_6105,N_5314,N_5526);
or U6106 (N_6106,N_5778,N_5303);
or U6107 (N_6107,N_5116,N_5274);
nand U6108 (N_6108,N_5272,N_5117);
and U6109 (N_6109,N_5963,N_5836);
and U6110 (N_6110,N_5231,N_5859);
nand U6111 (N_6111,N_5862,N_5853);
or U6112 (N_6112,N_5920,N_5580);
or U6113 (N_6113,N_5479,N_5721);
and U6114 (N_6114,N_5904,N_5991);
nor U6115 (N_6115,N_5123,N_5734);
and U6116 (N_6116,N_5978,N_5616);
xnor U6117 (N_6117,N_5713,N_5234);
nand U6118 (N_6118,N_5791,N_5007);
nor U6119 (N_6119,N_5815,N_5939);
nor U6120 (N_6120,N_5769,N_5565);
or U6121 (N_6121,N_5024,N_5411);
and U6122 (N_6122,N_5516,N_5676);
xor U6123 (N_6123,N_5277,N_5313);
nor U6124 (N_6124,N_5041,N_5169);
nor U6125 (N_6125,N_5463,N_5069);
and U6126 (N_6126,N_5298,N_5146);
nand U6127 (N_6127,N_5365,N_5878);
or U6128 (N_6128,N_5254,N_5459);
nor U6129 (N_6129,N_5935,N_5079);
nor U6130 (N_6130,N_5514,N_5308);
nor U6131 (N_6131,N_5268,N_5695);
nand U6132 (N_6132,N_5433,N_5792);
nand U6133 (N_6133,N_5488,N_5683);
and U6134 (N_6134,N_5742,N_5034);
and U6135 (N_6135,N_5098,N_5829);
nor U6136 (N_6136,N_5370,N_5059);
xor U6137 (N_6137,N_5235,N_5476);
and U6138 (N_6138,N_5506,N_5845);
nor U6139 (N_6139,N_5728,N_5371);
nor U6140 (N_6140,N_5648,N_5390);
nor U6141 (N_6141,N_5626,N_5508);
nand U6142 (N_6142,N_5211,N_5668);
nand U6143 (N_6143,N_5128,N_5316);
or U6144 (N_6144,N_5458,N_5635);
nor U6145 (N_6145,N_5923,N_5220);
and U6146 (N_6146,N_5470,N_5320);
nand U6147 (N_6147,N_5968,N_5967);
or U6148 (N_6148,N_5525,N_5178);
nand U6149 (N_6149,N_5180,N_5245);
nor U6150 (N_6150,N_5398,N_5375);
and U6151 (N_6151,N_5215,N_5011);
nor U6152 (N_6152,N_5223,N_5115);
nand U6153 (N_6153,N_5610,N_5445);
nor U6154 (N_6154,N_5515,N_5407);
nor U6155 (N_6155,N_5663,N_5745);
nand U6156 (N_6156,N_5617,N_5780);
and U6157 (N_6157,N_5622,N_5671);
and U6158 (N_6158,N_5554,N_5141);
nor U6159 (N_6159,N_5605,N_5015);
or U6160 (N_6160,N_5326,N_5413);
xnor U6161 (N_6161,N_5743,N_5114);
nor U6162 (N_6162,N_5552,N_5221);
nor U6163 (N_6163,N_5595,N_5287);
nor U6164 (N_6164,N_5395,N_5266);
nor U6165 (N_6165,N_5962,N_5425);
or U6166 (N_6166,N_5139,N_5161);
or U6167 (N_6167,N_5996,N_5964);
nor U6168 (N_6168,N_5132,N_5576);
nor U6169 (N_6169,N_5995,N_5304);
and U6170 (N_6170,N_5310,N_5631);
and U6171 (N_6171,N_5529,N_5073);
nand U6172 (N_6172,N_5280,N_5808);
or U6173 (N_6173,N_5189,N_5261);
nor U6174 (N_6174,N_5941,N_5945);
nor U6175 (N_6175,N_5888,N_5499);
and U6176 (N_6176,N_5898,N_5660);
nand U6177 (N_6177,N_5434,N_5501);
and U6178 (N_6178,N_5134,N_5085);
and U6179 (N_6179,N_5443,N_5909);
and U6180 (N_6180,N_5185,N_5672);
nand U6181 (N_6181,N_5330,N_5051);
nand U6182 (N_6182,N_5182,N_5926);
nor U6183 (N_6183,N_5159,N_5164);
nand U6184 (N_6184,N_5466,N_5607);
or U6185 (N_6185,N_5093,N_5794);
or U6186 (N_6186,N_5121,N_5857);
nor U6187 (N_6187,N_5451,N_5993);
and U6188 (N_6188,N_5184,N_5000);
nor U6189 (N_6189,N_5627,N_5267);
and U6190 (N_6190,N_5799,N_5301);
and U6191 (N_6191,N_5714,N_5746);
and U6192 (N_6192,N_5448,N_5910);
and U6193 (N_6193,N_5810,N_5827);
and U6194 (N_6194,N_5922,N_5854);
and U6195 (N_6195,N_5970,N_5982);
or U6196 (N_6196,N_5588,N_5581);
nor U6197 (N_6197,N_5812,N_5170);
or U6198 (N_6198,N_5549,N_5442);
and U6199 (N_6199,N_5373,N_5294);
nor U6200 (N_6200,N_5773,N_5500);
or U6201 (N_6201,N_5012,N_5847);
and U6202 (N_6202,N_5593,N_5761);
and U6203 (N_6203,N_5072,N_5199);
nand U6204 (N_6204,N_5487,N_5031);
or U6205 (N_6205,N_5571,N_5594);
and U6206 (N_6206,N_5202,N_5297);
or U6207 (N_6207,N_5225,N_5842);
xor U6208 (N_6208,N_5813,N_5844);
and U6209 (N_6209,N_5976,N_5715);
nor U6210 (N_6210,N_5239,N_5160);
nor U6211 (N_6211,N_5014,N_5357);
nor U6212 (N_6212,N_5331,N_5475);
or U6213 (N_6213,N_5193,N_5618);
nand U6214 (N_6214,N_5238,N_5436);
and U6215 (N_6215,N_5484,N_5795);
and U6216 (N_6216,N_5387,N_5296);
or U6217 (N_6217,N_5291,N_5464);
nor U6218 (N_6218,N_5786,N_5461);
nand U6219 (N_6219,N_5612,N_5517);
and U6220 (N_6220,N_5379,N_5271);
and U6221 (N_6221,N_5368,N_5988);
nand U6222 (N_6222,N_5557,N_5747);
and U6223 (N_6223,N_5559,N_5440);
or U6224 (N_6224,N_5546,N_5329);
nor U6225 (N_6225,N_5602,N_5636);
and U6226 (N_6226,N_5864,N_5203);
nor U6227 (N_6227,N_5358,N_5633);
nand U6228 (N_6228,N_5905,N_5347);
or U6229 (N_6229,N_5275,N_5881);
or U6230 (N_6230,N_5183,N_5283);
nand U6231 (N_6231,N_5781,N_5077);
and U6232 (N_6232,N_5566,N_5856);
nor U6233 (N_6233,N_5548,N_5720);
or U6234 (N_6234,N_5858,N_5596);
nor U6235 (N_6235,N_5820,N_5021);
or U6236 (N_6236,N_5348,N_5091);
or U6237 (N_6237,N_5523,N_5218);
nor U6238 (N_6238,N_5645,N_5641);
nor U6239 (N_6239,N_5729,N_5126);
nand U6240 (N_6240,N_5681,N_5374);
or U6241 (N_6241,N_5352,N_5009);
nand U6242 (N_6242,N_5697,N_5017);
nand U6243 (N_6243,N_5068,N_5896);
or U6244 (N_6244,N_5270,N_5070);
and U6245 (N_6245,N_5039,N_5026);
nor U6246 (N_6246,N_5273,N_5054);
nand U6247 (N_6247,N_5136,N_5513);
nand U6248 (N_6248,N_5553,N_5106);
nor U6249 (N_6249,N_5639,N_5748);
or U6250 (N_6250,N_5754,N_5033);
nand U6251 (N_6251,N_5776,N_5403);
nor U6252 (N_6252,N_5956,N_5197);
nand U6253 (N_6253,N_5613,N_5025);
nand U6254 (N_6254,N_5376,N_5994);
nor U6255 (N_6255,N_5414,N_5536);
nor U6256 (N_6256,N_5542,N_5226);
or U6257 (N_6257,N_5831,N_5295);
or U6258 (N_6258,N_5209,N_5638);
nand U6259 (N_6259,N_5597,N_5483);
nand U6260 (N_6260,N_5248,N_5416);
or U6261 (N_6261,N_5789,N_5119);
nor U6262 (N_6262,N_5958,N_5230);
nor U6263 (N_6263,N_5113,N_5140);
nor U6264 (N_6264,N_5758,N_5162);
and U6265 (N_6265,N_5046,N_5678);
nand U6266 (N_6266,N_5380,N_5288);
nor U6267 (N_6267,N_5564,N_5408);
nor U6268 (N_6268,N_5090,N_5866);
nand U6269 (N_6269,N_5176,N_5195);
nand U6270 (N_6270,N_5652,N_5490);
nand U6271 (N_6271,N_5598,N_5768);
nor U6272 (N_6272,N_5726,N_5875);
nand U6273 (N_6273,N_5860,N_5460);
and U6274 (N_6274,N_5435,N_5940);
nand U6275 (N_6275,N_5509,N_5575);
or U6276 (N_6276,N_5543,N_5237);
or U6277 (N_6277,N_5578,N_5210);
nand U6278 (N_6278,N_5003,N_5628);
and U6279 (N_6279,N_5955,N_5760);
nor U6280 (N_6280,N_5801,N_5022);
and U6281 (N_6281,N_5289,N_5504);
and U6282 (N_6282,N_5285,N_5756);
nand U6283 (N_6283,N_5590,N_5129);
nand U6284 (N_6284,N_5462,N_5049);
nand U6285 (N_6285,N_5147,N_5213);
or U6286 (N_6286,N_5651,N_5067);
and U6287 (N_6287,N_5749,N_5556);
and U6288 (N_6288,N_5886,N_5894);
nand U6289 (N_6289,N_5101,N_5196);
nand U6290 (N_6290,N_5739,N_5816);
and U6291 (N_6291,N_5361,N_5871);
or U6292 (N_6292,N_5686,N_5253);
or U6293 (N_6293,N_5491,N_5345);
or U6294 (N_6294,N_5724,N_5201);
or U6295 (N_6295,N_5130,N_5716);
nand U6296 (N_6296,N_5465,N_5432);
or U6297 (N_6297,N_5623,N_5530);
nand U6298 (N_6298,N_5227,N_5143);
or U6299 (N_6299,N_5276,N_5120);
and U6300 (N_6300,N_5111,N_5682);
nand U6301 (N_6301,N_5194,N_5646);
and U6302 (N_6302,N_5507,N_5438);
and U6303 (N_6303,N_5001,N_5561);
or U6304 (N_6304,N_5544,N_5125);
nand U6305 (N_6305,N_5450,N_5611);
xor U6306 (N_6306,N_5619,N_5665);
nor U6307 (N_6307,N_5744,N_5688);
nor U6308 (N_6308,N_5817,N_5579);
or U6309 (N_6309,N_5133,N_5891);
and U6310 (N_6310,N_5089,N_5719);
nor U6311 (N_6311,N_5779,N_5087);
or U6312 (N_6312,N_5493,N_5340);
and U6313 (N_6313,N_5673,N_5948);
and U6314 (N_6314,N_5382,N_5040);
nor U6315 (N_6315,N_5725,N_5381);
nand U6316 (N_6316,N_5803,N_5946);
nand U6317 (N_6317,N_5356,N_5030);
xor U6318 (N_6318,N_5452,N_5152);
and U6319 (N_6319,N_5108,N_5764);
nor U6320 (N_6320,N_5353,N_5305);
nor U6321 (N_6321,N_5583,N_5325);
nor U6322 (N_6322,N_5974,N_5192);
or U6323 (N_6323,N_5572,N_5949);
and U6324 (N_6324,N_5315,N_5770);
nand U6325 (N_6325,N_5625,N_5427);
nor U6326 (N_6326,N_5980,N_5444);
or U6327 (N_6327,N_5174,N_5750);
nand U6328 (N_6328,N_5456,N_5251);
nand U6329 (N_6329,N_5233,N_5082);
nor U6330 (N_6330,N_5914,N_5103);
or U6331 (N_6331,N_5343,N_5841);
or U6332 (N_6332,N_5539,N_5028);
and U6333 (N_6333,N_5535,N_5110);
and U6334 (N_6334,N_5518,N_5558);
nor U6335 (N_6335,N_5247,N_5906);
and U6336 (N_6336,N_5521,N_5938);
and U6337 (N_6337,N_5150,N_5877);
nor U6338 (N_6338,N_5629,N_5474);
or U6339 (N_6339,N_5532,N_5586);
or U6340 (N_6340,N_5707,N_5911);
nor U6341 (N_6341,N_5056,N_5981);
nand U6342 (N_6342,N_5095,N_5306);
or U6343 (N_6343,N_5969,N_5042);
or U6344 (N_6344,N_5989,N_5533);
nor U6345 (N_6345,N_5977,N_5188);
nand U6346 (N_6346,N_5389,N_5324);
or U6347 (N_6347,N_5839,N_5406);
nor U6348 (N_6348,N_5200,N_5047);
nand U6349 (N_6349,N_5587,N_5029);
nand U6350 (N_6350,N_5541,N_5538);
nor U6351 (N_6351,N_5284,N_5907);
xor U6352 (N_6352,N_5740,N_5772);
nand U6353 (N_6353,N_5229,N_5709);
nor U6354 (N_6354,N_5833,N_5402);
and U6355 (N_6355,N_5942,N_5903);
nor U6356 (N_6356,N_5807,N_5614);
and U6357 (N_6357,N_5927,N_5893);
nor U6358 (N_6358,N_5951,N_5242);
nand U6359 (N_6359,N_5870,N_5104);
and U6360 (N_6360,N_5172,N_5074);
nor U6361 (N_6361,N_5080,N_5181);
or U6362 (N_6362,N_5145,N_5489);
or U6363 (N_6363,N_5151,N_5138);
and U6364 (N_6364,N_5512,N_5100);
nor U6365 (N_6365,N_5765,N_5889);
nand U6366 (N_6366,N_5321,N_5788);
or U6367 (N_6367,N_5262,N_5924);
nand U6368 (N_6368,N_5805,N_5653);
or U6369 (N_6369,N_5852,N_5696);
nand U6370 (N_6370,N_5336,N_5346);
or U6371 (N_6371,N_5050,N_5873);
nor U6372 (N_6372,N_5410,N_5534);
xnor U6373 (N_6373,N_5472,N_5895);
and U6374 (N_6374,N_5171,N_5478);
and U6375 (N_6375,N_5259,N_5018);
or U6376 (N_6376,N_5179,N_5045);
xor U6377 (N_6377,N_5008,N_5044);
or U6378 (N_6378,N_5584,N_5354);
nor U6379 (N_6379,N_5224,N_5142);
and U6380 (N_6380,N_5094,N_5249);
nand U6381 (N_6381,N_5608,N_5861);
or U6382 (N_6382,N_5338,N_5704);
and U6383 (N_6383,N_5258,N_5198);
or U6384 (N_6384,N_5060,N_5667);
xnor U6385 (N_6385,N_5823,N_5703);
xor U6386 (N_6386,N_5733,N_5019);
or U6387 (N_6387,N_5759,N_5971);
nor U6388 (N_6388,N_5943,N_5004);
nor U6389 (N_6389,N_5168,N_5915);
nand U6390 (N_6390,N_5577,N_5048);
and U6391 (N_6391,N_5236,N_5790);
and U6392 (N_6392,N_5157,N_5053);
nor U6393 (N_6393,N_5423,N_5369);
nand U6394 (N_6394,N_5706,N_5494);
nor U6395 (N_6395,N_5165,N_5717);
or U6396 (N_6396,N_5965,N_5496);
nand U6397 (N_6397,N_5917,N_5755);
nand U6398 (N_6398,N_5328,N_5711);
and U6399 (N_6399,N_5486,N_5752);
nand U6400 (N_6400,N_5933,N_5061);
or U6401 (N_6401,N_5603,N_5762);
or U6402 (N_6402,N_5723,N_5701);
nand U6403 (N_6403,N_5342,N_5691);
nand U6404 (N_6404,N_5341,N_5333);
nor U6405 (N_6405,N_5632,N_5825);
or U6406 (N_6406,N_5929,N_5205);
and U6407 (N_6407,N_5052,N_5890);
and U6408 (N_6408,N_5624,N_5735);
and U6409 (N_6409,N_5107,N_5286);
nand U6410 (N_6410,N_5153,N_5293);
nand U6411 (N_6411,N_5774,N_5959);
nand U6412 (N_6412,N_5105,N_5206);
and U6413 (N_6413,N_5531,N_5960);
and U6414 (N_6414,N_5035,N_5899);
or U6415 (N_6415,N_5708,N_5317);
nor U6416 (N_6416,N_5582,N_5055);
or U6417 (N_6417,N_5670,N_5837);
or U6418 (N_6418,N_5383,N_5394);
nor U6419 (N_6419,N_5928,N_5846);
or U6420 (N_6420,N_5826,N_5377);
nand U6421 (N_6421,N_5811,N_5687);
and U6422 (N_6422,N_5620,N_5405);
nor U6423 (N_6423,N_5096,N_5351);
or U6424 (N_6424,N_5921,N_5838);
nand U6425 (N_6425,N_5796,N_5880);
nor U6426 (N_6426,N_5950,N_5363);
and U6427 (N_6427,N_5355,N_5243);
or U6428 (N_6428,N_5282,N_5585);
nand U6429 (N_6429,N_5640,N_5757);
nand U6430 (N_6430,N_5692,N_5473);
and U6431 (N_6431,N_5175,N_5281);
nor U6432 (N_6432,N_5944,N_5913);
nand U6433 (N_6433,N_5388,N_5937);
and U6434 (N_6434,N_5897,N_5421);
or U6435 (N_6435,N_5102,N_5718);
nand U6436 (N_6436,N_5863,N_5883);
and U6437 (N_6437,N_5983,N_5892);
and U6438 (N_6438,N_5083,N_5664);
nand U6439 (N_6439,N_5062,N_5984);
and U6440 (N_6440,N_5510,N_5010);
and U6441 (N_6441,N_5384,N_5973);
nor U6442 (N_6442,N_5250,N_5279);
and U6443 (N_6443,N_5606,N_5675);
or U6444 (N_6444,N_5900,N_5887);
and U6445 (N_6445,N_5409,N_5834);
nor U6446 (N_6446,N_5063,N_5885);
nand U6447 (N_6447,N_5023,N_5359);
or U6448 (N_6448,N_5481,N_5736);
nor U6449 (N_6449,N_5782,N_5078);
nand U6450 (N_6450,N_5738,N_5567);
nand U6451 (N_6451,N_5417,N_5058);
nand U6452 (N_6452,N_5323,N_5404);
nand U6453 (N_6453,N_5339,N_5453);
or U6454 (N_6454,N_5650,N_5840);
nand U6455 (N_6455,N_5449,N_5527);
or U6456 (N_6456,N_5732,N_5699);
nor U6457 (N_6457,N_5437,N_5422);
nand U6458 (N_6458,N_5038,N_5867);
or U6459 (N_6459,N_5216,N_5426);
nor U6460 (N_6460,N_5798,N_5643);
xor U6461 (N_6461,N_5002,N_5349);
nand U6462 (N_6462,N_5412,N_5855);
nor U6463 (N_6463,N_5037,N_5802);
nor U6464 (N_6464,N_5076,N_5835);
xor U6465 (N_6465,N_5865,N_5492);
and U6466 (N_6466,N_5397,N_5876);
nor U6467 (N_6467,N_5537,N_5337);
nor U6468 (N_6468,N_5241,N_5824);
nand U6469 (N_6469,N_5662,N_5666);
and U6470 (N_6470,N_5131,N_5560);
and U6471 (N_6471,N_5524,N_5647);
and U6472 (N_6472,N_5694,N_5999);
nand U6473 (N_6473,N_5882,N_5814);
nand U6474 (N_6474,N_5809,N_5149);
nor U6475 (N_6475,N_5902,N_5016);
nand U6476 (N_6476,N_5591,N_5290);
or U6477 (N_6477,N_5901,N_5644);
nor U6478 (N_6478,N_5784,N_5555);
nand U6479 (N_6479,N_5467,N_5600);
and U6480 (N_6480,N_5264,N_5777);
or U6481 (N_6481,N_5020,N_5191);
nor U6482 (N_6482,N_5783,N_5214);
nand U6483 (N_6483,N_5485,N_5367);
or U6484 (N_6484,N_5292,N_5257);
xnor U6485 (N_6485,N_5334,N_5925);
and U6486 (N_6486,N_5849,N_5468);
nor U6487 (N_6487,N_5430,N_5934);
nor U6488 (N_6488,N_5071,N_5818);
and U6489 (N_6489,N_5562,N_5589);
nor U6490 (N_6490,N_5066,N_5265);
nand U6491 (N_6491,N_5832,N_5621);
nand U6492 (N_6492,N_5806,N_5457);
and U6493 (N_6493,N_5109,N_5495);
nand U6494 (N_6494,N_5741,N_5975);
nor U6495 (N_6495,N_5155,N_5207);
and U6496 (N_6496,N_5961,N_5441);
and U6497 (N_6497,N_5657,N_5689);
nand U6498 (N_6498,N_5439,N_5391);
nand U6499 (N_6499,N_5177,N_5674);
or U6500 (N_6500,N_5670,N_5824);
and U6501 (N_6501,N_5762,N_5218);
and U6502 (N_6502,N_5840,N_5137);
nand U6503 (N_6503,N_5403,N_5486);
and U6504 (N_6504,N_5234,N_5279);
nand U6505 (N_6505,N_5521,N_5822);
nor U6506 (N_6506,N_5767,N_5080);
nor U6507 (N_6507,N_5970,N_5744);
nand U6508 (N_6508,N_5773,N_5508);
and U6509 (N_6509,N_5830,N_5566);
nand U6510 (N_6510,N_5837,N_5665);
or U6511 (N_6511,N_5598,N_5888);
nand U6512 (N_6512,N_5587,N_5292);
and U6513 (N_6513,N_5707,N_5975);
or U6514 (N_6514,N_5776,N_5481);
nand U6515 (N_6515,N_5749,N_5257);
nor U6516 (N_6516,N_5149,N_5676);
and U6517 (N_6517,N_5992,N_5041);
or U6518 (N_6518,N_5393,N_5974);
or U6519 (N_6519,N_5342,N_5154);
nand U6520 (N_6520,N_5173,N_5469);
nand U6521 (N_6521,N_5124,N_5907);
and U6522 (N_6522,N_5878,N_5403);
or U6523 (N_6523,N_5863,N_5055);
and U6524 (N_6524,N_5526,N_5562);
xnor U6525 (N_6525,N_5128,N_5073);
nor U6526 (N_6526,N_5959,N_5372);
nor U6527 (N_6527,N_5422,N_5467);
or U6528 (N_6528,N_5575,N_5154);
and U6529 (N_6529,N_5833,N_5290);
xnor U6530 (N_6530,N_5693,N_5256);
and U6531 (N_6531,N_5953,N_5687);
nor U6532 (N_6532,N_5996,N_5797);
nor U6533 (N_6533,N_5149,N_5044);
nor U6534 (N_6534,N_5479,N_5038);
nor U6535 (N_6535,N_5044,N_5582);
nand U6536 (N_6536,N_5048,N_5888);
nor U6537 (N_6537,N_5932,N_5808);
or U6538 (N_6538,N_5712,N_5490);
nand U6539 (N_6539,N_5258,N_5951);
and U6540 (N_6540,N_5096,N_5246);
or U6541 (N_6541,N_5773,N_5057);
nand U6542 (N_6542,N_5794,N_5253);
nand U6543 (N_6543,N_5407,N_5997);
nand U6544 (N_6544,N_5532,N_5906);
nand U6545 (N_6545,N_5473,N_5810);
nor U6546 (N_6546,N_5703,N_5811);
xnor U6547 (N_6547,N_5464,N_5162);
nand U6548 (N_6548,N_5520,N_5303);
nand U6549 (N_6549,N_5339,N_5575);
or U6550 (N_6550,N_5714,N_5873);
and U6551 (N_6551,N_5869,N_5177);
nor U6552 (N_6552,N_5007,N_5743);
nor U6553 (N_6553,N_5901,N_5736);
and U6554 (N_6554,N_5813,N_5070);
nor U6555 (N_6555,N_5335,N_5199);
and U6556 (N_6556,N_5181,N_5914);
or U6557 (N_6557,N_5089,N_5467);
and U6558 (N_6558,N_5639,N_5491);
nand U6559 (N_6559,N_5815,N_5860);
nand U6560 (N_6560,N_5655,N_5957);
nand U6561 (N_6561,N_5545,N_5829);
and U6562 (N_6562,N_5130,N_5094);
or U6563 (N_6563,N_5217,N_5697);
and U6564 (N_6564,N_5344,N_5229);
and U6565 (N_6565,N_5408,N_5766);
or U6566 (N_6566,N_5201,N_5795);
or U6567 (N_6567,N_5609,N_5631);
nor U6568 (N_6568,N_5405,N_5471);
nor U6569 (N_6569,N_5504,N_5772);
and U6570 (N_6570,N_5048,N_5104);
nand U6571 (N_6571,N_5141,N_5163);
or U6572 (N_6572,N_5291,N_5461);
or U6573 (N_6573,N_5098,N_5308);
nor U6574 (N_6574,N_5197,N_5133);
nor U6575 (N_6575,N_5013,N_5598);
or U6576 (N_6576,N_5589,N_5815);
and U6577 (N_6577,N_5490,N_5574);
nor U6578 (N_6578,N_5738,N_5328);
nor U6579 (N_6579,N_5659,N_5611);
nor U6580 (N_6580,N_5033,N_5293);
xor U6581 (N_6581,N_5409,N_5081);
nor U6582 (N_6582,N_5888,N_5294);
and U6583 (N_6583,N_5470,N_5277);
and U6584 (N_6584,N_5425,N_5535);
and U6585 (N_6585,N_5658,N_5752);
nand U6586 (N_6586,N_5134,N_5475);
nor U6587 (N_6587,N_5155,N_5759);
nand U6588 (N_6588,N_5623,N_5281);
or U6589 (N_6589,N_5503,N_5605);
nor U6590 (N_6590,N_5723,N_5893);
or U6591 (N_6591,N_5424,N_5508);
or U6592 (N_6592,N_5475,N_5139);
nand U6593 (N_6593,N_5155,N_5240);
nand U6594 (N_6594,N_5733,N_5072);
or U6595 (N_6595,N_5283,N_5443);
and U6596 (N_6596,N_5909,N_5264);
or U6597 (N_6597,N_5029,N_5330);
nand U6598 (N_6598,N_5089,N_5664);
or U6599 (N_6599,N_5776,N_5214);
and U6600 (N_6600,N_5311,N_5607);
nor U6601 (N_6601,N_5370,N_5351);
nand U6602 (N_6602,N_5459,N_5404);
and U6603 (N_6603,N_5832,N_5591);
and U6604 (N_6604,N_5052,N_5277);
nor U6605 (N_6605,N_5176,N_5678);
xnor U6606 (N_6606,N_5862,N_5437);
and U6607 (N_6607,N_5439,N_5642);
xor U6608 (N_6608,N_5226,N_5786);
and U6609 (N_6609,N_5194,N_5335);
and U6610 (N_6610,N_5239,N_5972);
and U6611 (N_6611,N_5074,N_5441);
nand U6612 (N_6612,N_5819,N_5789);
and U6613 (N_6613,N_5786,N_5504);
nand U6614 (N_6614,N_5181,N_5196);
or U6615 (N_6615,N_5244,N_5287);
nor U6616 (N_6616,N_5788,N_5928);
and U6617 (N_6617,N_5399,N_5087);
and U6618 (N_6618,N_5565,N_5761);
or U6619 (N_6619,N_5542,N_5421);
or U6620 (N_6620,N_5480,N_5507);
or U6621 (N_6621,N_5002,N_5094);
nand U6622 (N_6622,N_5564,N_5355);
nor U6623 (N_6623,N_5812,N_5077);
or U6624 (N_6624,N_5552,N_5476);
and U6625 (N_6625,N_5455,N_5721);
or U6626 (N_6626,N_5086,N_5487);
and U6627 (N_6627,N_5696,N_5180);
nand U6628 (N_6628,N_5274,N_5808);
nand U6629 (N_6629,N_5684,N_5476);
nor U6630 (N_6630,N_5279,N_5437);
nand U6631 (N_6631,N_5697,N_5852);
and U6632 (N_6632,N_5930,N_5612);
or U6633 (N_6633,N_5865,N_5011);
nand U6634 (N_6634,N_5767,N_5293);
nand U6635 (N_6635,N_5109,N_5600);
nand U6636 (N_6636,N_5314,N_5924);
nor U6637 (N_6637,N_5879,N_5389);
nor U6638 (N_6638,N_5373,N_5411);
and U6639 (N_6639,N_5311,N_5800);
nand U6640 (N_6640,N_5749,N_5550);
or U6641 (N_6641,N_5304,N_5315);
nor U6642 (N_6642,N_5336,N_5020);
nand U6643 (N_6643,N_5412,N_5194);
and U6644 (N_6644,N_5546,N_5070);
nand U6645 (N_6645,N_5816,N_5909);
nand U6646 (N_6646,N_5129,N_5687);
nor U6647 (N_6647,N_5661,N_5338);
or U6648 (N_6648,N_5679,N_5202);
nand U6649 (N_6649,N_5235,N_5004);
nor U6650 (N_6650,N_5018,N_5353);
or U6651 (N_6651,N_5177,N_5199);
or U6652 (N_6652,N_5649,N_5979);
nand U6653 (N_6653,N_5495,N_5118);
nor U6654 (N_6654,N_5674,N_5229);
nor U6655 (N_6655,N_5171,N_5881);
or U6656 (N_6656,N_5605,N_5056);
nor U6657 (N_6657,N_5701,N_5730);
xnor U6658 (N_6658,N_5625,N_5807);
nand U6659 (N_6659,N_5710,N_5099);
and U6660 (N_6660,N_5597,N_5224);
nor U6661 (N_6661,N_5302,N_5473);
nand U6662 (N_6662,N_5406,N_5436);
and U6663 (N_6663,N_5732,N_5733);
or U6664 (N_6664,N_5506,N_5693);
nor U6665 (N_6665,N_5307,N_5168);
or U6666 (N_6666,N_5098,N_5298);
nor U6667 (N_6667,N_5159,N_5652);
or U6668 (N_6668,N_5692,N_5097);
nor U6669 (N_6669,N_5014,N_5054);
nor U6670 (N_6670,N_5770,N_5052);
and U6671 (N_6671,N_5794,N_5954);
and U6672 (N_6672,N_5068,N_5671);
and U6673 (N_6673,N_5438,N_5154);
xor U6674 (N_6674,N_5871,N_5616);
nor U6675 (N_6675,N_5797,N_5526);
and U6676 (N_6676,N_5580,N_5493);
or U6677 (N_6677,N_5211,N_5872);
xnor U6678 (N_6678,N_5944,N_5516);
or U6679 (N_6679,N_5606,N_5226);
or U6680 (N_6680,N_5028,N_5989);
nor U6681 (N_6681,N_5926,N_5235);
nand U6682 (N_6682,N_5844,N_5929);
nor U6683 (N_6683,N_5519,N_5179);
and U6684 (N_6684,N_5038,N_5236);
nor U6685 (N_6685,N_5433,N_5724);
nand U6686 (N_6686,N_5445,N_5296);
nor U6687 (N_6687,N_5570,N_5149);
nand U6688 (N_6688,N_5424,N_5756);
and U6689 (N_6689,N_5090,N_5316);
and U6690 (N_6690,N_5552,N_5471);
and U6691 (N_6691,N_5138,N_5858);
nor U6692 (N_6692,N_5806,N_5764);
nand U6693 (N_6693,N_5223,N_5438);
nor U6694 (N_6694,N_5392,N_5129);
nand U6695 (N_6695,N_5617,N_5457);
nand U6696 (N_6696,N_5602,N_5881);
nand U6697 (N_6697,N_5261,N_5731);
nand U6698 (N_6698,N_5205,N_5940);
nor U6699 (N_6699,N_5703,N_5220);
nor U6700 (N_6700,N_5400,N_5851);
nand U6701 (N_6701,N_5349,N_5118);
nor U6702 (N_6702,N_5555,N_5363);
and U6703 (N_6703,N_5384,N_5388);
and U6704 (N_6704,N_5051,N_5541);
or U6705 (N_6705,N_5014,N_5547);
or U6706 (N_6706,N_5198,N_5166);
nand U6707 (N_6707,N_5746,N_5735);
and U6708 (N_6708,N_5295,N_5773);
or U6709 (N_6709,N_5124,N_5271);
nor U6710 (N_6710,N_5427,N_5209);
nor U6711 (N_6711,N_5036,N_5024);
xor U6712 (N_6712,N_5866,N_5509);
nand U6713 (N_6713,N_5987,N_5102);
and U6714 (N_6714,N_5800,N_5312);
nand U6715 (N_6715,N_5146,N_5935);
xnor U6716 (N_6716,N_5408,N_5703);
and U6717 (N_6717,N_5010,N_5350);
nor U6718 (N_6718,N_5907,N_5895);
nor U6719 (N_6719,N_5691,N_5972);
nand U6720 (N_6720,N_5556,N_5828);
nand U6721 (N_6721,N_5977,N_5553);
or U6722 (N_6722,N_5880,N_5427);
or U6723 (N_6723,N_5861,N_5014);
or U6724 (N_6724,N_5096,N_5558);
or U6725 (N_6725,N_5638,N_5565);
and U6726 (N_6726,N_5123,N_5437);
or U6727 (N_6727,N_5725,N_5891);
and U6728 (N_6728,N_5701,N_5836);
nand U6729 (N_6729,N_5907,N_5005);
or U6730 (N_6730,N_5703,N_5852);
and U6731 (N_6731,N_5784,N_5345);
or U6732 (N_6732,N_5556,N_5149);
nand U6733 (N_6733,N_5754,N_5496);
and U6734 (N_6734,N_5468,N_5660);
nand U6735 (N_6735,N_5969,N_5965);
and U6736 (N_6736,N_5608,N_5494);
nand U6737 (N_6737,N_5464,N_5941);
and U6738 (N_6738,N_5309,N_5816);
and U6739 (N_6739,N_5958,N_5597);
nor U6740 (N_6740,N_5652,N_5345);
nor U6741 (N_6741,N_5038,N_5778);
or U6742 (N_6742,N_5521,N_5080);
or U6743 (N_6743,N_5784,N_5192);
nor U6744 (N_6744,N_5941,N_5116);
nand U6745 (N_6745,N_5571,N_5450);
nand U6746 (N_6746,N_5876,N_5461);
nor U6747 (N_6747,N_5725,N_5813);
and U6748 (N_6748,N_5186,N_5329);
nor U6749 (N_6749,N_5406,N_5473);
nand U6750 (N_6750,N_5400,N_5218);
or U6751 (N_6751,N_5509,N_5018);
or U6752 (N_6752,N_5882,N_5093);
nor U6753 (N_6753,N_5968,N_5096);
nor U6754 (N_6754,N_5301,N_5380);
nor U6755 (N_6755,N_5634,N_5075);
and U6756 (N_6756,N_5880,N_5016);
nor U6757 (N_6757,N_5874,N_5644);
and U6758 (N_6758,N_5475,N_5876);
nand U6759 (N_6759,N_5865,N_5761);
nand U6760 (N_6760,N_5251,N_5294);
and U6761 (N_6761,N_5484,N_5605);
or U6762 (N_6762,N_5108,N_5684);
or U6763 (N_6763,N_5083,N_5110);
nor U6764 (N_6764,N_5166,N_5957);
or U6765 (N_6765,N_5299,N_5867);
or U6766 (N_6766,N_5826,N_5933);
and U6767 (N_6767,N_5857,N_5585);
and U6768 (N_6768,N_5070,N_5126);
and U6769 (N_6769,N_5561,N_5133);
nor U6770 (N_6770,N_5716,N_5767);
nand U6771 (N_6771,N_5072,N_5907);
or U6772 (N_6772,N_5424,N_5750);
and U6773 (N_6773,N_5472,N_5871);
and U6774 (N_6774,N_5845,N_5239);
or U6775 (N_6775,N_5160,N_5436);
nand U6776 (N_6776,N_5946,N_5016);
nand U6777 (N_6777,N_5350,N_5307);
nor U6778 (N_6778,N_5359,N_5496);
and U6779 (N_6779,N_5048,N_5084);
nor U6780 (N_6780,N_5062,N_5175);
xnor U6781 (N_6781,N_5722,N_5883);
nand U6782 (N_6782,N_5300,N_5431);
nor U6783 (N_6783,N_5029,N_5178);
or U6784 (N_6784,N_5876,N_5168);
or U6785 (N_6785,N_5653,N_5125);
nand U6786 (N_6786,N_5848,N_5405);
xor U6787 (N_6787,N_5540,N_5972);
or U6788 (N_6788,N_5949,N_5486);
or U6789 (N_6789,N_5432,N_5407);
nor U6790 (N_6790,N_5648,N_5188);
or U6791 (N_6791,N_5973,N_5024);
or U6792 (N_6792,N_5788,N_5940);
and U6793 (N_6793,N_5978,N_5802);
and U6794 (N_6794,N_5688,N_5280);
or U6795 (N_6795,N_5347,N_5584);
and U6796 (N_6796,N_5222,N_5418);
nand U6797 (N_6797,N_5924,N_5635);
nor U6798 (N_6798,N_5164,N_5606);
and U6799 (N_6799,N_5481,N_5225);
and U6800 (N_6800,N_5329,N_5209);
nand U6801 (N_6801,N_5397,N_5367);
and U6802 (N_6802,N_5712,N_5070);
nor U6803 (N_6803,N_5750,N_5215);
and U6804 (N_6804,N_5167,N_5902);
nor U6805 (N_6805,N_5232,N_5301);
nand U6806 (N_6806,N_5033,N_5736);
nand U6807 (N_6807,N_5621,N_5662);
nand U6808 (N_6808,N_5841,N_5451);
and U6809 (N_6809,N_5681,N_5336);
nand U6810 (N_6810,N_5656,N_5905);
and U6811 (N_6811,N_5345,N_5139);
or U6812 (N_6812,N_5511,N_5625);
and U6813 (N_6813,N_5495,N_5890);
nor U6814 (N_6814,N_5973,N_5096);
nand U6815 (N_6815,N_5207,N_5335);
or U6816 (N_6816,N_5020,N_5477);
nand U6817 (N_6817,N_5804,N_5015);
nand U6818 (N_6818,N_5754,N_5603);
nand U6819 (N_6819,N_5317,N_5030);
xnor U6820 (N_6820,N_5659,N_5475);
or U6821 (N_6821,N_5166,N_5146);
and U6822 (N_6822,N_5258,N_5056);
nand U6823 (N_6823,N_5271,N_5726);
nor U6824 (N_6824,N_5442,N_5810);
nand U6825 (N_6825,N_5848,N_5478);
nand U6826 (N_6826,N_5516,N_5422);
and U6827 (N_6827,N_5087,N_5872);
and U6828 (N_6828,N_5190,N_5121);
and U6829 (N_6829,N_5551,N_5312);
and U6830 (N_6830,N_5351,N_5674);
or U6831 (N_6831,N_5633,N_5605);
nand U6832 (N_6832,N_5791,N_5012);
nand U6833 (N_6833,N_5053,N_5489);
nand U6834 (N_6834,N_5536,N_5742);
and U6835 (N_6835,N_5062,N_5694);
and U6836 (N_6836,N_5324,N_5036);
or U6837 (N_6837,N_5745,N_5190);
nand U6838 (N_6838,N_5649,N_5801);
nor U6839 (N_6839,N_5852,N_5900);
or U6840 (N_6840,N_5332,N_5352);
nand U6841 (N_6841,N_5163,N_5071);
nand U6842 (N_6842,N_5061,N_5430);
and U6843 (N_6843,N_5825,N_5792);
and U6844 (N_6844,N_5688,N_5803);
and U6845 (N_6845,N_5054,N_5831);
and U6846 (N_6846,N_5232,N_5247);
and U6847 (N_6847,N_5626,N_5029);
or U6848 (N_6848,N_5589,N_5226);
and U6849 (N_6849,N_5642,N_5829);
nand U6850 (N_6850,N_5129,N_5596);
nand U6851 (N_6851,N_5910,N_5184);
xor U6852 (N_6852,N_5057,N_5833);
or U6853 (N_6853,N_5494,N_5574);
nand U6854 (N_6854,N_5307,N_5496);
nand U6855 (N_6855,N_5198,N_5243);
nand U6856 (N_6856,N_5920,N_5285);
or U6857 (N_6857,N_5307,N_5490);
nor U6858 (N_6858,N_5181,N_5550);
and U6859 (N_6859,N_5188,N_5036);
nor U6860 (N_6860,N_5295,N_5417);
nor U6861 (N_6861,N_5838,N_5181);
and U6862 (N_6862,N_5417,N_5450);
nand U6863 (N_6863,N_5856,N_5745);
and U6864 (N_6864,N_5406,N_5446);
and U6865 (N_6865,N_5826,N_5169);
nor U6866 (N_6866,N_5408,N_5552);
and U6867 (N_6867,N_5745,N_5204);
and U6868 (N_6868,N_5029,N_5465);
nor U6869 (N_6869,N_5720,N_5761);
and U6870 (N_6870,N_5642,N_5968);
and U6871 (N_6871,N_5241,N_5083);
and U6872 (N_6872,N_5487,N_5837);
and U6873 (N_6873,N_5247,N_5584);
nand U6874 (N_6874,N_5033,N_5419);
and U6875 (N_6875,N_5124,N_5115);
and U6876 (N_6876,N_5970,N_5295);
nor U6877 (N_6877,N_5866,N_5508);
nand U6878 (N_6878,N_5530,N_5818);
or U6879 (N_6879,N_5005,N_5824);
nor U6880 (N_6880,N_5740,N_5102);
nand U6881 (N_6881,N_5542,N_5344);
and U6882 (N_6882,N_5933,N_5449);
and U6883 (N_6883,N_5617,N_5615);
and U6884 (N_6884,N_5596,N_5676);
nor U6885 (N_6885,N_5357,N_5097);
or U6886 (N_6886,N_5715,N_5992);
nand U6887 (N_6887,N_5076,N_5496);
nand U6888 (N_6888,N_5354,N_5328);
nand U6889 (N_6889,N_5083,N_5266);
or U6890 (N_6890,N_5765,N_5547);
or U6891 (N_6891,N_5292,N_5504);
nand U6892 (N_6892,N_5747,N_5152);
or U6893 (N_6893,N_5344,N_5948);
nand U6894 (N_6894,N_5084,N_5731);
or U6895 (N_6895,N_5014,N_5169);
and U6896 (N_6896,N_5688,N_5593);
and U6897 (N_6897,N_5099,N_5492);
and U6898 (N_6898,N_5336,N_5442);
xnor U6899 (N_6899,N_5876,N_5167);
nor U6900 (N_6900,N_5090,N_5702);
and U6901 (N_6901,N_5665,N_5442);
nor U6902 (N_6902,N_5751,N_5190);
nand U6903 (N_6903,N_5909,N_5317);
nand U6904 (N_6904,N_5426,N_5965);
and U6905 (N_6905,N_5550,N_5769);
nor U6906 (N_6906,N_5748,N_5659);
or U6907 (N_6907,N_5143,N_5317);
nor U6908 (N_6908,N_5111,N_5223);
and U6909 (N_6909,N_5151,N_5168);
or U6910 (N_6910,N_5259,N_5981);
nor U6911 (N_6911,N_5817,N_5778);
or U6912 (N_6912,N_5448,N_5040);
nand U6913 (N_6913,N_5406,N_5748);
and U6914 (N_6914,N_5539,N_5284);
nand U6915 (N_6915,N_5814,N_5925);
nand U6916 (N_6916,N_5357,N_5902);
nand U6917 (N_6917,N_5854,N_5320);
or U6918 (N_6918,N_5834,N_5140);
and U6919 (N_6919,N_5400,N_5461);
nand U6920 (N_6920,N_5331,N_5425);
and U6921 (N_6921,N_5047,N_5226);
and U6922 (N_6922,N_5133,N_5592);
or U6923 (N_6923,N_5163,N_5924);
and U6924 (N_6924,N_5585,N_5165);
or U6925 (N_6925,N_5439,N_5510);
nor U6926 (N_6926,N_5419,N_5647);
or U6927 (N_6927,N_5746,N_5816);
or U6928 (N_6928,N_5867,N_5917);
or U6929 (N_6929,N_5503,N_5053);
and U6930 (N_6930,N_5040,N_5231);
or U6931 (N_6931,N_5001,N_5027);
nand U6932 (N_6932,N_5515,N_5405);
and U6933 (N_6933,N_5441,N_5059);
nor U6934 (N_6934,N_5363,N_5347);
and U6935 (N_6935,N_5043,N_5824);
nor U6936 (N_6936,N_5875,N_5275);
nand U6937 (N_6937,N_5957,N_5826);
and U6938 (N_6938,N_5736,N_5162);
nor U6939 (N_6939,N_5054,N_5304);
or U6940 (N_6940,N_5212,N_5265);
and U6941 (N_6941,N_5960,N_5686);
xor U6942 (N_6942,N_5053,N_5674);
or U6943 (N_6943,N_5856,N_5492);
and U6944 (N_6944,N_5043,N_5382);
and U6945 (N_6945,N_5736,N_5088);
or U6946 (N_6946,N_5880,N_5178);
and U6947 (N_6947,N_5914,N_5054);
nor U6948 (N_6948,N_5250,N_5367);
or U6949 (N_6949,N_5459,N_5412);
nand U6950 (N_6950,N_5121,N_5878);
and U6951 (N_6951,N_5149,N_5009);
or U6952 (N_6952,N_5887,N_5333);
nand U6953 (N_6953,N_5722,N_5470);
and U6954 (N_6954,N_5491,N_5581);
and U6955 (N_6955,N_5559,N_5305);
or U6956 (N_6956,N_5761,N_5251);
nor U6957 (N_6957,N_5890,N_5306);
nand U6958 (N_6958,N_5218,N_5151);
nand U6959 (N_6959,N_5055,N_5802);
and U6960 (N_6960,N_5015,N_5394);
and U6961 (N_6961,N_5764,N_5074);
nor U6962 (N_6962,N_5615,N_5690);
nand U6963 (N_6963,N_5325,N_5595);
nor U6964 (N_6964,N_5229,N_5023);
nor U6965 (N_6965,N_5723,N_5283);
and U6966 (N_6966,N_5326,N_5291);
or U6967 (N_6967,N_5870,N_5362);
or U6968 (N_6968,N_5953,N_5041);
or U6969 (N_6969,N_5274,N_5959);
and U6970 (N_6970,N_5272,N_5239);
and U6971 (N_6971,N_5848,N_5606);
or U6972 (N_6972,N_5609,N_5375);
nand U6973 (N_6973,N_5243,N_5622);
nand U6974 (N_6974,N_5243,N_5983);
or U6975 (N_6975,N_5408,N_5248);
nor U6976 (N_6976,N_5579,N_5173);
nor U6977 (N_6977,N_5286,N_5600);
nor U6978 (N_6978,N_5620,N_5450);
nand U6979 (N_6979,N_5532,N_5802);
and U6980 (N_6980,N_5288,N_5962);
nor U6981 (N_6981,N_5409,N_5013);
nand U6982 (N_6982,N_5588,N_5649);
or U6983 (N_6983,N_5515,N_5213);
nor U6984 (N_6984,N_5077,N_5756);
or U6985 (N_6985,N_5295,N_5833);
and U6986 (N_6986,N_5465,N_5504);
or U6987 (N_6987,N_5337,N_5089);
or U6988 (N_6988,N_5258,N_5767);
and U6989 (N_6989,N_5753,N_5519);
or U6990 (N_6990,N_5024,N_5998);
nand U6991 (N_6991,N_5632,N_5559);
nor U6992 (N_6992,N_5994,N_5944);
and U6993 (N_6993,N_5268,N_5795);
xnor U6994 (N_6994,N_5224,N_5184);
nand U6995 (N_6995,N_5278,N_5948);
nor U6996 (N_6996,N_5266,N_5529);
and U6997 (N_6997,N_5205,N_5017);
nor U6998 (N_6998,N_5982,N_5590);
and U6999 (N_6999,N_5711,N_5334);
or U7000 (N_7000,N_6829,N_6710);
and U7001 (N_7001,N_6661,N_6298);
nor U7002 (N_7002,N_6217,N_6989);
or U7003 (N_7003,N_6891,N_6443);
nand U7004 (N_7004,N_6343,N_6057);
or U7005 (N_7005,N_6130,N_6004);
nor U7006 (N_7006,N_6736,N_6475);
xnor U7007 (N_7007,N_6812,N_6421);
nor U7008 (N_7008,N_6066,N_6072);
nor U7009 (N_7009,N_6441,N_6593);
nor U7010 (N_7010,N_6694,N_6265);
nor U7011 (N_7011,N_6370,N_6769);
or U7012 (N_7012,N_6333,N_6880);
and U7013 (N_7013,N_6641,N_6925);
nand U7014 (N_7014,N_6949,N_6210);
nor U7015 (N_7015,N_6083,N_6259);
or U7016 (N_7016,N_6348,N_6323);
nor U7017 (N_7017,N_6454,N_6418);
and U7018 (N_7018,N_6584,N_6128);
nand U7019 (N_7019,N_6380,N_6852);
nand U7020 (N_7020,N_6818,N_6195);
or U7021 (N_7021,N_6539,N_6528);
and U7022 (N_7022,N_6378,N_6894);
or U7023 (N_7023,N_6470,N_6801);
nand U7024 (N_7024,N_6100,N_6885);
or U7025 (N_7025,N_6286,N_6342);
nand U7026 (N_7026,N_6501,N_6058);
nor U7027 (N_7027,N_6615,N_6937);
nand U7028 (N_7028,N_6336,N_6645);
or U7029 (N_7029,N_6510,N_6558);
nor U7030 (N_7030,N_6665,N_6244);
nand U7031 (N_7031,N_6858,N_6010);
and U7032 (N_7032,N_6236,N_6177);
and U7033 (N_7033,N_6837,N_6403);
nand U7034 (N_7034,N_6832,N_6126);
xor U7035 (N_7035,N_6803,N_6693);
or U7036 (N_7036,N_6912,N_6432);
or U7037 (N_7037,N_6131,N_6749);
nor U7038 (N_7038,N_6881,N_6563);
or U7039 (N_7039,N_6473,N_6082);
and U7040 (N_7040,N_6377,N_6133);
nand U7041 (N_7041,N_6318,N_6511);
nand U7042 (N_7042,N_6491,N_6260);
or U7043 (N_7043,N_6247,N_6033);
nand U7044 (N_7044,N_6022,N_6146);
nand U7045 (N_7045,N_6723,N_6172);
or U7046 (N_7046,N_6440,N_6412);
nor U7047 (N_7047,N_6163,N_6371);
nand U7048 (N_7048,N_6701,N_6479);
nand U7049 (N_7049,N_6225,N_6149);
or U7050 (N_7050,N_6631,N_6626);
or U7051 (N_7051,N_6923,N_6353);
and U7052 (N_7052,N_6625,N_6819);
and U7053 (N_7053,N_6814,N_6293);
and U7054 (N_7054,N_6411,N_6028);
nor U7055 (N_7055,N_6586,N_6215);
and U7056 (N_7056,N_6171,N_6173);
nand U7057 (N_7057,N_6638,N_6391);
and U7058 (N_7058,N_6277,N_6525);
nand U7059 (N_7059,N_6101,N_6901);
or U7060 (N_7060,N_6484,N_6587);
or U7061 (N_7061,N_6945,N_6692);
nor U7062 (N_7062,N_6597,N_6999);
nand U7063 (N_7063,N_6042,N_6205);
nand U7064 (N_7064,N_6299,N_6822);
nor U7065 (N_7065,N_6538,N_6129);
or U7066 (N_7066,N_6202,N_6482);
and U7067 (N_7067,N_6547,N_6246);
and U7068 (N_7068,N_6843,N_6888);
and U7069 (N_7069,N_6680,N_6513);
and U7070 (N_7070,N_6958,N_6493);
or U7071 (N_7071,N_6972,N_6982);
and U7072 (N_7072,N_6154,N_6867);
nand U7073 (N_7073,N_6959,N_6496);
or U7074 (N_7074,N_6352,N_6571);
nand U7075 (N_7075,N_6142,N_6086);
nand U7076 (N_7076,N_6598,N_6872);
and U7077 (N_7077,N_6366,N_6024);
nand U7078 (N_7078,N_6158,N_6316);
and U7079 (N_7079,N_6237,N_6091);
nand U7080 (N_7080,N_6870,N_6288);
nor U7081 (N_7081,N_6400,N_6752);
nand U7082 (N_7082,N_6595,N_6292);
nor U7083 (N_7083,N_6355,N_6477);
nor U7084 (N_7084,N_6678,N_6415);
or U7085 (N_7085,N_6178,N_6519);
or U7086 (N_7086,N_6255,N_6434);
or U7087 (N_7087,N_6253,N_6036);
or U7088 (N_7088,N_6204,N_6939);
and U7089 (N_7089,N_6241,N_6799);
nor U7090 (N_7090,N_6242,N_6324);
and U7091 (N_7091,N_6719,N_6811);
or U7092 (N_7092,N_6940,N_6676);
or U7093 (N_7093,N_6712,N_6809);
nand U7094 (N_7094,N_6789,N_6385);
xnor U7095 (N_7095,N_6214,N_6389);
and U7096 (N_7096,N_6974,N_6189);
or U7097 (N_7097,N_6798,N_6649);
or U7098 (N_7098,N_6349,N_6656);
and U7099 (N_7099,N_6627,N_6107);
nand U7100 (N_7100,N_6087,N_6469);
or U7101 (N_7101,N_6330,N_6369);
nand U7102 (N_7102,N_6950,N_6953);
nand U7103 (N_7103,N_6927,N_6280);
and U7104 (N_7104,N_6576,N_6766);
or U7105 (N_7105,N_6887,N_6849);
nor U7106 (N_7106,N_6367,N_6933);
nand U7107 (N_7107,N_6644,N_6695);
nand U7108 (N_7108,N_6635,N_6612);
and U7109 (N_7109,N_6398,N_6282);
nor U7110 (N_7110,N_6014,N_6805);
nand U7111 (N_7111,N_6754,N_6900);
nand U7112 (N_7112,N_6979,N_6393);
or U7113 (N_7113,N_6998,N_6851);
nand U7114 (N_7114,N_6170,N_6853);
xor U7115 (N_7115,N_6614,N_6660);
and U7116 (N_7116,N_6565,N_6860);
nand U7117 (N_7117,N_6793,N_6097);
and U7118 (N_7118,N_6842,N_6977);
or U7119 (N_7119,N_6567,N_6704);
or U7120 (N_7120,N_6362,N_6740);
and U7121 (N_7121,N_6971,N_6499);
and U7122 (N_7122,N_6351,N_6015);
and U7123 (N_7123,N_6404,N_6250);
or U7124 (N_7124,N_6850,N_6472);
and U7125 (N_7125,N_6579,N_6985);
or U7126 (N_7126,N_6762,N_6744);
or U7127 (N_7127,N_6630,N_6046);
nor U7128 (N_7128,N_6021,N_6976);
nand U7129 (N_7129,N_6673,N_6228);
nor U7130 (N_7130,N_6183,N_6655);
nand U7131 (N_7131,N_6588,N_6081);
nor U7132 (N_7132,N_6487,N_6148);
or U7133 (N_7133,N_6556,N_6456);
or U7134 (N_7134,N_6451,N_6186);
nor U7135 (N_7135,N_6585,N_6921);
or U7136 (N_7136,N_6827,N_6486);
nand U7137 (N_7137,N_6934,N_6428);
or U7138 (N_7138,N_6738,N_6117);
nand U7139 (N_7139,N_6011,N_6379);
nand U7140 (N_7140,N_6747,N_6720);
or U7141 (N_7141,N_6965,N_6657);
nand U7142 (N_7142,N_6908,N_6007);
and U7143 (N_7143,N_6709,N_6480);
nand U7144 (N_7144,N_6697,N_6700);
nand U7145 (N_7145,N_6254,N_6535);
nand U7146 (N_7146,N_6685,N_6788);
and U7147 (N_7147,N_6460,N_6957);
nor U7148 (N_7148,N_6981,N_6606);
nand U7149 (N_7149,N_6532,N_6941);
nor U7150 (N_7150,N_6537,N_6319);
or U7151 (N_7151,N_6840,N_6284);
and U7152 (N_7152,N_6450,N_6652);
nand U7153 (N_7153,N_6771,N_6116);
xor U7154 (N_7154,N_6229,N_6690);
nand U7155 (N_7155,N_6917,N_6753);
nand U7156 (N_7156,N_6063,N_6208);
and U7157 (N_7157,N_6844,N_6397);
nand U7158 (N_7158,N_6735,N_6806);
nor U7159 (N_7159,N_6031,N_6577);
and U7160 (N_7160,N_6203,N_6113);
or U7161 (N_7161,N_6702,N_6787);
or U7162 (N_7162,N_6359,N_6185);
or U7163 (N_7163,N_6703,N_6313);
nand U7164 (N_7164,N_6727,N_6037);
nand U7165 (N_7165,N_6119,N_6834);
nand U7166 (N_7166,N_6018,N_6152);
or U7167 (N_7167,N_6368,N_6764);
nand U7168 (N_7168,N_6325,N_6713);
or U7169 (N_7169,N_6734,N_6151);
nor U7170 (N_7170,N_6447,N_6760);
nor U7171 (N_7171,N_6121,N_6674);
and U7172 (N_7172,N_6725,N_6309);
nor U7173 (N_7173,N_6105,N_6032);
nor U7174 (N_7174,N_6137,N_6668);
nor U7175 (N_7175,N_6748,N_6497);
nor U7176 (N_7176,N_6162,N_6746);
and U7177 (N_7177,N_6636,N_6138);
nand U7178 (N_7178,N_6431,N_6180);
nor U7179 (N_7179,N_6967,N_6029);
and U7180 (N_7180,N_6104,N_6573);
nand U7181 (N_7181,N_6954,N_6426);
nor U7182 (N_7182,N_6707,N_6624);
or U7183 (N_7183,N_6817,N_6304);
and U7184 (N_7184,N_6591,N_6592);
nor U7185 (N_7185,N_6212,N_6670);
and U7186 (N_7186,N_6013,N_6562);
and U7187 (N_7187,N_6227,N_6845);
and U7188 (N_7188,N_6886,N_6874);
nor U7189 (N_7189,N_6653,N_6808);
nor U7190 (N_7190,N_6596,N_6303);
or U7191 (N_7191,N_6495,N_6581);
nor U7192 (N_7192,N_6948,N_6270);
nand U7193 (N_7193,N_6932,N_6669);
and U7194 (N_7194,N_6297,N_6308);
or U7195 (N_7195,N_6272,N_6181);
or U7196 (N_7196,N_6085,N_6341);
or U7197 (N_7197,N_6751,N_6914);
nand U7198 (N_7198,N_6448,N_6381);
nand U7199 (N_7199,N_6508,N_6252);
and U7200 (N_7200,N_6048,N_6728);
nand U7201 (N_7201,N_6768,N_6281);
nand U7202 (N_7202,N_6980,N_6759);
or U7203 (N_7203,N_6865,N_6618);
nor U7204 (N_7204,N_6446,N_6708);
or U7205 (N_7205,N_6603,N_6453);
xnor U7206 (N_7206,N_6120,N_6873);
and U7207 (N_7207,N_6098,N_6485);
and U7208 (N_7208,N_6039,N_6311);
nor U7209 (N_7209,N_6717,N_6836);
or U7210 (N_7210,N_6276,N_6060);
or U7211 (N_7211,N_6053,N_6111);
and U7212 (N_7212,N_6970,N_6966);
and U7213 (N_7213,N_6339,N_6758);
nand U7214 (N_7214,N_6005,N_6876);
xor U7215 (N_7215,N_6729,N_6190);
or U7216 (N_7216,N_6517,N_6640);
and U7217 (N_7217,N_6145,N_6468);
or U7218 (N_7218,N_6607,N_6350);
and U7219 (N_7219,N_6675,N_6092);
nor U7220 (N_7220,N_6034,N_6340);
nor U7221 (N_7221,N_6463,N_6582);
and U7222 (N_7222,N_6188,N_6975);
nand U7223 (N_7223,N_6893,N_6016);
or U7224 (N_7224,N_6429,N_6020);
nand U7225 (N_7225,N_6821,N_6781);
nand U7226 (N_7226,N_6983,N_6938);
or U7227 (N_7227,N_6964,N_6416);
nor U7228 (N_7228,N_6012,N_6155);
or U7229 (N_7229,N_6346,N_6520);
or U7230 (N_7230,N_6363,N_6838);
nand U7231 (N_7231,N_6796,N_6521);
and U7232 (N_7232,N_6273,N_6605);
nand U7233 (N_7233,N_6604,N_6364);
or U7234 (N_7234,N_6248,N_6540);
or U7235 (N_7235,N_6731,N_6628);
nor U7236 (N_7236,N_6667,N_6962);
or U7237 (N_7237,N_6399,N_6716);
and U7238 (N_7238,N_6159,N_6686);
nand U7239 (N_7239,N_6461,N_6220);
and U7240 (N_7240,N_6191,N_6533);
nor U7241 (N_7241,N_6909,N_6414);
nor U7242 (N_7242,N_6643,N_6462);
and U7243 (N_7243,N_6763,N_6095);
xnor U7244 (N_7244,N_6561,N_6001);
nand U7245 (N_7245,N_6386,N_6542);
nand U7246 (N_7246,N_6049,N_6489);
xor U7247 (N_7247,N_6507,N_6218);
nand U7248 (N_7248,N_6356,N_6772);
and U7249 (N_7249,N_6526,N_6407);
nor U7250 (N_7250,N_6541,N_6503);
nor U7251 (N_7251,N_6930,N_6813);
nor U7252 (N_7252,N_6358,N_6616);
and U7253 (N_7253,N_6310,N_6984);
or U7254 (N_7254,N_6935,N_6471);
nor U7255 (N_7255,N_6619,N_6402);
nand U7256 (N_7256,N_6884,N_6642);
and U7257 (N_7257,N_6164,N_6165);
nand U7258 (N_7258,N_6960,N_6854);
or U7259 (N_7259,N_6622,N_6928);
or U7260 (N_7260,N_6544,N_6094);
and U7261 (N_7261,N_6554,N_6848);
xor U7262 (N_7262,N_6677,N_6125);
and U7263 (N_7263,N_6384,N_6502);
and U7264 (N_7264,N_6687,N_6807);
nand U7265 (N_7265,N_6345,N_6417);
nand U7266 (N_7266,N_6682,N_6422);
and U7267 (N_7267,N_6207,N_6611);
nor U7268 (N_7268,N_6266,N_6846);
and U7269 (N_7269,N_6823,N_6936);
nand U7270 (N_7270,N_6509,N_6816);
nor U7271 (N_7271,N_6040,N_6841);
and U7272 (N_7272,N_6955,N_6500);
xnor U7273 (N_7273,N_6056,N_6051);
nand U7274 (N_7274,N_6742,N_6833);
nand U7275 (N_7275,N_6123,N_6196);
nand U7276 (N_7276,N_6903,N_6200);
and U7277 (N_7277,N_6904,N_6099);
or U7278 (N_7278,N_6257,N_6156);
nand U7279 (N_7279,N_6791,N_6911);
nand U7280 (N_7280,N_6770,N_6103);
and U7281 (N_7281,N_6394,N_6375);
and U7282 (N_7282,N_6439,N_6756);
and U7283 (N_7283,N_6483,N_6683);
nor U7284 (N_7284,N_6869,N_6739);
nand U7285 (N_7285,N_6376,N_6529);
nand U7286 (N_7286,N_6724,N_6944);
nand U7287 (N_7287,N_6179,N_6409);
and U7288 (N_7288,N_6922,N_6613);
and U7289 (N_7289,N_6327,N_6354);
or U7290 (N_7290,N_6522,N_6344);
nand U7291 (N_7291,N_6147,N_6637);
and U7292 (N_7292,N_6372,N_6546);
and U7293 (N_7293,N_6498,N_6919);
and U7294 (N_7294,N_6140,N_6564);
and U7295 (N_7295,N_6420,N_6224);
nor U7296 (N_7296,N_6124,N_6531);
nor U7297 (N_7297,N_6863,N_6289);
or U7298 (N_7298,N_6054,N_6396);
or U7299 (N_7299,N_6910,N_6251);
or U7300 (N_7300,N_6317,N_6608);
or U7301 (N_7301,N_6610,N_6599);
nor U7302 (N_7302,N_6868,N_6992);
and U7303 (N_7303,N_6824,N_6750);
and U7304 (N_7304,N_6335,N_6296);
nor U7305 (N_7305,N_6523,N_6698);
nor U7306 (N_7306,N_6390,N_6073);
nand U7307 (N_7307,N_6074,N_6861);
or U7308 (N_7308,N_6264,N_6688);
nand U7309 (N_7309,N_6830,N_6826);
and U7310 (N_7310,N_6524,N_6575);
nor U7311 (N_7311,N_6629,N_6465);
and U7312 (N_7312,N_6926,N_6786);
nand U7313 (N_7313,N_6895,N_6069);
and U7314 (N_7314,N_6176,N_6915);
nor U7315 (N_7315,N_6757,N_6552);
or U7316 (N_7316,N_6328,N_6516);
and U7317 (N_7317,N_6387,N_6182);
or U7318 (N_7318,N_6408,N_6942);
or U7319 (N_7319,N_6580,N_6589);
or U7320 (N_7320,N_6679,N_6263);
or U7321 (N_7321,N_6305,N_6433);
and U7322 (N_7322,N_6947,N_6570);
and U7323 (N_7323,N_6518,N_6543);
or U7324 (N_7324,N_6231,N_6916);
and U7325 (N_7325,N_6436,N_6550);
nand U7326 (N_7326,N_6150,N_6777);
nor U7327 (N_7327,N_6139,N_6043);
nand U7328 (N_7328,N_6184,N_6206);
or U7329 (N_7329,N_6361,N_6650);
nand U7330 (N_7330,N_6442,N_6783);
or U7331 (N_7331,N_6347,N_6108);
nor U7332 (N_7332,N_6968,N_6437);
nor U7333 (N_7333,N_6425,N_6249);
and U7334 (N_7334,N_6672,N_6291);
nor U7335 (N_7335,N_6088,N_6044);
and U7336 (N_7336,N_6157,N_6357);
or U7337 (N_7337,N_6952,N_6096);
or U7338 (N_7338,N_6135,N_6320);
or U7339 (N_7339,N_6951,N_6623);
nand U7340 (N_7340,N_6711,N_6035);
nor U7341 (N_7341,N_6153,N_6560);
and U7342 (N_7342,N_6905,N_6127);
or U7343 (N_7343,N_6855,N_6659);
nor U7344 (N_7344,N_6551,N_6134);
nor U7345 (N_7345,N_6654,N_6337);
and U7346 (N_7346,N_6267,N_6492);
or U7347 (N_7347,N_6019,N_6230);
or U7348 (N_7348,N_6555,N_6794);
and U7349 (N_7349,N_6071,N_6197);
and U7350 (N_7350,N_6000,N_6144);
and U7351 (N_7351,N_6233,N_6080);
and U7352 (N_7352,N_6785,N_6601);
nand U7353 (N_7353,N_6030,N_6114);
nand U7354 (N_7354,N_6681,N_6474);
or U7355 (N_7355,N_6706,N_6194);
nand U7356 (N_7356,N_6913,N_6864);
nand U7357 (N_7357,N_6285,N_6906);
nor U7358 (N_7358,N_6201,N_6295);
nor U7359 (N_7359,N_6279,N_6232);
and U7360 (N_7360,N_6223,N_6430);
nand U7361 (N_7361,N_6025,N_6988);
or U7362 (N_7362,N_6294,N_6553);
nor U7363 (N_7363,N_6234,N_6055);
and U7364 (N_7364,N_6780,N_6792);
or U7365 (N_7365,N_6856,N_6578);
or U7366 (N_7366,N_6920,N_6662);
nand U7367 (N_7367,N_6892,N_6963);
and U7368 (N_7368,N_6459,N_6222);
nand U7369 (N_7369,N_6767,N_6382);
nor U7370 (N_7370,N_6115,N_6102);
nor U7371 (N_7371,N_6847,N_6755);
nor U7372 (N_7372,N_6790,N_6275);
nand U7373 (N_7373,N_6026,N_6090);
nor U7374 (N_7374,N_6269,N_6600);
nor U7375 (N_7375,N_6240,N_6047);
or U7376 (N_7376,N_6061,N_6388);
and U7377 (N_7377,N_6997,N_6271);
and U7378 (N_7378,N_6978,N_6122);
nand U7379 (N_7379,N_6312,N_6326);
xnor U7380 (N_7380,N_6797,N_6219);
nor U7381 (N_7381,N_6986,N_6718);
or U7382 (N_7382,N_6689,N_6877);
and U7383 (N_7383,N_6765,N_6410);
and U7384 (N_7384,N_6245,N_6559);
nand U7385 (N_7385,N_6478,N_6365);
nor U7386 (N_7386,N_6902,N_6490);
nand U7387 (N_7387,N_6338,N_6078);
nand U7388 (N_7388,N_6070,N_6632);
nand U7389 (N_7389,N_6775,N_6721);
nor U7390 (N_7390,N_6776,N_6302);
and U7391 (N_7391,N_6737,N_6545);
nor U7392 (N_7392,N_6859,N_6332);
and U7393 (N_7393,N_6946,N_6109);
nor U7394 (N_7394,N_6435,N_6882);
or U7395 (N_7395,N_6574,N_6136);
or U7396 (N_7396,N_6160,N_6994);
or U7397 (N_7397,N_6699,N_6956);
and U7398 (N_7398,N_6169,N_6514);
xor U7399 (N_7399,N_6373,N_6003);
or U7400 (N_7400,N_6696,N_6590);
nand U7401 (N_7401,N_6866,N_6878);
or U7402 (N_7402,N_6527,N_6633);
nand U7403 (N_7403,N_6557,N_6722);
nand U7404 (N_7404,N_6106,N_6457);
or U7405 (N_7405,N_6889,N_6199);
nand U7406 (N_7406,N_6306,N_6449);
nand U7407 (N_7407,N_6494,N_6168);
nand U7408 (N_7408,N_6193,N_6455);
or U7409 (N_7409,N_6831,N_6795);
nor U7410 (N_7410,N_6617,N_6235);
nand U7411 (N_7411,N_6068,N_6321);
nand U7412 (N_7412,N_6782,N_6278);
nor U7413 (N_7413,N_6929,N_6084);
and U7414 (N_7414,N_6401,N_6990);
nor U7415 (N_7415,N_6209,N_6896);
and U7416 (N_7416,N_6079,N_6050);
and U7417 (N_7417,N_6262,N_6715);
or U7418 (N_7418,N_6481,N_6118);
xor U7419 (N_7419,N_6002,N_6009);
and U7420 (N_7420,N_6658,N_6283);
and U7421 (N_7421,N_6536,N_6256);
nand U7422 (N_7422,N_6871,N_6857);
and U7423 (N_7423,N_6452,N_6041);
nor U7424 (N_7424,N_6444,N_6213);
and U7425 (N_7425,N_6067,N_6879);
or U7426 (N_7426,N_6646,N_6969);
nand U7427 (N_7427,N_6467,N_6897);
and U7428 (N_7428,N_6052,N_6110);
nand U7429 (N_7429,N_6089,N_6476);
xor U7430 (N_7430,N_6395,N_6062);
or U7431 (N_7431,N_6568,N_6973);
nor U7432 (N_7432,N_6825,N_6093);
or U7433 (N_7433,N_6017,N_6261);
and U7434 (N_7434,N_6726,N_6875);
or U7435 (N_7435,N_6413,N_6334);
and U7436 (N_7436,N_6211,N_6761);
or U7437 (N_7437,N_6466,N_6027);
and U7438 (N_7438,N_6187,N_6300);
or U7439 (N_7439,N_6647,N_6383);
nor U7440 (N_7440,N_6360,N_6572);
and U7441 (N_7441,N_6828,N_6732);
nor U7442 (N_7442,N_6006,N_6268);
nor U7443 (N_7443,N_6112,N_6566);
nand U7444 (N_7444,N_6730,N_6512);
nor U7445 (N_7445,N_6705,N_6290);
or U7446 (N_7446,N_6991,N_6023);
nor U7447 (N_7447,N_6594,N_6175);
or U7448 (N_7448,N_6621,N_6405);
nor U7449 (N_7449,N_6045,N_6274);
nor U7450 (N_7450,N_6907,N_6810);
or U7451 (N_7451,N_6488,N_6663);
or U7452 (N_7452,N_6392,N_6943);
nand U7453 (N_7453,N_6198,N_6505);
and U7454 (N_7454,N_6374,N_6899);
nor U7455 (N_7455,N_6784,N_6075);
nor U7456 (N_7456,N_6424,N_6530);
nor U7457 (N_7457,N_6774,N_6008);
and U7458 (N_7458,N_6996,N_6548);
nor U7459 (N_7459,N_6504,N_6143);
nand U7460 (N_7460,N_6583,N_6639);
and U7461 (N_7461,N_6221,N_6569);
nand U7462 (N_7462,N_6314,N_6077);
nor U7463 (N_7463,N_6800,N_6666);
nor U7464 (N_7464,N_6515,N_6664);
or U7465 (N_7465,N_6243,N_6192);
nor U7466 (N_7466,N_6315,N_6835);
and U7467 (N_7467,N_6671,N_6406);
and U7468 (N_7468,N_6506,N_6331);
and U7469 (N_7469,N_6464,N_6065);
nor U7470 (N_7470,N_6995,N_6329);
or U7471 (N_7471,N_6301,N_6691);
nor U7472 (N_7472,N_6741,N_6820);
or U7473 (N_7473,N_6733,N_6174);
nand U7474 (N_7474,N_6549,N_6076);
nand U7475 (N_7475,N_6804,N_6534);
nor U7476 (N_7476,N_6802,N_6883);
and U7477 (N_7477,N_6898,N_6132);
nor U7478 (N_7478,N_6743,N_6961);
nand U7479 (N_7479,N_6166,N_6714);
and U7480 (N_7480,N_6064,N_6924);
or U7481 (N_7481,N_6161,N_6634);
and U7482 (N_7482,N_6918,N_6651);
and U7483 (N_7483,N_6322,N_6167);
nor U7484 (N_7484,N_6216,N_6423);
nand U7485 (N_7485,N_6419,N_6238);
nor U7486 (N_7486,N_6745,N_6779);
nand U7487 (N_7487,N_6890,N_6648);
and U7488 (N_7488,N_6239,N_6987);
or U7489 (N_7489,N_6038,N_6226);
nand U7490 (N_7490,N_6141,N_6307);
nand U7491 (N_7491,N_6438,N_6778);
xnor U7492 (N_7492,N_6931,N_6684);
or U7493 (N_7493,N_6258,N_6839);
nor U7494 (N_7494,N_6620,N_6815);
nand U7495 (N_7495,N_6773,N_6445);
nor U7496 (N_7496,N_6993,N_6059);
and U7497 (N_7497,N_6609,N_6427);
and U7498 (N_7498,N_6287,N_6602);
or U7499 (N_7499,N_6862,N_6458);
nand U7500 (N_7500,N_6024,N_6636);
nand U7501 (N_7501,N_6220,N_6419);
nor U7502 (N_7502,N_6608,N_6473);
nand U7503 (N_7503,N_6513,N_6598);
and U7504 (N_7504,N_6210,N_6843);
or U7505 (N_7505,N_6129,N_6489);
and U7506 (N_7506,N_6865,N_6177);
nor U7507 (N_7507,N_6167,N_6261);
and U7508 (N_7508,N_6362,N_6442);
nor U7509 (N_7509,N_6730,N_6822);
nand U7510 (N_7510,N_6556,N_6172);
and U7511 (N_7511,N_6568,N_6196);
nor U7512 (N_7512,N_6588,N_6088);
nor U7513 (N_7513,N_6662,N_6293);
and U7514 (N_7514,N_6190,N_6373);
and U7515 (N_7515,N_6907,N_6422);
or U7516 (N_7516,N_6137,N_6987);
nand U7517 (N_7517,N_6368,N_6706);
nor U7518 (N_7518,N_6679,N_6358);
or U7519 (N_7519,N_6335,N_6676);
or U7520 (N_7520,N_6731,N_6653);
or U7521 (N_7521,N_6789,N_6900);
nor U7522 (N_7522,N_6214,N_6550);
or U7523 (N_7523,N_6278,N_6040);
nand U7524 (N_7524,N_6293,N_6343);
and U7525 (N_7525,N_6390,N_6911);
nor U7526 (N_7526,N_6500,N_6349);
and U7527 (N_7527,N_6102,N_6178);
nand U7528 (N_7528,N_6614,N_6524);
or U7529 (N_7529,N_6417,N_6658);
or U7530 (N_7530,N_6764,N_6960);
or U7531 (N_7531,N_6075,N_6982);
or U7532 (N_7532,N_6750,N_6087);
nand U7533 (N_7533,N_6087,N_6006);
or U7534 (N_7534,N_6783,N_6311);
nor U7535 (N_7535,N_6398,N_6075);
nor U7536 (N_7536,N_6017,N_6829);
nand U7537 (N_7537,N_6163,N_6977);
and U7538 (N_7538,N_6279,N_6545);
nand U7539 (N_7539,N_6866,N_6686);
or U7540 (N_7540,N_6704,N_6526);
and U7541 (N_7541,N_6308,N_6823);
and U7542 (N_7542,N_6071,N_6433);
and U7543 (N_7543,N_6888,N_6926);
nor U7544 (N_7544,N_6178,N_6322);
or U7545 (N_7545,N_6365,N_6572);
nand U7546 (N_7546,N_6050,N_6275);
nor U7547 (N_7547,N_6819,N_6782);
nor U7548 (N_7548,N_6112,N_6774);
or U7549 (N_7549,N_6623,N_6713);
and U7550 (N_7550,N_6374,N_6817);
nor U7551 (N_7551,N_6910,N_6999);
and U7552 (N_7552,N_6770,N_6465);
nand U7553 (N_7553,N_6866,N_6011);
or U7554 (N_7554,N_6034,N_6999);
or U7555 (N_7555,N_6395,N_6397);
nand U7556 (N_7556,N_6855,N_6083);
nand U7557 (N_7557,N_6493,N_6003);
and U7558 (N_7558,N_6699,N_6753);
nor U7559 (N_7559,N_6047,N_6443);
or U7560 (N_7560,N_6568,N_6432);
nor U7561 (N_7561,N_6457,N_6258);
nand U7562 (N_7562,N_6361,N_6403);
and U7563 (N_7563,N_6871,N_6619);
nand U7564 (N_7564,N_6264,N_6873);
and U7565 (N_7565,N_6219,N_6868);
nand U7566 (N_7566,N_6734,N_6056);
and U7567 (N_7567,N_6635,N_6126);
nor U7568 (N_7568,N_6744,N_6149);
nor U7569 (N_7569,N_6157,N_6959);
nand U7570 (N_7570,N_6114,N_6600);
and U7571 (N_7571,N_6307,N_6061);
and U7572 (N_7572,N_6320,N_6825);
or U7573 (N_7573,N_6840,N_6833);
nor U7574 (N_7574,N_6923,N_6661);
and U7575 (N_7575,N_6282,N_6288);
nor U7576 (N_7576,N_6730,N_6664);
nor U7577 (N_7577,N_6395,N_6036);
or U7578 (N_7578,N_6840,N_6116);
or U7579 (N_7579,N_6139,N_6413);
nand U7580 (N_7580,N_6748,N_6411);
and U7581 (N_7581,N_6737,N_6091);
nor U7582 (N_7582,N_6037,N_6469);
nor U7583 (N_7583,N_6801,N_6160);
or U7584 (N_7584,N_6839,N_6438);
or U7585 (N_7585,N_6475,N_6413);
nor U7586 (N_7586,N_6939,N_6212);
nand U7587 (N_7587,N_6742,N_6683);
and U7588 (N_7588,N_6559,N_6800);
or U7589 (N_7589,N_6282,N_6293);
or U7590 (N_7590,N_6481,N_6187);
or U7591 (N_7591,N_6852,N_6893);
or U7592 (N_7592,N_6362,N_6385);
nor U7593 (N_7593,N_6909,N_6577);
and U7594 (N_7594,N_6235,N_6483);
or U7595 (N_7595,N_6376,N_6773);
nor U7596 (N_7596,N_6970,N_6115);
or U7597 (N_7597,N_6305,N_6763);
nor U7598 (N_7598,N_6847,N_6937);
nand U7599 (N_7599,N_6794,N_6498);
or U7600 (N_7600,N_6188,N_6632);
and U7601 (N_7601,N_6911,N_6601);
nor U7602 (N_7602,N_6493,N_6566);
nand U7603 (N_7603,N_6361,N_6593);
nand U7604 (N_7604,N_6408,N_6393);
or U7605 (N_7605,N_6937,N_6055);
and U7606 (N_7606,N_6853,N_6193);
or U7607 (N_7607,N_6997,N_6861);
or U7608 (N_7608,N_6309,N_6821);
nor U7609 (N_7609,N_6624,N_6093);
nand U7610 (N_7610,N_6249,N_6779);
and U7611 (N_7611,N_6122,N_6441);
nand U7612 (N_7612,N_6390,N_6645);
and U7613 (N_7613,N_6793,N_6464);
nand U7614 (N_7614,N_6875,N_6604);
nand U7615 (N_7615,N_6553,N_6026);
and U7616 (N_7616,N_6510,N_6903);
nand U7617 (N_7617,N_6087,N_6396);
or U7618 (N_7618,N_6946,N_6221);
nand U7619 (N_7619,N_6087,N_6434);
or U7620 (N_7620,N_6313,N_6923);
and U7621 (N_7621,N_6242,N_6979);
xor U7622 (N_7622,N_6774,N_6615);
xor U7623 (N_7623,N_6371,N_6059);
nand U7624 (N_7624,N_6188,N_6717);
or U7625 (N_7625,N_6312,N_6077);
nand U7626 (N_7626,N_6373,N_6517);
xnor U7627 (N_7627,N_6494,N_6134);
nor U7628 (N_7628,N_6300,N_6862);
nor U7629 (N_7629,N_6093,N_6966);
or U7630 (N_7630,N_6326,N_6952);
nor U7631 (N_7631,N_6045,N_6059);
and U7632 (N_7632,N_6653,N_6198);
nor U7633 (N_7633,N_6169,N_6883);
or U7634 (N_7634,N_6089,N_6759);
xor U7635 (N_7635,N_6437,N_6014);
nor U7636 (N_7636,N_6823,N_6715);
and U7637 (N_7637,N_6875,N_6118);
nand U7638 (N_7638,N_6003,N_6530);
and U7639 (N_7639,N_6772,N_6774);
and U7640 (N_7640,N_6490,N_6497);
nand U7641 (N_7641,N_6573,N_6665);
or U7642 (N_7642,N_6604,N_6139);
and U7643 (N_7643,N_6574,N_6838);
xnor U7644 (N_7644,N_6527,N_6668);
and U7645 (N_7645,N_6560,N_6158);
nor U7646 (N_7646,N_6099,N_6365);
nand U7647 (N_7647,N_6002,N_6491);
nand U7648 (N_7648,N_6429,N_6948);
nand U7649 (N_7649,N_6867,N_6404);
or U7650 (N_7650,N_6926,N_6717);
nand U7651 (N_7651,N_6183,N_6929);
xor U7652 (N_7652,N_6143,N_6448);
nand U7653 (N_7653,N_6797,N_6806);
nor U7654 (N_7654,N_6844,N_6638);
or U7655 (N_7655,N_6138,N_6580);
xor U7656 (N_7656,N_6020,N_6988);
nand U7657 (N_7657,N_6679,N_6443);
or U7658 (N_7658,N_6365,N_6653);
or U7659 (N_7659,N_6538,N_6789);
nor U7660 (N_7660,N_6982,N_6133);
or U7661 (N_7661,N_6100,N_6207);
nand U7662 (N_7662,N_6405,N_6860);
or U7663 (N_7663,N_6129,N_6289);
or U7664 (N_7664,N_6889,N_6208);
and U7665 (N_7665,N_6814,N_6335);
and U7666 (N_7666,N_6092,N_6493);
or U7667 (N_7667,N_6586,N_6819);
or U7668 (N_7668,N_6513,N_6160);
nand U7669 (N_7669,N_6592,N_6104);
nand U7670 (N_7670,N_6067,N_6616);
nor U7671 (N_7671,N_6153,N_6691);
or U7672 (N_7672,N_6937,N_6340);
nor U7673 (N_7673,N_6480,N_6392);
nor U7674 (N_7674,N_6101,N_6281);
nand U7675 (N_7675,N_6686,N_6569);
nor U7676 (N_7676,N_6976,N_6274);
nand U7677 (N_7677,N_6988,N_6496);
nor U7678 (N_7678,N_6098,N_6499);
or U7679 (N_7679,N_6386,N_6674);
nor U7680 (N_7680,N_6656,N_6083);
and U7681 (N_7681,N_6525,N_6567);
and U7682 (N_7682,N_6910,N_6477);
xor U7683 (N_7683,N_6561,N_6621);
or U7684 (N_7684,N_6820,N_6386);
and U7685 (N_7685,N_6788,N_6082);
nor U7686 (N_7686,N_6087,N_6103);
nor U7687 (N_7687,N_6899,N_6742);
and U7688 (N_7688,N_6037,N_6762);
nand U7689 (N_7689,N_6559,N_6250);
and U7690 (N_7690,N_6626,N_6750);
nor U7691 (N_7691,N_6345,N_6798);
and U7692 (N_7692,N_6859,N_6654);
nor U7693 (N_7693,N_6510,N_6895);
and U7694 (N_7694,N_6572,N_6748);
nor U7695 (N_7695,N_6356,N_6612);
and U7696 (N_7696,N_6855,N_6165);
nor U7697 (N_7697,N_6054,N_6809);
nand U7698 (N_7698,N_6069,N_6806);
nand U7699 (N_7699,N_6549,N_6068);
and U7700 (N_7700,N_6968,N_6864);
and U7701 (N_7701,N_6354,N_6544);
nand U7702 (N_7702,N_6460,N_6307);
nand U7703 (N_7703,N_6863,N_6451);
nand U7704 (N_7704,N_6359,N_6272);
nor U7705 (N_7705,N_6863,N_6083);
xnor U7706 (N_7706,N_6034,N_6822);
or U7707 (N_7707,N_6185,N_6150);
or U7708 (N_7708,N_6833,N_6685);
xnor U7709 (N_7709,N_6863,N_6670);
or U7710 (N_7710,N_6422,N_6281);
nor U7711 (N_7711,N_6754,N_6315);
or U7712 (N_7712,N_6351,N_6036);
nand U7713 (N_7713,N_6070,N_6557);
nor U7714 (N_7714,N_6769,N_6716);
nor U7715 (N_7715,N_6574,N_6651);
nor U7716 (N_7716,N_6786,N_6158);
nor U7717 (N_7717,N_6541,N_6556);
nand U7718 (N_7718,N_6805,N_6643);
nand U7719 (N_7719,N_6810,N_6743);
nand U7720 (N_7720,N_6339,N_6163);
or U7721 (N_7721,N_6046,N_6692);
and U7722 (N_7722,N_6544,N_6240);
nor U7723 (N_7723,N_6698,N_6119);
or U7724 (N_7724,N_6987,N_6303);
and U7725 (N_7725,N_6787,N_6084);
or U7726 (N_7726,N_6886,N_6328);
xnor U7727 (N_7727,N_6886,N_6500);
or U7728 (N_7728,N_6480,N_6953);
nor U7729 (N_7729,N_6669,N_6294);
or U7730 (N_7730,N_6842,N_6415);
nand U7731 (N_7731,N_6367,N_6856);
and U7732 (N_7732,N_6685,N_6840);
nor U7733 (N_7733,N_6050,N_6633);
nand U7734 (N_7734,N_6351,N_6196);
and U7735 (N_7735,N_6252,N_6350);
and U7736 (N_7736,N_6171,N_6225);
and U7737 (N_7737,N_6981,N_6182);
nor U7738 (N_7738,N_6379,N_6145);
nor U7739 (N_7739,N_6147,N_6876);
nor U7740 (N_7740,N_6881,N_6589);
nor U7741 (N_7741,N_6644,N_6169);
and U7742 (N_7742,N_6477,N_6983);
and U7743 (N_7743,N_6724,N_6276);
nor U7744 (N_7744,N_6637,N_6559);
and U7745 (N_7745,N_6173,N_6655);
nand U7746 (N_7746,N_6103,N_6064);
or U7747 (N_7747,N_6058,N_6529);
nand U7748 (N_7748,N_6781,N_6697);
and U7749 (N_7749,N_6036,N_6240);
and U7750 (N_7750,N_6756,N_6200);
or U7751 (N_7751,N_6288,N_6639);
or U7752 (N_7752,N_6976,N_6930);
and U7753 (N_7753,N_6102,N_6427);
nand U7754 (N_7754,N_6365,N_6446);
or U7755 (N_7755,N_6202,N_6710);
nand U7756 (N_7756,N_6621,N_6590);
and U7757 (N_7757,N_6514,N_6748);
nor U7758 (N_7758,N_6441,N_6385);
nand U7759 (N_7759,N_6363,N_6203);
nand U7760 (N_7760,N_6758,N_6963);
nand U7761 (N_7761,N_6868,N_6161);
nand U7762 (N_7762,N_6290,N_6641);
nand U7763 (N_7763,N_6799,N_6972);
nand U7764 (N_7764,N_6109,N_6674);
and U7765 (N_7765,N_6569,N_6678);
or U7766 (N_7766,N_6026,N_6016);
and U7767 (N_7767,N_6730,N_6703);
and U7768 (N_7768,N_6054,N_6490);
nand U7769 (N_7769,N_6439,N_6066);
nand U7770 (N_7770,N_6042,N_6932);
nand U7771 (N_7771,N_6620,N_6275);
nand U7772 (N_7772,N_6135,N_6224);
nor U7773 (N_7773,N_6368,N_6843);
nand U7774 (N_7774,N_6423,N_6281);
and U7775 (N_7775,N_6144,N_6334);
or U7776 (N_7776,N_6711,N_6574);
and U7777 (N_7777,N_6313,N_6721);
nor U7778 (N_7778,N_6263,N_6069);
nand U7779 (N_7779,N_6609,N_6635);
or U7780 (N_7780,N_6089,N_6192);
nand U7781 (N_7781,N_6437,N_6281);
or U7782 (N_7782,N_6390,N_6996);
or U7783 (N_7783,N_6284,N_6134);
and U7784 (N_7784,N_6003,N_6142);
or U7785 (N_7785,N_6037,N_6140);
and U7786 (N_7786,N_6270,N_6589);
nand U7787 (N_7787,N_6068,N_6726);
and U7788 (N_7788,N_6863,N_6882);
nor U7789 (N_7789,N_6317,N_6818);
and U7790 (N_7790,N_6086,N_6369);
nor U7791 (N_7791,N_6687,N_6490);
and U7792 (N_7792,N_6636,N_6966);
or U7793 (N_7793,N_6680,N_6023);
nor U7794 (N_7794,N_6308,N_6466);
nor U7795 (N_7795,N_6220,N_6485);
nand U7796 (N_7796,N_6811,N_6040);
nor U7797 (N_7797,N_6915,N_6110);
and U7798 (N_7798,N_6912,N_6767);
nor U7799 (N_7799,N_6895,N_6579);
or U7800 (N_7800,N_6926,N_6721);
and U7801 (N_7801,N_6346,N_6255);
nor U7802 (N_7802,N_6570,N_6747);
nand U7803 (N_7803,N_6808,N_6733);
nand U7804 (N_7804,N_6178,N_6662);
or U7805 (N_7805,N_6305,N_6146);
and U7806 (N_7806,N_6238,N_6766);
nor U7807 (N_7807,N_6978,N_6068);
nand U7808 (N_7808,N_6891,N_6974);
and U7809 (N_7809,N_6332,N_6987);
or U7810 (N_7810,N_6086,N_6501);
nand U7811 (N_7811,N_6676,N_6072);
and U7812 (N_7812,N_6730,N_6587);
and U7813 (N_7813,N_6321,N_6074);
nand U7814 (N_7814,N_6426,N_6046);
or U7815 (N_7815,N_6810,N_6479);
nor U7816 (N_7816,N_6098,N_6518);
xnor U7817 (N_7817,N_6429,N_6754);
or U7818 (N_7818,N_6881,N_6998);
nor U7819 (N_7819,N_6412,N_6633);
and U7820 (N_7820,N_6803,N_6739);
and U7821 (N_7821,N_6090,N_6267);
and U7822 (N_7822,N_6432,N_6908);
or U7823 (N_7823,N_6069,N_6072);
and U7824 (N_7824,N_6352,N_6019);
nor U7825 (N_7825,N_6569,N_6117);
nand U7826 (N_7826,N_6136,N_6008);
nor U7827 (N_7827,N_6486,N_6866);
or U7828 (N_7828,N_6672,N_6007);
and U7829 (N_7829,N_6068,N_6122);
nor U7830 (N_7830,N_6555,N_6473);
nor U7831 (N_7831,N_6597,N_6925);
nor U7832 (N_7832,N_6731,N_6218);
and U7833 (N_7833,N_6736,N_6734);
or U7834 (N_7834,N_6810,N_6845);
or U7835 (N_7835,N_6925,N_6112);
nor U7836 (N_7836,N_6796,N_6617);
or U7837 (N_7837,N_6302,N_6420);
nor U7838 (N_7838,N_6020,N_6102);
nor U7839 (N_7839,N_6826,N_6498);
nor U7840 (N_7840,N_6843,N_6100);
nor U7841 (N_7841,N_6271,N_6782);
nor U7842 (N_7842,N_6705,N_6339);
or U7843 (N_7843,N_6039,N_6303);
and U7844 (N_7844,N_6741,N_6593);
xnor U7845 (N_7845,N_6138,N_6956);
or U7846 (N_7846,N_6551,N_6888);
nand U7847 (N_7847,N_6734,N_6036);
and U7848 (N_7848,N_6645,N_6566);
nor U7849 (N_7849,N_6597,N_6231);
or U7850 (N_7850,N_6518,N_6778);
nor U7851 (N_7851,N_6087,N_6509);
and U7852 (N_7852,N_6201,N_6678);
xnor U7853 (N_7853,N_6909,N_6413);
nor U7854 (N_7854,N_6502,N_6585);
and U7855 (N_7855,N_6644,N_6633);
and U7856 (N_7856,N_6648,N_6052);
nand U7857 (N_7857,N_6532,N_6427);
and U7858 (N_7858,N_6552,N_6142);
nand U7859 (N_7859,N_6940,N_6467);
or U7860 (N_7860,N_6377,N_6786);
and U7861 (N_7861,N_6007,N_6856);
and U7862 (N_7862,N_6475,N_6006);
and U7863 (N_7863,N_6748,N_6521);
or U7864 (N_7864,N_6373,N_6764);
nor U7865 (N_7865,N_6987,N_6667);
nand U7866 (N_7866,N_6007,N_6753);
nand U7867 (N_7867,N_6472,N_6341);
or U7868 (N_7868,N_6198,N_6530);
or U7869 (N_7869,N_6659,N_6638);
and U7870 (N_7870,N_6456,N_6830);
nor U7871 (N_7871,N_6152,N_6069);
nand U7872 (N_7872,N_6655,N_6545);
nor U7873 (N_7873,N_6821,N_6610);
nand U7874 (N_7874,N_6698,N_6073);
nand U7875 (N_7875,N_6704,N_6817);
nor U7876 (N_7876,N_6405,N_6966);
and U7877 (N_7877,N_6343,N_6354);
nor U7878 (N_7878,N_6718,N_6633);
or U7879 (N_7879,N_6516,N_6023);
and U7880 (N_7880,N_6969,N_6070);
or U7881 (N_7881,N_6981,N_6403);
or U7882 (N_7882,N_6777,N_6047);
nand U7883 (N_7883,N_6886,N_6665);
nor U7884 (N_7884,N_6164,N_6881);
nor U7885 (N_7885,N_6320,N_6123);
nand U7886 (N_7886,N_6938,N_6581);
and U7887 (N_7887,N_6153,N_6880);
nand U7888 (N_7888,N_6193,N_6662);
and U7889 (N_7889,N_6518,N_6951);
nor U7890 (N_7890,N_6352,N_6583);
and U7891 (N_7891,N_6416,N_6686);
nor U7892 (N_7892,N_6495,N_6594);
nor U7893 (N_7893,N_6678,N_6323);
or U7894 (N_7894,N_6638,N_6541);
nand U7895 (N_7895,N_6358,N_6930);
and U7896 (N_7896,N_6373,N_6829);
nor U7897 (N_7897,N_6362,N_6054);
nand U7898 (N_7898,N_6949,N_6978);
nand U7899 (N_7899,N_6866,N_6419);
and U7900 (N_7900,N_6001,N_6756);
nor U7901 (N_7901,N_6244,N_6897);
nor U7902 (N_7902,N_6768,N_6505);
nand U7903 (N_7903,N_6396,N_6061);
nand U7904 (N_7904,N_6707,N_6213);
or U7905 (N_7905,N_6266,N_6597);
and U7906 (N_7906,N_6034,N_6578);
nor U7907 (N_7907,N_6201,N_6188);
nor U7908 (N_7908,N_6743,N_6189);
nand U7909 (N_7909,N_6304,N_6382);
and U7910 (N_7910,N_6131,N_6847);
nand U7911 (N_7911,N_6324,N_6770);
nand U7912 (N_7912,N_6386,N_6257);
nor U7913 (N_7913,N_6951,N_6725);
nor U7914 (N_7914,N_6787,N_6381);
xor U7915 (N_7915,N_6581,N_6810);
nand U7916 (N_7916,N_6187,N_6884);
nand U7917 (N_7917,N_6702,N_6206);
or U7918 (N_7918,N_6780,N_6230);
nand U7919 (N_7919,N_6885,N_6137);
or U7920 (N_7920,N_6090,N_6833);
nand U7921 (N_7921,N_6967,N_6660);
and U7922 (N_7922,N_6223,N_6073);
nor U7923 (N_7923,N_6178,N_6147);
or U7924 (N_7924,N_6293,N_6986);
or U7925 (N_7925,N_6954,N_6754);
nor U7926 (N_7926,N_6644,N_6497);
nor U7927 (N_7927,N_6834,N_6303);
and U7928 (N_7928,N_6637,N_6055);
and U7929 (N_7929,N_6124,N_6495);
or U7930 (N_7930,N_6559,N_6775);
and U7931 (N_7931,N_6712,N_6538);
or U7932 (N_7932,N_6103,N_6664);
nand U7933 (N_7933,N_6971,N_6920);
nor U7934 (N_7934,N_6089,N_6490);
and U7935 (N_7935,N_6282,N_6505);
and U7936 (N_7936,N_6205,N_6201);
or U7937 (N_7937,N_6146,N_6059);
and U7938 (N_7938,N_6288,N_6876);
nor U7939 (N_7939,N_6583,N_6967);
nor U7940 (N_7940,N_6956,N_6397);
nor U7941 (N_7941,N_6566,N_6882);
nand U7942 (N_7942,N_6447,N_6212);
or U7943 (N_7943,N_6289,N_6782);
nor U7944 (N_7944,N_6240,N_6698);
nor U7945 (N_7945,N_6550,N_6769);
or U7946 (N_7946,N_6445,N_6316);
and U7947 (N_7947,N_6278,N_6482);
xnor U7948 (N_7948,N_6749,N_6093);
nand U7949 (N_7949,N_6776,N_6438);
nor U7950 (N_7950,N_6539,N_6206);
nand U7951 (N_7951,N_6307,N_6306);
and U7952 (N_7952,N_6873,N_6802);
and U7953 (N_7953,N_6894,N_6009);
and U7954 (N_7954,N_6284,N_6897);
nor U7955 (N_7955,N_6815,N_6736);
and U7956 (N_7956,N_6909,N_6336);
and U7957 (N_7957,N_6174,N_6675);
or U7958 (N_7958,N_6173,N_6523);
nand U7959 (N_7959,N_6832,N_6790);
and U7960 (N_7960,N_6450,N_6824);
nand U7961 (N_7961,N_6667,N_6165);
and U7962 (N_7962,N_6697,N_6410);
nand U7963 (N_7963,N_6971,N_6735);
nand U7964 (N_7964,N_6560,N_6597);
nor U7965 (N_7965,N_6266,N_6128);
xor U7966 (N_7966,N_6800,N_6538);
or U7967 (N_7967,N_6917,N_6546);
or U7968 (N_7968,N_6318,N_6189);
and U7969 (N_7969,N_6622,N_6097);
nor U7970 (N_7970,N_6508,N_6549);
nand U7971 (N_7971,N_6321,N_6759);
nand U7972 (N_7972,N_6321,N_6803);
or U7973 (N_7973,N_6319,N_6152);
and U7974 (N_7974,N_6541,N_6665);
and U7975 (N_7975,N_6078,N_6672);
and U7976 (N_7976,N_6822,N_6783);
and U7977 (N_7977,N_6055,N_6448);
or U7978 (N_7978,N_6575,N_6198);
nand U7979 (N_7979,N_6446,N_6424);
and U7980 (N_7980,N_6650,N_6302);
or U7981 (N_7981,N_6170,N_6601);
or U7982 (N_7982,N_6506,N_6699);
nor U7983 (N_7983,N_6310,N_6036);
or U7984 (N_7984,N_6409,N_6766);
nand U7985 (N_7985,N_6674,N_6287);
or U7986 (N_7986,N_6378,N_6081);
nor U7987 (N_7987,N_6738,N_6541);
nor U7988 (N_7988,N_6765,N_6014);
or U7989 (N_7989,N_6193,N_6880);
and U7990 (N_7990,N_6154,N_6746);
nor U7991 (N_7991,N_6961,N_6544);
nor U7992 (N_7992,N_6893,N_6588);
nand U7993 (N_7993,N_6347,N_6462);
or U7994 (N_7994,N_6686,N_6296);
and U7995 (N_7995,N_6917,N_6449);
and U7996 (N_7996,N_6875,N_6670);
or U7997 (N_7997,N_6153,N_6100);
nor U7998 (N_7998,N_6417,N_6178);
and U7999 (N_7999,N_6777,N_6994);
nand U8000 (N_8000,N_7813,N_7481);
nand U8001 (N_8001,N_7843,N_7333);
and U8002 (N_8002,N_7307,N_7922);
and U8003 (N_8003,N_7953,N_7687);
nand U8004 (N_8004,N_7088,N_7279);
or U8005 (N_8005,N_7300,N_7766);
nor U8006 (N_8006,N_7486,N_7814);
and U8007 (N_8007,N_7151,N_7564);
or U8008 (N_8008,N_7132,N_7145);
or U8009 (N_8009,N_7835,N_7919);
or U8010 (N_8010,N_7556,N_7160);
and U8011 (N_8011,N_7857,N_7040);
nor U8012 (N_8012,N_7668,N_7441);
nand U8013 (N_8013,N_7029,N_7391);
or U8014 (N_8014,N_7815,N_7508);
nor U8015 (N_8015,N_7005,N_7312);
and U8016 (N_8016,N_7870,N_7460);
nand U8017 (N_8017,N_7008,N_7255);
or U8018 (N_8018,N_7253,N_7742);
nand U8019 (N_8019,N_7317,N_7389);
and U8020 (N_8020,N_7730,N_7530);
and U8021 (N_8021,N_7394,N_7130);
nand U8022 (N_8022,N_7174,N_7167);
nor U8023 (N_8023,N_7139,N_7271);
or U8024 (N_8024,N_7136,N_7940);
and U8025 (N_8025,N_7961,N_7753);
nand U8026 (N_8026,N_7349,N_7304);
or U8027 (N_8027,N_7283,N_7350);
nor U8028 (N_8028,N_7528,N_7869);
or U8029 (N_8029,N_7015,N_7746);
or U8030 (N_8030,N_7229,N_7945);
nand U8031 (N_8031,N_7363,N_7334);
nand U8032 (N_8032,N_7175,N_7625);
and U8033 (N_8033,N_7091,N_7912);
or U8034 (N_8034,N_7242,N_7803);
and U8035 (N_8035,N_7001,N_7704);
nand U8036 (N_8036,N_7303,N_7102);
nor U8037 (N_8037,N_7262,N_7387);
nand U8038 (N_8038,N_7951,N_7685);
or U8039 (N_8039,N_7631,N_7831);
or U8040 (N_8040,N_7010,N_7534);
nor U8041 (N_8041,N_7731,N_7608);
and U8042 (N_8042,N_7182,N_7849);
xor U8043 (N_8043,N_7112,N_7542);
and U8044 (N_8044,N_7234,N_7546);
or U8045 (N_8045,N_7434,N_7957);
or U8046 (N_8046,N_7222,N_7830);
or U8047 (N_8047,N_7764,N_7773);
and U8048 (N_8048,N_7641,N_7189);
or U8049 (N_8049,N_7527,N_7850);
nand U8050 (N_8050,N_7427,N_7258);
nor U8051 (N_8051,N_7886,N_7584);
nand U8052 (N_8052,N_7729,N_7034);
or U8053 (N_8053,N_7287,N_7899);
nor U8054 (N_8054,N_7269,N_7632);
nor U8055 (N_8055,N_7288,N_7038);
nor U8056 (N_8056,N_7747,N_7928);
and U8057 (N_8057,N_7547,N_7696);
or U8058 (N_8058,N_7586,N_7539);
or U8059 (N_8059,N_7430,N_7875);
nand U8060 (N_8060,N_7330,N_7716);
and U8061 (N_8061,N_7737,N_7021);
nor U8062 (N_8062,N_7932,N_7724);
or U8063 (N_8063,N_7738,N_7030);
and U8064 (N_8064,N_7995,N_7698);
xor U8065 (N_8065,N_7491,N_7763);
xnor U8066 (N_8066,N_7471,N_7210);
nor U8067 (N_8067,N_7465,N_7709);
and U8068 (N_8068,N_7461,N_7141);
nand U8069 (N_8069,N_7140,N_7101);
xor U8070 (N_8070,N_7109,N_7103);
nor U8071 (N_8071,N_7971,N_7553);
or U8072 (N_8072,N_7822,N_7464);
and U8073 (N_8073,N_7195,N_7640);
nor U8074 (N_8074,N_7075,N_7301);
or U8075 (N_8075,N_7986,N_7676);
xor U8076 (N_8076,N_7446,N_7201);
or U8077 (N_8077,N_7183,N_7874);
nand U8078 (N_8078,N_7117,N_7212);
or U8079 (N_8079,N_7431,N_7045);
and U8080 (N_8080,N_7209,N_7377);
nor U8081 (N_8081,N_7808,N_7261);
nor U8082 (N_8082,N_7052,N_7126);
or U8083 (N_8083,N_7617,N_7555);
and U8084 (N_8084,N_7416,N_7106);
nand U8085 (N_8085,N_7690,N_7149);
and U8086 (N_8086,N_7423,N_7090);
nand U8087 (N_8087,N_7295,N_7834);
nor U8088 (N_8088,N_7791,N_7326);
and U8089 (N_8089,N_7259,N_7517);
or U8090 (N_8090,N_7779,N_7550);
nand U8091 (N_8091,N_7935,N_7769);
nor U8092 (N_8092,N_7969,N_7384);
and U8093 (N_8093,N_7268,N_7845);
and U8094 (N_8094,N_7807,N_7054);
or U8095 (N_8095,N_7644,N_7913);
nor U8096 (N_8096,N_7891,N_7273);
nand U8097 (N_8097,N_7455,N_7442);
nor U8098 (N_8098,N_7655,N_7392);
nor U8099 (N_8099,N_7329,N_7415);
or U8100 (N_8100,N_7785,N_7852);
nand U8101 (N_8101,N_7395,N_7548);
nand U8102 (N_8102,N_7232,N_7732);
nand U8103 (N_8103,N_7828,N_7171);
nand U8104 (N_8104,N_7068,N_7858);
nor U8105 (N_8105,N_7993,N_7223);
nand U8106 (N_8106,N_7647,N_7179);
and U8107 (N_8107,N_7809,N_7777);
nand U8108 (N_8108,N_7457,N_7633);
xnor U8109 (N_8109,N_7203,N_7514);
nand U8110 (N_8110,N_7572,N_7386);
and U8111 (N_8111,N_7211,N_7235);
or U8112 (N_8112,N_7249,N_7656);
nand U8113 (N_8113,N_7135,N_7256);
nand U8114 (N_8114,N_7445,N_7600);
and U8115 (N_8115,N_7751,N_7247);
or U8116 (N_8116,N_7314,N_7675);
and U8117 (N_8117,N_7208,N_7161);
nor U8118 (N_8118,N_7615,N_7462);
and U8119 (N_8119,N_7535,N_7362);
or U8120 (N_8120,N_7991,N_7405);
and U8121 (N_8121,N_7509,N_7373);
nor U8122 (N_8122,N_7477,N_7400);
nand U8123 (N_8123,N_7162,N_7824);
nand U8124 (N_8124,N_7131,N_7770);
or U8125 (N_8125,N_7467,N_7342);
nor U8126 (N_8126,N_7799,N_7817);
or U8127 (N_8127,N_7097,N_7293);
or U8128 (N_8128,N_7420,N_7152);
or U8129 (N_8129,N_7598,N_7191);
and U8130 (N_8130,N_7516,N_7551);
and U8131 (N_8131,N_7390,N_7049);
nor U8132 (N_8132,N_7421,N_7325);
nor U8133 (N_8133,N_7634,N_7241);
xnor U8134 (N_8134,N_7449,N_7270);
nand U8135 (N_8135,N_7901,N_7336);
xor U8136 (N_8136,N_7958,N_7989);
and U8137 (N_8137,N_7645,N_7868);
or U8138 (N_8138,N_7368,N_7926);
nor U8139 (N_8139,N_7931,N_7627);
nand U8140 (N_8140,N_7257,N_7712);
nand U8141 (N_8141,N_7887,N_7309);
xor U8142 (N_8142,N_7401,N_7412);
nor U8143 (N_8143,N_7865,N_7847);
and U8144 (N_8144,N_7576,N_7890);
nand U8145 (N_8145,N_7708,N_7923);
or U8146 (N_8146,N_7359,N_7695);
and U8147 (N_8147,N_7670,N_7612);
nand U8148 (N_8148,N_7322,N_7299);
or U8149 (N_8149,N_7358,N_7002);
nor U8150 (N_8150,N_7818,N_7012);
nor U8151 (N_8151,N_7009,N_7474);
or U8152 (N_8152,N_7422,N_7673);
nand U8153 (N_8153,N_7419,N_7793);
or U8154 (N_8154,N_7978,N_7851);
nand U8155 (N_8155,N_7559,N_7137);
and U8156 (N_8156,N_7315,N_7050);
and U8157 (N_8157,N_7646,N_7078);
and U8158 (N_8158,N_7485,N_7607);
and U8159 (N_8159,N_7642,N_7761);
and U8160 (N_8160,N_7093,N_7024);
or U8161 (N_8161,N_7177,N_7736);
or U8162 (N_8162,N_7100,N_7072);
and U8163 (N_8163,N_7609,N_7525);
and U8164 (N_8164,N_7988,N_7910);
or U8165 (N_8165,N_7533,N_7678);
nand U8166 (N_8166,N_7251,N_7067);
nor U8167 (N_8167,N_7292,N_7193);
nor U8168 (N_8168,N_7264,N_7487);
nor U8169 (N_8169,N_7278,N_7904);
nand U8170 (N_8170,N_7768,N_7666);
or U8171 (N_8171,N_7410,N_7026);
nand U8172 (N_8172,N_7048,N_7894);
and U8173 (N_8173,N_7425,N_7114);
nand U8174 (N_8174,N_7744,N_7839);
and U8175 (N_8175,N_7066,N_7037);
nor U8176 (N_8176,N_7649,N_7150);
nor U8177 (N_8177,N_7417,N_7157);
nand U8178 (N_8178,N_7372,N_7680);
or U8179 (N_8179,N_7340,N_7291);
nand U8180 (N_8180,N_7702,N_7677);
and U8181 (N_8181,N_7099,N_7409);
nor U8182 (N_8182,N_7328,N_7244);
nand U8183 (N_8183,N_7041,N_7408);
or U8184 (N_8184,N_7490,N_7693);
nand U8185 (N_8185,N_7407,N_7217);
nor U8186 (N_8186,N_7492,N_7611);
or U8187 (N_8187,N_7082,N_7762);
nor U8188 (N_8188,N_7321,N_7780);
and U8189 (N_8189,N_7275,N_7842);
or U8190 (N_8190,N_7374,N_7892);
xor U8191 (N_8191,N_7393,N_7679);
nand U8192 (N_8192,N_7243,N_7519);
nor U8193 (N_8193,N_7713,N_7610);
or U8194 (N_8194,N_7236,N_7087);
nor U8195 (N_8195,N_7118,N_7888);
nor U8196 (N_8196,N_7345,N_7254);
or U8197 (N_8197,N_7844,N_7083);
and U8198 (N_8198,N_7697,N_7838);
and U8199 (N_8199,N_7129,N_7164);
or U8200 (N_8200,N_7233,N_7942);
nand U8201 (N_8201,N_7802,N_7186);
nor U8202 (N_8202,N_7571,N_7263);
nor U8203 (N_8203,N_7638,N_7128);
and U8204 (N_8204,N_7125,N_7765);
and U8205 (N_8205,N_7905,N_7031);
nor U8206 (N_8206,N_7825,N_7659);
nand U8207 (N_8207,N_7365,N_7495);
nand U8208 (N_8208,N_7783,N_7285);
and U8209 (N_8209,N_7418,N_7565);
and U8210 (N_8210,N_7216,N_7781);
nand U8211 (N_8211,N_7863,N_7938);
nand U8212 (N_8212,N_7743,N_7170);
nand U8213 (N_8213,N_7570,N_7884);
nor U8214 (N_8214,N_7504,N_7614);
nor U8215 (N_8215,N_7883,N_7811);
nor U8216 (N_8216,N_7033,N_7383);
nor U8217 (N_8217,N_7604,N_7798);
and U8218 (N_8218,N_7827,N_7250);
and U8219 (N_8219,N_7080,N_7823);
nor U8220 (N_8220,N_7399,N_7671);
nand U8221 (N_8221,N_7515,N_7156);
nand U8222 (N_8222,N_7710,N_7933);
nand U8223 (N_8223,N_7180,N_7380);
nand U8224 (N_8224,N_7804,N_7053);
and U8225 (N_8225,N_7214,N_7451);
or U8226 (N_8226,N_7829,N_7906);
xnor U8227 (N_8227,N_7227,N_7748);
nor U8228 (N_8228,N_7947,N_7726);
and U8229 (N_8229,N_7375,N_7626);
or U8230 (N_8230,N_7366,N_7665);
nand U8231 (N_8231,N_7480,N_7027);
and U8232 (N_8232,N_7206,N_7521);
nor U8233 (N_8233,N_7952,N_7893);
or U8234 (N_8234,N_7601,N_7602);
nand U8235 (N_8235,N_7154,N_7428);
nor U8236 (N_8236,N_7801,N_7028);
or U8237 (N_8237,N_7558,N_7582);
and U8238 (N_8238,N_7511,N_7122);
and U8239 (N_8239,N_7836,N_7281);
xor U8240 (N_8240,N_7364,N_7723);
and U8241 (N_8241,N_7406,N_7057);
and U8242 (N_8242,N_7098,N_7226);
or U8243 (N_8243,N_7651,N_7691);
nand U8244 (N_8244,N_7898,N_7841);
and U8245 (N_8245,N_7296,N_7606);
nor U8246 (N_8246,N_7153,N_7178);
and U8247 (N_8247,N_7854,N_7111);
xnor U8248 (N_8248,N_7867,N_7560);
and U8249 (N_8249,N_7290,N_7660);
nor U8250 (N_8250,N_7715,N_7204);
nand U8251 (N_8251,N_7864,N_7925);
or U8252 (N_8252,N_7541,N_7812);
and U8253 (N_8253,N_7348,N_7569);
nand U8254 (N_8254,N_7820,N_7004);
or U8255 (N_8255,N_7970,N_7603);
and U8256 (N_8256,N_7512,N_7484);
nand U8257 (N_8257,N_7897,N_7661);
and U8258 (N_8258,N_7219,N_7086);
and U8259 (N_8259,N_7774,N_7589);
or U8260 (N_8260,N_7503,N_7563);
nand U8261 (N_8261,N_7518,N_7635);
and U8262 (N_8262,N_7079,N_7058);
or U8263 (N_8263,N_7583,N_7821);
nand U8264 (N_8264,N_7096,N_7414);
nand U8265 (N_8265,N_7084,N_7963);
and U8266 (N_8266,N_7146,N_7192);
nor U8267 (N_8267,N_7018,N_7218);
nor U8268 (N_8268,N_7994,N_7056);
nor U8269 (N_8269,N_7934,N_7444);
nand U8270 (N_8270,N_7949,N_7733);
and U8271 (N_8271,N_7915,N_7432);
nor U8272 (N_8272,N_7168,N_7591);
or U8273 (N_8273,N_7650,N_7866);
or U8274 (N_8274,N_7950,N_7158);
nor U8275 (N_8275,N_7436,N_7784);
nor U8276 (N_8276,N_7960,N_7681);
nor U8277 (N_8277,N_7020,N_7238);
xor U8278 (N_8278,N_7277,N_7155);
or U8279 (N_8279,N_7344,N_7319);
or U8280 (N_8280,N_7187,N_7466);
and U8281 (N_8281,N_7682,N_7159);
nand U8282 (N_8282,N_7311,N_7717);
nor U8283 (N_8283,N_7134,N_7507);
nor U8284 (N_8284,N_7469,N_7795);
and U8285 (N_8285,N_7335,N_7361);
or U8286 (N_8286,N_7260,N_7876);
or U8287 (N_8287,N_7501,N_7061);
nor U8288 (N_8288,N_7976,N_7148);
or U8289 (N_8289,N_7190,N_7590);
or U8290 (N_8290,N_7964,N_7593);
and U8291 (N_8291,N_7699,N_7286);
nor U8292 (N_8292,N_7105,N_7943);
and U8293 (N_8293,N_7794,N_7166);
nand U8294 (N_8294,N_7755,N_7310);
or U8295 (N_8295,N_7683,N_7092);
nor U8296 (N_8296,N_7987,N_7313);
nand U8297 (N_8297,N_7974,N_7488);
or U8298 (N_8298,N_7356,N_7115);
nand U8299 (N_8299,N_7473,N_7044);
and U8300 (N_8300,N_7089,N_7231);
nor U8301 (N_8301,N_7578,N_7554);
nand U8302 (N_8302,N_7998,N_7071);
nand U8303 (N_8303,N_7107,N_7948);
nor U8304 (N_8304,N_7537,N_7388);
and U8305 (N_8305,N_7452,N_7902);
nand U8306 (N_8306,N_7318,N_7557);
xor U8307 (N_8307,N_7619,N_7701);
and U8308 (N_8308,N_7200,N_7714);
and U8309 (N_8309,N_7197,N_7921);
and U8310 (N_8310,N_7623,N_7246);
and U8311 (N_8311,N_7523,N_7536);
and U8312 (N_8312,N_7735,N_7526);
and U8313 (N_8313,N_7298,N_7120);
and U8314 (N_8314,N_7520,N_7032);
or U8315 (N_8315,N_7355,N_7853);
or U8316 (N_8316,N_7489,N_7580);
nor U8317 (N_8317,N_7230,N_7483);
nand U8318 (N_8318,N_7006,N_7767);
or U8319 (N_8319,N_7184,N_7700);
or U8320 (N_8320,N_7352,N_7116);
nor U8321 (N_8321,N_7705,N_7686);
and U8322 (N_8322,N_7694,N_7707);
or U8323 (N_8323,N_7215,N_7848);
and U8324 (N_8324,N_7142,N_7095);
and U8325 (N_8325,N_7720,N_7343);
nand U8326 (N_8326,N_7955,N_7076);
nor U8327 (N_8327,N_7522,N_7585);
nand U8328 (N_8328,N_7438,N_7065);
nand U8329 (N_8329,N_7968,N_7331);
or U8330 (N_8330,N_7003,N_7597);
and U8331 (N_8331,N_7920,N_7917);
and U8332 (N_8332,N_7975,N_7404);
or U8333 (N_8333,N_7346,N_7385);
nand U8334 (N_8334,N_7051,N_7579);
nand U8335 (N_8335,N_7143,N_7475);
nand U8336 (N_8336,N_7378,N_7741);
nor U8337 (N_8337,N_7039,N_7879);
or U8338 (N_8338,N_7792,N_7790);
nand U8339 (N_8339,N_7568,N_7306);
or U8340 (N_8340,N_7429,N_7629);
and U8341 (N_8341,N_7605,N_7983);
nand U8342 (N_8342,N_7104,N_7463);
nor U8343 (N_8343,N_7992,N_7133);
nand U8344 (N_8344,N_7454,N_7500);
nor U8345 (N_8345,N_7936,N_7688);
or U8346 (N_8346,N_7360,N_7188);
and U8347 (N_8347,N_7805,N_7482);
nor U8348 (N_8348,N_7035,N_7630);
or U8349 (N_8349,N_7648,N_7351);
and U8350 (N_8350,N_7787,N_7962);
and U8351 (N_8351,N_7739,N_7138);
or U8352 (N_8352,N_7036,N_7110);
nor U8353 (N_8353,N_7594,N_7213);
nor U8354 (N_8354,N_7435,N_7972);
and U8355 (N_8355,N_7956,N_7581);
nor U8356 (N_8356,N_7433,N_7069);
nand U8357 (N_8357,N_7176,N_7880);
nor U8358 (N_8358,N_7984,N_7398);
nand U8359 (N_8359,N_7144,N_7757);
xnor U8360 (N_8360,N_7081,N_7929);
or U8361 (N_8361,N_7924,N_7458);
or U8362 (N_8362,N_7448,N_7173);
nand U8363 (N_8363,N_7237,N_7621);
nand U8364 (N_8364,N_7728,N_7305);
or U8365 (N_8365,N_7513,N_7930);
and U8366 (N_8366,N_7672,N_7220);
and U8367 (N_8367,N_7810,N_7667);
nand U8368 (N_8368,N_7337,N_7706);
xor U8369 (N_8369,N_7121,N_7914);
or U8370 (N_8370,N_7561,N_7944);
nor U8371 (N_8371,N_7339,N_7245);
nor U8372 (N_8372,N_7725,N_7837);
and U8373 (N_8373,N_7977,N_7085);
nor U8374 (N_8374,N_7252,N_7896);
and U8375 (N_8375,N_7872,N_7443);
nand U8376 (N_8376,N_7575,N_7806);
nand U8377 (N_8377,N_7911,N_7341);
nor U8378 (N_8378,N_7240,N_7900);
or U8379 (N_8379,N_7124,N_7440);
and U8380 (N_8380,N_7022,N_7878);
nor U8381 (N_8381,N_7788,N_7055);
and U8382 (N_8382,N_7982,N_7544);
and U8383 (N_8383,N_7426,N_7996);
nand U8384 (N_8384,N_7367,N_7267);
xnor U8385 (N_8385,N_7711,N_7127);
nand U8386 (N_8386,N_7771,N_7637);
and U8387 (N_8387,N_7224,N_7778);
or U8388 (N_8388,N_7745,N_7577);
or U8389 (N_8389,N_7113,N_7221);
nand U8390 (N_8390,N_7357,N_7596);
nor U8391 (N_8391,N_7265,N_7618);
nor U8392 (N_8392,N_7199,N_7877);
nand U8393 (N_8393,N_7916,N_7013);
nand U8394 (N_8394,N_7980,N_7985);
and U8395 (N_8395,N_7439,N_7754);
nor U8396 (N_8396,N_7692,N_7043);
nand U8397 (N_8397,N_7636,N_7308);
nand U8398 (N_8398,N_7918,N_7562);
nor U8399 (N_8399,N_7062,N_7782);
or U8400 (N_8400,N_7510,N_7000);
nor U8401 (N_8401,N_7652,N_7064);
nand U8402 (N_8402,N_7228,N_7889);
nor U8403 (N_8403,N_7059,N_7468);
and U8404 (N_8404,N_7826,N_7871);
and U8405 (N_8405,N_7276,N_7007);
and U8406 (N_8406,N_7424,N_7639);
and U8407 (N_8407,N_7347,N_7239);
nand U8408 (N_8408,N_7025,N_7587);
and U8409 (N_8409,N_7371,N_7524);
nor U8410 (N_8410,N_7077,N_7496);
nor U8411 (N_8411,N_7840,N_7573);
nor U8412 (N_8412,N_7959,N_7756);
nor U8413 (N_8413,N_7941,N_7538);
nor U8414 (N_8414,N_7734,N_7658);
nand U8415 (N_8415,N_7499,N_7332);
or U8416 (N_8416,N_7786,N_7165);
nor U8417 (N_8417,N_7297,N_7074);
and U8418 (N_8418,N_7776,N_7816);
and U8419 (N_8419,N_7939,N_7272);
and U8420 (N_8420,N_7017,N_7860);
or U8421 (N_8421,N_7532,N_7727);
and U8422 (N_8422,N_7689,N_7722);
nor U8423 (N_8423,N_7397,N_7721);
nor U8424 (N_8424,N_7908,N_7459);
xnor U8425 (N_8425,N_7502,N_7479);
nand U8426 (N_8426,N_7796,N_7967);
nand U8427 (N_8427,N_7882,N_7859);
nor U8428 (N_8428,N_7396,N_7019);
nor U8429 (N_8429,N_7453,N_7966);
and U8430 (N_8430,N_7198,N_7316);
nor U8431 (N_8431,N_7997,N_7750);
nand U8432 (N_8432,N_7354,N_7379);
nand U8433 (N_8433,N_7531,N_7529);
and U8434 (N_8434,N_7494,N_7885);
nand U8435 (N_8435,N_7616,N_7772);
nand U8436 (N_8436,N_7194,N_7284);
nor U8437 (N_8437,N_7046,N_7289);
nand U8438 (N_8438,N_7280,N_7895);
and U8439 (N_8439,N_7505,N_7181);
or U8440 (N_8440,N_7937,N_7657);
xor U8441 (N_8441,N_7643,N_7094);
or U8442 (N_8442,N_7881,N_7909);
nor U8443 (N_8443,N_7664,N_7775);
or U8444 (N_8444,N_7819,N_7447);
or U8445 (N_8445,N_7758,N_7540);
or U8446 (N_8446,N_7476,N_7450);
or U8447 (N_8447,N_7833,N_7370);
or U8448 (N_8448,N_7628,N_7472);
and U8449 (N_8449,N_7123,N_7108);
or U8450 (N_8450,N_7752,N_7990);
and U8451 (N_8451,N_7663,N_7011);
or U8452 (N_8452,N_7413,N_7202);
nor U8453 (N_8453,N_7376,N_7759);
nand U8454 (N_8454,N_7954,N_7493);
nor U8455 (N_8455,N_7060,N_7903);
and U8456 (N_8456,N_7599,N_7327);
and U8457 (N_8457,N_7973,N_7662);
or U8458 (N_8458,N_7381,N_7979);
nand U8459 (N_8459,N_7543,N_7653);
and U8460 (N_8460,N_7574,N_7070);
and U8461 (N_8461,N_7566,N_7965);
or U8462 (N_8462,N_7927,N_7789);
or U8463 (N_8463,N_7620,N_7855);
or U8464 (N_8464,N_7592,N_7169);
nor U8465 (N_8465,N_7382,N_7498);
or U8466 (N_8466,N_7549,N_7402);
nand U8467 (N_8467,N_7172,N_7073);
and U8468 (N_8468,N_7225,N_7613);
nor U8469 (N_8469,N_7274,N_7797);
or U8470 (N_8470,N_7588,N_7014);
nor U8471 (N_8471,N_7196,N_7163);
xor U8472 (N_8472,N_7353,N_7832);
nor U8473 (N_8473,N_7023,N_7567);
nor U8474 (N_8474,N_7185,N_7497);
or U8475 (N_8475,N_7403,N_7946);
or U8476 (N_8476,N_7205,N_7147);
and U8477 (N_8477,N_7622,N_7981);
and U8478 (N_8478,N_7338,N_7478);
nor U8479 (N_8479,N_7800,N_7119);
nor U8480 (N_8480,N_7545,N_7719);
nand U8481 (N_8481,N_7042,N_7624);
nor U8482 (N_8482,N_7016,N_7456);
xnor U8483 (N_8483,N_7862,N_7674);
or U8484 (N_8484,N_7856,N_7302);
nand U8485 (N_8485,N_7740,N_7248);
nor U8486 (N_8486,N_7323,N_7266);
and U8487 (N_8487,N_7282,N_7907);
nor U8488 (N_8488,N_7873,N_7437);
xor U8489 (N_8489,N_7470,N_7669);
nor U8490 (N_8490,N_7749,N_7703);
nor U8491 (N_8491,N_7506,N_7411);
nand U8492 (N_8492,N_7063,N_7718);
nand U8493 (N_8493,N_7654,N_7324);
and U8494 (N_8494,N_7846,N_7320);
and U8495 (N_8495,N_7552,N_7684);
nor U8496 (N_8496,N_7369,N_7047);
nor U8497 (N_8497,N_7595,N_7999);
or U8498 (N_8498,N_7207,N_7294);
nor U8499 (N_8499,N_7861,N_7760);
or U8500 (N_8500,N_7968,N_7612);
nor U8501 (N_8501,N_7965,N_7314);
nor U8502 (N_8502,N_7664,N_7984);
nor U8503 (N_8503,N_7486,N_7557);
nor U8504 (N_8504,N_7928,N_7794);
nor U8505 (N_8505,N_7156,N_7286);
or U8506 (N_8506,N_7306,N_7125);
or U8507 (N_8507,N_7342,N_7326);
and U8508 (N_8508,N_7869,N_7707);
nor U8509 (N_8509,N_7648,N_7939);
or U8510 (N_8510,N_7055,N_7315);
or U8511 (N_8511,N_7228,N_7308);
nor U8512 (N_8512,N_7695,N_7074);
nand U8513 (N_8513,N_7427,N_7421);
and U8514 (N_8514,N_7877,N_7543);
and U8515 (N_8515,N_7558,N_7597);
xor U8516 (N_8516,N_7678,N_7781);
nor U8517 (N_8517,N_7321,N_7474);
nand U8518 (N_8518,N_7591,N_7766);
nor U8519 (N_8519,N_7523,N_7117);
nor U8520 (N_8520,N_7804,N_7894);
and U8521 (N_8521,N_7073,N_7839);
and U8522 (N_8522,N_7907,N_7731);
xnor U8523 (N_8523,N_7048,N_7615);
and U8524 (N_8524,N_7389,N_7777);
or U8525 (N_8525,N_7678,N_7996);
or U8526 (N_8526,N_7799,N_7646);
nand U8527 (N_8527,N_7500,N_7605);
nor U8528 (N_8528,N_7840,N_7534);
or U8529 (N_8529,N_7674,N_7146);
or U8530 (N_8530,N_7292,N_7476);
nor U8531 (N_8531,N_7669,N_7457);
and U8532 (N_8532,N_7245,N_7870);
and U8533 (N_8533,N_7118,N_7341);
nor U8534 (N_8534,N_7432,N_7408);
or U8535 (N_8535,N_7084,N_7613);
nor U8536 (N_8536,N_7152,N_7493);
nor U8537 (N_8537,N_7949,N_7978);
nor U8538 (N_8538,N_7821,N_7555);
nor U8539 (N_8539,N_7415,N_7048);
or U8540 (N_8540,N_7491,N_7258);
nor U8541 (N_8541,N_7145,N_7952);
nand U8542 (N_8542,N_7103,N_7508);
or U8543 (N_8543,N_7492,N_7721);
or U8544 (N_8544,N_7057,N_7288);
and U8545 (N_8545,N_7591,N_7163);
and U8546 (N_8546,N_7785,N_7492);
nor U8547 (N_8547,N_7666,N_7170);
and U8548 (N_8548,N_7752,N_7670);
nand U8549 (N_8549,N_7449,N_7549);
or U8550 (N_8550,N_7813,N_7543);
nand U8551 (N_8551,N_7384,N_7269);
and U8552 (N_8552,N_7003,N_7041);
and U8553 (N_8553,N_7207,N_7747);
nor U8554 (N_8554,N_7740,N_7641);
nand U8555 (N_8555,N_7873,N_7515);
or U8556 (N_8556,N_7334,N_7484);
and U8557 (N_8557,N_7611,N_7445);
and U8558 (N_8558,N_7375,N_7852);
and U8559 (N_8559,N_7318,N_7292);
nand U8560 (N_8560,N_7912,N_7585);
nor U8561 (N_8561,N_7301,N_7196);
or U8562 (N_8562,N_7028,N_7378);
nor U8563 (N_8563,N_7840,N_7505);
or U8564 (N_8564,N_7849,N_7675);
or U8565 (N_8565,N_7508,N_7819);
or U8566 (N_8566,N_7724,N_7026);
or U8567 (N_8567,N_7328,N_7026);
or U8568 (N_8568,N_7687,N_7045);
nand U8569 (N_8569,N_7873,N_7690);
or U8570 (N_8570,N_7972,N_7501);
or U8571 (N_8571,N_7205,N_7042);
nand U8572 (N_8572,N_7877,N_7888);
or U8573 (N_8573,N_7354,N_7693);
and U8574 (N_8574,N_7486,N_7178);
nor U8575 (N_8575,N_7059,N_7352);
or U8576 (N_8576,N_7624,N_7128);
and U8577 (N_8577,N_7442,N_7021);
or U8578 (N_8578,N_7871,N_7413);
or U8579 (N_8579,N_7402,N_7730);
and U8580 (N_8580,N_7363,N_7931);
or U8581 (N_8581,N_7713,N_7604);
or U8582 (N_8582,N_7137,N_7886);
nand U8583 (N_8583,N_7518,N_7197);
and U8584 (N_8584,N_7867,N_7559);
or U8585 (N_8585,N_7290,N_7007);
nand U8586 (N_8586,N_7325,N_7338);
nor U8587 (N_8587,N_7064,N_7494);
nand U8588 (N_8588,N_7461,N_7589);
nand U8589 (N_8589,N_7697,N_7662);
or U8590 (N_8590,N_7041,N_7826);
nor U8591 (N_8591,N_7609,N_7941);
or U8592 (N_8592,N_7267,N_7653);
and U8593 (N_8593,N_7522,N_7723);
or U8594 (N_8594,N_7383,N_7173);
nand U8595 (N_8595,N_7595,N_7908);
or U8596 (N_8596,N_7592,N_7116);
or U8597 (N_8597,N_7217,N_7173);
or U8598 (N_8598,N_7272,N_7952);
and U8599 (N_8599,N_7667,N_7710);
nor U8600 (N_8600,N_7965,N_7044);
nor U8601 (N_8601,N_7066,N_7710);
nor U8602 (N_8602,N_7998,N_7103);
or U8603 (N_8603,N_7547,N_7312);
or U8604 (N_8604,N_7026,N_7584);
nand U8605 (N_8605,N_7879,N_7835);
or U8606 (N_8606,N_7689,N_7178);
nor U8607 (N_8607,N_7273,N_7540);
xor U8608 (N_8608,N_7739,N_7600);
nor U8609 (N_8609,N_7566,N_7153);
nand U8610 (N_8610,N_7244,N_7432);
nand U8611 (N_8611,N_7066,N_7911);
and U8612 (N_8612,N_7575,N_7926);
nand U8613 (N_8613,N_7012,N_7550);
or U8614 (N_8614,N_7596,N_7898);
nor U8615 (N_8615,N_7771,N_7550);
nor U8616 (N_8616,N_7165,N_7715);
or U8617 (N_8617,N_7766,N_7812);
and U8618 (N_8618,N_7813,N_7513);
nand U8619 (N_8619,N_7936,N_7663);
nand U8620 (N_8620,N_7131,N_7024);
nand U8621 (N_8621,N_7428,N_7512);
or U8622 (N_8622,N_7429,N_7402);
nor U8623 (N_8623,N_7094,N_7076);
nand U8624 (N_8624,N_7033,N_7035);
nor U8625 (N_8625,N_7041,N_7090);
nand U8626 (N_8626,N_7238,N_7920);
nor U8627 (N_8627,N_7126,N_7368);
nand U8628 (N_8628,N_7612,N_7131);
nor U8629 (N_8629,N_7764,N_7122);
or U8630 (N_8630,N_7014,N_7542);
and U8631 (N_8631,N_7183,N_7205);
or U8632 (N_8632,N_7736,N_7597);
and U8633 (N_8633,N_7263,N_7092);
nand U8634 (N_8634,N_7681,N_7627);
nand U8635 (N_8635,N_7652,N_7344);
nand U8636 (N_8636,N_7883,N_7768);
and U8637 (N_8637,N_7025,N_7367);
or U8638 (N_8638,N_7791,N_7184);
nand U8639 (N_8639,N_7195,N_7608);
or U8640 (N_8640,N_7304,N_7983);
and U8641 (N_8641,N_7298,N_7474);
nor U8642 (N_8642,N_7160,N_7416);
nand U8643 (N_8643,N_7059,N_7573);
nand U8644 (N_8644,N_7877,N_7890);
nor U8645 (N_8645,N_7770,N_7672);
nor U8646 (N_8646,N_7139,N_7697);
and U8647 (N_8647,N_7603,N_7046);
nand U8648 (N_8648,N_7821,N_7744);
and U8649 (N_8649,N_7567,N_7579);
and U8650 (N_8650,N_7039,N_7504);
nor U8651 (N_8651,N_7834,N_7276);
and U8652 (N_8652,N_7286,N_7324);
nor U8653 (N_8653,N_7333,N_7121);
nor U8654 (N_8654,N_7200,N_7381);
nor U8655 (N_8655,N_7045,N_7030);
and U8656 (N_8656,N_7258,N_7972);
and U8657 (N_8657,N_7822,N_7876);
nand U8658 (N_8658,N_7749,N_7351);
and U8659 (N_8659,N_7845,N_7680);
and U8660 (N_8660,N_7856,N_7596);
xnor U8661 (N_8661,N_7223,N_7192);
nand U8662 (N_8662,N_7437,N_7872);
nor U8663 (N_8663,N_7817,N_7730);
and U8664 (N_8664,N_7843,N_7063);
or U8665 (N_8665,N_7144,N_7950);
and U8666 (N_8666,N_7851,N_7839);
nand U8667 (N_8667,N_7354,N_7845);
or U8668 (N_8668,N_7500,N_7876);
and U8669 (N_8669,N_7304,N_7002);
or U8670 (N_8670,N_7710,N_7513);
nand U8671 (N_8671,N_7618,N_7799);
nand U8672 (N_8672,N_7346,N_7662);
nand U8673 (N_8673,N_7161,N_7322);
or U8674 (N_8674,N_7322,N_7160);
and U8675 (N_8675,N_7507,N_7916);
nand U8676 (N_8676,N_7059,N_7053);
nand U8677 (N_8677,N_7084,N_7725);
nor U8678 (N_8678,N_7683,N_7378);
or U8679 (N_8679,N_7908,N_7609);
nand U8680 (N_8680,N_7948,N_7567);
nor U8681 (N_8681,N_7346,N_7113);
and U8682 (N_8682,N_7579,N_7936);
nor U8683 (N_8683,N_7465,N_7735);
nand U8684 (N_8684,N_7253,N_7567);
or U8685 (N_8685,N_7769,N_7558);
nand U8686 (N_8686,N_7789,N_7497);
or U8687 (N_8687,N_7168,N_7682);
nand U8688 (N_8688,N_7401,N_7873);
nand U8689 (N_8689,N_7734,N_7945);
or U8690 (N_8690,N_7564,N_7137);
nand U8691 (N_8691,N_7515,N_7475);
or U8692 (N_8692,N_7675,N_7137);
and U8693 (N_8693,N_7575,N_7525);
nor U8694 (N_8694,N_7656,N_7694);
nand U8695 (N_8695,N_7024,N_7550);
nor U8696 (N_8696,N_7648,N_7975);
and U8697 (N_8697,N_7640,N_7842);
nand U8698 (N_8698,N_7536,N_7922);
or U8699 (N_8699,N_7519,N_7607);
nor U8700 (N_8700,N_7375,N_7337);
or U8701 (N_8701,N_7720,N_7303);
nor U8702 (N_8702,N_7462,N_7487);
or U8703 (N_8703,N_7276,N_7577);
and U8704 (N_8704,N_7961,N_7815);
nor U8705 (N_8705,N_7214,N_7330);
and U8706 (N_8706,N_7106,N_7438);
nand U8707 (N_8707,N_7690,N_7657);
nand U8708 (N_8708,N_7359,N_7691);
nand U8709 (N_8709,N_7565,N_7262);
nand U8710 (N_8710,N_7967,N_7382);
nand U8711 (N_8711,N_7350,N_7255);
nand U8712 (N_8712,N_7661,N_7701);
and U8713 (N_8713,N_7594,N_7010);
nand U8714 (N_8714,N_7995,N_7186);
or U8715 (N_8715,N_7396,N_7917);
nand U8716 (N_8716,N_7859,N_7159);
nand U8717 (N_8717,N_7462,N_7054);
and U8718 (N_8718,N_7286,N_7770);
and U8719 (N_8719,N_7699,N_7599);
nor U8720 (N_8720,N_7091,N_7829);
nand U8721 (N_8721,N_7242,N_7963);
and U8722 (N_8722,N_7777,N_7586);
or U8723 (N_8723,N_7905,N_7352);
and U8724 (N_8724,N_7994,N_7941);
nand U8725 (N_8725,N_7540,N_7205);
nor U8726 (N_8726,N_7857,N_7771);
nor U8727 (N_8727,N_7776,N_7401);
or U8728 (N_8728,N_7171,N_7422);
nor U8729 (N_8729,N_7032,N_7210);
and U8730 (N_8730,N_7016,N_7265);
and U8731 (N_8731,N_7984,N_7392);
and U8732 (N_8732,N_7779,N_7610);
and U8733 (N_8733,N_7678,N_7072);
nand U8734 (N_8734,N_7315,N_7094);
nand U8735 (N_8735,N_7438,N_7484);
nand U8736 (N_8736,N_7603,N_7786);
or U8737 (N_8737,N_7551,N_7752);
nand U8738 (N_8738,N_7191,N_7541);
or U8739 (N_8739,N_7735,N_7323);
xnor U8740 (N_8740,N_7703,N_7913);
nor U8741 (N_8741,N_7392,N_7150);
and U8742 (N_8742,N_7349,N_7852);
xor U8743 (N_8743,N_7157,N_7617);
or U8744 (N_8744,N_7286,N_7924);
or U8745 (N_8745,N_7670,N_7807);
nor U8746 (N_8746,N_7917,N_7990);
nand U8747 (N_8747,N_7585,N_7876);
nand U8748 (N_8748,N_7075,N_7282);
nor U8749 (N_8749,N_7200,N_7464);
and U8750 (N_8750,N_7963,N_7687);
nand U8751 (N_8751,N_7801,N_7985);
and U8752 (N_8752,N_7161,N_7987);
or U8753 (N_8753,N_7494,N_7531);
and U8754 (N_8754,N_7829,N_7017);
or U8755 (N_8755,N_7524,N_7386);
nand U8756 (N_8756,N_7496,N_7699);
and U8757 (N_8757,N_7979,N_7287);
and U8758 (N_8758,N_7235,N_7187);
or U8759 (N_8759,N_7437,N_7854);
nor U8760 (N_8760,N_7063,N_7611);
and U8761 (N_8761,N_7670,N_7620);
and U8762 (N_8762,N_7945,N_7510);
and U8763 (N_8763,N_7036,N_7740);
and U8764 (N_8764,N_7042,N_7509);
nand U8765 (N_8765,N_7015,N_7393);
nand U8766 (N_8766,N_7464,N_7821);
or U8767 (N_8767,N_7149,N_7372);
nand U8768 (N_8768,N_7620,N_7268);
nor U8769 (N_8769,N_7059,N_7072);
nor U8770 (N_8770,N_7715,N_7249);
and U8771 (N_8771,N_7210,N_7653);
nand U8772 (N_8772,N_7985,N_7616);
and U8773 (N_8773,N_7928,N_7945);
and U8774 (N_8774,N_7387,N_7482);
nand U8775 (N_8775,N_7700,N_7477);
nor U8776 (N_8776,N_7908,N_7091);
nor U8777 (N_8777,N_7173,N_7295);
nor U8778 (N_8778,N_7898,N_7991);
nor U8779 (N_8779,N_7839,N_7471);
or U8780 (N_8780,N_7273,N_7872);
nand U8781 (N_8781,N_7363,N_7856);
nor U8782 (N_8782,N_7586,N_7626);
or U8783 (N_8783,N_7632,N_7085);
nand U8784 (N_8784,N_7099,N_7613);
nand U8785 (N_8785,N_7834,N_7166);
or U8786 (N_8786,N_7844,N_7816);
or U8787 (N_8787,N_7295,N_7849);
nor U8788 (N_8788,N_7931,N_7011);
nor U8789 (N_8789,N_7445,N_7290);
nor U8790 (N_8790,N_7453,N_7094);
xor U8791 (N_8791,N_7631,N_7483);
or U8792 (N_8792,N_7116,N_7058);
nand U8793 (N_8793,N_7691,N_7988);
nor U8794 (N_8794,N_7608,N_7185);
and U8795 (N_8795,N_7768,N_7164);
nand U8796 (N_8796,N_7647,N_7305);
nor U8797 (N_8797,N_7906,N_7208);
xnor U8798 (N_8798,N_7958,N_7590);
nor U8799 (N_8799,N_7134,N_7761);
or U8800 (N_8800,N_7540,N_7406);
and U8801 (N_8801,N_7163,N_7602);
and U8802 (N_8802,N_7092,N_7757);
and U8803 (N_8803,N_7476,N_7168);
or U8804 (N_8804,N_7259,N_7503);
nor U8805 (N_8805,N_7294,N_7409);
and U8806 (N_8806,N_7207,N_7350);
nand U8807 (N_8807,N_7588,N_7840);
and U8808 (N_8808,N_7753,N_7727);
and U8809 (N_8809,N_7480,N_7781);
nor U8810 (N_8810,N_7207,N_7455);
nand U8811 (N_8811,N_7354,N_7411);
and U8812 (N_8812,N_7232,N_7498);
nor U8813 (N_8813,N_7180,N_7955);
nor U8814 (N_8814,N_7355,N_7745);
xor U8815 (N_8815,N_7313,N_7598);
xnor U8816 (N_8816,N_7184,N_7857);
nor U8817 (N_8817,N_7881,N_7190);
nor U8818 (N_8818,N_7248,N_7273);
and U8819 (N_8819,N_7652,N_7620);
and U8820 (N_8820,N_7620,N_7683);
and U8821 (N_8821,N_7235,N_7693);
xor U8822 (N_8822,N_7765,N_7722);
nor U8823 (N_8823,N_7367,N_7487);
nand U8824 (N_8824,N_7525,N_7186);
and U8825 (N_8825,N_7150,N_7317);
nor U8826 (N_8826,N_7119,N_7453);
or U8827 (N_8827,N_7469,N_7929);
and U8828 (N_8828,N_7178,N_7390);
nor U8829 (N_8829,N_7974,N_7299);
or U8830 (N_8830,N_7507,N_7891);
nor U8831 (N_8831,N_7457,N_7250);
or U8832 (N_8832,N_7352,N_7584);
or U8833 (N_8833,N_7276,N_7436);
nor U8834 (N_8834,N_7363,N_7524);
nand U8835 (N_8835,N_7886,N_7031);
and U8836 (N_8836,N_7222,N_7223);
nor U8837 (N_8837,N_7918,N_7579);
xor U8838 (N_8838,N_7412,N_7549);
and U8839 (N_8839,N_7320,N_7592);
nand U8840 (N_8840,N_7872,N_7494);
nand U8841 (N_8841,N_7540,N_7341);
and U8842 (N_8842,N_7618,N_7769);
or U8843 (N_8843,N_7320,N_7754);
nor U8844 (N_8844,N_7574,N_7408);
nor U8845 (N_8845,N_7976,N_7510);
nand U8846 (N_8846,N_7513,N_7236);
and U8847 (N_8847,N_7514,N_7346);
and U8848 (N_8848,N_7679,N_7610);
or U8849 (N_8849,N_7449,N_7604);
nand U8850 (N_8850,N_7084,N_7352);
nor U8851 (N_8851,N_7780,N_7844);
or U8852 (N_8852,N_7444,N_7345);
xor U8853 (N_8853,N_7948,N_7851);
or U8854 (N_8854,N_7622,N_7575);
and U8855 (N_8855,N_7557,N_7094);
nand U8856 (N_8856,N_7284,N_7822);
nor U8857 (N_8857,N_7837,N_7947);
and U8858 (N_8858,N_7506,N_7094);
nand U8859 (N_8859,N_7192,N_7134);
and U8860 (N_8860,N_7526,N_7728);
nor U8861 (N_8861,N_7874,N_7788);
and U8862 (N_8862,N_7467,N_7563);
or U8863 (N_8863,N_7776,N_7325);
or U8864 (N_8864,N_7381,N_7893);
nor U8865 (N_8865,N_7570,N_7178);
nor U8866 (N_8866,N_7480,N_7617);
nand U8867 (N_8867,N_7466,N_7141);
and U8868 (N_8868,N_7537,N_7357);
or U8869 (N_8869,N_7284,N_7300);
nor U8870 (N_8870,N_7213,N_7210);
nor U8871 (N_8871,N_7435,N_7185);
and U8872 (N_8872,N_7458,N_7221);
nand U8873 (N_8873,N_7947,N_7154);
and U8874 (N_8874,N_7959,N_7679);
nand U8875 (N_8875,N_7662,N_7153);
and U8876 (N_8876,N_7889,N_7359);
or U8877 (N_8877,N_7115,N_7768);
nand U8878 (N_8878,N_7975,N_7270);
nand U8879 (N_8879,N_7723,N_7246);
or U8880 (N_8880,N_7175,N_7474);
nand U8881 (N_8881,N_7538,N_7638);
or U8882 (N_8882,N_7854,N_7395);
or U8883 (N_8883,N_7209,N_7875);
nor U8884 (N_8884,N_7105,N_7122);
nand U8885 (N_8885,N_7389,N_7028);
nand U8886 (N_8886,N_7864,N_7363);
nor U8887 (N_8887,N_7475,N_7114);
nand U8888 (N_8888,N_7510,N_7591);
and U8889 (N_8889,N_7328,N_7271);
and U8890 (N_8890,N_7723,N_7026);
or U8891 (N_8891,N_7884,N_7508);
nand U8892 (N_8892,N_7294,N_7304);
nor U8893 (N_8893,N_7867,N_7554);
nand U8894 (N_8894,N_7923,N_7333);
nor U8895 (N_8895,N_7485,N_7288);
nor U8896 (N_8896,N_7596,N_7437);
nor U8897 (N_8897,N_7264,N_7500);
nand U8898 (N_8898,N_7814,N_7947);
nor U8899 (N_8899,N_7750,N_7763);
nor U8900 (N_8900,N_7836,N_7524);
nand U8901 (N_8901,N_7709,N_7613);
or U8902 (N_8902,N_7782,N_7010);
or U8903 (N_8903,N_7317,N_7041);
and U8904 (N_8904,N_7757,N_7163);
nor U8905 (N_8905,N_7101,N_7750);
and U8906 (N_8906,N_7456,N_7378);
and U8907 (N_8907,N_7945,N_7754);
or U8908 (N_8908,N_7961,N_7609);
nor U8909 (N_8909,N_7102,N_7050);
nand U8910 (N_8910,N_7198,N_7510);
or U8911 (N_8911,N_7004,N_7735);
nor U8912 (N_8912,N_7612,N_7643);
nor U8913 (N_8913,N_7267,N_7216);
nand U8914 (N_8914,N_7141,N_7131);
nand U8915 (N_8915,N_7442,N_7692);
and U8916 (N_8916,N_7600,N_7166);
nor U8917 (N_8917,N_7491,N_7292);
or U8918 (N_8918,N_7618,N_7123);
nor U8919 (N_8919,N_7225,N_7957);
or U8920 (N_8920,N_7882,N_7571);
or U8921 (N_8921,N_7018,N_7013);
nor U8922 (N_8922,N_7525,N_7000);
or U8923 (N_8923,N_7366,N_7157);
nor U8924 (N_8924,N_7079,N_7216);
and U8925 (N_8925,N_7393,N_7404);
nand U8926 (N_8926,N_7401,N_7949);
nor U8927 (N_8927,N_7607,N_7880);
nand U8928 (N_8928,N_7213,N_7450);
or U8929 (N_8929,N_7531,N_7258);
nor U8930 (N_8930,N_7962,N_7699);
or U8931 (N_8931,N_7542,N_7879);
or U8932 (N_8932,N_7561,N_7392);
nor U8933 (N_8933,N_7449,N_7445);
and U8934 (N_8934,N_7725,N_7627);
or U8935 (N_8935,N_7331,N_7198);
or U8936 (N_8936,N_7700,N_7284);
nand U8937 (N_8937,N_7944,N_7522);
or U8938 (N_8938,N_7122,N_7049);
and U8939 (N_8939,N_7465,N_7647);
or U8940 (N_8940,N_7837,N_7473);
nor U8941 (N_8941,N_7347,N_7893);
nor U8942 (N_8942,N_7594,N_7031);
nor U8943 (N_8943,N_7749,N_7456);
or U8944 (N_8944,N_7454,N_7347);
and U8945 (N_8945,N_7812,N_7923);
or U8946 (N_8946,N_7025,N_7803);
and U8947 (N_8947,N_7217,N_7465);
nand U8948 (N_8948,N_7299,N_7339);
nand U8949 (N_8949,N_7050,N_7476);
or U8950 (N_8950,N_7305,N_7800);
nor U8951 (N_8951,N_7917,N_7965);
xor U8952 (N_8952,N_7000,N_7793);
or U8953 (N_8953,N_7895,N_7730);
and U8954 (N_8954,N_7246,N_7552);
and U8955 (N_8955,N_7021,N_7450);
nor U8956 (N_8956,N_7941,N_7351);
nor U8957 (N_8957,N_7337,N_7960);
and U8958 (N_8958,N_7289,N_7218);
and U8959 (N_8959,N_7769,N_7180);
nor U8960 (N_8960,N_7492,N_7679);
nor U8961 (N_8961,N_7557,N_7632);
xor U8962 (N_8962,N_7742,N_7633);
or U8963 (N_8963,N_7358,N_7459);
nor U8964 (N_8964,N_7800,N_7071);
nor U8965 (N_8965,N_7774,N_7491);
nand U8966 (N_8966,N_7120,N_7673);
nor U8967 (N_8967,N_7082,N_7447);
and U8968 (N_8968,N_7759,N_7457);
nor U8969 (N_8969,N_7888,N_7408);
xor U8970 (N_8970,N_7489,N_7789);
or U8971 (N_8971,N_7889,N_7465);
nand U8972 (N_8972,N_7676,N_7435);
or U8973 (N_8973,N_7027,N_7061);
and U8974 (N_8974,N_7857,N_7757);
nand U8975 (N_8975,N_7857,N_7059);
nand U8976 (N_8976,N_7170,N_7222);
or U8977 (N_8977,N_7545,N_7322);
nand U8978 (N_8978,N_7246,N_7841);
nand U8979 (N_8979,N_7092,N_7588);
nor U8980 (N_8980,N_7417,N_7690);
or U8981 (N_8981,N_7074,N_7654);
nand U8982 (N_8982,N_7024,N_7470);
or U8983 (N_8983,N_7989,N_7427);
or U8984 (N_8984,N_7015,N_7675);
or U8985 (N_8985,N_7102,N_7169);
and U8986 (N_8986,N_7590,N_7359);
or U8987 (N_8987,N_7759,N_7196);
nor U8988 (N_8988,N_7299,N_7961);
nand U8989 (N_8989,N_7125,N_7819);
nand U8990 (N_8990,N_7693,N_7142);
and U8991 (N_8991,N_7348,N_7021);
or U8992 (N_8992,N_7693,N_7968);
or U8993 (N_8993,N_7105,N_7545);
and U8994 (N_8994,N_7424,N_7708);
nor U8995 (N_8995,N_7495,N_7704);
xnor U8996 (N_8996,N_7870,N_7518);
xnor U8997 (N_8997,N_7880,N_7267);
and U8998 (N_8998,N_7360,N_7023);
nor U8999 (N_8999,N_7233,N_7144);
and U9000 (N_9000,N_8616,N_8299);
nand U9001 (N_9001,N_8589,N_8413);
or U9002 (N_9002,N_8747,N_8549);
nand U9003 (N_9003,N_8551,N_8343);
or U9004 (N_9004,N_8916,N_8587);
and U9005 (N_9005,N_8316,N_8466);
nand U9006 (N_9006,N_8910,N_8679);
nor U9007 (N_9007,N_8186,N_8775);
and U9008 (N_9008,N_8215,N_8245);
nand U9009 (N_9009,N_8352,N_8820);
nand U9010 (N_9010,N_8975,N_8986);
nand U9011 (N_9011,N_8298,N_8686);
or U9012 (N_9012,N_8485,N_8395);
or U9013 (N_9013,N_8458,N_8711);
nor U9014 (N_9014,N_8491,N_8596);
or U9015 (N_9015,N_8782,N_8535);
nor U9016 (N_9016,N_8946,N_8571);
xor U9017 (N_9017,N_8236,N_8635);
and U9018 (N_9018,N_8366,N_8423);
or U9019 (N_9019,N_8618,N_8005);
and U9020 (N_9020,N_8893,N_8852);
nor U9021 (N_9021,N_8225,N_8894);
and U9022 (N_9022,N_8147,N_8454);
and U9023 (N_9023,N_8895,N_8884);
nor U9024 (N_9024,N_8375,N_8054);
nand U9025 (N_9025,N_8151,N_8414);
or U9026 (N_9026,N_8733,N_8603);
nor U9027 (N_9027,N_8218,N_8953);
and U9028 (N_9028,N_8987,N_8611);
nand U9029 (N_9029,N_8036,N_8842);
or U9030 (N_9030,N_8488,N_8398);
or U9031 (N_9031,N_8950,N_8079);
nand U9032 (N_9032,N_8082,N_8256);
or U9033 (N_9033,N_8633,N_8802);
nor U9034 (N_9034,N_8695,N_8780);
and U9035 (N_9035,N_8273,N_8154);
nand U9036 (N_9036,N_8709,N_8443);
and U9037 (N_9037,N_8383,N_8740);
nand U9038 (N_9038,N_8873,N_8922);
and U9039 (N_9039,N_8905,N_8216);
nand U9040 (N_9040,N_8815,N_8113);
nor U9041 (N_9041,N_8762,N_8008);
nor U9042 (N_9042,N_8965,N_8866);
nand U9043 (N_9043,N_8687,N_8801);
nand U9044 (N_9044,N_8087,N_8704);
nand U9045 (N_9045,N_8201,N_8029);
and U9046 (N_9046,N_8561,N_8532);
nand U9047 (N_9047,N_8536,N_8149);
or U9048 (N_9048,N_8558,N_8967);
nand U9049 (N_9049,N_8097,N_8858);
or U9050 (N_9050,N_8572,N_8930);
or U9051 (N_9051,N_8690,N_8527);
nor U9052 (N_9052,N_8867,N_8503);
or U9053 (N_9053,N_8988,N_8684);
or U9054 (N_9054,N_8031,N_8470);
and U9055 (N_9055,N_8850,N_8391);
nand U9056 (N_9056,N_8416,N_8301);
nor U9057 (N_9057,N_8244,N_8026);
or U9058 (N_9058,N_8058,N_8311);
nor U9059 (N_9059,N_8292,N_8737);
nor U9060 (N_9060,N_8289,N_8754);
or U9061 (N_9061,N_8796,N_8533);
nor U9062 (N_9062,N_8806,N_8593);
nand U9063 (N_9063,N_8789,N_8662);
nand U9064 (N_9064,N_8957,N_8075);
nor U9065 (N_9065,N_8497,N_8411);
xnor U9066 (N_9066,N_8260,N_8857);
nor U9067 (N_9067,N_8328,N_8592);
and U9068 (N_9068,N_8211,N_8584);
xor U9069 (N_9069,N_8230,N_8804);
and U9070 (N_9070,N_8148,N_8076);
nor U9071 (N_9071,N_8390,N_8727);
and U9072 (N_9072,N_8247,N_8233);
or U9073 (N_9073,N_8351,N_8604);
and U9074 (N_9074,N_8983,N_8537);
nor U9075 (N_9075,N_8045,N_8656);
nor U9076 (N_9076,N_8899,N_8904);
or U9077 (N_9077,N_8146,N_8280);
nand U9078 (N_9078,N_8315,N_8102);
nor U9079 (N_9079,N_8481,N_8406);
nor U9080 (N_9080,N_8544,N_8548);
nor U9081 (N_9081,N_8430,N_8150);
nor U9082 (N_9082,N_8312,N_8510);
and U9083 (N_9083,N_8600,N_8321);
and U9084 (N_9084,N_8823,N_8606);
nor U9085 (N_9085,N_8732,N_8438);
and U9086 (N_9086,N_8122,N_8407);
nor U9087 (N_9087,N_8977,N_8250);
or U9088 (N_9088,N_8277,N_8614);
nand U9089 (N_9089,N_8174,N_8234);
or U9090 (N_9090,N_8098,N_8972);
nor U9091 (N_9091,N_8799,N_8169);
or U9092 (N_9092,N_8581,N_8420);
or U9093 (N_9093,N_8748,N_8719);
or U9094 (N_9094,N_8519,N_8278);
and U9095 (N_9095,N_8943,N_8396);
nor U9096 (N_9096,N_8582,N_8750);
nand U9097 (N_9097,N_8124,N_8263);
or U9098 (N_9098,N_8018,N_8118);
or U9099 (N_9099,N_8106,N_8619);
nand U9100 (N_9100,N_8394,N_8402);
nand U9101 (N_9101,N_8172,N_8261);
or U9102 (N_9102,N_8157,N_8735);
and U9103 (N_9103,N_8586,N_8878);
and U9104 (N_9104,N_8089,N_8410);
or U9105 (N_9105,N_8528,N_8376);
nand U9106 (N_9106,N_8545,N_8185);
or U9107 (N_9107,N_8210,N_8104);
xor U9108 (N_9108,N_8502,N_8770);
nand U9109 (N_9109,N_8346,N_8962);
nor U9110 (N_9110,N_8012,N_8513);
and U9111 (N_9111,N_8196,N_8999);
nand U9112 (N_9112,N_8574,N_8274);
nor U9113 (N_9113,N_8083,N_8693);
or U9114 (N_9114,N_8968,N_8412);
and U9115 (N_9115,N_8178,N_8550);
nand U9116 (N_9116,N_8359,N_8035);
and U9117 (N_9117,N_8307,N_8966);
xnor U9118 (N_9118,N_8153,N_8064);
nand U9119 (N_9119,N_8672,N_8267);
or U9120 (N_9120,N_8349,N_8745);
and U9121 (N_9121,N_8973,N_8477);
nor U9122 (N_9122,N_8941,N_8652);
or U9123 (N_9123,N_8074,N_8241);
nand U9124 (N_9124,N_8167,N_8275);
nor U9125 (N_9125,N_8291,N_8816);
or U9126 (N_9126,N_8744,N_8025);
xor U9127 (N_9127,N_8379,N_8556);
and U9128 (N_9128,N_8863,N_8632);
and U9129 (N_9129,N_8761,N_8634);
nor U9130 (N_9130,N_8129,N_8070);
nand U9131 (N_9131,N_8115,N_8627);
nand U9132 (N_9132,N_8720,N_8363);
or U9133 (N_9133,N_8387,N_8791);
or U9134 (N_9134,N_8339,N_8168);
or U9135 (N_9135,N_8807,N_8907);
nand U9136 (N_9136,N_8004,N_8998);
nor U9137 (N_9137,N_8325,N_8355);
and U9138 (N_9138,N_8476,N_8963);
nor U9139 (N_9139,N_8200,N_8979);
or U9140 (N_9140,N_8824,N_8373);
nor U9141 (N_9141,N_8692,N_8874);
and U9142 (N_9142,N_8710,N_8023);
nor U9143 (N_9143,N_8771,N_8577);
or U9144 (N_9144,N_8594,N_8994);
and U9145 (N_9145,N_8993,N_8794);
or U9146 (N_9146,N_8439,N_8235);
or U9147 (N_9147,N_8175,N_8348);
nand U9148 (N_9148,N_8790,N_8431);
or U9149 (N_9149,N_8781,N_8859);
or U9150 (N_9150,N_8678,N_8334);
and U9151 (N_9151,N_8223,N_8371);
and U9152 (N_9152,N_8840,N_8897);
nand U9153 (N_9153,N_8116,N_8085);
nor U9154 (N_9154,N_8323,N_8248);
and U9155 (N_9155,N_8259,N_8769);
nor U9156 (N_9156,N_8182,N_8521);
or U9157 (N_9157,N_8564,N_8404);
nor U9158 (N_9158,N_8433,N_8500);
nand U9159 (N_9159,N_8934,N_8475);
nand U9160 (N_9160,N_8156,N_8989);
nand U9161 (N_9161,N_8798,N_8034);
or U9162 (N_9162,N_8320,N_8547);
nor U9163 (N_9163,N_8708,N_8162);
nand U9164 (N_9164,N_8607,N_8161);
and U9165 (N_9165,N_8380,N_8332);
and U9166 (N_9166,N_8206,N_8341);
nor U9167 (N_9167,N_8610,N_8296);
nor U9168 (N_9168,N_8197,N_8123);
and U9169 (N_9169,N_8903,N_8658);
nor U9170 (N_9170,N_8960,N_8069);
nand U9171 (N_9171,N_8764,N_8835);
and U9172 (N_9172,N_8474,N_8163);
nand U9173 (N_9173,N_8177,N_8357);
nor U9174 (N_9174,N_8847,N_8049);
nand U9175 (N_9175,N_8920,N_8121);
nor U9176 (N_9176,N_8871,N_8496);
nor U9177 (N_9177,N_8746,N_8655);
and U9178 (N_9178,N_8898,N_8117);
nor U9179 (N_9179,N_8531,N_8974);
or U9180 (N_9180,N_8539,N_8336);
and U9181 (N_9181,N_8570,N_8212);
or U9182 (N_9182,N_8872,N_8130);
or U9183 (N_9183,N_8468,N_8636);
nor U9184 (N_9184,N_8942,N_8674);
nand U9185 (N_9185,N_8501,N_8489);
and U9186 (N_9186,N_8016,N_8073);
nand U9187 (N_9187,N_8252,N_8314);
nand U9188 (N_9188,N_8313,N_8830);
nor U9189 (N_9189,N_8715,N_8429);
or U9190 (N_9190,N_8759,N_8567);
and U9191 (N_9191,N_8462,N_8668);
nor U9192 (N_9192,N_8961,N_8653);
or U9193 (N_9193,N_8703,N_8140);
xnor U9194 (N_9194,N_8927,N_8426);
and U9195 (N_9195,N_8845,N_8659);
or U9196 (N_9196,N_8812,N_8626);
or U9197 (N_9197,N_8015,N_8081);
and U9198 (N_9198,N_8958,N_8839);
nand U9199 (N_9199,N_8243,N_8555);
nand U9200 (N_9200,N_8494,N_8698);
and U9201 (N_9201,N_8131,N_8482);
nand U9202 (N_9202,N_8728,N_8694);
nor U9203 (N_9203,N_8204,N_8006);
and U9204 (N_9204,N_8415,N_8400);
xor U9205 (N_9205,N_8524,N_8763);
and U9206 (N_9206,N_8734,N_8552);
nor U9207 (N_9207,N_8623,N_8188);
and U9208 (N_9208,N_8887,N_8939);
nor U9209 (N_9209,N_8249,N_8829);
nand U9210 (N_9210,N_8997,N_8526);
nor U9211 (N_9211,N_8721,N_8766);
or U9212 (N_9212,N_8370,N_8566);
or U9213 (N_9213,N_8417,N_8714);
nand U9214 (N_9214,N_8933,N_8160);
nor U9215 (N_9215,N_8155,N_8803);
or U9216 (N_9216,N_8257,N_8183);
nand U9217 (N_9217,N_8682,N_8788);
and U9218 (N_9218,N_8621,N_8848);
nor U9219 (N_9219,N_8324,N_8518);
nor U9220 (N_9220,N_8890,N_8663);
and U9221 (N_9221,N_8385,N_8622);
nand U9222 (N_9222,N_8392,N_8691);
and U9223 (N_9223,N_8194,N_8624);
nor U9224 (N_9224,N_8882,N_8354);
and U9225 (N_9225,N_8459,N_8209);
nand U9226 (N_9226,N_8309,N_8645);
or U9227 (N_9227,N_8638,N_8595);
or U9228 (N_9228,N_8152,N_8718);
nand U9229 (N_9229,N_8199,N_8393);
xnor U9230 (N_9230,N_8198,N_8498);
or U9231 (N_9231,N_8976,N_8101);
nor U9232 (N_9232,N_8514,N_8099);
or U9233 (N_9233,N_8043,N_8573);
nand U9234 (N_9234,N_8646,N_8487);
nand U9235 (N_9235,N_8418,N_8050);
and U9236 (N_9236,N_8327,N_8995);
and U9237 (N_9237,N_8001,N_8294);
and U9238 (N_9238,N_8569,N_8749);
nor U9239 (N_9239,N_8819,N_8650);
or U9240 (N_9240,N_8377,N_8702);
and U9241 (N_9241,N_8795,N_8176);
and U9242 (N_9242,N_8926,N_8836);
xnor U9243 (N_9243,N_8062,N_8925);
nand U9244 (N_9244,N_8495,N_8456);
or U9245 (N_9245,N_8724,N_8892);
nor U9246 (N_9246,N_8827,N_8665);
nand U9247 (N_9247,N_8705,N_8367);
and U9248 (N_9248,N_8512,N_8868);
and U9249 (N_9249,N_8128,N_8560);
nor U9250 (N_9250,N_8061,N_8282);
nor U9251 (N_9251,N_8068,N_8078);
nand U9252 (N_9252,N_8660,N_8885);
nand U9253 (N_9253,N_8723,N_8755);
nand U9254 (N_9254,N_8208,N_8304);
and U9255 (N_9255,N_8013,N_8171);
xnor U9256 (N_9256,N_8369,N_8180);
nand U9257 (N_9257,N_8597,N_8543);
nor U9258 (N_9258,N_8165,N_8254);
nand U9259 (N_9259,N_8598,N_8287);
and U9260 (N_9260,N_8114,N_8628);
nand U9261 (N_9261,N_8649,N_8669);
nand U9262 (N_9262,N_8347,N_8010);
nand U9263 (N_9263,N_8664,N_8120);
and U9264 (N_9264,N_8279,N_8881);
or U9265 (N_9265,N_8787,N_8612);
nor U9266 (N_9266,N_8530,N_8936);
nor U9267 (N_9267,N_8838,N_8318);
or U9268 (N_9268,N_8461,N_8760);
nand U9269 (N_9269,N_8805,N_8909);
or U9270 (N_9270,N_8056,N_8181);
or U9271 (N_9271,N_8810,N_8337);
or U9272 (N_9272,N_8063,N_8699);
nand U9273 (N_9273,N_8319,N_8242);
and U9274 (N_9274,N_8333,N_8195);
nor U9275 (N_9275,N_8455,N_8040);
or U9276 (N_9276,N_8486,N_8768);
and U9277 (N_9277,N_8000,N_8493);
or U9278 (N_9278,N_8266,N_8164);
nand U9279 (N_9279,N_8639,N_8913);
nor U9280 (N_9280,N_8880,N_8701);
xnor U9281 (N_9281,N_8362,N_8436);
or U9282 (N_9282,N_8350,N_8896);
and U9283 (N_9283,N_8024,N_8969);
nor U9284 (N_9284,N_8403,N_8931);
or U9285 (N_9285,N_8657,N_8384);
nand U9286 (N_9286,N_8011,N_8305);
or U9287 (N_9287,N_8110,N_8478);
or U9288 (N_9288,N_8583,N_8588);
and U9289 (N_9289,N_8725,N_8090);
or U9290 (N_9290,N_8870,N_8978);
and U9291 (N_9291,N_8844,N_8515);
nand U9292 (N_9292,N_8615,N_8877);
and U9293 (N_9293,N_8901,N_8281);
or U9294 (N_9294,N_8007,N_8297);
nand U9295 (N_9295,N_8435,N_8509);
nand U9296 (N_9296,N_8300,N_8224);
nand U9297 (N_9297,N_8631,N_8405);
and U9298 (N_9298,N_8875,N_8504);
and U9299 (N_9299,N_8908,N_8271);
nand U9300 (N_9300,N_8219,N_8322);
or U9301 (N_9301,N_8849,N_8340);
and U9302 (N_9302,N_8428,N_8317);
or U9303 (N_9303,N_8134,N_8139);
nor U9304 (N_9304,N_8792,N_8751);
or U9305 (N_9305,N_8706,N_8401);
nor U9306 (N_9306,N_8832,N_8358);
nand U9307 (N_9307,N_8105,N_8712);
nor U9308 (N_9308,N_8951,N_8540);
or U9309 (N_9309,N_8166,N_8879);
nand U9310 (N_9310,N_8753,N_8643);
nand U9311 (N_9311,N_8862,N_8368);
or U9312 (N_9312,N_8902,N_8522);
or U9313 (N_9313,N_8467,N_8579);
and U9314 (N_9314,N_8553,N_8173);
nand U9315 (N_9315,N_8575,N_8688);
nand U9316 (N_9316,N_8856,N_8921);
or U9317 (N_9317,N_8345,N_8463);
nand U9318 (N_9318,N_8421,N_8091);
and U9319 (N_9319,N_8092,N_8772);
nor U9320 (N_9320,N_8232,N_8743);
or U9321 (N_9321,N_8060,N_8947);
nand U9322 (N_9322,N_8372,N_8542);
or U9323 (N_9323,N_8479,N_8184);
or U9324 (N_9324,N_8065,N_8356);
or U9325 (N_9325,N_8932,N_8742);
or U9326 (N_9326,N_8591,N_8814);
xnor U9327 (N_9327,N_8044,N_8047);
nand U9328 (N_9328,N_8825,N_8629);
and U9329 (N_9329,N_8251,N_8834);
or U9330 (N_9330,N_8937,N_8538);
and U9331 (N_9331,N_8285,N_8473);
and U9332 (N_9332,N_8096,N_8042);
nand U9333 (N_9333,N_8364,N_8517);
nand U9334 (N_9334,N_8217,N_8440);
nand U9335 (N_9335,N_8716,N_8889);
or U9336 (N_9336,N_8483,N_8142);
nand U9337 (N_9337,N_8959,N_8021);
nand U9338 (N_9338,N_8697,N_8460);
and U9339 (N_9339,N_8471,N_8644);
nand U9340 (N_9340,N_8888,N_8264);
and U9341 (N_9341,N_8620,N_8765);
xnor U9342 (N_9342,N_8290,N_8295);
nand U9343 (N_9343,N_8253,N_8984);
nor U9344 (N_9344,N_8864,N_8828);
or U9345 (N_9345,N_8135,N_8143);
and U9346 (N_9346,N_8944,N_8783);
and U9347 (N_9347,N_8924,N_8095);
and U9348 (N_9348,N_8675,N_8344);
and U9349 (N_9349,N_8919,N_8565);
nor U9350 (N_9350,N_8239,N_8084);
nor U9351 (N_9351,N_8757,N_8302);
nor U9352 (N_9352,N_8205,N_8109);
nor U9353 (N_9353,N_8949,N_8214);
and U9354 (N_9354,N_8837,N_8956);
and U9355 (N_9355,N_8971,N_8237);
nand U9356 (N_9356,N_8310,N_8666);
nor U9357 (N_9357,N_8507,N_8141);
or U9358 (N_9358,N_8055,N_8258);
nand U9359 (N_9359,N_8052,N_8231);
nand U9360 (N_9360,N_8576,N_8111);
or U9361 (N_9361,N_8683,N_8525);
nand U9362 (N_9362,N_8144,N_8809);
xor U9363 (N_9363,N_8918,N_8752);
or U9364 (N_9364,N_8326,N_8048);
nor U9365 (N_9365,N_8038,N_8992);
and U9366 (N_9366,N_8826,N_8952);
and U9367 (N_9367,N_8179,N_8381);
nand U9368 (N_9368,N_8399,N_8935);
nand U9369 (N_9369,N_8793,N_8094);
or U9370 (N_9370,N_8424,N_8917);
nor U9371 (N_9371,N_8030,N_8923);
nand U9372 (N_9372,N_8457,N_8677);
and U9373 (N_9373,N_8453,N_8027);
nor U9374 (N_9374,N_8599,N_8738);
xor U9375 (N_9375,N_8767,N_8991);
nand U9376 (N_9376,N_8067,N_8990);
or U9377 (N_9377,N_8255,N_8818);
and U9378 (N_9378,N_8448,N_8409);
and U9379 (N_9379,N_8444,N_8900);
or U9380 (N_9380,N_8730,N_8563);
or U9381 (N_9381,N_8227,N_8861);
nor U9382 (N_9382,N_8817,N_8189);
and U9383 (N_9383,N_8492,N_8821);
nor U9384 (N_9384,N_8568,N_8003);
or U9385 (N_9385,N_8865,N_8108);
and U9386 (N_9386,N_8700,N_8883);
nand U9387 (N_9387,N_8159,N_8360);
nand U9388 (N_9388,N_8107,N_8511);
and U9389 (N_9389,N_8246,N_8193);
and U9390 (N_9390,N_8331,N_8833);
nor U9391 (N_9391,N_8386,N_8422);
and U9392 (N_9392,N_8449,N_8046);
nor U9393 (N_9393,N_8057,N_8886);
xnor U9394 (N_9394,N_8221,N_8022);
nor U9395 (N_9395,N_8203,N_8126);
nor U9396 (N_9396,N_8707,N_8964);
nand U9397 (N_9397,N_8546,N_8676);
and U9398 (N_9398,N_8681,N_8613);
and U9399 (N_9399,N_8434,N_8673);
nand U9400 (N_9400,N_8685,N_8080);
and U9401 (N_9401,N_8726,N_8736);
nand U9402 (N_9402,N_8869,N_8112);
nand U9403 (N_9403,N_8945,N_8608);
nor U9404 (N_9404,N_8397,N_8602);
nand U9405 (N_9405,N_8929,N_8970);
or U9406 (N_9406,N_8138,N_8329);
nor U9407 (N_9407,N_8262,N_8088);
or U9408 (N_9408,N_8276,N_8441);
nand U9409 (N_9409,N_8388,N_8283);
or U9410 (N_9410,N_8132,N_8284);
nand U9411 (N_9411,N_8306,N_8541);
or U9412 (N_9412,N_8671,N_8051);
and U9413 (N_9413,N_8938,N_8450);
nor U9414 (N_9414,N_8982,N_8797);
and U9415 (N_9415,N_8265,N_8077);
nor U9416 (N_9416,N_8948,N_8758);
or U9417 (N_9417,N_8041,N_8037);
or U9418 (N_9418,N_8020,N_8286);
or U9419 (N_9419,N_8667,N_8446);
nand U9420 (N_9420,N_8293,N_8469);
or U9421 (N_9421,N_8033,N_8137);
nor U9422 (N_9422,N_8442,N_8019);
nand U9423 (N_9423,N_8554,N_8637);
and U9424 (N_9424,N_8119,N_8559);
and U9425 (N_9425,N_8776,N_8335);
and U9426 (N_9426,N_8860,N_8854);
nor U9427 (N_9427,N_8911,N_8580);
and U9428 (N_9428,N_8912,N_8220);
nand U9429 (N_9429,N_8985,N_8072);
or U9430 (N_9430,N_8464,N_8557);
or U9431 (N_9431,N_8831,N_8202);
or U9432 (N_9432,N_8427,N_8419);
and U9433 (N_9433,N_8190,N_8374);
and U9434 (N_9434,N_8272,N_8891);
nand U9435 (N_9435,N_8841,N_8981);
nand U9436 (N_9436,N_8661,N_8389);
and U9437 (N_9437,N_8851,N_8640);
and U9438 (N_9438,N_8689,N_8382);
nor U9439 (N_9439,N_8071,N_8445);
nand U9440 (N_9440,N_8145,N_8808);
nor U9441 (N_9441,N_8562,N_8432);
and U9442 (N_9442,N_8523,N_8773);
or U9443 (N_9443,N_8534,N_8158);
or U9444 (N_9444,N_8187,N_8066);
nor U9445 (N_9445,N_8009,N_8813);
and U9446 (N_9446,N_8954,N_8601);
and U9447 (N_9447,N_8270,N_8213);
or U9448 (N_9448,N_8756,N_8032);
nor U9449 (N_9449,N_8028,N_8609);
nor U9450 (N_9450,N_8437,N_8303);
nand U9451 (N_9451,N_8505,N_8955);
nor U9452 (N_9452,N_8452,N_8447);
or U9453 (N_9453,N_8451,N_8353);
or U9454 (N_9454,N_8785,N_8800);
or U9455 (N_9455,N_8465,N_8876);
nand U9456 (N_9456,N_8741,N_8739);
nand U9457 (N_9457,N_8651,N_8378);
or U9458 (N_9458,N_8647,N_8811);
or U9459 (N_9459,N_8338,N_8654);
or U9460 (N_9460,N_8641,N_8617);
and U9461 (N_9461,N_8713,N_8940);
nand U9462 (N_9462,N_8059,N_8717);
xor U9463 (N_9463,N_8774,N_8170);
and U9464 (N_9464,N_8914,N_8529);
and U9465 (N_9465,N_8670,N_8490);
nor U9466 (N_9466,N_8731,N_8779);
or U9467 (N_9467,N_8928,N_8002);
or U9468 (N_9468,N_8625,N_8228);
and U9469 (N_9469,N_8365,N_8226);
and U9470 (N_9470,N_8268,N_8222);
or U9471 (N_9471,N_8778,N_8240);
xnor U9472 (N_9472,N_8125,N_8472);
and U9473 (N_9473,N_8207,N_8330);
or U9474 (N_9474,N_8996,N_8093);
nand U9475 (N_9475,N_8127,N_8648);
and U9476 (N_9476,N_8642,N_8846);
nor U9477 (N_9477,N_8590,N_8499);
xnor U9478 (N_9478,N_8915,N_8269);
nor U9479 (N_9479,N_8086,N_8843);
or U9480 (N_9480,N_8136,N_8906);
nand U9481 (N_9481,N_8014,N_8508);
and U9482 (N_9482,N_8822,N_8605);
or U9483 (N_9483,N_8238,N_8484);
or U9484 (N_9484,N_8361,N_8229);
and U9485 (N_9485,N_8425,N_8786);
and U9486 (N_9486,N_8191,N_8777);
or U9487 (N_9487,N_8980,N_8288);
and U9488 (N_9488,N_8722,N_8133);
and U9489 (N_9489,N_8630,N_8516);
nand U9490 (N_9490,N_8520,N_8784);
nand U9491 (N_9491,N_8585,N_8408);
nand U9492 (N_9492,N_8308,N_8480);
nor U9493 (N_9493,N_8342,N_8680);
nand U9494 (N_9494,N_8100,N_8053);
nor U9495 (N_9495,N_8192,N_8017);
nand U9496 (N_9496,N_8855,N_8506);
and U9497 (N_9497,N_8853,N_8039);
nand U9498 (N_9498,N_8578,N_8103);
nand U9499 (N_9499,N_8696,N_8729);
and U9500 (N_9500,N_8468,N_8236);
and U9501 (N_9501,N_8075,N_8099);
or U9502 (N_9502,N_8178,N_8312);
or U9503 (N_9503,N_8763,N_8730);
nor U9504 (N_9504,N_8011,N_8109);
nand U9505 (N_9505,N_8330,N_8953);
nand U9506 (N_9506,N_8223,N_8718);
nor U9507 (N_9507,N_8121,N_8501);
and U9508 (N_9508,N_8394,N_8406);
nor U9509 (N_9509,N_8050,N_8838);
nand U9510 (N_9510,N_8894,N_8469);
and U9511 (N_9511,N_8660,N_8066);
nand U9512 (N_9512,N_8807,N_8659);
and U9513 (N_9513,N_8573,N_8858);
nor U9514 (N_9514,N_8654,N_8430);
and U9515 (N_9515,N_8610,N_8439);
or U9516 (N_9516,N_8297,N_8838);
xnor U9517 (N_9517,N_8869,N_8550);
nor U9518 (N_9518,N_8424,N_8293);
or U9519 (N_9519,N_8659,N_8135);
nor U9520 (N_9520,N_8509,N_8559);
and U9521 (N_9521,N_8715,N_8926);
nor U9522 (N_9522,N_8718,N_8245);
nand U9523 (N_9523,N_8149,N_8129);
nand U9524 (N_9524,N_8573,N_8484);
or U9525 (N_9525,N_8690,N_8699);
or U9526 (N_9526,N_8238,N_8492);
and U9527 (N_9527,N_8751,N_8294);
nor U9528 (N_9528,N_8775,N_8041);
nor U9529 (N_9529,N_8241,N_8373);
nor U9530 (N_9530,N_8637,N_8595);
or U9531 (N_9531,N_8869,N_8997);
or U9532 (N_9532,N_8589,N_8310);
nand U9533 (N_9533,N_8600,N_8404);
and U9534 (N_9534,N_8602,N_8669);
nand U9535 (N_9535,N_8551,N_8727);
and U9536 (N_9536,N_8908,N_8037);
and U9537 (N_9537,N_8218,N_8239);
nand U9538 (N_9538,N_8239,N_8800);
or U9539 (N_9539,N_8540,N_8238);
or U9540 (N_9540,N_8838,N_8800);
nand U9541 (N_9541,N_8564,N_8117);
nand U9542 (N_9542,N_8547,N_8072);
and U9543 (N_9543,N_8690,N_8971);
nor U9544 (N_9544,N_8961,N_8272);
nor U9545 (N_9545,N_8317,N_8667);
nand U9546 (N_9546,N_8984,N_8117);
or U9547 (N_9547,N_8920,N_8698);
nor U9548 (N_9548,N_8838,N_8852);
and U9549 (N_9549,N_8692,N_8974);
nor U9550 (N_9550,N_8818,N_8779);
and U9551 (N_9551,N_8091,N_8244);
nor U9552 (N_9552,N_8468,N_8960);
nor U9553 (N_9553,N_8254,N_8483);
nand U9554 (N_9554,N_8024,N_8840);
or U9555 (N_9555,N_8527,N_8558);
nand U9556 (N_9556,N_8754,N_8150);
nor U9557 (N_9557,N_8873,N_8257);
nand U9558 (N_9558,N_8080,N_8046);
and U9559 (N_9559,N_8568,N_8886);
nand U9560 (N_9560,N_8538,N_8665);
or U9561 (N_9561,N_8500,N_8182);
and U9562 (N_9562,N_8330,N_8011);
nor U9563 (N_9563,N_8113,N_8790);
xor U9564 (N_9564,N_8042,N_8697);
or U9565 (N_9565,N_8370,N_8309);
xor U9566 (N_9566,N_8783,N_8768);
or U9567 (N_9567,N_8883,N_8586);
or U9568 (N_9568,N_8735,N_8255);
and U9569 (N_9569,N_8253,N_8947);
nor U9570 (N_9570,N_8671,N_8191);
and U9571 (N_9571,N_8216,N_8669);
nand U9572 (N_9572,N_8442,N_8262);
nand U9573 (N_9573,N_8064,N_8433);
nor U9574 (N_9574,N_8347,N_8428);
or U9575 (N_9575,N_8947,N_8756);
and U9576 (N_9576,N_8766,N_8005);
nand U9577 (N_9577,N_8409,N_8413);
nand U9578 (N_9578,N_8877,N_8152);
nor U9579 (N_9579,N_8082,N_8073);
nor U9580 (N_9580,N_8583,N_8853);
nand U9581 (N_9581,N_8260,N_8061);
nor U9582 (N_9582,N_8722,N_8848);
or U9583 (N_9583,N_8488,N_8263);
nand U9584 (N_9584,N_8596,N_8176);
xor U9585 (N_9585,N_8804,N_8664);
nand U9586 (N_9586,N_8365,N_8012);
or U9587 (N_9587,N_8262,N_8312);
nand U9588 (N_9588,N_8162,N_8165);
xor U9589 (N_9589,N_8055,N_8925);
nor U9590 (N_9590,N_8237,N_8092);
and U9591 (N_9591,N_8959,N_8942);
nor U9592 (N_9592,N_8168,N_8385);
nand U9593 (N_9593,N_8583,N_8130);
nand U9594 (N_9594,N_8372,N_8229);
or U9595 (N_9595,N_8487,N_8160);
nor U9596 (N_9596,N_8216,N_8315);
nor U9597 (N_9597,N_8878,N_8153);
and U9598 (N_9598,N_8106,N_8659);
or U9599 (N_9599,N_8716,N_8289);
or U9600 (N_9600,N_8346,N_8773);
and U9601 (N_9601,N_8023,N_8727);
or U9602 (N_9602,N_8688,N_8043);
nor U9603 (N_9603,N_8210,N_8993);
or U9604 (N_9604,N_8415,N_8730);
and U9605 (N_9605,N_8255,N_8177);
and U9606 (N_9606,N_8530,N_8201);
nor U9607 (N_9607,N_8740,N_8137);
nand U9608 (N_9608,N_8355,N_8420);
nor U9609 (N_9609,N_8031,N_8370);
nor U9610 (N_9610,N_8024,N_8328);
and U9611 (N_9611,N_8205,N_8518);
or U9612 (N_9612,N_8192,N_8096);
nor U9613 (N_9613,N_8392,N_8968);
nor U9614 (N_9614,N_8808,N_8182);
or U9615 (N_9615,N_8867,N_8147);
nor U9616 (N_9616,N_8397,N_8311);
nor U9617 (N_9617,N_8945,N_8544);
and U9618 (N_9618,N_8005,N_8255);
and U9619 (N_9619,N_8313,N_8272);
nor U9620 (N_9620,N_8061,N_8403);
and U9621 (N_9621,N_8993,N_8097);
nor U9622 (N_9622,N_8141,N_8366);
or U9623 (N_9623,N_8301,N_8187);
nand U9624 (N_9624,N_8065,N_8464);
or U9625 (N_9625,N_8802,N_8053);
nor U9626 (N_9626,N_8171,N_8078);
xnor U9627 (N_9627,N_8968,N_8342);
nand U9628 (N_9628,N_8412,N_8525);
nand U9629 (N_9629,N_8875,N_8541);
nand U9630 (N_9630,N_8158,N_8460);
nand U9631 (N_9631,N_8884,N_8539);
or U9632 (N_9632,N_8000,N_8158);
and U9633 (N_9633,N_8985,N_8941);
nand U9634 (N_9634,N_8432,N_8789);
nand U9635 (N_9635,N_8087,N_8798);
or U9636 (N_9636,N_8626,N_8509);
nand U9637 (N_9637,N_8962,N_8452);
or U9638 (N_9638,N_8418,N_8962);
and U9639 (N_9639,N_8285,N_8566);
nand U9640 (N_9640,N_8319,N_8477);
nor U9641 (N_9641,N_8258,N_8026);
nor U9642 (N_9642,N_8800,N_8880);
or U9643 (N_9643,N_8228,N_8058);
nor U9644 (N_9644,N_8834,N_8841);
nor U9645 (N_9645,N_8416,N_8429);
and U9646 (N_9646,N_8475,N_8054);
or U9647 (N_9647,N_8781,N_8551);
nand U9648 (N_9648,N_8561,N_8979);
nand U9649 (N_9649,N_8974,N_8003);
and U9650 (N_9650,N_8341,N_8474);
or U9651 (N_9651,N_8336,N_8942);
and U9652 (N_9652,N_8804,N_8729);
xor U9653 (N_9653,N_8687,N_8594);
and U9654 (N_9654,N_8575,N_8307);
or U9655 (N_9655,N_8623,N_8445);
nand U9656 (N_9656,N_8211,N_8176);
nor U9657 (N_9657,N_8570,N_8824);
and U9658 (N_9658,N_8735,N_8960);
or U9659 (N_9659,N_8994,N_8035);
nand U9660 (N_9660,N_8962,N_8823);
nand U9661 (N_9661,N_8408,N_8902);
nand U9662 (N_9662,N_8940,N_8357);
nand U9663 (N_9663,N_8374,N_8586);
nand U9664 (N_9664,N_8097,N_8881);
nand U9665 (N_9665,N_8434,N_8527);
nand U9666 (N_9666,N_8207,N_8938);
nand U9667 (N_9667,N_8062,N_8663);
nor U9668 (N_9668,N_8094,N_8753);
nand U9669 (N_9669,N_8812,N_8280);
nor U9670 (N_9670,N_8471,N_8934);
nor U9671 (N_9671,N_8517,N_8724);
nor U9672 (N_9672,N_8051,N_8673);
or U9673 (N_9673,N_8073,N_8989);
or U9674 (N_9674,N_8582,N_8050);
nor U9675 (N_9675,N_8589,N_8314);
nand U9676 (N_9676,N_8490,N_8585);
or U9677 (N_9677,N_8325,N_8422);
and U9678 (N_9678,N_8603,N_8282);
nor U9679 (N_9679,N_8716,N_8396);
and U9680 (N_9680,N_8942,N_8538);
and U9681 (N_9681,N_8648,N_8849);
or U9682 (N_9682,N_8642,N_8069);
or U9683 (N_9683,N_8433,N_8424);
nand U9684 (N_9684,N_8162,N_8175);
and U9685 (N_9685,N_8247,N_8805);
or U9686 (N_9686,N_8149,N_8958);
nand U9687 (N_9687,N_8964,N_8107);
and U9688 (N_9688,N_8366,N_8151);
xor U9689 (N_9689,N_8153,N_8474);
xnor U9690 (N_9690,N_8456,N_8711);
nor U9691 (N_9691,N_8939,N_8878);
xnor U9692 (N_9692,N_8197,N_8756);
and U9693 (N_9693,N_8674,N_8155);
nand U9694 (N_9694,N_8938,N_8853);
nand U9695 (N_9695,N_8815,N_8987);
or U9696 (N_9696,N_8842,N_8003);
nor U9697 (N_9697,N_8361,N_8596);
nand U9698 (N_9698,N_8052,N_8523);
or U9699 (N_9699,N_8475,N_8349);
nand U9700 (N_9700,N_8431,N_8007);
or U9701 (N_9701,N_8433,N_8890);
and U9702 (N_9702,N_8121,N_8958);
and U9703 (N_9703,N_8303,N_8976);
nand U9704 (N_9704,N_8111,N_8779);
or U9705 (N_9705,N_8577,N_8110);
and U9706 (N_9706,N_8667,N_8904);
nand U9707 (N_9707,N_8173,N_8562);
and U9708 (N_9708,N_8267,N_8576);
nor U9709 (N_9709,N_8202,N_8124);
nand U9710 (N_9710,N_8403,N_8103);
xor U9711 (N_9711,N_8941,N_8902);
nand U9712 (N_9712,N_8691,N_8185);
and U9713 (N_9713,N_8916,N_8657);
and U9714 (N_9714,N_8016,N_8175);
xnor U9715 (N_9715,N_8398,N_8836);
nor U9716 (N_9716,N_8262,N_8432);
nor U9717 (N_9717,N_8968,N_8847);
or U9718 (N_9718,N_8230,N_8347);
and U9719 (N_9719,N_8526,N_8202);
or U9720 (N_9720,N_8618,N_8720);
and U9721 (N_9721,N_8089,N_8728);
nand U9722 (N_9722,N_8651,N_8647);
or U9723 (N_9723,N_8676,N_8165);
nor U9724 (N_9724,N_8083,N_8239);
nor U9725 (N_9725,N_8449,N_8967);
and U9726 (N_9726,N_8014,N_8858);
nand U9727 (N_9727,N_8158,N_8899);
or U9728 (N_9728,N_8778,N_8139);
or U9729 (N_9729,N_8137,N_8560);
nor U9730 (N_9730,N_8484,N_8762);
and U9731 (N_9731,N_8794,N_8079);
and U9732 (N_9732,N_8380,N_8182);
nor U9733 (N_9733,N_8897,N_8842);
nand U9734 (N_9734,N_8003,N_8324);
or U9735 (N_9735,N_8741,N_8547);
or U9736 (N_9736,N_8112,N_8558);
nand U9737 (N_9737,N_8923,N_8711);
nand U9738 (N_9738,N_8232,N_8268);
or U9739 (N_9739,N_8914,N_8112);
and U9740 (N_9740,N_8941,N_8885);
nor U9741 (N_9741,N_8726,N_8123);
nand U9742 (N_9742,N_8746,N_8806);
nand U9743 (N_9743,N_8830,N_8106);
or U9744 (N_9744,N_8266,N_8007);
or U9745 (N_9745,N_8634,N_8262);
and U9746 (N_9746,N_8697,N_8906);
nor U9747 (N_9747,N_8524,N_8692);
nand U9748 (N_9748,N_8962,N_8961);
nand U9749 (N_9749,N_8910,N_8847);
nor U9750 (N_9750,N_8644,N_8740);
or U9751 (N_9751,N_8785,N_8528);
nor U9752 (N_9752,N_8374,N_8512);
nor U9753 (N_9753,N_8446,N_8488);
and U9754 (N_9754,N_8291,N_8558);
or U9755 (N_9755,N_8249,N_8094);
xor U9756 (N_9756,N_8208,N_8772);
or U9757 (N_9757,N_8478,N_8496);
or U9758 (N_9758,N_8808,N_8488);
or U9759 (N_9759,N_8999,N_8488);
nand U9760 (N_9760,N_8975,N_8191);
and U9761 (N_9761,N_8969,N_8092);
or U9762 (N_9762,N_8657,N_8721);
or U9763 (N_9763,N_8511,N_8994);
and U9764 (N_9764,N_8574,N_8598);
and U9765 (N_9765,N_8894,N_8307);
nand U9766 (N_9766,N_8951,N_8678);
or U9767 (N_9767,N_8796,N_8891);
and U9768 (N_9768,N_8196,N_8146);
or U9769 (N_9769,N_8181,N_8609);
nand U9770 (N_9770,N_8944,N_8606);
or U9771 (N_9771,N_8745,N_8009);
nor U9772 (N_9772,N_8434,N_8414);
and U9773 (N_9773,N_8875,N_8730);
nand U9774 (N_9774,N_8506,N_8260);
nor U9775 (N_9775,N_8515,N_8869);
or U9776 (N_9776,N_8615,N_8429);
nand U9777 (N_9777,N_8315,N_8292);
nand U9778 (N_9778,N_8425,N_8479);
or U9779 (N_9779,N_8987,N_8076);
and U9780 (N_9780,N_8322,N_8952);
and U9781 (N_9781,N_8955,N_8264);
nand U9782 (N_9782,N_8854,N_8557);
nand U9783 (N_9783,N_8413,N_8014);
and U9784 (N_9784,N_8165,N_8036);
or U9785 (N_9785,N_8468,N_8659);
and U9786 (N_9786,N_8096,N_8689);
and U9787 (N_9787,N_8205,N_8234);
or U9788 (N_9788,N_8344,N_8457);
and U9789 (N_9789,N_8625,N_8403);
and U9790 (N_9790,N_8808,N_8505);
nor U9791 (N_9791,N_8030,N_8893);
and U9792 (N_9792,N_8897,N_8760);
nor U9793 (N_9793,N_8054,N_8583);
and U9794 (N_9794,N_8964,N_8853);
and U9795 (N_9795,N_8787,N_8015);
nor U9796 (N_9796,N_8722,N_8883);
and U9797 (N_9797,N_8361,N_8312);
xnor U9798 (N_9798,N_8402,N_8196);
nand U9799 (N_9799,N_8999,N_8397);
or U9800 (N_9800,N_8614,N_8625);
or U9801 (N_9801,N_8394,N_8586);
nor U9802 (N_9802,N_8723,N_8879);
or U9803 (N_9803,N_8010,N_8869);
nor U9804 (N_9804,N_8587,N_8691);
or U9805 (N_9805,N_8162,N_8526);
and U9806 (N_9806,N_8336,N_8801);
nor U9807 (N_9807,N_8995,N_8434);
nor U9808 (N_9808,N_8513,N_8162);
or U9809 (N_9809,N_8743,N_8369);
nor U9810 (N_9810,N_8236,N_8208);
or U9811 (N_9811,N_8353,N_8404);
nand U9812 (N_9812,N_8787,N_8892);
nor U9813 (N_9813,N_8581,N_8382);
or U9814 (N_9814,N_8748,N_8410);
nor U9815 (N_9815,N_8167,N_8805);
and U9816 (N_9816,N_8886,N_8132);
nand U9817 (N_9817,N_8815,N_8613);
and U9818 (N_9818,N_8461,N_8852);
nor U9819 (N_9819,N_8497,N_8786);
xnor U9820 (N_9820,N_8163,N_8975);
xnor U9821 (N_9821,N_8711,N_8289);
and U9822 (N_9822,N_8115,N_8212);
and U9823 (N_9823,N_8768,N_8925);
nand U9824 (N_9824,N_8534,N_8576);
and U9825 (N_9825,N_8109,N_8789);
or U9826 (N_9826,N_8067,N_8340);
or U9827 (N_9827,N_8467,N_8419);
nor U9828 (N_9828,N_8884,N_8775);
and U9829 (N_9829,N_8720,N_8135);
nor U9830 (N_9830,N_8396,N_8449);
and U9831 (N_9831,N_8632,N_8175);
nand U9832 (N_9832,N_8170,N_8146);
nand U9833 (N_9833,N_8175,N_8892);
and U9834 (N_9834,N_8971,N_8540);
or U9835 (N_9835,N_8041,N_8035);
and U9836 (N_9836,N_8463,N_8473);
and U9837 (N_9837,N_8957,N_8554);
or U9838 (N_9838,N_8578,N_8690);
nor U9839 (N_9839,N_8078,N_8347);
xnor U9840 (N_9840,N_8324,N_8709);
or U9841 (N_9841,N_8216,N_8657);
nand U9842 (N_9842,N_8695,N_8964);
nor U9843 (N_9843,N_8013,N_8027);
nor U9844 (N_9844,N_8453,N_8956);
nand U9845 (N_9845,N_8906,N_8370);
or U9846 (N_9846,N_8176,N_8064);
and U9847 (N_9847,N_8745,N_8259);
nor U9848 (N_9848,N_8667,N_8664);
and U9849 (N_9849,N_8247,N_8604);
and U9850 (N_9850,N_8573,N_8078);
xnor U9851 (N_9851,N_8490,N_8308);
nor U9852 (N_9852,N_8081,N_8705);
or U9853 (N_9853,N_8428,N_8216);
nand U9854 (N_9854,N_8836,N_8291);
or U9855 (N_9855,N_8664,N_8714);
and U9856 (N_9856,N_8224,N_8882);
nor U9857 (N_9857,N_8607,N_8334);
and U9858 (N_9858,N_8892,N_8923);
and U9859 (N_9859,N_8050,N_8009);
nor U9860 (N_9860,N_8990,N_8438);
and U9861 (N_9861,N_8033,N_8322);
or U9862 (N_9862,N_8580,N_8456);
or U9863 (N_9863,N_8764,N_8699);
nand U9864 (N_9864,N_8358,N_8564);
nor U9865 (N_9865,N_8312,N_8703);
nor U9866 (N_9866,N_8097,N_8746);
and U9867 (N_9867,N_8871,N_8361);
nor U9868 (N_9868,N_8111,N_8656);
xor U9869 (N_9869,N_8768,N_8203);
or U9870 (N_9870,N_8266,N_8184);
nor U9871 (N_9871,N_8052,N_8417);
nor U9872 (N_9872,N_8034,N_8863);
or U9873 (N_9873,N_8368,N_8515);
and U9874 (N_9874,N_8226,N_8876);
nand U9875 (N_9875,N_8415,N_8535);
nor U9876 (N_9876,N_8343,N_8788);
or U9877 (N_9877,N_8076,N_8500);
or U9878 (N_9878,N_8984,N_8945);
or U9879 (N_9879,N_8384,N_8165);
or U9880 (N_9880,N_8199,N_8433);
nor U9881 (N_9881,N_8338,N_8941);
nor U9882 (N_9882,N_8139,N_8361);
or U9883 (N_9883,N_8174,N_8491);
or U9884 (N_9884,N_8877,N_8562);
nor U9885 (N_9885,N_8818,N_8118);
nor U9886 (N_9886,N_8570,N_8075);
nor U9887 (N_9887,N_8982,N_8310);
nand U9888 (N_9888,N_8068,N_8566);
or U9889 (N_9889,N_8573,N_8184);
nand U9890 (N_9890,N_8110,N_8735);
and U9891 (N_9891,N_8727,N_8525);
or U9892 (N_9892,N_8622,N_8659);
and U9893 (N_9893,N_8622,N_8965);
nand U9894 (N_9894,N_8376,N_8280);
nor U9895 (N_9895,N_8060,N_8697);
and U9896 (N_9896,N_8819,N_8042);
and U9897 (N_9897,N_8462,N_8385);
nor U9898 (N_9898,N_8095,N_8571);
and U9899 (N_9899,N_8309,N_8768);
nor U9900 (N_9900,N_8774,N_8674);
or U9901 (N_9901,N_8932,N_8715);
nor U9902 (N_9902,N_8032,N_8725);
nor U9903 (N_9903,N_8063,N_8945);
and U9904 (N_9904,N_8610,N_8072);
or U9905 (N_9905,N_8845,N_8613);
or U9906 (N_9906,N_8796,N_8835);
and U9907 (N_9907,N_8978,N_8575);
nor U9908 (N_9908,N_8938,N_8912);
and U9909 (N_9909,N_8711,N_8497);
or U9910 (N_9910,N_8376,N_8208);
nor U9911 (N_9911,N_8606,N_8575);
nor U9912 (N_9912,N_8873,N_8806);
nand U9913 (N_9913,N_8513,N_8188);
nand U9914 (N_9914,N_8111,N_8843);
and U9915 (N_9915,N_8966,N_8913);
or U9916 (N_9916,N_8409,N_8318);
nor U9917 (N_9917,N_8155,N_8501);
or U9918 (N_9918,N_8476,N_8229);
nor U9919 (N_9919,N_8818,N_8185);
nor U9920 (N_9920,N_8164,N_8662);
xor U9921 (N_9921,N_8725,N_8785);
and U9922 (N_9922,N_8097,N_8196);
and U9923 (N_9923,N_8459,N_8696);
and U9924 (N_9924,N_8793,N_8708);
or U9925 (N_9925,N_8690,N_8499);
nor U9926 (N_9926,N_8861,N_8073);
or U9927 (N_9927,N_8599,N_8646);
nand U9928 (N_9928,N_8946,N_8714);
or U9929 (N_9929,N_8591,N_8835);
nand U9930 (N_9930,N_8326,N_8422);
and U9931 (N_9931,N_8341,N_8268);
nor U9932 (N_9932,N_8561,N_8436);
or U9933 (N_9933,N_8941,N_8333);
and U9934 (N_9934,N_8667,N_8698);
and U9935 (N_9935,N_8349,N_8241);
or U9936 (N_9936,N_8681,N_8247);
xnor U9937 (N_9937,N_8293,N_8056);
or U9938 (N_9938,N_8515,N_8768);
nand U9939 (N_9939,N_8698,N_8031);
nand U9940 (N_9940,N_8169,N_8851);
and U9941 (N_9941,N_8448,N_8622);
nor U9942 (N_9942,N_8537,N_8216);
nand U9943 (N_9943,N_8326,N_8844);
nand U9944 (N_9944,N_8904,N_8967);
and U9945 (N_9945,N_8380,N_8638);
or U9946 (N_9946,N_8779,N_8025);
nor U9947 (N_9947,N_8261,N_8902);
and U9948 (N_9948,N_8009,N_8366);
nand U9949 (N_9949,N_8371,N_8993);
or U9950 (N_9950,N_8214,N_8115);
nand U9951 (N_9951,N_8144,N_8243);
nor U9952 (N_9952,N_8767,N_8489);
or U9953 (N_9953,N_8739,N_8309);
nand U9954 (N_9954,N_8984,N_8198);
and U9955 (N_9955,N_8537,N_8427);
nand U9956 (N_9956,N_8695,N_8603);
nor U9957 (N_9957,N_8661,N_8954);
nand U9958 (N_9958,N_8945,N_8264);
nor U9959 (N_9959,N_8064,N_8382);
and U9960 (N_9960,N_8928,N_8769);
nor U9961 (N_9961,N_8643,N_8862);
or U9962 (N_9962,N_8910,N_8850);
nor U9963 (N_9963,N_8206,N_8491);
and U9964 (N_9964,N_8286,N_8818);
nor U9965 (N_9965,N_8540,N_8470);
nor U9966 (N_9966,N_8899,N_8055);
or U9967 (N_9967,N_8153,N_8888);
and U9968 (N_9968,N_8048,N_8171);
nor U9969 (N_9969,N_8190,N_8040);
xor U9970 (N_9970,N_8033,N_8709);
and U9971 (N_9971,N_8995,N_8545);
xor U9972 (N_9972,N_8924,N_8545);
and U9973 (N_9973,N_8412,N_8654);
or U9974 (N_9974,N_8838,N_8605);
nor U9975 (N_9975,N_8255,N_8354);
nand U9976 (N_9976,N_8431,N_8362);
nor U9977 (N_9977,N_8338,N_8033);
nand U9978 (N_9978,N_8310,N_8318);
nand U9979 (N_9979,N_8430,N_8662);
xor U9980 (N_9980,N_8134,N_8782);
nor U9981 (N_9981,N_8883,N_8075);
nand U9982 (N_9982,N_8764,N_8155);
nor U9983 (N_9983,N_8360,N_8394);
or U9984 (N_9984,N_8990,N_8493);
or U9985 (N_9985,N_8483,N_8375);
nand U9986 (N_9986,N_8849,N_8883);
nor U9987 (N_9987,N_8510,N_8561);
nor U9988 (N_9988,N_8078,N_8449);
nand U9989 (N_9989,N_8264,N_8589);
or U9990 (N_9990,N_8242,N_8877);
xor U9991 (N_9991,N_8660,N_8977);
nand U9992 (N_9992,N_8318,N_8541);
and U9993 (N_9993,N_8288,N_8368);
and U9994 (N_9994,N_8341,N_8724);
nand U9995 (N_9995,N_8733,N_8823);
nand U9996 (N_9996,N_8349,N_8488);
nand U9997 (N_9997,N_8714,N_8907);
nor U9998 (N_9998,N_8231,N_8002);
or U9999 (N_9999,N_8406,N_8509);
and UO_0 (O_0,N_9037,N_9325);
nor UO_1 (O_1,N_9696,N_9440);
nand UO_2 (O_2,N_9835,N_9523);
and UO_3 (O_3,N_9115,N_9788);
and UO_4 (O_4,N_9389,N_9890);
and UO_5 (O_5,N_9393,N_9051);
or UO_6 (O_6,N_9940,N_9023);
nand UO_7 (O_7,N_9375,N_9084);
or UO_8 (O_8,N_9821,N_9799);
nand UO_9 (O_9,N_9823,N_9424);
nor UO_10 (O_10,N_9842,N_9625);
or UO_11 (O_11,N_9483,N_9571);
or UO_12 (O_12,N_9584,N_9118);
nor UO_13 (O_13,N_9709,N_9364);
nand UO_14 (O_14,N_9630,N_9260);
and UO_15 (O_15,N_9242,N_9038);
and UO_16 (O_16,N_9882,N_9144);
and UO_17 (O_17,N_9870,N_9559);
or UO_18 (O_18,N_9666,N_9908);
nand UO_19 (O_19,N_9831,N_9427);
nor UO_20 (O_20,N_9861,N_9984);
nand UO_21 (O_21,N_9694,N_9490);
xor UO_22 (O_22,N_9172,N_9922);
nor UO_23 (O_23,N_9065,N_9949);
or UO_24 (O_24,N_9638,N_9508);
and UO_25 (O_25,N_9879,N_9824);
nand UO_26 (O_26,N_9288,N_9199);
nand UO_27 (O_27,N_9676,N_9374);
and UO_28 (O_28,N_9511,N_9255);
or UO_29 (O_29,N_9329,N_9649);
nand UO_30 (O_30,N_9756,N_9425);
nor UO_31 (O_31,N_9281,N_9341);
nor UO_32 (O_32,N_9970,N_9647);
or UO_33 (O_33,N_9176,N_9175);
xor UO_34 (O_34,N_9955,N_9719);
or UO_35 (O_35,N_9104,N_9088);
nand UO_36 (O_36,N_9365,N_9860);
nor UO_37 (O_37,N_9189,N_9096);
or UO_38 (O_38,N_9867,N_9204);
or UO_39 (O_39,N_9733,N_9310);
or UO_40 (O_40,N_9520,N_9320);
nand UO_41 (O_41,N_9943,N_9106);
nor UO_42 (O_42,N_9330,N_9463);
nand UO_43 (O_43,N_9053,N_9928);
or UO_44 (O_44,N_9566,N_9976);
and UO_45 (O_45,N_9752,N_9293);
nand UO_46 (O_46,N_9224,N_9459);
or UO_47 (O_47,N_9070,N_9800);
nand UO_48 (O_48,N_9911,N_9685);
nand UO_49 (O_49,N_9311,N_9679);
nand UO_50 (O_50,N_9141,N_9889);
nor UO_51 (O_51,N_9136,N_9094);
nor UO_52 (O_52,N_9658,N_9631);
nand UO_53 (O_53,N_9677,N_9160);
and UO_54 (O_54,N_9642,N_9818);
and UO_55 (O_55,N_9482,N_9801);
nand UO_56 (O_56,N_9188,N_9367);
or UO_57 (O_57,N_9624,N_9787);
xnor UO_58 (O_58,N_9004,N_9877);
nand UO_59 (O_59,N_9468,N_9057);
nor UO_60 (O_60,N_9689,N_9186);
nand UO_61 (O_61,N_9539,N_9639);
or UO_62 (O_62,N_9282,N_9525);
or UO_63 (O_63,N_9028,N_9110);
nand UO_64 (O_64,N_9581,N_9011);
or UO_65 (O_65,N_9122,N_9612);
nor UO_66 (O_66,N_9589,N_9198);
and UO_67 (O_67,N_9243,N_9034);
and UO_68 (O_68,N_9682,N_9797);
nor UO_69 (O_69,N_9662,N_9058);
or UO_70 (O_70,N_9864,N_9267);
nor UO_71 (O_71,N_9646,N_9203);
and UO_72 (O_72,N_9193,N_9181);
nor UO_73 (O_73,N_9335,N_9415);
nand UO_74 (O_74,N_9572,N_9368);
nand UO_75 (O_75,N_9904,N_9405);
nand UO_76 (O_76,N_9985,N_9085);
nand UO_77 (O_77,N_9099,N_9822);
nand UO_78 (O_78,N_9875,N_9771);
nor UO_79 (O_79,N_9066,N_9361);
xnor UO_80 (O_80,N_9245,N_9447);
nand UO_81 (O_81,N_9516,N_9116);
and UO_82 (O_82,N_9919,N_9829);
and UO_83 (O_83,N_9497,N_9806);
or UO_84 (O_84,N_9628,N_9924);
nand UO_85 (O_85,N_9072,N_9419);
and UO_86 (O_86,N_9741,N_9794);
or UO_87 (O_87,N_9276,N_9734);
nand UO_88 (O_88,N_9993,N_9074);
or UO_89 (O_89,N_9180,N_9123);
or UO_90 (O_90,N_9443,N_9640);
nand UO_91 (O_91,N_9183,N_9167);
xnor UO_92 (O_92,N_9636,N_9207);
nand UO_93 (O_93,N_9754,N_9804);
and UO_94 (O_94,N_9888,N_9112);
nor UO_95 (O_95,N_9700,N_9915);
or UO_96 (O_96,N_9323,N_9645);
nor UO_97 (O_97,N_9796,N_9237);
nand UO_98 (O_98,N_9776,N_9306);
nand UO_99 (O_99,N_9934,N_9151);
and UO_100 (O_100,N_9397,N_9248);
or UO_101 (O_101,N_9385,N_9359);
nand UO_102 (O_102,N_9878,N_9891);
nand UO_103 (O_103,N_9960,N_9579);
and UO_104 (O_104,N_9377,N_9309);
nand UO_105 (O_105,N_9973,N_9708);
nor UO_106 (O_106,N_9716,N_9978);
and UO_107 (O_107,N_9035,N_9608);
and UO_108 (O_108,N_9456,N_9544);
and UO_109 (O_109,N_9462,N_9880);
nor UO_110 (O_110,N_9674,N_9495);
and UO_111 (O_111,N_9120,N_9308);
nor UO_112 (O_112,N_9568,N_9277);
nor UO_113 (O_113,N_9580,N_9554);
xor UO_114 (O_114,N_9097,N_9270);
nor UO_115 (O_115,N_9262,N_9812);
nor UO_116 (O_116,N_9157,N_9143);
nand UO_117 (O_117,N_9721,N_9827);
nor UO_118 (O_118,N_9912,N_9672);
and UO_119 (O_119,N_9760,N_9078);
and UO_120 (O_120,N_9974,N_9531);
or UO_121 (O_121,N_9863,N_9016);
or UO_122 (O_122,N_9938,N_9394);
nand UO_123 (O_123,N_9107,N_9898);
and UO_124 (O_124,N_9986,N_9965);
nand UO_125 (O_125,N_9656,N_9913);
nor UO_126 (O_126,N_9856,N_9504);
or UO_127 (O_127,N_9522,N_9414);
and UO_128 (O_128,N_9363,N_9486);
and UO_129 (O_129,N_9464,N_9844);
nand UO_130 (O_130,N_9944,N_9914);
nand UO_131 (O_131,N_9980,N_9475);
nor UO_132 (O_132,N_9130,N_9613);
nand UO_133 (O_133,N_9697,N_9062);
and UO_134 (O_134,N_9644,N_9266);
nor UO_135 (O_135,N_9594,N_9576);
nor UO_136 (O_136,N_9603,N_9211);
or UO_137 (O_137,N_9014,N_9948);
nand UO_138 (O_138,N_9421,N_9318);
and UO_139 (O_139,N_9221,N_9931);
nor UO_140 (O_140,N_9187,N_9457);
or UO_141 (O_141,N_9530,N_9047);
nor UO_142 (O_142,N_9748,N_9905);
and UO_143 (O_143,N_9100,N_9396);
and UO_144 (O_144,N_9710,N_9304);
or UO_145 (O_145,N_9049,N_9635);
nor UO_146 (O_146,N_9972,N_9811);
or UO_147 (O_147,N_9843,N_9022);
or UO_148 (O_148,N_9356,N_9027);
nor UO_149 (O_149,N_9460,N_9481);
nand UO_150 (O_150,N_9869,N_9032);
nor UO_151 (O_151,N_9585,N_9010);
nor UO_152 (O_152,N_9437,N_9269);
nor UO_153 (O_153,N_9968,N_9372);
or UO_154 (O_154,N_9769,N_9055);
or UO_155 (O_155,N_9213,N_9046);
and UO_156 (O_156,N_9258,N_9466);
nand UO_157 (O_157,N_9202,N_9279);
nor UO_158 (O_158,N_9533,N_9815);
and UO_159 (O_159,N_9668,N_9006);
nand UO_160 (O_160,N_9707,N_9409);
nor UO_161 (O_161,N_9814,N_9471);
or UO_162 (O_162,N_9527,N_9252);
and UO_163 (O_163,N_9966,N_9127);
and UO_164 (O_164,N_9229,N_9453);
or UO_165 (O_165,N_9836,N_9515);
nor UO_166 (O_166,N_9852,N_9287);
and UO_167 (O_167,N_9597,N_9586);
and UO_168 (O_168,N_9764,N_9902);
nand UO_169 (O_169,N_9219,N_9770);
and UO_170 (O_170,N_9506,N_9775);
or UO_171 (O_171,N_9126,N_9681);
nand UO_172 (O_172,N_9015,N_9434);
nor UO_173 (O_173,N_9050,N_9461);
or UO_174 (O_174,N_9355,N_9979);
and UO_175 (O_175,N_9897,N_9614);
nand UO_176 (O_176,N_9623,N_9975);
and UO_177 (O_177,N_9268,N_9163);
or UO_178 (O_178,N_9598,N_9412);
nand UO_179 (O_179,N_9688,N_9587);
or UO_180 (O_180,N_9013,N_9737);
and UO_181 (O_181,N_9387,N_9289);
and UO_182 (O_182,N_9762,N_9782);
or UO_183 (O_183,N_9534,N_9247);
nand UO_184 (O_184,N_9191,N_9487);
or UO_185 (O_185,N_9362,N_9197);
and UO_186 (O_186,N_9432,N_9670);
nor UO_187 (O_187,N_9458,N_9551);
nand UO_188 (O_188,N_9535,N_9493);
and UO_189 (O_189,N_9491,N_9655);
nor UO_190 (O_190,N_9315,N_9406);
or UO_191 (O_191,N_9484,N_9041);
nor UO_192 (O_192,N_9798,N_9717);
nand UO_193 (O_193,N_9786,N_9847);
or UO_194 (O_194,N_9778,N_9546);
nand UO_195 (O_195,N_9871,N_9570);
and UO_196 (O_196,N_9828,N_9500);
and UO_197 (O_197,N_9164,N_9449);
nand UO_198 (O_198,N_9060,N_9736);
or UO_199 (O_199,N_9654,N_9059);
or UO_200 (O_200,N_9723,N_9729);
nor UO_201 (O_201,N_9956,N_9184);
and UO_202 (O_202,N_9226,N_9599);
nand UO_203 (O_203,N_9780,N_9900);
nand UO_204 (O_204,N_9839,N_9773);
or UO_205 (O_205,N_9650,N_9138);
xnor UO_206 (O_206,N_9606,N_9711);
nor UO_207 (O_207,N_9052,N_9868);
nand UO_208 (O_208,N_9350,N_9926);
and UO_209 (O_209,N_9008,N_9557);
nor UO_210 (O_210,N_9702,N_9933);
or UO_211 (O_211,N_9166,N_9317);
nor UO_212 (O_212,N_9299,N_9125);
and UO_213 (O_213,N_9954,N_9404);
nand UO_214 (O_214,N_9210,N_9101);
or UO_215 (O_215,N_9673,N_9837);
and UO_216 (O_216,N_9273,N_9684);
or UO_217 (O_217,N_9917,N_9018);
nor UO_218 (O_218,N_9067,N_9600);
nor UO_219 (O_219,N_9918,N_9390);
nand UO_220 (O_220,N_9542,N_9333);
nand UO_221 (O_221,N_9946,N_9496);
or UO_222 (O_222,N_9841,N_9007);
nand UO_223 (O_223,N_9177,N_9507);
and UO_224 (O_224,N_9033,N_9391);
nand UO_225 (O_225,N_9338,N_9884);
xor UO_226 (O_226,N_9724,N_9667);
nand UO_227 (O_227,N_9371,N_9292);
and UO_228 (O_228,N_9766,N_9692);
or UO_229 (O_229,N_9698,N_9064);
nor UO_230 (O_230,N_9784,N_9617);
nand UO_231 (O_231,N_9077,N_9147);
nor UO_232 (O_232,N_9230,N_9509);
and UO_233 (O_233,N_9963,N_9321);
or UO_234 (O_234,N_9567,N_9632);
or UO_235 (O_235,N_9114,N_9379);
nand UO_236 (O_236,N_9300,N_9240);
and UO_237 (O_237,N_9524,N_9537);
or UO_238 (O_238,N_9081,N_9809);
nand UO_239 (O_239,N_9403,N_9967);
nor UO_240 (O_240,N_9235,N_9858);
nor UO_241 (O_241,N_9234,N_9030);
nor UO_242 (O_242,N_9098,N_9997);
and UO_243 (O_243,N_9873,N_9703);
nand UO_244 (O_244,N_9561,N_9439);
and UO_245 (O_245,N_9961,N_9959);
or UO_246 (O_246,N_9855,N_9326);
or UO_247 (O_247,N_9992,N_9382);
nor UO_248 (O_248,N_9146,N_9169);
or UO_249 (O_249,N_9383,N_9358);
nand UO_250 (O_250,N_9607,N_9284);
nand UO_251 (O_251,N_9344,N_9020);
nand UO_252 (O_252,N_9349,N_9170);
nand UO_253 (O_253,N_9781,N_9222);
nand UO_254 (O_254,N_9789,N_9669);
nand UO_255 (O_255,N_9653,N_9885);
nand UO_256 (O_256,N_9423,N_9932);
and UO_257 (O_257,N_9339,N_9261);
nand UO_258 (O_258,N_9331,N_9302);
or UO_259 (O_259,N_9121,N_9386);
or UO_260 (O_260,N_9582,N_9357);
or UO_261 (O_261,N_9347,N_9793);
nor UO_262 (O_262,N_9381,N_9410);
nor UO_263 (O_263,N_9366,N_9024);
nor UO_264 (O_264,N_9953,N_9431);
nand UO_265 (O_265,N_9887,N_9563);
and UO_266 (O_266,N_9264,N_9162);
nand UO_267 (O_267,N_9605,N_9592);
nand UO_268 (O_268,N_9610,N_9615);
and UO_269 (O_269,N_9907,N_9091);
nand UO_270 (O_270,N_9250,N_9036);
nand UO_271 (O_271,N_9705,N_9133);
and UO_272 (O_272,N_9817,N_9865);
nand UO_273 (O_273,N_9555,N_9351);
nor UO_274 (O_274,N_9813,N_9611);
and UO_275 (O_275,N_9556,N_9805);
and UO_276 (O_276,N_9549,N_9082);
nand UO_277 (O_277,N_9178,N_9562);
and UO_278 (O_278,N_9452,N_9505);
nand UO_279 (O_279,N_9045,N_9923);
and UO_280 (O_280,N_9271,N_9701);
and UO_281 (O_281,N_9179,N_9820);
nor UO_282 (O_282,N_9513,N_9489);
or UO_283 (O_283,N_9429,N_9407);
or UO_284 (O_284,N_9763,N_9512);
nor UO_285 (O_285,N_9352,N_9012);
or UO_286 (O_286,N_9738,N_9989);
or UO_287 (O_287,N_9426,N_9095);
nor UO_288 (O_288,N_9275,N_9850);
or UO_289 (O_289,N_9477,N_9981);
nor UO_290 (O_290,N_9117,N_9641);
and UO_291 (O_291,N_9661,N_9758);
nand UO_292 (O_292,N_9233,N_9470);
nor UO_293 (O_293,N_9777,N_9947);
nand UO_294 (O_294,N_9529,N_9241);
or UO_295 (O_295,N_9872,N_9768);
or UO_296 (O_296,N_9353,N_9238);
nor UO_297 (O_297,N_9990,N_9680);
and UO_298 (O_298,N_9455,N_9274);
and UO_299 (O_299,N_9343,N_9201);
and UO_300 (O_300,N_9663,N_9671);
nor UO_301 (O_301,N_9704,N_9939);
and UO_302 (O_302,N_9420,N_9054);
nor UO_303 (O_303,N_9772,N_9039);
or UO_304 (O_304,N_9294,N_9411);
or UO_305 (O_305,N_9526,N_9278);
xor UO_306 (O_306,N_9450,N_9153);
nor UO_307 (O_307,N_9291,N_9678);
and UO_308 (O_308,N_9548,N_9753);
nor UO_309 (O_309,N_9693,N_9982);
nand UO_310 (O_310,N_9009,N_9208);
or UO_311 (O_311,N_9312,N_9699);
nand UO_312 (O_312,N_9626,N_9727);
or UO_313 (O_313,N_9886,N_9790);
and UO_314 (O_314,N_9418,N_9435);
and UO_315 (O_315,N_9079,N_9750);
and UO_316 (O_316,N_9853,N_9690);
nor UO_317 (O_317,N_9659,N_9916);
nand UO_318 (O_318,N_9925,N_9190);
or UO_319 (O_319,N_9192,N_9892);
or UO_320 (O_320,N_9936,N_9392);
and UO_321 (O_321,N_9388,N_9259);
nor UO_322 (O_322,N_9519,N_9545);
nor UO_323 (O_323,N_9174,N_9467);
nand UO_324 (O_324,N_9073,N_9298);
and UO_325 (O_325,N_9433,N_9595);
or UO_326 (O_326,N_9182,N_9552);
nor UO_327 (O_327,N_9223,N_9373);
nor UO_328 (O_328,N_9416,N_9706);
or UO_329 (O_329,N_9340,N_9652);
and UO_330 (O_330,N_9845,N_9851);
nand UO_331 (O_331,N_9596,N_9730);
or UO_332 (O_332,N_9921,N_9825);
and UO_333 (O_333,N_9360,N_9958);
and UO_334 (O_334,N_9307,N_9543);
nor UO_335 (O_335,N_9422,N_9591);
or UO_336 (O_336,N_9135,N_9929);
and UO_337 (O_337,N_9324,N_9951);
nor UO_338 (O_338,N_9622,N_9017);
nand UO_339 (O_339,N_9538,N_9109);
and UO_340 (O_340,N_9846,N_9089);
and UO_341 (O_341,N_9171,N_9795);
xnor UO_342 (O_342,N_9807,N_9345);
or UO_343 (O_343,N_9840,N_9774);
or UO_344 (O_344,N_9732,N_9480);
nand UO_345 (O_345,N_9301,N_9492);
nor UO_346 (O_346,N_9942,N_9217);
xnor UO_347 (O_347,N_9742,N_9558);
nor UO_348 (O_348,N_9792,N_9231);
or UO_349 (O_349,N_9128,N_9194);
nor UO_350 (O_350,N_9528,N_9560);
nor UO_351 (O_351,N_9994,N_9239);
or UO_352 (O_352,N_9148,N_9687);
and UO_353 (O_353,N_9521,N_9895);
nor UO_354 (O_354,N_9498,N_9479);
or UO_355 (O_355,N_9142,N_9369);
and UO_356 (O_356,N_9803,N_9080);
nand UO_357 (O_357,N_9297,N_9451);
nand UO_358 (O_358,N_9152,N_9857);
nor UO_359 (O_359,N_9783,N_9718);
nand UO_360 (O_360,N_9485,N_9316);
and UO_361 (O_361,N_9588,N_9236);
nor UO_362 (O_362,N_9124,N_9745);
or UO_363 (O_363,N_9140,N_9149);
and UO_364 (O_364,N_9952,N_9573);
nand UO_365 (O_365,N_9998,N_9314);
nor UO_366 (O_366,N_9195,N_9132);
nor UO_367 (O_367,N_9618,N_9883);
or UO_368 (O_368,N_9826,N_9962);
and UO_369 (O_369,N_9629,N_9810);
nor UO_370 (O_370,N_9903,N_9686);
nor UO_371 (O_371,N_9728,N_9042);
and UO_372 (O_372,N_9621,N_9637);
or UO_373 (O_373,N_9150,N_9044);
and UO_374 (O_374,N_9322,N_9747);
and UO_375 (O_375,N_9665,N_9735);
or UO_376 (O_376,N_9465,N_9071);
nor UO_377 (O_377,N_9894,N_9547);
nand UO_378 (O_378,N_9000,N_9802);
nor UO_379 (O_379,N_9725,N_9145);
nor UO_380 (O_380,N_9501,N_9739);
or UO_381 (O_381,N_9092,N_9832);
nor UO_382 (O_382,N_9478,N_9876);
or UO_383 (O_383,N_9971,N_9937);
and UO_384 (O_384,N_9859,N_9510);
and UO_385 (O_385,N_9108,N_9996);
and UO_386 (O_386,N_9265,N_9327);
nor UO_387 (O_387,N_9206,N_9575);
nand UO_388 (O_388,N_9830,N_9244);
or UO_389 (O_389,N_9577,N_9755);
nor UO_390 (O_390,N_9767,N_9906);
nor UO_391 (O_391,N_9950,N_9816);
nand UO_392 (O_392,N_9969,N_9473);
nor UO_393 (O_393,N_9909,N_9712);
nand UO_394 (O_394,N_9838,N_9541);
or UO_395 (O_395,N_9228,N_9025);
nand UO_396 (O_396,N_9848,N_9720);
nor UO_397 (O_397,N_9232,N_9417);
nand UO_398 (O_398,N_9634,N_9664);
nor UO_399 (O_399,N_9643,N_9168);
or UO_400 (O_400,N_9158,N_9384);
nand UO_401 (O_401,N_9910,N_9165);
or UO_402 (O_402,N_9866,N_9348);
and UO_403 (O_403,N_9332,N_9209);
nor UO_404 (O_404,N_9616,N_9779);
nor UO_405 (O_405,N_9602,N_9263);
or UO_406 (O_406,N_9683,N_9319);
or UO_407 (O_407,N_9313,N_9137);
or UO_408 (O_408,N_9633,N_9590);
or UO_409 (O_409,N_9593,N_9651);
nand UO_410 (O_410,N_9283,N_9048);
nor UO_411 (O_411,N_9249,N_9200);
nor UO_412 (O_412,N_9469,N_9791);
nand UO_413 (O_413,N_9401,N_9286);
or UO_414 (O_414,N_9494,N_9001);
nor UO_415 (O_415,N_9402,N_9173);
and UO_416 (O_416,N_9977,N_9454);
and UO_417 (O_417,N_9380,N_9376);
xor UO_418 (O_418,N_9087,N_9517);
or UO_419 (O_419,N_9003,N_9019);
nand UO_420 (O_420,N_9988,N_9161);
nand UO_421 (O_421,N_9881,N_9395);
nor UO_422 (O_422,N_9086,N_9159);
or UO_423 (O_423,N_9285,N_9808);
and UO_424 (O_424,N_9896,N_9413);
nand UO_425 (O_425,N_9550,N_9026);
or UO_426 (O_426,N_9819,N_9225);
xor UO_427 (O_427,N_9695,N_9731);
and UO_428 (O_428,N_9514,N_9021);
nor UO_429 (O_429,N_9246,N_9214);
or UO_430 (O_430,N_9995,N_9290);
nor UO_431 (O_431,N_9983,N_9218);
nor UO_432 (O_432,N_9499,N_9744);
xor UO_433 (O_433,N_9991,N_9893);
xnor UO_434 (O_434,N_9657,N_9354);
nor UO_435 (O_435,N_9532,N_9675);
or UO_436 (O_436,N_9185,N_9609);
nand UO_437 (O_437,N_9031,N_9305);
xor UO_438 (O_438,N_9927,N_9215);
or UO_439 (O_439,N_9503,N_9296);
nor UO_440 (O_440,N_9272,N_9156);
or UO_441 (O_441,N_9619,N_9399);
nor UO_442 (O_442,N_9620,N_9400);
and UO_443 (O_443,N_9761,N_9063);
or UO_444 (O_444,N_9029,N_9251);
nor UO_445 (O_445,N_9834,N_9999);
and UO_446 (O_446,N_9196,N_9930);
and UO_447 (O_447,N_9920,N_9069);
nand UO_448 (O_448,N_9303,N_9005);
nor UO_449 (O_449,N_9536,N_9205);
nand UO_450 (O_450,N_9154,N_9061);
and UO_451 (O_451,N_9257,N_9564);
nand UO_452 (O_452,N_9901,N_9119);
nor UO_453 (O_453,N_9220,N_9691);
or UO_454 (O_454,N_9722,N_9227);
xnor UO_455 (O_455,N_9139,N_9448);
nand UO_456 (O_456,N_9987,N_9862);
xnor UO_457 (O_457,N_9103,N_9334);
nand UO_458 (O_458,N_9518,N_9441);
nand UO_459 (O_459,N_9076,N_9346);
and UO_460 (O_460,N_9212,N_9488);
or UO_461 (O_461,N_9743,N_9134);
nor UO_462 (O_462,N_9874,N_9428);
nand UO_463 (O_463,N_9740,N_9056);
and UO_464 (O_464,N_9408,N_9833);
nor UO_465 (O_465,N_9444,N_9849);
nand UO_466 (O_466,N_9155,N_9131);
nand UO_467 (O_467,N_9714,N_9604);
and UO_468 (O_468,N_9785,N_9726);
or UO_469 (O_469,N_9445,N_9254);
nor UO_470 (O_470,N_9553,N_9751);
xnor UO_471 (O_471,N_9083,N_9660);
or UO_472 (O_472,N_9601,N_9713);
or UO_473 (O_473,N_9578,N_9336);
nand UO_474 (O_474,N_9102,N_9105);
and UO_475 (O_475,N_9746,N_9964);
and UO_476 (O_476,N_9945,N_9093);
nand UO_477 (O_477,N_9436,N_9370);
nand UO_478 (O_478,N_9090,N_9438);
nand UO_479 (O_479,N_9935,N_9957);
xnor UO_480 (O_480,N_9899,N_9715);
or UO_481 (O_481,N_9342,N_9129);
or UO_482 (O_482,N_9759,N_9474);
nor UO_483 (O_483,N_9068,N_9648);
and UO_484 (O_484,N_9337,N_9111);
nand UO_485 (O_485,N_9398,N_9765);
and UO_486 (O_486,N_9280,N_9757);
nor UO_487 (O_487,N_9583,N_9442);
nand UO_488 (O_488,N_9941,N_9043);
or UO_489 (O_489,N_9040,N_9854);
nand UO_490 (O_490,N_9295,N_9476);
and UO_491 (O_491,N_9378,N_9502);
or UO_492 (O_492,N_9216,N_9574);
or UO_493 (O_493,N_9565,N_9256);
nor UO_494 (O_494,N_9446,N_9472);
or UO_495 (O_495,N_9075,N_9627);
and UO_496 (O_496,N_9113,N_9749);
nand UO_497 (O_497,N_9328,N_9569);
nand UO_498 (O_498,N_9253,N_9002);
nand UO_499 (O_499,N_9540,N_9430);
nand UO_500 (O_500,N_9576,N_9786);
nor UO_501 (O_501,N_9581,N_9489);
and UO_502 (O_502,N_9785,N_9988);
nand UO_503 (O_503,N_9245,N_9839);
nor UO_504 (O_504,N_9735,N_9159);
or UO_505 (O_505,N_9625,N_9027);
and UO_506 (O_506,N_9077,N_9350);
and UO_507 (O_507,N_9719,N_9342);
nand UO_508 (O_508,N_9278,N_9221);
and UO_509 (O_509,N_9612,N_9731);
or UO_510 (O_510,N_9464,N_9338);
xnor UO_511 (O_511,N_9383,N_9077);
nor UO_512 (O_512,N_9757,N_9413);
or UO_513 (O_513,N_9761,N_9615);
nor UO_514 (O_514,N_9187,N_9602);
nand UO_515 (O_515,N_9682,N_9454);
or UO_516 (O_516,N_9015,N_9717);
or UO_517 (O_517,N_9254,N_9862);
or UO_518 (O_518,N_9170,N_9152);
nand UO_519 (O_519,N_9349,N_9459);
nand UO_520 (O_520,N_9780,N_9635);
or UO_521 (O_521,N_9840,N_9198);
nand UO_522 (O_522,N_9116,N_9566);
xnor UO_523 (O_523,N_9126,N_9760);
or UO_524 (O_524,N_9493,N_9064);
or UO_525 (O_525,N_9950,N_9799);
nand UO_526 (O_526,N_9297,N_9520);
nor UO_527 (O_527,N_9476,N_9275);
nand UO_528 (O_528,N_9031,N_9487);
nor UO_529 (O_529,N_9449,N_9136);
nor UO_530 (O_530,N_9060,N_9050);
and UO_531 (O_531,N_9154,N_9962);
and UO_532 (O_532,N_9218,N_9022);
nor UO_533 (O_533,N_9862,N_9509);
nor UO_534 (O_534,N_9712,N_9325);
or UO_535 (O_535,N_9577,N_9397);
or UO_536 (O_536,N_9520,N_9914);
or UO_537 (O_537,N_9400,N_9363);
nand UO_538 (O_538,N_9288,N_9009);
nand UO_539 (O_539,N_9357,N_9954);
or UO_540 (O_540,N_9379,N_9516);
nand UO_541 (O_541,N_9844,N_9858);
nand UO_542 (O_542,N_9597,N_9344);
or UO_543 (O_543,N_9131,N_9200);
or UO_544 (O_544,N_9869,N_9113);
or UO_545 (O_545,N_9023,N_9010);
or UO_546 (O_546,N_9715,N_9319);
nand UO_547 (O_547,N_9734,N_9601);
and UO_548 (O_548,N_9705,N_9377);
nor UO_549 (O_549,N_9265,N_9869);
and UO_550 (O_550,N_9363,N_9882);
nor UO_551 (O_551,N_9078,N_9644);
nor UO_552 (O_552,N_9160,N_9292);
nand UO_553 (O_553,N_9651,N_9444);
and UO_554 (O_554,N_9473,N_9793);
or UO_555 (O_555,N_9066,N_9428);
xor UO_556 (O_556,N_9446,N_9966);
nor UO_557 (O_557,N_9759,N_9276);
nand UO_558 (O_558,N_9822,N_9042);
nand UO_559 (O_559,N_9137,N_9309);
and UO_560 (O_560,N_9498,N_9478);
nand UO_561 (O_561,N_9627,N_9496);
and UO_562 (O_562,N_9985,N_9590);
and UO_563 (O_563,N_9900,N_9646);
and UO_564 (O_564,N_9968,N_9453);
or UO_565 (O_565,N_9031,N_9028);
and UO_566 (O_566,N_9648,N_9167);
xnor UO_567 (O_567,N_9202,N_9081);
or UO_568 (O_568,N_9105,N_9871);
nor UO_569 (O_569,N_9322,N_9637);
nand UO_570 (O_570,N_9548,N_9914);
nand UO_571 (O_571,N_9862,N_9858);
and UO_572 (O_572,N_9418,N_9224);
or UO_573 (O_573,N_9258,N_9817);
nor UO_574 (O_574,N_9801,N_9537);
nand UO_575 (O_575,N_9287,N_9203);
or UO_576 (O_576,N_9915,N_9613);
nor UO_577 (O_577,N_9626,N_9919);
and UO_578 (O_578,N_9081,N_9448);
and UO_579 (O_579,N_9481,N_9416);
and UO_580 (O_580,N_9805,N_9812);
and UO_581 (O_581,N_9033,N_9894);
and UO_582 (O_582,N_9970,N_9775);
nand UO_583 (O_583,N_9256,N_9822);
or UO_584 (O_584,N_9780,N_9319);
nand UO_585 (O_585,N_9897,N_9888);
nor UO_586 (O_586,N_9187,N_9550);
nand UO_587 (O_587,N_9020,N_9949);
xor UO_588 (O_588,N_9242,N_9883);
and UO_589 (O_589,N_9914,N_9329);
and UO_590 (O_590,N_9877,N_9339);
and UO_591 (O_591,N_9630,N_9439);
xnor UO_592 (O_592,N_9618,N_9895);
and UO_593 (O_593,N_9671,N_9232);
and UO_594 (O_594,N_9084,N_9540);
nand UO_595 (O_595,N_9558,N_9571);
nor UO_596 (O_596,N_9664,N_9707);
xor UO_597 (O_597,N_9097,N_9386);
or UO_598 (O_598,N_9232,N_9602);
or UO_599 (O_599,N_9574,N_9914);
and UO_600 (O_600,N_9461,N_9588);
nand UO_601 (O_601,N_9654,N_9736);
nand UO_602 (O_602,N_9294,N_9361);
nand UO_603 (O_603,N_9815,N_9505);
and UO_604 (O_604,N_9352,N_9055);
or UO_605 (O_605,N_9971,N_9187);
and UO_606 (O_606,N_9478,N_9255);
and UO_607 (O_607,N_9983,N_9862);
or UO_608 (O_608,N_9203,N_9321);
and UO_609 (O_609,N_9355,N_9930);
nor UO_610 (O_610,N_9846,N_9555);
or UO_611 (O_611,N_9698,N_9995);
nor UO_612 (O_612,N_9775,N_9046);
or UO_613 (O_613,N_9249,N_9326);
nand UO_614 (O_614,N_9783,N_9114);
nand UO_615 (O_615,N_9608,N_9747);
and UO_616 (O_616,N_9044,N_9694);
and UO_617 (O_617,N_9647,N_9579);
and UO_618 (O_618,N_9107,N_9917);
nor UO_619 (O_619,N_9494,N_9416);
nor UO_620 (O_620,N_9247,N_9451);
nand UO_621 (O_621,N_9445,N_9011);
or UO_622 (O_622,N_9288,N_9557);
nand UO_623 (O_623,N_9450,N_9364);
nand UO_624 (O_624,N_9030,N_9721);
nor UO_625 (O_625,N_9582,N_9024);
nor UO_626 (O_626,N_9062,N_9080);
and UO_627 (O_627,N_9663,N_9245);
or UO_628 (O_628,N_9694,N_9025);
and UO_629 (O_629,N_9550,N_9571);
and UO_630 (O_630,N_9290,N_9164);
nand UO_631 (O_631,N_9027,N_9568);
or UO_632 (O_632,N_9270,N_9979);
nand UO_633 (O_633,N_9170,N_9419);
nand UO_634 (O_634,N_9730,N_9440);
nand UO_635 (O_635,N_9179,N_9277);
and UO_636 (O_636,N_9208,N_9462);
or UO_637 (O_637,N_9419,N_9322);
xnor UO_638 (O_638,N_9231,N_9492);
and UO_639 (O_639,N_9540,N_9528);
and UO_640 (O_640,N_9308,N_9063);
or UO_641 (O_641,N_9806,N_9932);
nand UO_642 (O_642,N_9416,N_9949);
and UO_643 (O_643,N_9817,N_9410);
nand UO_644 (O_644,N_9340,N_9709);
or UO_645 (O_645,N_9881,N_9434);
nand UO_646 (O_646,N_9096,N_9995);
or UO_647 (O_647,N_9467,N_9551);
nand UO_648 (O_648,N_9406,N_9954);
and UO_649 (O_649,N_9476,N_9112);
or UO_650 (O_650,N_9306,N_9988);
nand UO_651 (O_651,N_9988,N_9680);
nor UO_652 (O_652,N_9263,N_9907);
nor UO_653 (O_653,N_9159,N_9464);
nor UO_654 (O_654,N_9939,N_9398);
xnor UO_655 (O_655,N_9060,N_9973);
nor UO_656 (O_656,N_9570,N_9462);
nor UO_657 (O_657,N_9254,N_9407);
nor UO_658 (O_658,N_9598,N_9468);
xnor UO_659 (O_659,N_9129,N_9943);
nor UO_660 (O_660,N_9453,N_9276);
nand UO_661 (O_661,N_9274,N_9661);
or UO_662 (O_662,N_9841,N_9770);
nor UO_663 (O_663,N_9632,N_9865);
and UO_664 (O_664,N_9028,N_9981);
or UO_665 (O_665,N_9376,N_9350);
nor UO_666 (O_666,N_9858,N_9576);
or UO_667 (O_667,N_9703,N_9383);
nor UO_668 (O_668,N_9955,N_9440);
or UO_669 (O_669,N_9666,N_9231);
or UO_670 (O_670,N_9347,N_9753);
nor UO_671 (O_671,N_9478,N_9487);
nand UO_672 (O_672,N_9460,N_9874);
and UO_673 (O_673,N_9889,N_9038);
or UO_674 (O_674,N_9233,N_9090);
and UO_675 (O_675,N_9184,N_9663);
nand UO_676 (O_676,N_9836,N_9252);
nand UO_677 (O_677,N_9170,N_9377);
and UO_678 (O_678,N_9962,N_9477);
nand UO_679 (O_679,N_9344,N_9719);
and UO_680 (O_680,N_9704,N_9586);
nand UO_681 (O_681,N_9003,N_9436);
or UO_682 (O_682,N_9630,N_9398);
or UO_683 (O_683,N_9684,N_9193);
or UO_684 (O_684,N_9217,N_9926);
nor UO_685 (O_685,N_9933,N_9865);
nor UO_686 (O_686,N_9837,N_9235);
and UO_687 (O_687,N_9475,N_9175);
and UO_688 (O_688,N_9172,N_9610);
and UO_689 (O_689,N_9083,N_9872);
xor UO_690 (O_690,N_9296,N_9769);
nand UO_691 (O_691,N_9157,N_9688);
and UO_692 (O_692,N_9110,N_9608);
or UO_693 (O_693,N_9499,N_9375);
and UO_694 (O_694,N_9556,N_9036);
nor UO_695 (O_695,N_9120,N_9218);
and UO_696 (O_696,N_9670,N_9127);
xnor UO_697 (O_697,N_9057,N_9738);
xnor UO_698 (O_698,N_9831,N_9496);
nor UO_699 (O_699,N_9009,N_9602);
and UO_700 (O_700,N_9324,N_9731);
nand UO_701 (O_701,N_9442,N_9060);
and UO_702 (O_702,N_9170,N_9011);
nor UO_703 (O_703,N_9286,N_9714);
nand UO_704 (O_704,N_9957,N_9522);
and UO_705 (O_705,N_9434,N_9489);
and UO_706 (O_706,N_9063,N_9642);
and UO_707 (O_707,N_9194,N_9743);
nand UO_708 (O_708,N_9955,N_9050);
or UO_709 (O_709,N_9931,N_9968);
nor UO_710 (O_710,N_9392,N_9940);
nand UO_711 (O_711,N_9929,N_9571);
or UO_712 (O_712,N_9414,N_9272);
or UO_713 (O_713,N_9532,N_9365);
nand UO_714 (O_714,N_9670,N_9964);
nor UO_715 (O_715,N_9432,N_9387);
nor UO_716 (O_716,N_9435,N_9233);
nor UO_717 (O_717,N_9143,N_9386);
nand UO_718 (O_718,N_9514,N_9546);
nor UO_719 (O_719,N_9674,N_9822);
and UO_720 (O_720,N_9455,N_9361);
and UO_721 (O_721,N_9037,N_9544);
nor UO_722 (O_722,N_9390,N_9597);
nor UO_723 (O_723,N_9175,N_9371);
or UO_724 (O_724,N_9256,N_9121);
and UO_725 (O_725,N_9246,N_9135);
nor UO_726 (O_726,N_9712,N_9358);
and UO_727 (O_727,N_9128,N_9541);
nand UO_728 (O_728,N_9557,N_9884);
nor UO_729 (O_729,N_9169,N_9232);
nor UO_730 (O_730,N_9354,N_9633);
and UO_731 (O_731,N_9934,N_9014);
or UO_732 (O_732,N_9306,N_9520);
nor UO_733 (O_733,N_9872,N_9713);
and UO_734 (O_734,N_9427,N_9042);
nand UO_735 (O_735,N_9720,N_9377);
nor UO_736 (O_736,N_9976,N_9022);
and UO_737 (O_737,N_9885,N_9919);
and UO_738 (O_738,N_9245,N_9872);
nor UO_739 (O_739,N_9543,N_9082);
and UO_740 (O_740,N_9935,N_9164);
nand UO_741 (O_741,N_9953,N_9248);
nor UO_742 (O_742,N_9670,N_9717);
or UO_743 (O_743,N_9687,N_9037);
and UO_744 (O_744,N_9979,N_9047);
and UO_745 (O_745,N_9720,N_9009);
and UO_746 (O_746,N_9494,N_9376);
nor UO_747 (O_747,N_9116,N_9892);
and UO_748 (O_748,N_9981,N_9492);
nor UO_749 (O_749,N_9012,N_9077);
nand UO_750 (O_750,N_9817,N_9092);
nor UO_751 (O_751,N_9178,N_9154);
or UO_752 (O_752,N_9299,N_9008);
nand UO_753 (O_753,N_9071,N_9652);
nand UO_754 (O_754,N_9306,N_9419);
and UO_755 (O_755,N_9301,N_9620);
nor UO_756 (O_756,N_9230,N_9536);
or UO_757 (O_757,N_9412,N_9681);
nor UO_758 (O_758,N_9294,N_9210);
or UO_759 (O_759,N_9030,N_9589);
or UO_760 (O_760,N_9773,N_9081);
and UO_761 (O_761,N_9918,N_9865);
or UO_762 (O_762,N_9253,N_9381);
and UO_763 (O_763,N_9182,N_9115);
and UO_764 (O_764,N_9043,N_9002);
nand UO_765 (O_765,N_9036,N_9989);
nand UO_766 (O_766,N_9391,N_9404);
and UO_767 (O_767,N_9568,N_9316);
or UO_768 (O_768,N_9536,N_9544);
nand UO_769 (O_769,N_9574,N_9718);
nor UO_770 (O_770,N_9519,N_9851);
nand UO_771 (O_771,N_9943,N_9224);
nor UO_772 (O_772,N_9223,N_9581);
and UO_773 (O_773,N_9731,N_9208);
or UO_774 (O_774,N_9923,N_9472);
and UO_775 (O_775,N_9161,N_9317);
or UO_776 (O_776,N_9615,N_9011);
and UO_777 (O_777,N_9634,N_9462);
nand UO_778 (O_778,N_9085,N_9765);
or UO_779 (O_779,N_9356,N_9758);
and UO_780 (O_780,N_9740,N_9070);
or UO_781 (O_781,N_9543,N_9645);
nor UO_782 (O_782,N_9623,N_9238);
or UO_783 (O_783,N_9834,N_9734);
or UO_784 (O_784,N_9601,N_9850);
or UO_785 (O_785,N_9304,N_9888);
nand UO_786 (O_786,N_9200,N_9762);
or UO_787 (O_787,N_9417,N_9043);
and UO_788 (O_788,N_9342,N_9179);
nor UO_789 (O_789,N_9488,N_9497);
nor UO_790 (O_790,N_9680,N_9861);
and UO_791 (O_791,N_9309,N_9936);
or UO_792 (O_792,N_9189,N_9284);
and UO_793 (O_793,N_9551,N_9131);
nand UO_794 (O_794,N_9889,N_9981);
nor UO_795 (O_795,N_9823,N_9843);
or UO_796 (O_796,N_9625,N_9191);
and UO_797 (O_797,N_9238,N_9732);
and UO_798 (O_798,N_9884,N_9803);
nor UO_799 (O_799,N_9725,N_9885);
nor UO_800 (O_800,N_9907,N_9933);
nand UO_801 (O_801,N_9793,N_9949);
nand UO_802 (O_802,N_9520,N_9955);
nand UO_803 (O_803,N_9077,N_9888);
xnor UO_804 (O_804,N_9010,N_9695);
or UO_805 (O_805,N_9130,N_9535);
and UO_806 (O_806,N_9891,N_9694);
and UO_807 (O_807,N_9964,N_9848);
nor UO_808 (O_808,N_9623,N_9239);
nor UO_809 (O_809,N_9860,N_9728);
and UO_810 (O_810,N_9648,N_9296);
xnor UO_811 (O_811,N_9413,N_9242);
and UO_812 (O_812,N_9322,N_9672);
or UO_813 (O_813,N_9796,N_9002);
nor UO_814 (O_814,N_9726,N_9940);
or UO_815 (O_815,N_9081,N_9799);
and UO_816 (O_816,N_9270,N_9258);
nand UO_817 (O_817,N_9965,N_9131);
and UO_818 (O_818,N_9175,N_9471);
nand UO_819 (O_819,N_9805,N_9694);
nand UO_820 (O_820,N_9130,N_9310);
or UO_821 (O_821,N_9547,N_9615);
nor UO_822 (O_822,N_9389,N_9735);
or UO_823 (O_823,N_9620,N_9359);
or UO_824 (O_824,N_9106,N_9305);
nand UO_825 (O_825,N_9732,N_9596);
xor UO_826 (O_826,N_9787,N_9693);
or UO_827 (O_827,N_9872,N_9215);
nor UO_828 (O_828,N_9796,N_9967);
nor UO_829 (O_829,N_9053,N_9580);
nand UO_830 (O_830,N_9383,N_9472);
nand UO_831 (O_831,N_9719,N_9358);
or UO_832 (O_832,N_9042,N_9178);
or UO_833 (O_833,N_9620,N_9826);
or UO_834 (O_834,N_9168,N_9981);
nand UO_835 (O_835,N_9872,N_9124);
nand UO_836 (O_836,N_9959,N_9499);
nor UO_837 (O_837,N_9193,N_9209);
or UO_838 (O_838,N_9867,N_9318);
nand UO_839 (O_839,N_9546,N_9916);
nor UO_840 (O_840,N_9772,N_9319);
nor UO_841 (O_841,N_9689,N_9084);
and UO_842 (O_842,N_9389,N_9321);
or UO_843 (O_843,N_9258,N_9568);
and UO_844 (O_844,N_9723,N_9772);
and UO_845 (O_845,N_9568,N_9911);
nor UO_846 (O_846,N_9545,N_9860);
and UO_847 (O_847,N_9546,N_9019);
and UO_848 (O_848,N_9428,N_9909);
or UO_849 (O_849,N_9269,N_9110);
or UO_850 (O_850,N_9699,N_9891);
nor UO_851 (O_851,N_9678,N_9297);
nand UO_852 (O_852,N_9991,N_9007);
or UO_853 (O_853,N_9832,N_9353);
nor UO_854 (O_854,N_9889,N_9508);
nand UO_855 (O_855,N_9007,N_9981);
and UO_856 (O_856,N_9719,N_9946);
nand UO_857 (O_857,N_9335,N_9117);
and UO_858 (O_858,N_9822,N_9547);
and UO_859 (O_859,N_9562,N_9946);
and UO_860 (O_860,N_9821,N_9745);
nand UO_861 (O_861,N_9479,N_9202);
nand UO_862 (O_862,N_9072,N_9659);
or UO_863 (O_863,N_9490,N_9867);
nand UO_864 (O_864,N_9789,N_9907);
nand UO_865 (O_865,N_9504,N_9316);
and UO_866 (O_866,N_9853,N_9599);
or UO_867 (O_867,N_9914,N_9543);
nor UO_868 (O_868,N_9766,N_9902);
or UO_869 (O_869,N_9709,N_9553);
xnor UO_870 (O_870,N_9276,N_9943);
and UO_871 (O_871,N_9363,N_9039);
nand UO_872 (O_872,N_9972,N_9470);
and UO_873 (O_873,N_9283,N_9752);
nor UO_874 (O_874,N_9136,N_9290);
or UO_875 (O_875,N_9324,N_9855);
and UO_876 (O_876,N_9274,N_9736);
nor UO_877 (O_877,N_9657,N_9348);
or UO_878 (O_878,N_9721,N_9870);
and UO_879 (O_879,N_9774,N_9913);
nor UO_880 (O_880,N_9112,N_9513);
nand UO_881 (O_881,N_9682,N_9688);
nand UO_882 (O_882,N_9205,N_9584);
nand UO_883 (O_883,N_9038,N_9476);
nor UO_884 (O_884,N_9576,N_9305);
nor UO_885 (O_885,N_9336,N_9016);
and UO_886 (O_886,N_9454,N_9013);
nand UO_887 (O_887,N_9908,N_9147);
nand UO_888 (O_888,N_9611,N_9366);
nor UO_889 (O_889,N_9213,N_9540);
or UO_890 (O_890,N_9880,N_9993);
nor UO_891 (O_891,N_9086,N_9962);
xor UO_892 (O_892,N_9851,N_9460);
xnor UO_893 (O_893,N_9102,N_9087);
nand UO_894 (O_894,N_9123,N_9858);
or UO_895 (O_895,N_9110,N_9831);
nor UO_896 (O_896,N_9088,N_9818);
and UO_897 (O_897,N_9802,N_9442);
nor UO_898 (O_898,N_9721,N_9136);
or UO_899 (O_899,N_9870,N_9427);
nor UO_900 (O_900,N_9438,N_9080);
and UO_901 (O_901,N_9438,N_9756);
nand UO_902 (O_902,N_9190,N_9429);
and UO_903 (O_903,N_9346,N_9722);
or UO_904 (O_904,N_9762,N_9218);
nor UO_905 (O_905,N_9701,N_9284);
nand UO_906 (O_906,N_9142,N_9505);
or UO_907 (O_907,N_9005,N_9797);
or UO_908 (O_908,N_9555,N_9721);
and UO_909 (O_909,N_9360,N_9303);
or UO_910 (O_910,N_9481,N_9940);
and UO_911 (O_911,N_9168,N_9708);
and UO_912 (O_912,N_9221,N_9656);
nand UO_913 (O_913,N_9713,N_9848);
or UO_914 (O_914,N_9539,N_9840);
and UO_915 (O_915,N_9561,N_9759);
nand UO_916 (O_916,N_9226,N_9360);
and UO_917 (O_917,N_9429,N_9629);
and UO_918 (O_918,N_9630,N_9018);
nor UO_919 (O_919,N_9536,N_9400);
nor UO_920 (O_920,N_9032,N_9640);
and UO_921 (O_921,N_9377,N_9392);
nor UO_922 (O_922,N_9787,N_9803);
or UO_923 (O_923,N_9966,N_9499);
or UO_924 (O_924,N_9775,N_9412);
and UO_925 (O_925,N_9415,N_9729);
and UO_926 (O_926,N_9022,N_9784);
and UO_927 (O_927,N_9186,N_9703);
nor UO_928 (O_928,N_9867,N_9755);
and UO_929 (O_929,N_9890,N_9374);
nand UO_930 (O_930,N_9147,N_9742);
nor UO_931 (O_931,N_9604,N_9879);
and UO_932 (O_932,N_9818,N_9168);
nand UO_933 (O_933,N_9212,N_9531);
nand UO_934 (O_934,N_9226,N_9618);
or UO_935 (O_935,N_9655,N_9451);
and UO_936 (O_936,N_9657,N_9166);
nor UO_937 (O_937,N_9116,N_9769);
and UO_938 (O_938,N_9329,N_9067);
nand UO_939 (O_939,N_9425,N_9074);
nand UO_940 (O_940,N_9364,N_9896);
or UO_941 (O_941,N_9919,N_9177);
or UO_942 (O_942,N_9166,N_9288);
or UO_943 (O_943,N_9595,N_9221);
and UO_944 (O_944,N_9144,N_9499);
or UO_945 (O_945,N_9485,N_9528);
or UO_946 (O_946,N_9037,N_9661);
nor UO_947 (O_947,N_9591,N_9875);
and UO_948 (O_948,N_9372,N_9062);
or UO_949 (O_949,N_9032,N_9407);
or UO_950 (O_950,N_9867,N_9074);
nor UO_951 (O_951,N_9241,N_9963);
nand UO_952 (O_952,N_9492,N_9787);
or UO_953 (O_953,N_9301,N_9002);
nand UO_954 (O_954,N_9509,N_9628);
xor UO_955 (O_955,N_9417,N_9559);
nand UO_956 (O_956,N_9695,N_9245);
and UO_957 (O_957,N_9050,N_9185);
or UO_958 (O_958,N_9984,N_9968);
nand UO_959 (O_959,N_9862,N_9612);
nor UO_960 (O_960,N_9689,N_9694);
and UO_961 (O_961,N_9711,N_9187);
nand UO_962 (O_962,N_9463,N_9102);
or UO_963 (O_963,N_9038,N_9126);
nor UO_964 (O_964,N_9508,N_9853);
nor UO_965 (O_965,N_9534,N_9935);
nor UO_966 (O_966,N_9309,N_9926);
nand UO_967 (O_967,N_9394,N_9268);
nor UO_968 (O_968,N_9023,N_9759);
nor UO_969 (O_969,N_9589,N_9063);
and UO_970 (O_970,N_9784,N_9196);
and UO_971 (O_971,N_9114,N_9776);
and UO_972 (O_972,N_9986,N_9707);
nor UO_973 (O_973,N_9446,N_9492);
nand UO_974 (O_974,N_9179,N_9520);
or UO_975 (O_975,N_9241,N_9032);
nand UO_976 (O_976,N_9468,N_9325);
and UO_977 (O_977,N_9055,N_9419);
or UO_978 (O_978,N_9834,N_9560);
nor UO_979 (O_979,N_9792,N_9373);
nand UO_980 (O_980,N_9748,N_9713);
nand UO_981 (O_981,N_9942,N_9888);
nand UO_982 (O_982,N_9406,N_9916);
or UO_983 (O_983,N_9616,N_9483);
nand UO_984 (O_984,N_9785,N_9235);
and UO_985 (O_985,N_9071,N_9833);
or UO_986 (O_986,N_9108,N_9844);
nor UO_987 (O_987,N_9228,N_9918);
nand UO_988 (O_988,N_9495,N_9583);
nor UO_989 (O_989,N_9495,N_9659);
or UO_990 (O_990,N_9042,N_9729);
and UO_991 (O_991,N_9875,N_9577);
and UO_992 (O_992,N_9981,N_9706);
nand UO_993 (O_993,N_9447,N_9101);
or UO_994 (O_994,N_9956,N_9046);
or UO_995 (O_995,N_9646,N_9664);
nand UO_996 (O_996,N_9773,N_9971);
and UO_997 (O_997,N_9630,N_9135);
nor UO_998 (O_998,N_9861,N_9353);
or UO_999 (O_999,N_9055,N_9705);
nand UO_1000 (O_1000,N_9135,N_9389);
and UO_1001 (O_1001,N_9557,N_9236);
nand UO_1002 (O_1002,N_9610,N_9707);
and UO_1003 (O_1003,N_9915,N_9068);
nor UO_1004 (O_1004,N_9997,N_9651);
and UO_1005 (O_1005,N_9350,N_9550);
and UO_1006 (O_1006,N_9441,N_9371);
or UO_1007 (O_1007,N_9749,N_9336);
nand UO_1008 (O_1008,N_9280,N_9943);
or UO_1009 (O_1009,N_9407,N_9803);
nor UO_1010 (O_1010,N_9662,N_9928);
nand UO_1011 (O_1011,N_9805,N_9428);
and UO_1012 (O_1012,N_9665,N_9492);
and UO_1013 (O_1013,N_9155,N_9997);
or UO_1014 (O_1014,N_9401,N_9810);
nand UO_1015 (O_1015,N_9373,N_9168);
and UO_1016 (O_1016,N_9366,N_9640);
nor UO_1017 (O_1017,N_9868,N_9505);
nor UO_1018 (O_1018,N_9373,N_9875);
and UO_1019 (O_1019,N_9153,N_9295);
nor UO_1020 (O_1020,N_9357,N_9808);
or UO_1021 (O_1021,N_9279,N_9713);
nor UO_1022 (O_1022,N_9012,N_9153);
nand UO_1023 (O_1023,N_9813,N_9362);
and UO_1024 (O_1024,N_9786,N_9946);
or UO_1025 (O_1025,N_9485,N_9129);
or UO_1026 (O_1026,N_9921,N_9420);
or UO_1027 (O_1027,N_9325,N_9347);
or UO_1028 (O_1028,N_9358,N_9359);
nor UO_1029 (O_1029,N_9122,N_9186);
and UO_1030 (O_1030,N_9874,N_9205);
nor UO_1031 (O_1031,N_9460,N_9132);
or UO_1032 (O_1032,N_9085,N_9928);
nor UO_1033 (O_1033,N_9326,N_9717);
and UO_1034 (O_1034,N_9319,N_9110);
xor UO_1035 (O_1035,N_9670,N_9603);
or UO_1036 (O_1036,N_9987,N_9713);
and UO_1037 (O_1037,N_9792,N_9168);
or UO_1038 (O_1038,N_9810,N_9682);
nor UO_1039 (O_1039,N_9534,N_9952);
nor UO_1040 (O_1040,N_9016,N_9949);
and UO_1041 (O_1041,N_9863,N_9340);
nor UO_1042 (O_1042,N_9843,N_9160);
and UO_1043 (O_1043,N_9464,N_9626);
or UO_1044 (O_1044,N_9288,N_9418);
nand UO_1045 (O_1045,N_9411,N_9018);
or UO_1046 (O_1046,N_9930,N_9971);
or UO_1047 (O_1047,N_9992,N_9773);
nor UO_1048 (O_1048,N_9203,N_9882);
or UO_1049 (O_1049,N_9656,N_9231);
or UO_1050 (O_1050,N_9271,N_9861);
nand UO_1051 (O_1051,N_9777,N_9976);
or UO_1052 (O_1052,N_9786,N_9267);
nand UO_1053 (O_1053,N_9612,N_9660);
and UO_1054 (O_1054,N_9066,N_9319);
nand UO_1055 (O_1055,N_9391,N_9760);
and UO_1056 (O_1056,N_9671,N_9393);
nor UO_1057 (O_1057,N_9656,N_9303);
and UO_1058 (O_1058,N_9529,N_9256);
nand UO_1059 (O_1059,N_9148,N_9498);
nand UO_1060 (O_1060,N_9012,N_9687);
nand UO_1061 (O_1061,N_9434,N_9282);
and UO_1062 (O_1062,N_9636,N_9815);
or UO_1063 (O_1063,N_9263,N_9509);
nand UO_1064 (O_1064,N_9398,N_9884);
nand UO_1065 (O_1065,N_9870,N_9744);
nor UO_1066 (O_1066,N_9279,N_9753);
nand UO_1067 (O_1067,N_9530,N_9478);
nor UO_1068 (O_1068,N_9396,N_9469);
and UO_1069 (O_1069,N_9983,N_9617);
nor UO_1070 (O_1070,N_9596,N_9854);
or UO_1071 (O_1071,N_9027,N_9687);
nand UO_1072 (O_1072,N_9368,N_9025);
nand UO_1073 (O_1073,N_9979,N_9104);
nor UO_1074 (O_1074,N_9107,N_9763);
or UO_1075 (O_1075,N_9262,N_9723);
nand UO_1076 (O_1076,N_9138,N_9695);
and UO_1077 (O_1077,N_9938,N_9130);
nor UO_1078 (O_1078,N_9184,N_9415);
and UO_1079 (O_1079,N_9422,N_9998);
nand UO_1080 (O_1080,N_9008,N_9949);
nor UO_1081 (O_1081,N_9432,N_9433);
nand UO_1082 (O_1082,N_9882,N_9916);
nand UO_1083 (O_1083,N_9781,N_9180);
nor UO_1084 (O_1084,N_9841,N_9743);
nor UO_1085 (O_1085,N_9230,N_9319);
and UO_1086 (O_1086,N_9148,N_9285);
nor UO_1087 (O_1087,N_9937,N_9263);
or UO_1088 (O_1088,N_9584,N_9694);
nand UO_1089 (O_1089,N_9175,N_9691);
nand UO_1090 (O_1090,N_9742,N_9428);
nor UO_1091 (O_1091,N_9106,N_9516);
or UO_1092 (O_1092,N_9567,N_9621);
or UO_1093 (O_1093,N_9742,N_9881);
xnor UO_1094 (O_1094,N_9538,N_9358);
or UO_1095 (O_1095,N_9653,N_9537);
or UO_1096 (O_1096,N_9863,N_9431);
nor UO_1097 (O_1097,N_9332,N_9166);
and UO_1098 (O_1098,N_9326,N_9095);
and UO_1099 (O_1099,N_9353,N_9199);
xnor UO_1100 (O_1100,N_9420,N_9357);
nand UO_1101 (O_1101,N_9410,N_9578);
nand UO_1102 (O_1102,N_9339,N_9495);
nor UO_1103 (O_1103,N_9043,N_9311);
nand UO_1104 (O_1104,N_9509,N_9535);
nand UO_1105 (O_1105,N_9189,N_9628);
or UO_1106 (O_1106,N_9174,N_9213);
nand UO_1107 (O_1107,N_9135,N_9750);
or UO_1108 (O_1108,N_9176,N_9612);
xnor UO_1109 (O_1109,N_9499,N_9456);
nand UO_1110 (O_1110,N_9146,N_9626);
or UO_1111 (O_1111,N_9539,N_9640);
or UO_1112 (O_1112,N_9964,N_9235);
nand UO_1113 (O_1113,N_9727,N_9072);
and UO_1114 (O_1114,N_9799,N_9520);
or UO_1115 (O_1115,N_9810,N_9817);
nand UO_1116 (O_1116,N_9384,N_9025);
or UO_1117 (O_1117,N_9410,N_9150);
nor UO_1118 (O_1118,N_9042,N_9845);
and UO_1119 (O_1119,N_9623,N_9424);
or UO_1120 (O_1120,N_9258,N_9609);
and UO_1121 (O_1121,N_9391,N_9683);
nor UO_1122 (O_1122,N_9094,N_9118);
nand UO_1123 (O_1123,N_9929,N_9277);
and UO_1124 (O_1124,N_9444,N_9367);
and UO_1125 (O_1125,N_9168,N_9705);
nand UO_1126 (O_1126,N_9751,N_9107);
nand UO_1127 (O_1127,N_9737,N_9606);
or UO_1128 (O_1128,N_9697,N_9347);
or UO_1129 (O_1129,N_9931,N_9569);
nand UO_1130 (O_1130,N_9297,N_9595);
xor UO_1131 (O_1131,N_9985,N_9332);
nand UO_1132 (O_1132,N_9758,N_9421);
nor UO_1133 (O_1133,N_9871,N_9347);
and UO_1134 (O_1134,N_9093,N_9191);
or UO_1135 (O_1135,N_9579,N_9633);
and UO_1136 (O_1136,N_9652,N_9680);
or UO_1137 (O_1137,N_9922,N_9473);
nand UO_1138 (O_1138,N_9433,N_9405);
or UO_1139 (O_1139,N_9387,N_9368);
and UO_1140 (O_1140,N_9002,N_9423);
and UO_1141 (O_1141,N_9075,N_9470);
or UO_1142 (O_1142,N_9565,N_9659);
nand UO_1143 (O_1143,N_9351,N_9382);
and UO_1144 (O_1144,N_9321,N_9164);
nor UO_1145 (O_1145,N_9884,N_9253);
nand UO_1146 (O_1146,N_9635,N_9722);
nor UO_1147 (O_1147,N_9117,N_9415);
and UO_1148 (O_1148,N_9021,N_9306);
nand UO_1149 (O_1149,N_9628,N_9691);
and UO_1150 (O_1150,N_9888,N_9489);
or UO_1151 (O_1151,N_9606,N_9267);
nor UO_1152 (O_1152,N_9246,N_9534);
nand UO_1153 (O_1153,N_9167,N_9599);
and UO_1154 (O_1154,N_9672,N_9410);
or UO_1155 (O_1155,N_9849,N_9501);
or UO_1156 (O_1156,N_9068,N_9266);
or UO_1157 (O_1157,N_9486,N_9237);
xnor UO_1158 (O_1158,N_9866,N_9500);
nand UO_1159 (O_1159,N_9423,N_9823);
and UO_1160 (O_1160,N_9184,N_9570);
nand UO_1161 (O_1161,N_9473,N_9666);
xnor UO_1162 (O_1162,N_9127,N_9280);
nor UO_1163 (O_1163,N_9476,N_9747);
nor UO_1164 (O_1164,N_9558,N_9953);
and UO_1165 (O_1165,N_9912,N_9110);
or UO_1166 (O_1166,N_9318,N_9216);
nand UO_1167 (O_1167,N_9335,N_9329);
or UO_1168 (O_1168,N_9780,N_9497);
and UO_1169 (O_1169,N_9236,N_9579);
xnor UO_1170 (O_1170,N_9274,N_9758);
nand UO_1171 (O_1171,N_9977,N_9641);
and UO_1172 (O_1172,N_9666,N_9642);
nor UO_1173 (O_1173,N_9140,N_9399);
and UO_1174 (O_1174,N_9307,N_9970);
and UO_1175 (O_1175,N_9298,N_9496);
nor UO_1176 (O_1176,N_9282,N_9854);
nand UO_1177 (O_1177,N_9785,N_9532);
and UO_1178 (O_1178,N_9996,N_9038);
and UO_1179 (O_1179,N_9027,N_9008);
and UO_1180 (O_1180,N_9312,N_9053);
nor UO_1181 (O_1181,N_9865,N_9980);
nand UO_1182 (O_1182,N_9530,N_9624);
and UO_1183 (O_1183,N_9458,N_9329);
nor UO_1184 (O_1184,N_9482,N_9640);
nand UO_1185 (O_1185,N_9965,N_9193);
or UO_1186 (O_1186,N_9769,N_9364);
or UO_1187 (O_1187,N_9392,N_9087);
nor UO_1188 (O_1188,N_9493,N_9607);
or UO_1189 (O_1189,N_9723,N_9530);
and UO_1190 (O_1190,N_9751,N_9181);
or UO_1191 (O_1191,N_9761,N_9629);
nor UO_1192 (O_1192,N_9920,N_9339);
and UO_1193 (O_1193,N_9051,N_9691);
or UO_1194 (O_1194,N_9181,N_9447);
nand UO_1195 (O_1195,N_9843,N_9822);
and UO_1196 (O_1196,N_9579,N_9849);
or UO_1197 (O_1197,N_9475,N_9470);
or UO_1198 (O_1198,N_9960,N_9154);
and UO_1199 (O_1199,N_9683,N_9719);
or UO_1200 (O_1200,N_9420,N_9499);
nand UO_1201 (O_1201,N_9838,N_9878);
nand UO_1202 (O_1202,N_9352,N_9098);
or UO_1203 (O_1203,N_9724,N_9317);
nand UO_1204 (O_1204,N_9291,N_9386);
nand UO_1205 (O_1205,N_9393,N_9383);
or UO_1206 (O_1206,N_9024,N_9254);
nand UO_1207 (O_1207,N_9449,N_9341);
nand UO_1208 (O_1208,N_9936,N_9987);
or UO_1209 (O_1209,N_9570,N_9108);
or UO_1210 (O_1210,N_9383,N_9495);
xor UO_1211 (O_1211,N_9932,N_9440);
and UO_1212 (O_1212,N_9187,N_9184);
and UO_1213 (O_1213,N_9631,N_9761);
nor UO_1214 (O_1214,N_9999,N_9862);
nand UO_1215 (O_1215,N_9683,N_9653);
nor UO_1216 (O_1216,N_9168,N_9565);
nor UO_1217 (O_1217,N_9576,N_9193);
nor UO_1218 (O_1218,N_9763,N_9995);
nor UO_1219 (O_1219,N_9490,N_9186);
nor UO_1220 (O_1220,N_9135,N_9794);
or UO_1221 (O_1221,N_9333,N_9623);
nor UO_1222 (O_1222,N_9258,N_9209);
nor UO_1223 (O_1223,N_9715,N_9959);
or UO_1224 (O_1224,N_9599,N_9213);
or UO_1225 (O_1225,N_9274,N_9721);
and UO_1226 (O_1226,N_9142,N_9278);
or UO_1227 (O_1227,N_9315,N_9863);
or UO_1228 (O_1228,N_9939,N_9848);
nand UO_1229 (O_1229,N_9884,N_9746);
or UO_1230 (O_1230,N_9699,N_9576);
nand UO_1231 (O_1231,N_9592,N_9923);
nand UO_1232 (O_1232,N_9591,N_9312);
and UO_1233 (O_1233,N_9180,N_9094);
or UO_1234 (O_1234,N_9323,N_9940);
nor UO_1235 (O_1235,N_9634,N_9285);
or UO_1236 (O_1236,N_9094,N_9318);
nor UO_1237 (O_1237,N_9791,N_9787);
or UO_1238 (O_1238,N_9095,N_9697);
nor UO_1239 (O_1239,N_9400,N_9263);
or UO_1240 (O_1240,N_9263,N_9773);
nand UO_1241 (O_1241,N_9532,N_9931);
nand UO_1242 (O_1242,N_9201,N_9475);
nand UO_1243 (O_1243,N_9267,N_9307);
and UO_1244 (O_1244,N_9258,N_9999);
nor UO_1245 (O_1245,N_9750,N_9323);
nor UO_1246 (O_1246,N_9659,N_9373);
nor UO_1247 (O_1247,N_9309,N_9560);
nand UO_1248 (O_1248,N_9792,N_9812);
nand UO_1249 (O_1249,N_9655,N_9390);
nand UO_1250 (O_1250,N_9581,N_9316);
and UO_1251 (O_1251,N_9542,N_9389);
nand UO_1252 (O_1252,N_9645,N_9080);
nor UO_1253 (O_1253,N_9542,N_9467);
xnor UO_1254 (O_1254,N_9922,N_9288);
nand UO_1255 (O_1255,N_9007,N_9222);
nand UO_1256 (O_1256,N_9645,N_9250);
nor UO_1257 (O_1257,N_9022,N_9607);
or UO_1258 (O_1258,N_9961,N_9758);
and UO_1259 (O_1259,N_9575,N_9373);
or UO_1260 (O_1260,N_9842,N_9137);
and UO_1261 (O_1261,N_9745,N_9610);
nand UO_1262 (O_1262,N_9319,N_9293);
xnor UO_1263 (O_1263,N_9782,N_9665);
nand UO_1264 (O_1264,N_9049,N_9339);
nor UO_1265 (O_1265,N_9558,N_9686);
xor UO_1266 (O_1266,N_9073,N_9673);
nand UO_1267 (O_1267,N_9235,N_9147);
nand UO_1268 (O_1268,N_9110,N_9163);
or UO_1269 (O_1269,N_9016,N_9927);
nor UO_1270 (O_1270,N_9010,N_9218);
nor UO_1271 (O_1271,N_9594,N_9596);
or UO_1272 (O_1272,N_9077,N_9959);
or UO_1273 (O_1273,N_9922,N_9743);
or UO_1274 (O_1274,N_9811,N_9645);
nand UO_1275 (O_1275,N_9707,N_9681);
and UO_1276 (O_1276,N_9498,N_9829);
and UO_1277 (O_1277,N_9100,N_9891);
or UO_1278 (O_1278,N_9149,N_9933);
and UO_1279 (O_1279,N_9264,N_9663);
and UO_1280 (O_1280,N_9533,N_9067);
nand UO_1281 (O_1281,N_9937,N_9372);
and UO_1282 (O_1282,N_9960,N_9346);
or UO_1283 (O_1283,N_9234,N_9863);
nor UO_1284 (O_1284,N_9405,N_9541);
nor UO_1285 (O_1285,N_9526,N_9128);
nor UO_1286 (O_1286,N_9021,N_9338);
nand UO_1287 (O_1287,N_9534,N_9900);
nand UO_1288 (O_1288,N_9996,N_9162);
nor UO_1289 (O_1289,N_9988,N_9386);
or UO_1290 (O_1290,N_9311,N_9473);
or UO_1291 (O_1291,N_9402,N_9605);
or UO_1292 (O_1292,N_9205,N_9880);
nand UO_1293 (O_1293,N_9671,N_9662);
or UO_1294 (O_1294,N_9589,N_9285);
and UO_1295 (O_1295,N_9548,N_9820);
nor UO_1296 (O_1296,N_9790,N_9396);
and UO_1297 (O_1297,N_9607,N_9750);
nand UO_1298 (O_1298,N_9702,N_9155);
and UO_1299 (O_1299,N_9231,N_9848);
nand UO_1300 (O_1300,N_9317,N_9351);
nand UO_1301 (O_1301,N_9027,N_9857);
nor UO_1302 (O_1302,N_9361,N_9589);
nor UO_1303 (O_1303,N_9872,N_9930);
and UO_1304 (O_1304,N_9814,N_9776);
nand UO_1305 (O_1305,N_9935,N_9721);
or UO_1306 (O_1306,N_9620,N_9682);
and UO_1307 (O_1307,N_9504,N_9462);
nor UO_1308 (O_1308,N_9601,N_9482);
nor UO_1309 (O_1309,N_9350,N_9954);
nor UO_1310 (O_1310,N_9798,N_9193);
xnor UO_1311 (O_1311,N_9501,N_9116);
nand UO_1312 (O_1312,N_9676,N_9484);
nor UO_1313 (O_1313,N_9767,N_9587);
and UO_1314 (O_1314,N_9903,N_9809);
and UO_1315 (O_1315,N_9245,N_9466);
nand UO_1316 (O_1316,N_9638,N_9704);
and UO_1317 (O_1317,N_9529,N_9709);
nand UO_1318 (O_1318,N_9198,N_9848);
and UO_1319 (O_1319,N_9057,N_9283);
nor UO_1320 (O_1320,N_9086,N_9593);
and UO_1321 (O_1321,N_9718,N_9243);
nand UO_1322 (O_1322,N_9718,N_9013);
nand UO_1323 (O_1323,N_9336,N_9260);
nor UO_1324 (O_1324,N_9645,N_9406);
nor UO_1325 (O_1325,N_9514,N_9616);
and UO_1326 (O_1326,N_9259,N_9659);
nor UO_1327 (O_1327,N_9287,N_9836);
nand UO_1328 (O_1328,N_9129,N_9976);
nor UO_1329 (O_1329,N_9986,N_9216);
or UO_1330 (O_1330,N_9438,N_9234);
and UO_1331 (O_1331,N_9178,N_9212);
xor UO_1332 (O_1332,N_9199,N_9801);
nor UO_1333 (O_1333,N_9700,N_9957);
nand UO_1334 (O_1334,N_9061,N_9704);
or UO_1335 (O_1335,N_9333,N_9649);
nor UO_1336 (O_1336,N_9830,N_9837);
nor UO_1337 (O_1337,N_9321,N_9277);
nand UO_1338 (O_1338,N_9919,N_9149);
and UO_1339 (O_1339,N_9233,N_9156);
nor UO_1340 (O_1340,N_9098,N_9059);
nand UO_1341 (O_1341,N_9682,N_9054);
and UO_1342 (O_1342,N_9000,N_9569);
and UO_1343 (O_1343,N_9033,N_9979);
nand UO_1344 (O_1344,N_9238,N_9131);
nand UO_1345 (O_1345,N_9643,N_9418);
and UO_1346 (O_1346,N_9970,N_9337);
nor UO_1347 (O_1347,N_9376,N_9665);
nor UO_1348 (O_1348,N_9778,N_9188);
nand UO_1349 (O_1349,N_9091,N_9327);
and UO_1350 (O_1350,N_9074,N_9653);
or UO_1351 (O_1351,N_9309,N_9823);
or UO_1352 (O_1352,N_9003,N_9808);
or UO_1353 (O_1353,N_9094,N_9358);
and UO_1354 (O_1354,N_9528,N_9285);
nor UO_1355 (O_1355,N_9706,N_9334);
nand UO_1356 (O_1356,N_9613,N_9387);
and UO_1357 (O_1357,N_9431,N_9392);
or UO_1358 (O_1358,N_9097,N_9268);
or UO_1359 (O_1359,N_9021,N_9590);
nand UO_1360 (O_1360,N_9901,N_9956);
and UO_1361 (O_1361,N_9326,N_9670);
or UO_1362 (O_1362,N_9147,N_9464);
nand UO_1363 (O_1363,N_9044,N_9464);
and UO_1364 (O_1364,N_9000,N_9770);
nand UO_1365 (O_1365,N_9583,N_9537);
nand UO_1366 (O_1366,N_9462,N_9379);
nand UO_1367 (O_1367,N_9430,N_9057);
and UO_1368 (O_1368,N_9990,N_9929);
nor UO_1369 (O_1369,N_9654,N_9627);
nand UO_1370 (O_1370,N_9198,N_9909);
nand UO_1371 (O_1371,N_9278,N_9671);
nor UO_1372 (O_1372,N_9747,N_9475);
and UO_1373 (O_1373,N_9458,N_9399);
nor UO_1374 (O_1374,N_9238,N_9846);
and UO_1375 (O_1375,N_9608,N_9447);
or UO_1376 (O_1376,N_9985,N_9078);
nand UO_1377 (O_1377,N_9300,N_9880);
and UO_1378 (O_1378,N_9230,N_9648);
nand UO_1379 (O_1379,N_9149,N_9176);
or UO_1380 (O_1380,N_9988,N_9135);
and UO_1381 (O_1381,N_9881,N_9190);
or UO_1382 (O_1382,N_9979,N_9865);
and UO_1383 (O_1383,N_9922,N_9221);
nor UO_1384 (O_1384,N_9506,N_9156);
nand UO_1385 (O_1385,N_9675,N_9537);
and UO_1386 (O_1386,N_9119,N_9072);
nand UO_1387 (O_1387,N_9961,N_9326);
nor UO_1388 (O_1388,N_9456,N_9411);
nand UO_1389 (O_1389,N_9316,N_9121);
nor UO_1390 (O_1390,N_9121,N_9726);
and UO_1391 (O_1391,N_9318,N_9396);
nor UO_1392 (O_1392,N_9271,N_9422);
nand UO_1393 (O_1393,N_9602,N_9492);
nor UO_1394 (O_1394,N_9640,N_9293);
nor UO_1395 (O_1395,N_9509,N_9982);
nor UO_1396 (O_1396,N_9919,N_9706);
or UO_1397 (O_1397,N_9801,N_9730);
nor UO_1398 (O_1398,N_9117,N_9299);
nand UO_1399 (O_1399,N_9147,N_9845);
and UO_1400 (O_1400,N_9272,N_9084);
or UO_1401 (O_1401,N_9239,N_9584);
and UO_1402 (O_1402,N_9712,N_9275);
nand UO_1403 (O_1403,N_9534,N_9221);
nor UO_1404 (O_1404,N_9693,N_9209);
nand UO_1405 (O_1405,N_9277,N_9947);
and UO_1406 (O_1406,N_9262,N_9449);
or UO_1407 (O_1407,N_9285,N_9489);
and UO_1408 (O_1408,N_9097,N_9574);
nor UO_1409 (O_1409,N_9108,N_9460);
nor UO_1410 (O_1410,N_9571,N_9849);
xor UO_1411 (O_1411,N_9940,N_9087);
nor UO_1412 (O_1412,N_9571,N_9783);
or UO_1413 (O_1413,N_9451,N_9172);
nand UO_1414 (O_1414,N_9841,N_9086);
nand UO_1415 (O_1415,N_9632,N_9198);
nor UO_1416 (O_1416,N_9952,N_9492);
nor UO_1417 (O_1417,N_9990,N_9953);
or UO_1418 (O_1418,N_9199,N_9661);
nand UO_1419 (O_1419,N_9193,N_9330);
nor UO_1420 (O_1420,N_9973,N_9075);
and UO_1421 (O_1421,N_9457,N_9985);
nor UO_1422 (O_1422,N_9013,N_9421);
nand UO_1423 (O_1423,N_9272,N_9151);
or UO_1424 (O_1424,N_9371,N_9231);
or UO_1425 (O_1425,N_9206,N_9449);
and UO_1426 (O_1426,N_9203,N_9694);
nand UO_1427 (O_1427,N_9551,N_9593);
and UO_1428 (O_1428,N_9621,N_9444);
or UO_1429 (O_1429,N_9907,N_9069);
and UO_1430 (O_1430,N_9798,N_9570);
nand UO_1431 (O_1431,N_9832,N_9300);
or UO_1432 (O_1432,N_9379,N_9989);
nand UO_1433 (O_1433,N_9609,N_9158);
or UO_1434 (O_1434,N_9202,N_9419);
or UO_1435 (O_1435,N_9614,N_9462);
nand UO_1436 (O_1436,N_9658,N_9820);
nand UO_1437 (O_1437,N_9250,N_9334);
nand UO_1438 (O_1438,N_9830,N_9117);
or UO_1439 (O_1439,N_9224,N_9899);
or UO_1440 (O_1440,N_9890,N_9485);
xnor UO_1441 (O_1441,N_9249,N_9234);
nor UO_1442 (O_1442,N_9817,N_9597);
nand UO_1443 (O_1443,N_9438,N_9521);
nand UO_1444 (O_1444,N_9187,N_9787);
nor UO_1445 (O_1445,N_9510,N_9788);
and UO_1446 (O_1446,N_9928,N_9493);
or UO_1447 (O_1447,N_9946,N_9931);
nand UO_1448 (O_1448,N_9069,N_9125);
or UO_1449 (O_1449,N_9666,N_9803);
nand UO_1450 (O_1450,N_9752,N_9251);
nand UO_1451 (O_1451,N_9680,N_9791);
nand UO_1452 (O_1452,N_9950,N_9536);
or UO_1453 (O_1453,N_9962,N_9592);
nand UO_1454 (O_1454,N_9597,N_9906);
and UO_1455 (O_1455,N_9453,N_9397);
nand UO_1456 (O_1456,N_9557,N_9565);
or UO_1457 (O_1457,N_9217,N_9451);
nand UO_1458 (O_1458,N_9430,N_9669);
or UO_1459 (O_1459,N_9639,N_9638);
nand UO_1460 (O_1460,N_9395,N_9161);
nor UO_1461 (O_1461,N_9214,N_9371);
nand UO_1462 (O_1462,N_9850,N_9003);
or UO_1463 (O_1463,N_9949,N_9326);
and UO_1464 (O_1464,N_9503,N_9873);
nor UO_1465 (O_1465,N_9437,N_9808);
xor UO_1466 (O_1466,N_9189,N_9960);
or UO_1467 (O_1467,N_9409,N_9019);
nor UO_1468 (O_1468,N_9965,N_9245);
or UO_1469 (O_1469,N_9498,N_9887);
and UO_1470 (O_1470,N_9973,N_9849);
nand UO_1471 (O_1471,N_9939,N_9056);
or UO_1472 (O_1472,N_9860,N_9302);
nor UO_1473 (O_1473,N_9844,N_9461);
nand UO_1474 (O_1474,N_9711,N_9695);
nand UO_1475 (O_1475,N_9158,N_9914);
or UO_1476 (O_1476,N_9825,N_9959);
nor UO_1477 (O_1477,N_9289,N_9516);
nand UO_1478 (O_1478,N_9770,N_9071);
nand UO_1479 (O_1479,N_9245,N_9576);
nor UO_1480 (O_1480,N_9435,N_9497);
xor UO_1481 (O_1481,N_9143,N_9051);
nand UO_1482 (O_1482,N_9686,N_9596);
nor UO_1483 (O_1483,N_9885,N_9279);
nor UO_1484 (O_1484,N_9769,N_9900);
xor UO_1485 (O_1485,N_9692,N_9768);
or UO_1486 (O_1486,N_9376,N_9628);
nand UO_1487 (O_1487,N_9808,N_9281);
or UO_1488 (O_1488,N_9001,N_9675);
nand UO_1489 (O_1489,N_9441,N_9385);
or UO_1490 (O_1490,N_9707,N_9823);
nor UO_1491 (O_1491,N_9250,N_9257);
nand UO_1492 (O_1492,N_9072,N_9004);
xor UO_1493 (O_1493,N_9378,N_9351);
and UO_1494 (O_1494,N_9028,N_9781);
nand UO_1495 (O_1495,N_9902,N_9006);
and UO_1496 (O_1496,N_9726,N_9271);
nand UO_1497 (O_1497,N_9028,N_9456);
and UO_1498 (O_1498,N_9521,N_9035);
and UO_1499 (O_1499,N_9913,N_9972);
endmodule