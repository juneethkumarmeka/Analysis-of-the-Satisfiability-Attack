module basic_2500_25000_3000_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1037,In_1973);
nor U1 (N_1,In_113,In_528);
or U2 (N_2,In_2404,In_1960);
and U3 (N_3,In_940,In_402);
xor U4 (N_4,In_1748,In_2283);
nor U5 (N_5,In_480,In_237);
or U6 (N_6,In_589,In_1836);
xnor U7 (N_7,In_814,In_1891);
and U8 (N_8,In_678,In_972);
xnor U9 (N_9,In_2254,In_349);
nand U10 (N_10,In_609,In_1187);
xor U11 (N_11,In_837,In_2305);
nand U12 (N_12,In_1223,In_2288);
or U13 (N_13,In_1715,In_364);
or U14 (N_14,In_771,In_1309);
nand U15 (N_15,In_1705,In_71);
xor U16 (N_16,In_177,In_1350);
or U17 (N_17,In_756,In_335);
or U18 (N_18,In_2338,In_2136);
nand U19 (N_19,In_639,In_321);
and U20 (N_20,In_252,In_592);
nand U21 (N_21,In_384,In_2481);
or U22 (N_22,In_632,In_1781);
and U23 (N_23,In_1754,In_788);
nand U24 (N_24,In_1125,In_1961);
xor U25 (N_25,In_1261,In_1074);
or U26 (N_26,In_685,In_1731);
nand U27 (N_27,In_731,In_1712);
or U28 (N_28,In_919,In_442);
nor U29 (N_29,In_2449,In_1281);
and U30 (N_30,In_2215,In_1813);
nand U31 (N_31,In_2155,In_623);
and U32 (N_32,In_1943,In_2133);
or U33 (N_33,In_664,In_2034);
nor U34 (N_34,In_1292,In_819);
xor U35 (N_35,In_1686,In_93);
or U36 (N_36,In_412,In_2320);
nand U37 (N_37,In_2201,In_2248);
xnor U38 (N_38,In_850,In_726);
nor U39 (N_39,In_966,In_1010);
nor U40 (N_40,In_2251,In_408);
xor U41 (N_41,In_253,In_1041);
nand U42 (N_42,In_1232,In_2377);
xor U43 (N_43,In_943,In_2071);
nand U44 (N_44,In_1559,In_27);
nor U45 (N_45,In_330,In_1695);
nand U46 (N_46,In_1287,In_1931);
nand U47 (N_47,In_1468,In_1122);
xor U48 (N_48,In_2121,In_400);
nor U49 (N_49,In_211,In_1057);
or U50 (N_50,In_968,In_1410);
or U51 (N_51,In_719,In_957);
or U52 (N_52,In_1824,In_512);
or U53 (N_53,In_259,In_1828);
xnor U54 (N_54,In_1167,In_714);
xnor U55 (N_55,In_845,In_1180);
xor U56 (N_56,In_668,In_1782);
nand U57 (N_57,In_1012,In_8);
xor U58 (N_58,In_1371,In_1690);
and U59 (N_59,In_1124,In_1692);
xor U60 (N_60,In_513,In_974);
or U61 (N_61,In_1336,In_1434);
nor U62 (N_62,In_546,In_126);
nor U63 (N_63,In_2087,In_1738);
or U64 (N_64,In_2203,In_580);
nand U65 (N_65,In_427,In_646);
xor U66 (N_66,In_597,In_1302);
and U67 (N_67,In_1583,In_204);
and U68 (N_68,In_2126,In_1854);
nand U69 (N_69,In_212,In_161);
and U70 (N_70,In_110,In_306);
nand U71 (N_71,In_2359,In_2086);
and U72 (N_72,In_175,In_2441);
xor U73 (N_73,In_1369,In_1719);
nand U74 (N_74,In_1778,In_2055);
nor U75 (N_75,In_461,In_802);
xor U76 (N_76,In_1386,In_1967);
xor U77 (N_77,In_2080,In_2222);
or U78 (N_78,In_1558,In_2276);
nand U79 (N_79,In_1638,In_1421);
or U80 (N_80,In_2308,In_2156);
xor U81 (N_81,In_949,In_6);
or U82 (N_82,In_2267,In_923);
xnor U83 (N_83,In_1619,In_1581);
or U84 (N_84,In_2069,In_1955);
nand U85 (N_85,In_122,In_1405);
and U86 (N_86,In_1349,In_550);
nor U87 (N_87,In_622,In_2163);
nor U88 (N_88,In_1779,In_1197);
nand U89 (N_89,In_258,In_455);
or U90 (N_90,In_2202,In_41);
nand U91 (N_91,In_1228,In_2082);
xor U92 (N_92,In_1427,In_55);
nor U93 (N_93,In_1680,In_792);
xor U94 (N_94,In_2037,In_1681);
or U95 (N_95,In_453,In_395);
and U96 (N_96,In_1864,In_1173);
nand U97 (N_97,In_389,In_119);
and U98 (N_98,In_883,In_1353);
or U99 (N_99,In_2102,In_1075);
or U100 (N_100,In_228,In_1594);
nand U101 (N_101,In_1825,In_1776);
xor U102 (N_102,In_2366,In_1062);
and U103 (N_103,In_2002,In_820);
or U104 (N_104,In_356,In_429);
xor U105 (N_105,In_1480,In_963);
nand U106 (N_106,In_3,In_1602);
and U107 (N_107,In_519,In_1841);
or U108 (N_108,In_488,In_1551);
xor U109 (N_109,In_1015,In_1721);
or U110 (N_110,In_1821,In_2416);
nand U111 (N_111,In_897,In_1513);
nor U112 (N_112,In_2260,In_1615);
and U113 (N_113,In_1000,In_1377);
nand U114 (N_114,In_1839,In_137);
nor U115 (N_115,In_88,In_2218);
xor U116 (N_116,In_2384,In_2068);
or U117 (N_117,In_2399,In_1083);
nor U118 (N_118,In_1224,In_699);
or U119 (N_119,In_232,In_367);
and U120 (N_120,In_1519,In_1208);
xnor U121 (N_121,In_366,In_905);
xnor U122 (N_122,In_2499,In_274);
nand U123 (N_123,In_2483,In_344);
or U124 (N_124,In_1479,In_2357);
nor U125 (N_125,In_2165,In_502);
and U126 (N_126,In_1734,In_1425);
and U127 (N_127,In_1874,In_929);
or U128 (N_128,In_870,In_1267);
xor U129 (N_129,In_2411,In_2100);
xor U130 (N_130,In_2137,In_1308);
and U131 (N_131,In_1586,In_1411);
or U132 (N_132,In_1934,In_340);
and U133 (N_133,In_993,In_1959);
xor U134 (N_134,In_2261,In_842);
xor U135 (N_135,In_1073,In_1913);
or U136 (N_136,In_2461,In_267);
or U137 (N_137,In_992,In_1942);
nand U138 (N_138,In_254,In_420);
or U139 (N_139,In_1110,In_30);
or U140 (N_140,In_1424,In_2348);
xnor U141 (N_141,In_207,In_680);
nor U142 (N_142,In_62,In_1743);
nand U143 (N_143,In_1021,In_2041);
nand U144 (N_144,In_1490,In_939);
nor U145 (N_145,In_464,In_876);
or U146 (N_146,In_755,In_983);
or U147 (N_147,In_2056,In_459);
xor U148 (N_148,In_1507,In_2178);
or U149 (N_149,In_1851,In_106);
and U150 (N_150,In_573,In_1911);
nand U151 (N_151,In_68,In_28);
xor U152 (N_152,In_1295,In_1626);
nor U153 (N_153,In_1044,In_1254);
nor U154 (N_154,In_77,In_2373);
or U155 (N_155,In_1355,In_305);
or U156 (N_156,In_1667,In_1593);
nor U157 (N_157,In_835,In_1755);
nor U158 (N_158,In_2414,In_324);
or U159 (N_159,In_593,In_2021);
nand U160 (N_160,In_2060,In_2187);
xor U161 (N_161,In_1890,In_1387);
and U162 (N_162,In_2290,In_670);
xor U163 (N_163,In_524,In_2031);
or U164 (N_164,In_343,In_1226);
nor U165 (N_165,In_1177,In_426);
nand U166 (N_166,In_1248,In_261);
nor U167 (N_167,In_749,In_1130);
nand U168 (N_168,In_208,In_31);
and U169 (N_169,In_798,In_849);
xnor U170 (N_170,In_1493,In_348);
nand U171 (N_171,In_894,In_411);
and U172 (N_172,In_1843,In_1138);
nor U173 (N_173,In_1750,In_659);
nand U174 (N_174,In_1987,In_688);
and U175 (N_175,In_2192,In_369);
nand U176 (N_176,In_1118,In_2264);
and U177 (N_177,In_283,In_2333);
nor U178 (N_178,In_241,In_56);
xnor U179 (N_179,In_1277,In_909);
nor U180 (N_180,In_1040,In_1168);
nor U181 (N_181,In_1025,In_1429);
xnor U182 (N_182,In_1689,In_767);
nor U183 (N_183,In_672,In_2332);
nand U184 (N_184,In_826,In_1810);
nor U185 (N_185,In_1893,In_1347);
nor U186 (N_186,In_1321,In_158);
or U187 (N_187,In_482,In_987);
nand U188 (N_188,In_1724,In_147);
xor U189 (N_189,In_2387,In_575);
and U190 (N_190,In_1670,In_2164);
nor U191 (N_191,In_1898,In_79);
xnor U192 (N_192,In_1601,In_2470);
or U193 (N_193,In_1213,In_2197);
nand U194 (N_194,In_1956,In_1241);
nand U195 (N_195,In_1158,In_2105);
and U196 (N_196,In_1568,In_930);
and U197 (N_197,In_221,In_124);
or U198 (N_198,In_2392,In_631);
and U199 (N_199,In_1034,In_698);
or U200 (N_200,In_2048,In_82);
or U201 (N_201,In_772,In_388);
or U202 (N_202,In_1869,In_841);
and U203 (N_203,In_1103,In_2174);
or U204 (N_204,In_227,In_2094);
and U205 (N_205,In_421,In_709);
nor U206 (N_206,In_1844,In_2045);
or U207 (N_207,In_1749,In_332);
xor U208 (N_208,In_1744,In_2406);
nor U209 (N_209,In_2370,In_2117);
nand U210 (N_210,In_173,In_80);
nand U211 (N_211,In_583,In_1319);
nand U212 (N_212,In_499,In_722);
or U213 (N_213,In_893,In_2317);
nor U214 (N_214,In_982,In_149);
nor U215 (N_215,In_1327,In_878);
nor U216 (N_216,In_2463,In_1328);
nor U217 (N_217,In_2272,In_1669);
or U218 (N_218,In_687,In_1150);
or U219 (N_219,In_66,In_277);
and U220 (N_220,In_1787,In_747);
xor U221 (N_221,In_885,In_667);
nand U222 (N_222,In_1508,In_2408);
xor U223 (N_223,In_1487,In_1381);
nand U224 (N_224,In_2281,In_1720);
nand U225 (N_225,In_245,In_636);
nor U226 (N_226,In_675,In_118);
xnor U227 (N_227,In_1345,In_638);
and U228 (N_228,In_40,In_2020);
or U229 (N_229,In_1462,In_2437);
nor U230 (N_230,In_1294,In_785);
or U231 (N_231,In_168,In_407);
or U232 (N_232,In_469,In_1078);
xnor U233 (N_233,In_1183,In_1391);
nor U234 (N_234,In_202,In_1780);
or U235 (N_235,In_591,In_23);
or U236 (N_236,In_1968,In_311);
nor U237 (N_237,In_391,In_2232);
or U238 (N_238,In_222,In_69);
or U239 (N_239,In_1947,In_1099);
nand U240 (N_240,In_2091,In_256);
nand U241 (N_241,In_2444,In_316);
nor U242 (N_242,In_579,In_1298);
xor U243 (N_243,In_1323,In_445);
xnor U244 (N_244,In_120,In_1885);
xnor U245 (N_245,In_800,In_2167);
nor U246 (N_246,In_1026,In_536);
nand U247 (N_247,In_1660,In_1702);
nor U248 (N_248,In_936,In_2497);
nand U249 (N_249,In_1278,In_669);
or U250 (N_250,In_840,In_1629);
nand U251 (N_251,In_2149,In_1783);
nand U252 (N_252,In_135,In_1856);
nor U253 (N_253,In_2030,In_1239);
or U254 (N_254,In_1330,In_242);
or U255 (N_255,In_879,In_2017);
xor U256 (N_256,In_1300,In_2081);
nand U257 (N_257,In_361,In_1106);
nor U258 (N_258,In_776,In_1011);
or U259 (N_259,In_1486,In_18);
nand U260 (N_260,In_737,In_960);
nand U261 (N_261,In_833,In_1972);
and U262 (N_262,In_501,In_1991);
or U263 (N_263,In_2024,In_17);
or U264 (N_264,In_1404,In_365);
or U265 (N_265,In_1694,In_529);
and U266 (N_266,In_1446,In_736);
xnor U267 (N_267,In_2393,In_1896);
xor U268 (N_268,In_188,In_1904);
or U269 (N_269,In_1467,In_1286);
nor U270 (N_270,In_45,In_1693);
nand U271 (N_271,In_882,In_1220);
and U272 (N_272,In_2007,In_1614);
nand U273 (N_273,In_1521,In_1948);
nand U274 (N_274,In_1642,In_2230);
xor U275 (N_275,In_434,In_1364);
nor U276 (N_276,In_818,In_1113);
xnor U277 (N_277,In_2401,In_808);
nand U278 (N_278,In_2327,In_1799);
or U279 (N_279,In_652,In_465);
or U280 (N_280,In_333,In_2181);
or U281 (N_281,In_545,In_514);
or U282 (N_282,In_797,In_2095);
nor U283 (N_283,In_2005,In_108);
and U284 (N_284,In_1403,In_401);
and U285 (N_285,In_1495,In_1093);
or U286 (N_286,In_19,In_537);
or U287 (N_287,In_1950,In_708);
and U288 (N_288,In_1316,In_656);
or U289 (N_289,In_1580,In_662);
xor U290 (N_290,In_724,In_1033);
nor U291 (N_291,In_9,In_1662);
and U292 (N_292,In_2278,In_1822);
nand U293 (N_293,In_1472,In_1152);
xor U294 (N_294,In_326,In_1528);
or U295 (N_295,In_1582,In_2072);
xor U296 (N_296,In_780,In_1756);
nor U297 (N_297,In_2343,In_2249);
nor U298 (N_298,In_1354,In_991);
nand U299 (N_299,In_191,In_1491);
nand U300 (N_300,In_2452,In_1589);
xnor U301 (N_301,In_1798,In_1982);
or U302 (N_302,In_466,In_1023);
xnor U303 (N_303,In_2376,In_2205);
or U304 (N_304,In_1055,In_1489);
nand U305 (N_305,In_1204,In_677);
or U306 (N_306,In_1202,In_1613);
and U307 (N_307,In_1661,In_1951);
and U308 (N_308,In_294,In_980);
or U309 (N_309,In_2443,In_2211);
and U310 (N_310,In_1696,In_1352);
nand U311 (N_311,In_1623,In_811);
and U312 (N_312,In_2438,In_189);
nor U313 (N_313,In_1385,In_504);
nand U314 (N_314,In_125,In_888);
or U315 (N_315,In_60,In_1820);
nor U316 (N_316,In_1996,In_713);
or U317 (N_317,In_1886,In_336);
nor U318 (N_318,In_1708,In_1677);
nor U319 (N_319,In_872,In_2315);
xor U320 (N_320,In_594,In_1251);
and U321 (N_321,In_1710,In_1243);
nand U322 (N_322,In_2270,In_2077);
nand U323 (N_323,In_2235,In_1101);
nand U324 (N_324,In_12,In_902);
nand U325 (N_325,In_1532,In_1926);
nor U326 (N_326,In_740,In_1557);
nand U327 (N_327,In_2294,In_1178);
nor U328 (N_328,In_1198,In_239);
nor U329 (N_329,In_1440,In_72);
xnor U330 (N_330,In_406,In_603);
xor U331 (N_331,In_509,In_1238);
xnor U332 (N_332,In_1684,In_1092);
xor U333 (N_333,In_1999,In_543);
and U334 (N_334,In_347,In_1672);
nor U335 (N_335,In_1542,In_1064);
or U336 (N_336,In_26,In_1496);
nor U337 (N_337,In_1587,In_1830);
and U338 (N_338,In_1272,In_1408);
nand U339 (N_339,In_1443,In_1648);
xor U340 (N_340,In_2492,In_1870);
nand U341 (N_341,In_2400,In_718);
xnor U342 (N_342,In_1920,In_186);
and U343 (N_343,In_831,In_2336);
xnor U344 (N_344,In_43,In_1400);
nand U345 (N_345,In_1423,In_457);
nor U346 (N_346,In_1668,In_733);
and U347 (N_347,In_5,In_2447);
or U348 (N_348,In_959,In_2469);
nand U349 (N_349,In_1604,In_1505);
nand U350 (N_350,In_2368,In_54);
and U351 (N_351,In_1522,In_376);
xnor U352 (N_352,In_1133,In_1195);
and U353 (N_353,In_2029,In_1222);
xor U354 (N_354,In_16,In_477);
or U355 (N_355,In_2291,In_2292);
nor U356 (N_356,In_2114,In_157);
or U357 (N_357,In_2243,In_2151);
xnor U358 (N_358,In_1290,In_1988);
and U359 (N_359,In_64,In_900);
xnor U360 (N_360,In_103,In_2382);
and U361 (N_361,In_694,In_353);
nand U362 (N_362,In_20,In_2341);
nor U363 (N_363,In_1359,In_843);
nor U364 (N_364,In_78,In_1791);
and U365 (N_365,In_2398,In_1556);
or U366 (N_366,In_2494,In_2426);
or U367 (N_367,In_196,In_385);
and U368 (N_368,In_1571,In_2093);
or U369 (N_369,In_1873,In_2284);
xor U370 (N_370,In_1895,In_190);
xnor U371 (N_371,In_586,In_1182);
or U372 (N_372,In_2191,In_1861);
nor U373 (N_373,In_2138,In_2049);
xnor U374 (N_374,In_437,In_976);
and U375 (N_375,In_1827,In_607);
and U376 (N_376,In_2258,In_1714);
nor U377 (N_377,In_1435,In_1995);
and U378 (N_378,In_390,In_763);
nand U379 (N_379,In_192,In_1089);
nor U380 (N_380,In_910,In_525);
and U381 (N_381,In_2495,In_1052);
and U382 (N_382,In_438,In_1084);
nor U383 (N_383,In_1009,In_73);
xor U384 (N_384,In_2364,In_2141);
or U385 (N_385,In_1624,In_2360);
nand U386 (N_386,In_517,In_279);
xor U387 (N_387,In_1794,In_1190);
and U388 (N_388,In_418,In_2177);
nor U389 (N_389,In_285,In_1249);
nand U390 (N_390,In_2491,In_229);
xnor U391 (N_391,In_2006,In_1742);
nor U392 (N_392,In_1665,In_1883);
xor U393 (N_393,In_620,In_289);
nor U394 (N_394,In_263,In_2166);
or U395 (N_395,In_1230,In_1166);
nor U396 (N_396,In_1806,In_999);
nor U397 (N_397,In_1657,In_1284);
or U398 (N_398,In_781,In_2090);
nor U399 (N_399,In_906,In_1946);
xor U400 (N_400,In_1017,In_219);
nor U401 (N_401,In_2172,In_2078);
nor U402 (N_402,In_1482,In_853);
and U403 (N_403,In_2282,In_1941);
or U404 (N_404,In_2342,In_2073);
nor U405 (N_405,In_585,In_1266);
or U406 (N_406,In_1407,In_1797);
xnor U407 (N_407,In_490,In_1918);
and U408 (N_408,In_1372,In_1728);
nand U409 (N_409,In_10,In_1157);
and U410 (N_410,In_946,In_322);
nand U411 (N_411,In_979,In_49);
nor U412 (N_412,In_1514,In_2128);
nor U413 (N_413,In_150,In_1108);
or U414 (N_414,In_292,In_544);
nor U415 (N_415,In_2119,In_1175);
xnor U416 (N_416,In_1699,In_1531);
nor U417 (N_417,In_1126,In_565);
nand U418 (N_418,In_2208,In_1717);
and U419 (N_419,In_1739,In_554);
nand U420 (N_420,In_38,In_1520);
nand U421 (N_421,In_1161,In_588);
and U422 (N_422,In_732,In_935);
and U423 (N_423,In_1792,In_1484);
xnor U424 (N_424,In_1838,In_495);
nand U425 (N_425,In_2050,In_1339);
xnor U426 (N_426,In_2225,In_1053);
xor U427 (N_427,In_1014,In_1595);
xnor U428 (N_428,In_937,In_1216);
and U429 (N_429,In_2245,In_1303);
and U430 (N_430,In_1597,In_1135);
xnor U431 (N_431,In_1028,In_281);
nand U432 (N_432,In_712,In_2259);
nor U433 (N_433,In_269,In_2036);
and U434 (N_434,In_2388,In_2003);
nand U435 (N_435,In_1983,In_1509);
nor U436 (N_436,In_2280,In_505);
nor U437 (N_437,In_762,In_1549);
and U438 (N_438,In_904,In_2240);
nand U439 (N_439,In_2433,In_127);
and U440 (N_440,In_107,In_984);
nor U441 (N_441,In_1397,In_658);
or U442 (N_442,In_1603,In_2262);
xor U443 (N_443,In_961,In_508);
xor U444 (N_444,In_859,In_1240);
nor U445 (N_445,In_1718,In_1971);
and U446 (N_446,In_485,In_750);
and U447 (N_447,In_2033,In_1132);
xor U448 (N_448,In_2120,In_1301);
or U449 (N_449,In_1588,In_1585);
nor U450 (N_450,In_558,In_1450);
nor U451 (N_451,In_526,In_2250);
nand U452 (N_452,In_1121,In_1373);
nor U453 (N_453,In_264,In_2421);
and U454 (N_454,In_665,In_1970);
or U455 (N_455,In_2186,In_1401);
nand U456 (N_456,In_782,In_35);
and U457 (N_457,In_2277,In_950);
nand U458 (N_458,In_1072,In_2429);
or U459 (N_459,In_1343,In_2233);
xor U460 (N_460,In_2346,In_1264);
nand U461 (N_461,In_410,In_572);
or U462 (N_462,In_569,In_634);
nand U463 (N_463,In_1250,In_230);
xor U464 (N_464,In_1409,In_1376);
xnor U465 (N_465,In_2140,In_628);
nor U466 (N_466,In_1566,In_381);
and U467 (N_467,In_924,In_337);
or U468 (N_468,In_2383,In_2214);
xor U469 (N_469,In_2372,In_661);
xor U470 (N_470,In_1676,In_1650);
or U471 (N_471,In_2046,In_2083);
nor U472 (N_472,In_187,In_2409);
nand U473 (N_473,In_1765,In_2475);
xor U474 (N_474,In_1674,In_1170);
or U475 (N_475,In_1392,In_216);
or U476 (N_476,In_602,In_1819);
xor U477 (N_477,In_2389,In_1324);
or U478 (N_478,In_926,In_822);
or U479 (N_479,In_1811,In_439);
and U480 (N_480,In_610,In_1527);
or U481 (N_481,In_873,In_1077);
nand U482 (N_482,In_1143,In_303);
nand U483 (N_483,In_2035,In_1818);
nand U484 (N_484,In_1937,In_777);
nor U485 (N_485,In_738,In_25);
and U486 (N_486,In_483,In_810);
nand U487 (N_487,In_57,In_2079);
nand U488 (N_488,In_355,In_1771);
or U489 (N_489,In_338,In_2206);
nor U490 (N_490,In_481,In_880);
nand U491 (N_491,In_916,In_1939);
nor U492 (N_492,In_836,In_971);
or U493 (N_493,In_540,In_94);
nand U494 (N_494,In_1727,In_394);
and U495 (N_495,In_2395,In_1070);
xnor U496 (N_496,In_1945,In_1767);
and U497 (N_497,In_1001,In_1453);
or U498 (N_498,In_886,In_799);
xnor U499 (N_499,In_1837,In_1685);
nand U500 (N_500,N_42,In_2394);
nor U501 (N_501,In_342,In_1428);
nor U502 (N_502,In_1981,In_458);
nand U503 (N_503,In_1459,In_1733);
nand U504 (N_504,N_243,In_50);
nor U505 (N_505,In_531,In_2468);
and U506 (N_506,In_1115,N_323);
or U507 (N_507,In_2183,N_412);
nor U508 (N_508,In_1541,In_341);
xor U509 (N_509,In_1430,In_1884);
nand U510 (N_510,In_2011,In_2115);
or U511 (N_511,In_2440,In_1047);
and U512 (N_512,In_1100,In_1437);
nor U513 (N_513,In_858,In_1735);
or U514 (N_514,N_211,In_1760);
nand U515 (N_515,In_1156,In_1706);
or U516 (N_516,In_2358,In_2051);
and U517 (N_517,N_56,In_1418);
and U518 (N_518,In_102,In_890);
nand U519 (N_519,N_363,N_423);
xor U520 (N_520,In_616,In_2);
and U521 (N_521,In_1338,In_1829);
and U522 (N_522,In_302,In_964);
and U523 (N_523,In_1789,In_1850);
nor U524 (N_524,In_2353,In_2303);
nor U525 (N_525,In_817,N_199);
nor U526 (N_526,In_194,N_272);
and U527 (N_527,In_271,In_416);
and U528 (N_528,In_2378,In_1620);
or U529 (N_529,In_2484,N_207);
nand U530 (N_530,N_409,In_1050);
nand U531 (N_531,N_415,N_105);
or U532 (N_532,In_472,In_1914);
and U533 (N_533,N_310,In_1503);
nor U534 (N_534,In_1848,In_611);
or U535 (N_535,N_165,In_2018);
xnor U536 (N_536,In_1570,In_300);
nor U537 (N_537,In_443,In_46);
nor U538 (N_538,N_133,In_1512);
and U539 (N_539,In_1761,N_224);
or U540 (N_540,In_1652,In_598);
nor U541 (N_541,In_2247,N_392);
or U542 (N_542,In_276,In_223);
nand U543 (N_543,In_1304,N_301);
nor U544 (N_544,In_2350,N_97);
xor U545 (N_545,In_334,In_1060);
nor U546 (N_546,In_2042,In_200);
and U547 (N_547,N_221,In_2344);
nor U548 (N_548,In_539,In_627);
xor U549 (N_549,In_1107,In_2176);
and U550 (N_550,In_463,N_20);
nand U551 (N_551,N_354,In_774);
nor U552 (N_552,In_2299,In_1452);
nor U553 (N_553,In_595,N_201);
nor U554 (N_554,In_325,N_167);
nor U555 (N_555,In_1625,In_2144);
nor U556 (N_556,In_2423,N_3);
nor U557 (N_557,In_1233,In_1833);
nand U558 (N_558,In_265,In_1881);
xnor U559 (N_559,In_869,In_467);
or U560 (N_560,In_1803,In_1888);
nor U561 (N_561,In_2489,In_2058);
nand U562 (N_562,In_1105,In_96);
nor U563 (N_563,In_1574,In_922);
nand U564 (N_564,In_2412,In_2200);
and U565 (N_565,N_187,In_91);
xnor U566 (N_566,N_256,In_1131);
and U567 (N_567,In_2418,In_1659);
nor U568 (N_568,N_36,N_64);
and U569 (N_569,In_1584,In_2061);
xnor U570 (N_570,N_285,In_1431);
xor U571 (N_571,In_314,In_22);
xnor U572 (N_572,In_1986,In_679);
or U573 (N_573,In_1499,In_1517);
xor U574 (N_574,In_487,In_1600);
xnor U575 (N_575,In_1227,N_485);
nand U576 (N_576,In_527,In_1311);
nand U577 (N_577,In_604,In_1565);
and U578 (N_578,In_116,In_169);
nor U579 (N_579,In_1917,In_1039);
xor U580 (N_580,N_442,In_1540);
nor U581 (N_581,In_981,N_449);
nand U582 (N_582,N_0,N_185);
xor U583 (N_583,In_2237,N_210);
and U584 (N_584,N_459,N_261);
or U585 (N_585,In_1313,In_655);
nand U586 (N_586,In_2179,N_460);
and U587 (N_587,In_240,In_1500);
nor U588 (N_588,In_1270,In_440);
nand U589 (N_589,N_315,In_1933);
or U590 (N_590,N_8,In_1206);
xnor U591 (N_591,In_1494,In_1530);
xnor U592 (N_592,In_2269,In_2180);
and U593 (N_593,In_61,In_889);
nand U594 (N_594,In_1315,In_1253);
and U595 (N_595,In_34,In_185);
nor U596 (N_596,In_2076,N_231);
and U597 (N_597,N_481,In_994);
nor U598 (N_598,In_1877,N_330);
xnor U599 (N_599,In_1548,N_457);
nand U600 (N_600,N_447,In_419);
xor U601 (N_601,In_475,N_414);
nor U602 (N_602,In_1894,N_403);
nor U603 (N_603,In_1691,In_1066);
and U604 (N_604,In_556,In_1433);
xnor U605 (N_605,In_1814,N_52);
nand U606 (N_606,N_421,In_114);
or U607 (N_607,N_296,N_129);
nand U608 (N_608,In_117,N_338);
and U609 (N_609,In_2147,N_398);
xor U610 (N_610,In_2474,In_666);
or U611 (N_611,In_1938,In_761);
or U612 (N_612,N_401,In_266);
or U613 (N_613,In_1097,N_66);
or U614 (N_614,N_440,N_488);
and U615 (N_615,In_1518,N_132);
xor U616 (N_616,N_117,In_1636);
or U617 (N_617,N_308,N_395);
nor U618 (N_618,In_2356,In_233);
xnor U619 (N_619,N_139,In_804);
nand U620 (N_620,N_441,N_342);
nand U621 (N_621,In_1564,N_275);
or U622 (N_622,In_248,In_1279);
or U623 (N_623,In_1142,N_375);
nor U624 (N_624,In_2103,N_183);
xor U625 (N_625,In_217,In_145);
xor U626 (N_626,In_637,In_1181);
or U627 (N_627,In_2098,In_1709);
nor U628 (N_628,In_2339,In_2301);
nand U629 (N_629,In_2159,In_99);
and U630 (N_630,In_478,In_1906);
xor U631 (N_631,N_19,N_383);
nand U632 (N_632,In_1139,In_681);
and U633 (N_633,In_693,In_1465);
or U634 (N_634,In_468,In_1402);
nand U635 (N_635,In_1562,In_1332);
or U636 (N_636,In_2325,In_1800);
xnor U637 (N_637,N_326,In_561);
and U638 (N_638,In_1005,In_1217);
or U639 (N_639,In_2170,In_1088);
nand U640 (N_640,In_1802,N_492);
nand U641 (N_641,In_881,In_877);
nor U642 (N_642,In_1919,In_995);
nor U643 (N_643,N_4,N_232);
and U644 (N_644,In_899,In_1231);
nor U645 (N_645,In_2130,N_404);
or U646 (N_646,In_1022,N_450);
nor U647 (N_647,In_619,In_1741);
and U648 (N_648,In_2085,In_250);
nor U649 (N_649,In_278,In_605);
xor U650 (N_650,N_408,In_741);
and U651 (N_651,In_1697,In_2451);
nor U652 (N_652,In_2212,N_65);
nand U653 (N_653,In_1713,In_1823);
and U654 (N_654,In_1704,N_76);
or U655 (N_655,In_1857,In_14);
and U656 (N_656,In_92,In_1020);
or U657 (N_657,In_1590,In_2467);
nor U658 (N_658,In_1700,In_1067);
nor U659 (N_659,In_199,N_95);
or U660 (N_660,N_252,In_1362);
xor U661 (N_661,In_538,In_553);
nor U662 (N_662,N_156,In_128);
nor U663 (N_663,In_225,In_1129);
xnor U664 (N_664,In_312,In_42);
xnor U665 (N_665,In_866,In_2287);
or U666 (N_666,In_1363,In_1447);
nor U667 (N_667,In_816,In_288);
or U668 (N_668,In_948,N_493);
xnor U669 (N_669,In_1137,N_100);
nor U670 (N_670,In_486,In_67);
nor U671 (N_671,In_1179,In_346);
or U672 (N_672,N_116,In_758);
nand U673 (N_673,In_783,In_1348);
or U674 (N_674,N_146,N_314);
xnor U675 (N_675,N_295,N_51);
or U676 (N_676,In_2227,In_805);
nor U677 (N_677,In_1605,In_1974);
xnor U678 (N_678,In_2420,In_198);
nor U679 (N_679,N_118,In_1809);
or U680 (N_680,In_1905,In_1234);
xnor U681 (N_681,In_645,In_703);
nand U682 (N_682,In_462,In_2074);
and U683 (N_683,In_2298,In_2464);
nor U684 (N_684,In_1096,In_1688);
nor U685 (N_685,N_328,In_2096);
xor U686 (N_686,In_846,In_1003);
nor U687 (N_687,In_617,N_390);
xor U688 (N_688,N_159,In_1116);
nand U689 (N_689,In_1098,In_723);
or U690 (N_690,In_1305,N_486);
and U691 (N_691,In_2381,N_271);
xnor U692 (N_692,In_1176,In_1640);
xnor U693 (N_693,N_74,In_2015);
or U694 (N_694,In_1120,In_1144);
or U695 (N_695,In_2252,N_389);
or U696 (N_696,In_2488,In_1080);
nor U697 (N_697,In_1259,N_294);
or U698 (N_698,N_287,In_716);
nor U699 (N_699,In_1639,In_2157);
xnor U700 (N_700,N_202,N_175);
or U701 (N_701,In_1008,In_915);
nand U702 (N_702,In_907,N_145);
nor U703 (N_703,In_2062,In_1141);
and U704 (N_704,N_22,N_130);
and U705 (N_705,In_1544,N_428);
or U706 (N_706,In_1845,In_2221);
and U707 (N_707,N_290,N_439);
and U708 (N_708,In_1795,In_729);
or U709 (N_709,In_642,N_173);
and U710 (N_710,In_1865,N_142);
nor U711 (N_711,In_707,In_2161);
xor U712 (N_712,N_433,N_335);
and U713 (N_713,In_1535,In_1730);
nor U714 (N_714,N_140,In_1966);
or U715 (N_715,N_343,In_1117);
xnor U716 (N_716,In_2446,In_1289);
and U717 (N_717,In_506,In_139);
and U718 (N_718,In_2226,In_21);
nor U719 (N_719,In_1337,In_405);
nand U720 (N_720,N_240,In_65);
xnor U721 (N_721,In_1112,In_520);
or U722 (N_722,In_615,N_371);
nand U723 (N_723,N_1,N_300);
and U724 (N_724,N_49,In_1383);
or U725 (N_725,In_2485,N_276);
xnor U726 (N_726,In_1165,N_54);
or U727 (N_727,In_1412,In_496);
nor U728 (N_728,N_6,In_766);
nand U729 (N_729,In_184,In_151);
and U730 (N_730,In_162,In_769);
nor U731 (N_731,In_2472,N_196);
nand U732 (N_732,In_1262,In_700);
or U733 (N_733,In_1758,In_430);
xnor U734 (N_734,N_413,N_364);
xor U735 (N_735,In_373,In_542);
xnor U736 (N_736,N_124,N_362);
nand U737 (N_737,In_1526,In_861);
or U738 (N_738,N_346,In_865);
nand U739 (N_739,In_1203,In_1866);
or U740 (N_740,In_1189,In_452);
and U741 (N_741,In_476,In_2022);
xnor U742 (N_742,In_786,N_244);
or U743 (N_743,In_474,In_1333);
nor U744 (N_744,In_83,In_952);
or U745 (N_745,N_127,In_931);
nand U746 (N_746,In_2219,In_1759);
nor U747 (N_747,N_416,In_1038);
or U748 (N_748,In_422,N_192);
and U749 (N_749,N_289,In_2456);
nand U750 (N_750,In_813,N_205);
xor U751 (N_751,N_250,In_164);
xnor U752 (N_752,N_102,In_1444);
or U753 (N_753,In_1366,In_1398);
xnor U754 (N_754,In_441,In_297);
or U755 (N_755,N_253,In_887);
nand U756 (N_756,In_2297,N_238);
xor U757 (N_757,In_2386,In_121);
nand U758 (N_758,In_363,In_327);
nand U759 (N_759,N_111,In_1335);
nand U760 (N_760,In_2038,In_548);
and U761 (N_761,In_576,In_1921);
xnor U762 (N_762,In_768,N_128);
or U763 (N_763,N_360,In_1331);
or U764 (N_764,N_291,In_2135);
and U765 (N_765,In_534,In_1326);
and U766 (N_766,N_226,In_1420);
nor U767 (N_767,In_1504,N_47);
nor U768 (N_768,In_89,N_24);
nor U769 (N_769,N_464,In_1832);
and U770 (N_770,N_327,In_2337);
xor U771 (N_771,N_61,In_2313);
or U772 (N_772,N_147,In_1643);
or U773 (N_773,In_815,N_170);
nand U774 (N_774,In_996,N_265);
nand U775 (N_775,In_1030,In_13);
xor U776 (N_776,In_1641,In_1745);
nand U777 (N_777,In_1325,In_1086);
and U778 (N_778,In_1065,In_52);
xor U779 (N_779,N_482,In_852);
nor U780 (N_780,In_1457,In_1477);
nand U781 (N_781,In_567,In_2334);
or U782 (N_782,In_1048,In_2318);
xnor U783 (N_783,In_1609,In_1031);
and U784 (N_784,In_612,N_163);
nand U785 (N_785,N_427,In_2439);
xnor U786 (N_786,N_366,In_2016);
nand U787 (N_787,In_721,In_1678);
nor U788 (N_788,In_757,In_2362);
xnor U789 (N_789,In_1506,In_1024);
or U790 (N_790,In_2168,In_1346);
nand U791 (N_791,In_1058,In_1976);
nor U792 (N_792,In_1269,In_1901);
nor U793 (N_793,N_99,In_1984);
or U794 (N_794,In_129,In_1852);
or U795 (N_795,In_1498,In_1907);
xnor U796 (N_796,N_425,In_855);
nand U797 (N_797,In_1575,In_1395);
xor U798 (N_798,In_85,In_1651);
and U799 (N_799,In_2108,N_472);
xnor U800 (N_800,In_1273,In_1368);
nor U801 (N_801,N_350,In_867);
nand U802 (N_802,In_727,In_2052);
and U803 (N_803,N_358,In_2146);
or U804 (N_804,In_1764,In_1769);
nor U805 (N_805,N_153,N_138);
or U806 (N_806,In_789,In_2027);
or U807 (N_807,In_201,N_94);
xnor U808 (N_808,In_1722,N_131);
and U809 (N_809,In_2175,In_142);
or U810 (N_810,In_2145,In_132);
and U811 (N_811,In_1962,In_1529);
nand U812 (N_812,In_1215,In_874);
nor U813 (N_813,N_25,In_309);
nor U814 (N_814,N_432,N_206);
nor U815 (N_815,N_230,In_1645);
xor U816 (N_816,In_706,N_179);
nor U817 (N_817,In_1862,In_1853);
and U818 (N_818,In_689,In_825);
nand U819 (N_819,In_577,In_1944);
or U820 (N_820,N_334,In_100);
xor U821 (N_821,In_1687,N_467);
and U822 (N_822,N_496,In_2448);
nand U823 (N_823,In_2417,In_1119);
and U824 (N_824,N_103,In_398);
or U825 (N_825,In_2216,In_715);
or U826 (N_826,In_456,N_325);
or U827 (N_827,In_249,In_1930);
and U828 (N_828,In_160,N_166);
and U829 (N_829,N_473,In_1929);
xor U830 (N_830,In_1598,In_1111);
xor U831 (N_831,N_286,In_671);
nor U832 (N_832,In_1439,N_209);
xnor U833 (N_833,In_510,In_1079);
and U834 (N_834,In_1653,In_2396);
nor U835 (N_835,In_1644,In_2312);
and U836 (N_836,In_1171,N_197);
and U837 (N_837,In_1461,In_1627);
or U838 (N_838,N_53,In_1293);
and U839 (N_839,In_746,N_10);
and U840 (N_840,In_24,N_181);
and U841 (N_841,In_2352,In_2142);
xor U842 (N_842,In_286,In_1436);
xor U843 (N_843,In_255,N_58);
nor U844 (N_844,N_266,In_683);
nor U845 (N_845,N_426,In_1476);
nor U846 (N_846,In_570,In_2189);
and U847 (N_847,In_1545,In_796);
xor U848 (N_848,N_303,In_84);
xor U849 (N_849,In_1729,In_1631);
xor U850 (N_850,N_461,In_1666);
or U851 (N_851,In_1236,In_691);
or U852 (N_852,N_44,In_1469);
nand U853 (N_853,In_357,In_2023);
nand U854 (N_854,In_2428,In_2026);
nand U855 (N_855,N_466,In_578);
nor U856 (N_856,In_1637,In_2019);
or U857 (N_857,In_115,In_1940);
or U858 (N_858,In_47,In_2465);
and U859 (N_859,N_284,In_1235);
nor U860 (N_860,In_318,N_137);
and U861 (N_861,In_734,N_370);
nand U862 (N_862,N_498,N_487);
or U863 (N_863,In_760,In_484);
or U864 (N_864,In_1188,In_105);
and U865 (N_865,In_862,In_209);
nand U866 (N_866,In_414,N_106);
xor U867 (N_867,In_444,In_1554);
nor U868 (N_868,In_1867,In_742);
nand U869 (N_869,In_1547,In_1275);
and U870 (N_870,In_1912,In_280);
nor U871 (N_871,N_304,In_1384);
nor U872 (N_872,N_50,In_53);
nand U873 (N_873,In_751,N_236);
or U874 (N_874,In_2289,N_424);
nor U875 (N_875,In_1925,In_315);
and U876 (N_876,In_1567,N_107);
or U877 (N_877,In_516,In_2182);
or U878 (N_878,In_1796,In_370);
xnor U879 (N_879,In_1546,In_235);
nor U880 (N_880,N_302,In_1817);
nor U881 (N_881,N_444,In_1474);
xnor U882 (N_882,N_38,N_422);
xnor U883 (N_883,N_406,In_1897);
nor U884 (N_884,In_1379,In_2379);
nand U885 (N_885,In_97,In_36);
xor U886 (N_886,In_901,In_2311);
and U887 (N_887,In_989,In_1193);
nand U888 (N_888,In_1076,In_15);
nand U889 (N_889,In_1964,N_478);
nand U890 (N_890,In_2242,In_807);
xor U891 (N_891,N_476,In_479);
xnor U892 (N_892,In_582,In_571);
or U893 (N_893,In_1244,In_424);
xor U894 (N_894,In_134,N_15);
nor U895 (N_895,In_1994,In_339);
nor U896 (N_896,In_1145,In_1725);
nand U897 (N_897,In_1628,In_2039);
and U898 (N_898,In_1035,N_313);
or U899 (N_899,In_967,In_63);
xor U900 (N_900,In_997,N_222);
nor U901 (N_901,In_913,In_945);
nor U902 (N_902,In_2132,In_2106);
and U903 (N_903,N_320,In_1225);
and U904 (N_904,In_682,In_1785);
xor U905 (N_905,In_613,In_2371);
nor U906 (N_906,N_434,In_752);
nor U907 (N_907,In_1572,In_1773);
nand U908 (N_908,In_1200,In_1085);
nand U909 (N_909,In_450,N_195);
nand U910 (N_910,In_2153,In_140);
and U911 (N_911,In_549,In_148);
or U912 (N_912,In_257,N_430);
or U913 (N_913,In_375,N_471);
xor U914 (N_914,N_489,N_341);
and U915 (N_915,In_1868,In_2273);
and U916 (N_916,In_70,In_446);
or U917 (N_917,N_233,In_1902);
and U918 (N_918,In_1646,In_1859);
nor U919 (N_919,In_744,N_158);
xnor U920 (N_920,In_76,In_179);
nor U921 (N_921,N_263,In_2476);
nor U922 (N_922,In_2340,In_778);
nand U923 (N_923,N_193,In_745);
and U924 (N_924,In_2331,In_1634);
nor U925 (N_925,In_530,In_2246);
and U926 (N_926,In_2012,N_160);
nor U927 (N_927,N_438,In_1344);
and U928 (N_928,In_951,In_1419);
nand U929 (N_929,N_151,In_1630);
or U930 (N_930,In_511,In_911);
or U931 (N_931,In_51,In_2143);
nand U932 (N_932,In_1831,In_2010);
xnor U933 (N_933,N_136,N_39);
xor U934 (N_934,N_497,In_1515);
nor U935 (N_935,N_121,In_1550);
or U936 (N_936,In_684,In_2171);
xnor U937 (N_937,In_2152,In_1104);
xnor U938 (N_938,In_2390,In_1807);
nand U939 (N_939,In_1422,In_1682);
nor U940 (N_940,In_739,In_2410);
nand U941 (N_941,In_282,In_1985);
nor U942 (N_942,In_1257,In_2223);
nor U943 (N_943,N_495,In_2148);
nor U944 (N_944,In_2413,In_2099);
nor U945 (N_945,N_483,In_2496);
nor U946 (N_946,N_355,In_133);
or U947 (N_947,In_651,In_728);
and U948 (N_948,In_1063,In_1740);
nor U949 (N_949,In_2088,In_1958);
xor U950 (N_950,N_91,N_186);
and U951 (N_951,N_446,In_379);
and U952 (N_952,N_259,In_323);
xor U953 (N_953,N_45,In_801);
nand U954 (N_954,In_428,In_2044);
or U955 (N_955,In_969,In_635);
or U956 (N_956,In_1592,In_1815);
xnor U957 (N_957,In_978,In_1256);
and U958 (N_958,In_1356,In_2124);
nor U959 (N_959,In_155,In_1882);
and U960 (N_960,In_630,In_1016);
or U961 (N_961,N_216,In_203);
xnor U962 (N_962,In_1185,In_136);
xnor U963 (N_963,In_112,In_1516);
nand U964 (N_964,In_1618,N_292);
and U965 (N_965,N_148,In_1752);
xor U966 (N_966,In_75,N_46);
or U967 (N_967,In_2014,N_268);
nand U968 (N_968,N_469,N_387);
nor U969 (N_969,In_643,In_1900);
nor U970 (N_970,In_1707,N_68);
and U971 (N_971,In_2498,In_2217);
nor U972 (N_972,In_29,In_1483);
or U973 (N_973,N_316,In_1596);
or U974 (N_974,N_78,In_2238);
or U975 (N_975,In_1957,In_1963);
and U976 (N_976,N_200,In_1164);
or U977 (N_977,In_2043,In_301);
xor U978 (N_978,In_1671,N_356);
nor U979 (N_979,In_555,In_371);
nand U980 (N_980,N_96,In_2231);
xnor U981 (N_981,N_270,In_1997);
xnor U982 (N_982,In_2040,In_138);
or U983 (N_983,In_270,N_63);
nor U984 (N_984,N_384,In_857);
xor U985 (N_985,In_86,In_764);
nand U986 (N_986,N_247,In_1296);
xnor U987 (N_987,In_1438,In_1061);
or U988 (N_988,In_1808,In_431);
nand U989 (N_989,In_2047,In_2190);
nor U990 (N_990,N_135,In_1342);
nand U991 (N_991,In_1612,N_351);
nor U992 (N_992,N_69,N_171);
nor U993 (N_993,In_1329,In_2116);
nor U994 (N_994,In_986,In_1775);
or U995 (N_995,In_1378,In_1094);
nor U996 (N_996,In_2028,In_74);
or U997 (N_997,In_2196,In_1977);
or U998 (N_998,In_2109,In_928);
xnor U999 (N_999,In_1576,In_1056);
xor U1000 (N_1000,In_205,N_697);
xor U1001 (N_1001,N_720,In_1282);
nor U1002 (N_1002,In_557,In_1455);
or U1003 (N_1003,In_2415,N_623);
nand U1004 (N_1004,N_722,In_1842);
and U1005 (N_1005,In_717,N_608);
nand U1006 (N_1006,N_919,N_747);
nand U1007 (N_1007,N_738,N_393);
or U1008 (N_1008,In_965,N_721);
nor U1009 (N_1009,In_600,N_77);
nor U1010 (N_1010,In_1109,In_1711);
xnor U1011 (N_1011,In_2118,In_875);
and U1012 (N_1012,N_735,In_298);
xor U1013 (N_1013,N_982,In_748);
xnor U1014 (N_1014,In_2323,N_27);
nor U1015 (N_1015,N_357,N_348);
nor U1016 (N_1016,N_905,N_776);
or U1017 (N_1017,N_685,In_914);
xnor U1018 (N_1018,N_775,N_614);
xnor U1019 (N_1019,In_990,N_992);
nor U1020 (N_1020,N_853,In_2224);
or U1021 (N_1021,In_696,In_1561);
nor U1022 (N_1022,N_612,N_784);
or U1023 (N_1023,N_758,N_517);
and U1024 (N_1024,In_144,In_378);
nand U1025 (N_1025,N_693,N_182);
xor U1026 (N_1026,In_2466,In_2380);
nor U1027 (N_1027,In_1365,In_828);
nand U1028 (N_1028,In_1382,N_576);
nor U1029 (N_1029,In_2477,N_981);
and U1030 (N_1030,In_1878,In_2304);
or U1031 (N_1031,In_1307,N_840);
or U1032 (N_1032,N_764,In_834);
and U1033 (N_1033,In_690,In_521);
or U1034 (N_1034,In_1018,In_1762);
xnor U1035 (N_1035,In_2473,In_1871);
xor U1036 (N_1036,In_523,In_489);
xnor U1037 (N_1037,In_2204,In_1553);
nor U1038 (N_1038,N_709,In_299);
nand U1039 (N_1039,In_1426,N_983);
or U1040 (N_1040,N_376,N_9);
or U1041 (N_1041,In_1573,N_499);
or U1042 (N_1042,N_746,N_803);
xnor U1043 (N_1043,In_2185,In_2263);
nor U1044 (N_1044,N_324,In_2445);
nand U1045 (N_1045,In_1524,N_896);
or U1046 (N_1046,N_698,In_551);
nor U1047 (N_1047,In_1610,In_1998);
and U1048 (N_1048,In_1019,In_1051);
or U1049 (N_1049,N_543,N_322);
or U1050 (N_1050,In_1297,In_295);
nand U1051 (N_1051,In_2268,In_1563);
and U1052 (N_1052,N_592,N_752);
xor U1053 (N_1053,In_2351,N_934);
xnor U1054 (N_1054,N_959,In_868);
nand U1055 (N_1055,N_914,In_1258);
or U1056 (N_1056,N_152,In_2001);
xor U1057 (N_1057,In_392,In_1899);
nor U1058 (N_1058,In_2057,In_934);
xor U1059 (N_1059,In_2275,N_966);
nor U1060 (N_1060,N_180,N_506);
xnor U1061 (N_1061,In_1492,In_226);
nand U1062 (N_1062,In_2234,N_680);
and U1063 (N_1063,In_101,In_1880);
xor U1064 (N_1064,In_1608,In_1046);
xnor U1065 (N_1065,In_1497,N_386);
and U1066 (N_1066,In_1858,In_1415);
nand U1067 (N_1067,In_1675,In_1969);
or U1068 (N_1068,In_1194,N_306);
xnor U1069 (N_1069,In_1916,N_579);
nor U1070 (N_1070,N_832,N_643);
or U1071 (N_1071,N_807,N_655);
nor U1072 (N_1072,N_906,In_871);
xnor U1073 (N_1073,In_730,N_177);
and U1074 (N_1074,N_388,In_1255);
nand U1075 (N_1075,N_400,N_804);
and U1076 (N_1076,In_1647,N_7);
or U1077 (N_1077,N_670,In_1212);
nor U1078 (N_1078,N_321,In_1632);
nand U1079 (N_1079,N_379,In_838);
nor U1080 (N_1080,In_1134,In_1793);
or U1081 (N_1081,In_181,In_587);
or U1082 (N_1082,In_1140,N_730);
xnor U1083 (N_1083,N_18,In_795);
nor U1084 (N_1084,N_436,N_453);
nand U1085 (N_1085,N_668,N_921);
xor U1086 (N_1086,N_108,N_14);
xor U1087 (N_1087,In_1863,N_604);
or U1088 (N_1088,N_845,In_417);
or U1089 (N_1089,In_2453,N_550);
nor U1090 (N_1090,N_548,N_767);
xor U1091 (N_1091,N_35,N_353);
xnor U1092 (N_1092,In_59,N_590);
and U1093 (N_1093,N_652,In_1159);
nor U1094 (N_1094,In_1394,N_277);
and U1095 (N_1095,In_2065,N_560);
or U1096 (N_1096,N_766,In_2127);
xor U1097 (N_1097,In_2434,In_206);
nand U1098 (N_1098,In_152,In_830);
xor U1099 (N_1099,In_956,In_938);
xor U1100 (N_1100,In_1449,In_1683);
and U1101 (N_1101,N_797,N_134);
or U1102 (N_1102,N_529,In_1478);
or U1103 (N_1103,In_1537,N_794);
nand U1104 (N_1104,N_28,N_513);
xnor U1105 (N_1105,N_671,N_542);
or U1106 (N_1106,In_832,N_318);
nand U1107 (N_1107,In_1622,N_336);
xor U1108 (N_1108,In_2113,N_834);
or U1109 (N_1109,N_369,In_293);
and U1110 (N_1110,In_494,N_971);
nor U1111 (N_1111,N_331,In_2427);
nor U1112 (N_1112,In_1155,N_955);
nand U1113 (N_1113,N_616,N_228);
and U1114 (N_1114,N_569,N_815);
xnor U1115 (N_1115,In_1199,N_556);
nand U1116 (N_1116,N_41,N_635);
xnor U1117 (N_1117,In_2158,N_16);
and U1118 (N_1118,In_1442,In_1790);
nor U1119 (N_1119,N_915,N_637);
xor U1120 (N_1120,N_559,N_11);
nand U1121 (N_1121,N_726,In_1357);
or U1122 (N_1122,N_239,N_667);
and U1123 (N_1123,In_146,N_407);
or U1124 (N_1124,In_380,In_599);
and U1125 (N_1125,In_947,N_282);
and U1126 (N_1126,N_194,In_803);
or U1127 (N_1127,In_608,N_920);
nand U1128 (N_1128,In_1701,N_880);
nor U1129 (N_1129,N_164,In_1042);
nor U1130 (N_1130,N_659,N_23);
nand U1131 (N_1131,N_970,N_565);
and U1132 (N_1132,N_742,In_650);
nand U1133 (N_1133,In_260,N_765);
and U1134 (N_1134,N_823,N_88);
nand U1135 (N_1135,N_748,N_241);
or U1136 (N_1136,N_123,In_2239);
or U1137 (N_1137,N_311,In_1043);
or U1138 (N_1138,N_507,N_973);
nand U1139 (N_1139,In_159,N_777);
nor U1140 (N_1140,N_562,In_2054);
and U1141 (N_1141,N_694,N_257);
xor U1142 (N_1142,N_681,In_697);
xnor U1143 (N_1143,N_227,N_307);
xnor U1144 (N_1144,N_938,In_2256);
nor U1145 (N_1145,N_533,In_1768);
nor U1146 (N_1146,In_1448,N_339);
or U1147 (N_1147,In_1927,N_620);
and U1148 (N_1148,In_644,N_452);
xor U1149 (N_1149,In_2067,In_2013);
nand U1150 (N_1150,N_429,N_312);
xor U1151 (N_1151,N_377,N_660);
nor U1152 (N_1152,In_973,N_969);
and U1153 (N_1153,N_855,In_2129);
xnor U1154 (N_1154,N_741,N_885);
nand U1155 (N_1155,In_1069,N_817);
nor U1156 (N_1156,In_1835,In_1306);
nor U1157 (N_1157,In_130,In_2478);
or U1158 (N_1158,In_568,N_254);
or U1159 (N_1159,In_1784,In_1470);
nand U1160 (N_1160,In_141,N_26);
nor U1161 (N_1161,In_2302,In_345);
nor U1162 (N_1162,In_2053,N_684);
xor U1163 (N_1163,N_624,In_58);
or U1164 (N_1164,In_2255,N_229);
or U1165 (N_1165,In_48,In_1737);
xor U1166 (N_1166,In_1351,N_273);
nand U1167 (N_1167,N_524,In_541);
and U1168 (N_1168,N_126,N_979);
nand U1169 (N_1169,N_848,N_781);
or U1170 (N_1170,In_351,N_699);
and U1171 (N_1171,In_393,In_1174);
or U1172 (N_1172,In_941,In_1396);
and U1173 (N_1173,N_947,In_2457);
nor U1174 (N_1174,N_782,In_1840);
nor U1175 (N_1175,N_965,N_262);
xor U1176 (N_1176,N_898,N_154);
and U1177 (N_1177,In_2084,N_778);
nor U1178 (N_1178,N_999,In_844);
xor U1179 (N_1179,In_1360,In_1172);
and U1180 (N_1180,In_1965,In_1534);
or U1181 (N_1181,N_79,In_2123);
or U1182 (N_1182,In_1816,N_603);
xnor U1183 (N_1183,N_625,N_639);
or U1184 (N_1184,In_328,N_902);
xnor U1185 (N_1185,In_1923,N_858);
xor U1186 (N_1186,In_560,N_223);
nand U1187 (N_1187,In_2131,In_32);
or U1188 (N_1188,N_892,N_673);
nor U1189 (N_1189,In_626,N_913);
xnor U1190 (N_1190,N_208,In_33);
xnor U1191 (N_1191,N_928,In_1252);
and U1192 (N_1192,In_711,N_869);
and U1193 (N_1193,N_234,N_93);
nor U1194 (N_1194,In_649,In_787);
nor U1195 (N_1195,In_2244,In_2300);
nor U1196 (N_1196,N_645,In_1192);
and U1197 (N_1197,N_372,N_618);
nor U1198 (N_1198,In_2107,N_829);
nor U1199 (N_1199,In_1656,N_930);
xor U1200 (N_1200,N_198,N_456);
nand U1201 (N_1201,In_1184,In_1148);
or U1202 (N_1202,In_214,In_2059);
or U1203 (N_1203,In_1621,In_2407);
and U1204 (N_1204,In_1414,N_566);
nand U1205 (N_1205,In_1219,N_155);
or U1206 (N_1206,In_1454,In_1146);
nor U1207 (N_1207,N_367,N_235);
nor U1208 (N_1208,N_883,N_801);
or U1209 (N_1209,In_1777,In_1432);
nand U1210 (N_1210,In_2361,N_585);
and U1211 (N_1211,N_831,In_933);
and U1212 (N_1212,In_399,In_329);
and U1213 (N_1213,N_281,N_75);
xnor U1214 (N_1214,In_1501,N_873);
nand U1215 (N_1215,In_1464,N_864);
and U1216 (N_1216,N_633,In_1786);
or U1217 (N_1217,N_783,In_633);
and U1218 (N_1218,In_1341,N_991);
or U1219 (N_1219,In_2486,N_544);
nand U1220 (N_1220,N_458,In_503);
nor U1221 (N_1221,N_944,N_705);
xor U1222 (N_1222,N_675,In_606);
xor U1223 (N_1223,N_551,N_770);
xnor U1224 (N_1224,N_329,N_588);
or U1225 (N_1225,N_711,In_2310);
or U1226 (N_1226,N_691,In_1451);
nor U1227 (N_1227,N_477,In_2367);
xor U1228 (N_1228,In_131,In_704);
xnor U1229 (N_1229,In_37,N_836);
nand U1230 (N_1230,In_224,N_534);
nand U1231 (N_1231,In_676,N_634);
nand U1232 (N_1232,N_70,N_820);
nor U1233 (N_1233,In_449,In_1191);
and U1234 (N_1234,In_1952,N_217);
and U1235 (N_1235,In_360,N_237);
nand U1236 (N_1236,In_1186,N_710);
or U1237 (N_1237,In_2480,N_954);
nor U1238 (N_1238,N_610,In_2154);
and U1239 (N_1239,In_320,In_1751);
xor U1240 (N_1240,N_851,N_808);
nand U1241 (N_1241,In_1209,N_184);
or U1242 (N_1242,N_736,N_215);
xnor U1243 (N_1243,In_2330,In_1274);
nor U1244 (N_1244,In_2265,In_436);
and U1245 (N_1245,In_1265,In_2424);
or U1246 (N_1246,N_526,In_1935);
xnor U1247 (N_1247,N_98,In_2405);
and U1248 (N_1248,N_798,N_886);
nand U1249 (N_1249,N_475,N_859);
or U1250 (N_1250,N_615,In_1980);
or U1251 (N_1251,In_95,In_273);
xnor U1252 (N_1252,In_460,In_4);
and U1253 (N_1253,In_735,N_702);
or U1254 (N_1254,In_182,N_664);
and U1255 (N_1255,In_1949,In_1237);
and U1256 (N_1256,N_586,In_2139);
nand U1257 (N_1257,In_590,N_31);
or U1258 (N_1258,N_391,N_712);
nor U1259 (N_1259,N_714,In_2160);
xor U1260 (N_1260,N_941,N_964);
and U1261 (N_1261,In_1445,In_1317);
and U1262 (N_1262,N_950,N_723);
or U1263 (N_1263,In_1616,N_110);
nor U1264 (N_1264,N_825,N_37);
and U1265 (N_1265,N_649,N_884);
nand U1266 (N_1266,In_368,In_896);
nor U1267 (N_1267,In_1283,N_528);
nand U1268 (N_1268,In_1374,In_1475);
and U1269 (N_1269,N_508,N_933);
nor U1270 (N_1270,In_1288,In_2369);
or U1271 (N_1271,In_2066,In_629);
nor U1272 (N_1272,N_169,In_847);
and U1273 (N_1273,In_272,In_1932);
nand U1274 (N_1274,N_800,N_986);
xor U1275 (N_1275,In_470,In_2000);
or U1276 (N_1276,N_953,In_705);
nand U1277 (N_1277,In_1679,In_1389);
nand U1278 (N_1278,N_267,N_852);
or U1279 (N_1279,N_812,N_935);
nor U1280 (N_1280,N_305,In_2319);
or U1281 (N_1281,In_1320,In_584);
or U1282 (N_1282,N_490,N_299);
xnor U1283 (N_1283,In_435,N_220);
nor U1284 (N_1284,In_1889,In_1993);
and U1285 (N_1285,In_2101,In_397);
nand U1286 (N_1286,N_857,N_512);
or U1287 (N_1287,N_629,In_839);
nor U1288 (N_1288,N_665,N_465);
xnor U1289 (N_1289,In_673,N_990);
nand U1290 (N_1290,N_753,N_862);
and U1291 (N_1291,In_925,N_822);
nand U1292 (N_1292,N_443,N_703);
nand U1293 (N_1293,N_337,N_246);
and U1294 (N_1294,In_2274,In_409);
or U1295 (N_1295,N_575,In_1543);
xor U1296 (N_1296,In_793,In_944);
or U1297 (N_1297,In_454,N_73);
nand U1298 (N_1298,N_658,N_359);
or U1299 (N_1299,In_2375,N_587);
or U1300 (N_1300,N_638,N_448);
nand U1301 (N_1301,In_244,In_895);
xor U1302 (N_1302,N_708,In_2324);
or U1303 (N_1303,N_577,In_618);
or U1304 (N_1304,In_1607,N_30);
nand U1305 (N_1305,In_310,In_1312);
and U1306 (N_1306,In_1673,In_425);
or U1307 (N_1307,In_377,N_651);
xnor U1308 (N_1308,N_686,N_793);
nor U1309 (N_1309,N_850,N_662);
nor U1310 (N_1310,N_397,N_455);
and U1311 (N_1311,N_502,In_2009);
xor U1312 (N_1312,In_183,N_922);
xor U1313 (N_1313,In_1887,N_500);
nor U1314 (N_1314,N_162,In_87);
and U1315 (N_1315,N_841,In_2314);
nand U1316 (N_1316,N_863,In_2422);
xor U1317 (N_1317,In_809,In_2450);
or U1318 (N_1318,In_2442,N_945);
xor U1319 (N_1319,In_2220,In_354);
xnor U1320 (N_1320,In_2064,In_153);
nand U1321 (N_1321,N_809,In_1322);
xor U1322 (N_1322,In_1205,In_660);
nand U1323 (N_1323,In_1210,N_994);
xnor U1324 (N_1324,In_2150,In_358);
and U1325 (N_1325,N_641,N_656);
or U1326 (N_1326,In_98,In_657);
or U1327 (N_1327,In_1804,In_498);
xnor U1328 (N_1328,In_296,N_925);
nor U1329 (N_1329,N_535,In_2328);
xnor U1330 (N_1330,N_203,In_448);
nand U1331 (N_1331,N_87,In_1915);
and U1332 (N_1332,N_737,N_996);
nand U1333 (N_1333,N_597,In_674);
and U1334 (N_1334,In_2419,In_2025);
nor U1335 (N_1335,N_917,In_178);
nand U1336 (N_1336,N_849,N_71);
xor U1337 (N_1337,N_189,In_854);
xnor U1338 (N_1338,N_90,N_805);
nand U1339 (N_1339,In_908,N_125);
and U1340 (N_1340,N_437,In_104);
nor U1341 (N_1341,In_2213,N_530);
xnor U1342 (N_1342,N_689,In_304);
nor U1343 (N_1343,In_1703,In_1082);
xnor U1344 (N_1344,N_525,In_596);
or U1345 (N_1345,N_600,N_547);
nor U1346 (N_1346,N_672,N_901);
and U1347 (N_1347,In_2335,In_891);
and U1348 (N_1348,N_679,In_1314);
and U1349 (N_1349,In_2322,In_2487);
nor U1350 (N_1350,In_753,In_1910);
and U1351 (N_1351,N_875,In_784);
xnor U1352 (N_1352,N_821,N_283);
nand U1353 (N_1353,N_62,N_120);
and U1354 (N_1354,N_549,N_647);
xor U1355 (N_1355,In_1358,In_1552);
nor U1356 (N_1356,In_2326,In_231);
xnor U1357 (N_1357,N_595,In_1726);
xor U1358 (N_1358,In_2293,In_176);
or U1359 (N_1359,In_382,N_580);
or U1360 (N_1360,In_1908,In_653);
xor U1361 (N_1361,N_468,N_317);
nor U1362 (N_1362,In_686,N_509);
xnor U1363 (N_1363,In_898,In_942);
nand U1364 (N_1364,In_988,In_220);
and U1365 (N_1365,In_1271,In_284);
nand U1366 (N_1366,N_792,N_17);
and U1367 (N_1367,In_1723,In_1847);
nand U1368 (N_1368,In_2459,In_2309);
nor U1369 (N_1369,In_2236,N_814);
and U1370 (N_1370,In_1875,In_44);
or U1371 (N_1371,N_724,In_215);
xor U1372 (N_1372,N_813,In_1247);
nand U1373 (N_1373,N_687,In_954);
nand U1374 (N_1374,N_688,N_420);
or U1375 (N_1375,In_1846,In_291);
nand U1376 (N_1376,N_879,N_48);
or U1377 (N_1377,N_732,In_2279);
or U1378 (N_1378,In_2257,In_1826);
nand U1379 (N_1379,N_92,In_1569);
and U1380 (N_1380,N_854,In_2329);
xor U1381 (N_1381,In_533,N_890);
nor U1382 (N_1382,N_995,In_1510);
nor U1383 (N_1383,N_718,N_977);
nand U1384 (N_1384,N_957,N_773);
nor U1385 (N_1385,In_2089,N_532);
nor U1386 (N_1386,N_876,In_654);
or U1387 (N_1387,In_1211,N_122);
or U1388 (N_1388,N_827,N_690);
nand U1389 (N_1389,In_1698,In_1310);
and U1390 (N_1390,In_432,In_1903);
xor U1391 (N_1391,In_563,N_594);
nor U1392 (N_1392,In_1375,N_774);
nor U1393 (N_1393,In_624,N_622);
nand U1394 (N_1394,In_507,N_895);
and U1395 (N_1395,N_60,In_352);
xor U1396 (N_1396,In_1280,N_12);
xor U1397 (N_1397,N_539,N_653);
and U1398 (N_1398,N_826,In_331);
nor U1399 (N_1399,N_860,In_710);
nand U1400 (N_1400,In_2385,N_527);
or U1401 (N_1401,In_574,N_806);
xor U1402 (N_1402,In_743,In_1664);
and U1403 (N_1403,N_696,In_1245);
nand U1404 (N_1404,In_1538,In_918);
or U1405 (N_1405,N_949,In_2402);
xor U1406 (N_1406,N_59,N_631);
and U1407 (N_1407,In_2266,N_274);
or U1408 (N_1408,N_279,N_251);
nand U1409 (N_1409,N_918,N_997);
and U1410 (N_1410,N_214,N_931);
and U1411 (N_1411,N_779,N_319);
nor U1412 (N_1412,In_396,N_932);
or U1413 (N_1413,In_824,In_1007);
or U1414 (N_1414,In_1617,N_57);
nand U1415 (N_1415,In_2482,In_1147);
xor U1416 (N_1416,In_1036,N_378);
or U1417 (N_1417,N_757,In_953);
nand U1418 (N_1418,In_1268,N_772);
nor U1419 (N_1419,N_611,N_976);
and U1420 (N_1420,In_932,In_566);
and U1421 (N_1421,N_790,In_1413);
and U1422 (N_1422,In_1466,In_1246);
nor U1423 (N_1423,In_2347,N_522);
xnor U1424 (N_1424,In_111,N_993);
nand U1425 (N_1425,In_1655,In_955);
or U1426 (N_1426,In_2134,N_908);
or U1427 (N_1427,N_204,N_787);
and U1428 (N_1428,N_789,N_161);
or U1429 (N_1429,N_411,In_2345);
and U1430 (N_1430,In_1090,N_143);
or U1431 (N_1431,N_480,N_715);
or U1432 (N_1432,In_1770,N_553);
nor U1433 (N_1433,N_245,In_1162);
or U1434 (N_1434,N_743,N_558);
and U1435 (N_1435,In_123,In_1218);
or U1436 (N_1436,N_264,In_2321);
or U1437 (N_1437,In_1473,N_844);
and U1438 (N_1438,In_143,N_646);
xor U1439 (N_1439,In_1536,In_195);
nor U1440 (N_1440,In_1805,N_474);
xnor U1441 (N_1441,In_977,N_750);
nand U1442 (N_1442,N_974,In_1276);
xor U1443 (N_1443,N_141,In_2490);
nor U1444 (N_1444,In_491,N_511);
nand U1445 (N_1445,N_978,N_462);
xnor U1446 (N_1446,N_677,N_86);
and U1447 (N_1447,N_581,In_958);
nor U1448 (N_1448,In_1207,In_701);
xor U1449 (N_1449,N_734,In_1654);
and U1450 (N_1450,N_150,N_674);
nor U1451 (N_1451,In_7,In_154);
xor U1452 (N_1452,N_309,N_619);
or U1453 (N_1453,In_1318,N_510);
nand U1454 (N_1454,In_720,N_418);
xor U1455 (N_1455,In_90,In_246);
xnor U1456 (N_1456,N_961,N_663);
nand U1457 (N_1457,N_695,N_749);
or U1458 (N_1458,In_562,In_621);
nand U1459 (N_1459,In_625,In_998);
xor U1460 (N_1460,In_1027,N_762);
xnor U1461 (N_1461,In_1953,In_163);
xor U1462 (N_1462,N_942,In_497);
nor U1463 (N_1463,N_630,In_1989);
or U1464 (N_1464,In_1128,In_2460);
or U1465 (N_1465,In_725,N_591);
nand U1466 (N_1466,In_404,N_607);
xor U1467 (N_1467,In_1992,In_1788);
nor U1468 (N_1468,N_642,In_471);
nand U1469 (N_1469,N_636,N_903);
and U1470 (N_1470,In_1006,N_541);
nand U1471 (N_1471,In_829,N_828);
nand U1472 (N_1472,In_581,N_865);
xor U1473 (N_1473,In_2194,In_1417);
or U1474 (N_1474,N_707,In_1954);
nand U1475 (N_1475,In_236,N_819);
or U1476 (N_1476,In_2397,N_796);
xnor U1477 (N_1477,In_2199,In_1095);
nor U1478 (N_1478,N_989,N_72);
nand U1479 (N_1479,N_768,In_197);
or U1480 (N_1480,In_2354,In_2122);
or U1481 (N_1481,N_288,N_984);
nand U1482 (N_1482,In_1463,N_190);
xor U1483 (N_1483,In_2455,In_823);
nand U1484 (N_1484,N_861,N_669);
nor U1485 (N_1485,N_34,In_2195);
or U1486 (N_1486,N_786,N_531);
nor U1487 (N_1487,In_2316,N_682);
nand U1488 (N_1488,N_894,In_1488);
xor U1489 (N_1489,In_1753,In_2173);
nand U1490 (N_1490,N_503,In_912);
xor U1491 (N_1491,In_166,N_373);
nand U1492 (N_1492,In_1441,In_2431);
nand U1493 (N_1493,In_663,N_212);
xor U1494 (N_1494,N_728,N_347);
or U1495 (N_1495,N_399,N_740);
nor U1496 (N_1496,In_433,N_188);
and U1497 (N_1497,In_1196,N_333);
xnor U1498 (N_1498,N_887,In_2063);
or U1499 (N_1499,In_156,In_1834);
and U1500 (N_1500,N_1295,N_1300);
or U1501 (N_1501,N_1195,N_1151);
or U1502 (N_1502,N_1335,N_1353);
nor U1503 (N_1503,In_1013,In_2104);
nand U1504 (N_1504,N_515,In_1399);
and U1505 (N_1505,N_1379,N_1334);
and U1506 (N_1506,N_345,In_290);
xor U1507 (N_1507,N_84,N_1114);
nor U1508 (N_1508,In_1221,N_1152);
nor U1509 (N_1509,In_790,N_1368);
nor U1510 (N_1510,N_573,N_1265);
nor U1511 (N_1511,N_951,In_1114);
and U1512 (N_1512,In_1029,N_1383);
nor U1513 (N_1513,In_532,N_1243);
nand U1514 (N_1514,N_5,N_937);
nand U1515 (N_1515,N_1349,N_1274);
nand U1516 (N_1516,N_1450,In_1772);
nor U1517 (N_1517,N_1036,N_1468);
nand U1518 (N_1518,N_1141,N_871);
xor U1519 (N_1519,In_2228,N_1382);
and U1520 (N_1520,N_385,N_260);
and U1521 (N_1521,In_2075,N_1213);
or U1522 (N_1522,In_1746,N_419);
nand U1523 (N_1523,N_1312,N_1046);
nor U1524 (N_1524,N_1239,In_860);
xor U1525 (N_1525,N_1488,N_1138);
nor U1526 (N_1526,In_601,In_1533);
or U1527 (N_1527,N_628,In_251);
or U1528 (N_1528,N_1048,N_1369);
or U1529 (N_1529,In_641,N_719);
xor U1530 (N_1530,N_1282,N_916);
and U1531 (N_1531,N_365,N_998);
or U1532 (N_1532,In_1071,N_936);
or U1533 (N_1533,N_1310,N_112);
nor U1534 (N_1534,N_1035,N_1412);
and U1535 (N_1535,N_1007,N_874);
nor U1536 (N_1536,N_1279,N_1253);
and U1537 (N_1537,N_1381,N_1256);
xnor U1538 (N_1538,In_564,In_2430);
or U1539 (N_1539,In_920,N_1340);
and U1540 (N_1540,N_1144,N_1042);
nor U1541 (N_1541,N_1434,N_598);
nand U1542 (N_1542,N_1156,In_2296);
xnor U1543 (N_1543,N_1497,In_238);
xnor U1544 (N_1544,N_700,N_1415);
xor U1545 (N_1545,N_1483,N_1180);
nand U1546 (N_1546,N_1175,In_848);
nand U1547 (N_1547,N_1084,N_899);
xor U1548 (N_1548,In_319,N_838);
nand U1549 (N_1549,N_1031,N_225);
nor U1550 (N_1550,In_2241,In_1242);
nand U1551 (N_1551,In_473,N_1390);
and U1552 (N_1552,In_213,N_1408);
and U1553 (N_1553,N_1283,N_1398);
or U1554 (N_1554,N_856,N_818);
and U1555 (N_1555,N_1191,N_744);
or U1556 (N_1556,N_1484,In_773);
xor U1557 (N_1557,N_1323,N_1214);
nand U1558 (N_1558,N_1366,N_1370);
or U1559 (N_1559,N_1392,In_2207);
or U1560 (N_1560,N_280,N_1225);
xnor U1561 (N_1561,N_1402,N_1316);
xnor U1562 (N_1562,N_1314,N_1104);
xnor U1563 (N_1563,In_927,N_1227);
nand U1564 (N_1564,N_1343,N_1017);
nor U1565 (N_1565,N_1166,In_1068);
nand U1566 (N_1566,N_1161,N_816);
nand U1567 (N_1567,N_1301,N_1016);
or U1568 (N_1568,N_248,In_1716);
or U1569 (N_1569,In_648,In_2295);
and U1570 (N_1570,N_1427,N_1192);
nor U1571 (N_1571,N_1159,N_650);
nand U1572 (N_1572,In_2193,N_540);
and U1573 (N_1573,N_1413,N_1018);
and U1574 (N_1574,N_1297,N_1055);
and U1575 (N_1575,N_1117,In_359);
and U1576 (N_1576,N_1322,N_1240);
and U1577 (N_1577,N_956,N_1187);
nand U1578 (N_1578,N_1226,N_1206);
nor U1579 (N_1579,N_1439,In_1471);
nor U1580 (N_1580,N_596,N_1403);
nand U1581 (N_1581,N_13,In_515);
and U1582 (N_1582,N_1025,In_1611);
nand U1583 (N_1583,N_1241,N_910);
or U1584 (N_1584,N_176,In_985);
xnor U1585 (N_1585,N_1496,N_1249);
xor U1586 (N_1586,In_856,N_1423);
xor U1587 (N_1587,N_1090,N_1426);
nor U1588 (N_1588,In_2285,In_492);
nor U1589 (N_1589,In_170,N_82);
and U1590 (N_1590,In_791,N_1372);
nor U1591 (N_1591,N_1285,N_1129);
or U1592 (N_1592,N_1456,N_1385);
and U1593 (N_1593,N_1454,N_1131);
nor U1594 (N_1594,N_1096,N_754);
nand U1595 (N_1595,N_114,N_297);
nand U1596 (N_1596,In_415,N_666);
and U1597 (N_1597,N_725,N_1184);
nand U1598 (N_1598,N_1126,N_1167);
nand U1599 (N_1599,N_1203,In_1390);
xor U1600 (N_1600,N_1302,N_940);
xor U1601 (N_1601,N_1190,In_317);
nand U1602 (N_1602,N_1215,In_1);
xnor U1603 (N_1603,N_1150,N_269);
and U1604 (N_1604,N_1123,N_1264);
xor U1605 (N_1605,N_1286,N_1238);
xnor U1606 (N_1606,N_1064,N_1027);
or U1607 (N_1607,In_2210,N_1363);
nor U1608 (N_1608,In_770,N_927);
xnor U1609 (N_1609,In_413,N_1470);
xor U1610 (N_1610,In_1153,N_1002);
nand U1611 (N_1611,In_2355,N_1038);
or U1612 (N_1612,N_1458,N_298);
nand U1613 (N_1613,N_644,N_1433);
nand U1614 (N_1614,N_1331,N_1041);
or U1615 (N_1615,In_1263,N_1185);
nor U1616 (N_1616,N_1278,N_1079);
nand U1617 (N_1617,N_1047,N_1223);
nor U1618 (N_1618,N_1115,N_1262);
nand U1619 (N_1619,N_1396,N_601);
nand U1620 (N_1620,In_1928,N_1077);
nand U1621 (N_1621,In_884,In_1539);
xnor U1622 (N_1622,In_851,N_1447);
xnor U1623 (N_1623,N_891,In_1460);
or U1624 (N_1624,N_1134,N_1008);
nor U1625 (N_1625,In_1340,N_972);
xor U1626 (N_1626,In_1855,N_1030);
nor U1627 (N_1627,N_1113,In_863);
and U1628 (N_1628,N_1009,N_837);
or U1629 (N_1629,N_1270,In_827);
xor U1630 (N_1630,In_1872,N_83);
and U1631 (N_1631,N_788,In_1577);
or U1632 (N_1632,N_657,N_868);
or U1633 (N_1633,N_1380,N_1014);
and U1634 (N_1634,In_1732,N_410);
nand U1635 (N_1635,In_2032,In_247);
nor U1636 (N_1636,N_174,In_765);
or U1637 (N_1637,N_846,In_1370);
and U1638 (N_1638,N_1248,N_1122);
or U1639 (N_1639,N_1208,In_1299);
nor U1640 (N_1640,N_1168,N_713);
or U1641 (N_1641,In_2253,N_1091);
or U1642 (N_1642,N_1435,N_1393);
and U1643 (N_1643,N_939,N_717);
nand U1644 (N_1644,In_1975,In_1334);
xor U1645 (N_1645,N_952,N_332);
and U1646 (N_1646,N_479,In_1633);
nand U1647 (N_1647,In_2435,N_1204);
or U1648 (N_1648,In_262,N_1162);
nor U1649 (N_1649,N_494,N_948);
or U1650 (N_1650,N_988,N_1088);
or U1651 (N_1651,N_1222,N_1350);
and U1652 (N_1652,In_167,N_613);
nand U1653 (N_1653,In_1747,N_1217);
nor U1654 (N_1654,N_568,N_1207);
nand U1655 (N_1655,N_882,N_763);
or U1656 (N_1656,N_368,N_1266);
and U1657 (N_1657,In_2403,In_1002);
and U1658 (N_1658,In_1201,N_1453);
or U1659 (N_1659,N_1327,N_888);
or U1660 (N_1660,In_2184,N_89);
nor U1661 (N_1661,N_1358,N_1148);
nand U1662 (N_1662,In_1879,N_249);
nand U1663 (N_1663,In_1032,N_1319);
nand U1664 (N_1664,N_554,N_1232);
nor U1665 (N_1665,In_1736,N_1345);
nand U1666 (N_1666,N_985,N_811);
xor U1667 (N_1667,In_2479,N_381);
nor U1668 (N_1668,N_115,In_2188);
xnor U1669 (N_1669,N_405,N_599);
or U1670 (N_1670,N_1315,In_2363);
nand U1671 (N_1671,N_1102,N_1260);
and U1672 (N_1672,N_1058,N_463);
or U1673 (N_1673,N_578,N_564);
xnor U1674 (N_1674,N_1044,In_2365);
nor U1675 (N_1675,N_1015,N_835);
and U1676 (N_1676,N_640,N_1013);
xnor U1677 (N_1677,N_85,In_1892);
and U1678 (N_1678,N_1012,In_1285);
nor U1679 (N_1679,N_824,N_1119);
nand U1680 (N_1680,N_1201,N_537);
nor U1681 (N_1681,In_362,N_1086);
nand U1682 (N_1682,N_561,N_1306);
nand U1683 (N_1683,N_960,In_702);
nand U1684 (N_1684,In_1511,In_2307);
and U1685 (N_1685,In_1004,In_1774);
or U1686 (N_1686,N_1491,N_1377);
xor U1687 (N_1687,N_1029,N_1205);
and U1688 (N_1688,N_1135,In_1291);
or U1689 (N_1689,In_1406,N_1494);
nand U1690 (N_1690,N_1062,N_1471);
nand U1691 (N_1691,In_962,N_1033);
and U1692 (N_1692,In_794,N_878);
nand U1693 (N_1693,N_538,N_877);
xor U1694 (N_1694,N_904,N_1263);
nand U1695 (N_1695,N_617,N_1328);
nand U1696 (N_1696,In_2162,N_1420);
nand U1697 (N_1697,N_733,N_1125);
nand U1698 (N_1698,N_1364,N_1354);
and U1699 (N_1699,In_2271,In_647);
nor U1700 (N_1700,N_1330,N_1188);
nor U1701 (N_1701,In_1909,N_1045);
and U1702 (N_1702,N_574,N_1024);
nand U1703 (N_1703,In_1481,N_980);
and U1704 (N_1704,N_1053,In_275);
xnor U1705 (N_1705,N_1318,N_1236);
xor U1706 (N_1706,In_1635,N_1388);
xnor U1707 (N_1707,N_907,N_80);
xor U1708 (N_1708,N_1284,N_1107);
or U1709 (N_1709,N_1493,In_1936);
and U1710 (N_1710,N_1485,In_1763);
nor U1711 (N_1711,N_769,N_1277);
and U1712 (N_1712,N_1212,N_1242);
and U1713 (N_1713,N_1425,N_866);
nor U1714 (N_1714,N_1394,N_1313);
xor U1715 (N_1715,In_1136,N_1006);
and U1716 (N_1716,N_1083,N_1442);
or U1717 (N_1717,N_1010,In_1102);
nand U1718 (N_1718,N_1040,N_1216);
nand U1719 (N_1719,N_1076,N_1210);
nor U1720 (N_1720,N_1228,N_1399);
xnor U1721 (N_1721,In_754,N_484);
nor U1722 (N_1722,In_1149,N_1416);
nand U1723 (N_1723,N_1428,N_1257);
and U1724 (N_1724,N_536,N_1486);
nor U1725 (N_1725,In_387,N_1136);
or U1726 (N_1726,In_1380,N_1178);
xnor U1727 (N_1727,N_1418,N_1164);
xnor U1728 (N_1728,N_514,N_1132);
nand U1729 (N_1729,N_584,N_1034);
nand U1730 (N_1730,N_968,N_771);
nor U1731 (N_1731,N_1237,N_760);
or U1732 (N_1732,In_2391,In_174);
and U1733 (N_1733,N_1170,N_1234);
nand U1734 (N_1734,N_491,N_1250);
and U1735 (N_1735,In_1979,N_1365);
nand U1736 (N_1736,In_2004,N_1360);
or U1737 (N_1737,N_1071,N_1443);
nand U1738 (N_1738,N_1095,N_1085);
nor U1739 (N_1739,N_1255,N_1305);
nor U1740 (N_1740,N_1474,N_454);
and U1741 (N_1741,N_1142,N_1063);
nand U1742 (N_1742,In_1458,N_1112);
xnor U1743 (N_1743,N_1224,N_1384);
or U1744 (N_1744,N_1352,N_1371);
or U1745 (N_1745,N_1281,N_1499);
xor U1746 (N_1746,In_374,N_678);
nand U1747 (N_1747,N_1252,N_1329);
xor U1748 (N_1748,N_435,N_1109);
and U1749 (N_1749,In_917,In_1560);
and U1750 (N_1750,N_1124,N_109);
nor U1751 (N_1751,In_1081,In_372);
nand U1752 (N_1752,N_756,N_648);
nor U1753 (N_1753,N_1481,N_1120);
nand U1754 (N_1754,N_1169,N_1182);
or U1755 (N_1755,N_33,N_661);
nor U1756 (N_1756,N_1022,N_67);
xor U1757 (N_1757,N_191,In_81);
and U1758 (N_1758,N_830,N_1066);
or U1759 (N_1759,In_493,N_802);
nor U1760 (N_1760,N_791,In_1922);
xnor U1761 (N_1761,N_518,In_2425);
and U1762 (N_1762,N_1023,N_278);
or U1763 (N_1763,N_785,N_1149);
nand U1764 (N_1764,N_157,N_104);
nand U1765 (N_1765,N_521,N_1139);
and U1766 (N_1766,N_606,N_520);
xnor U1767 (N_1767,In_451,N_727);
or U1768 (N_1768,N_731,In_775);
and U1769 (N_1769,N_1419,N_987);
and U1770 (N_1770,N_1163,In_2374);
and U1771 (N_1771,N_759,N_352);
xor U1772 (N_1772,N_626,N_1089);
or U1773 (N_1773,N_1056,N_1268);
xor U1774 (N_1774,N_1137,N_609);
and U1775 (N_1775,N_1276,In_1091);
nor U1776 (N_1776,In_892,In_1054);
or U1777 (N_1777,N_1078,N_1183);
or U1778 (N_1778,N_1397,N_605);
or U1779 (N_1779,N_361,N_394);
or U1780 (N_1780,N_1462,N_519);
and U1781 (N_1781,N_1376,N_1037);
or U1782 (N_1782,N_1356,N_1275);
and U1783 (N_1783,N_847,N_43);
nor U1784 (N_1784,N_912,N_1005);
and U1785 (N_1785,In_1801,In_1523);
nor U1786 (N_1786,N_1431,N_843);
and U1787 (N_1787,N_1118,N_557);
nand U1788 (N_1788,N_1097,In_1990);
or U1789 (N_1789,In_180,N_745);
and U1790 (N_1790,N_1438,In_2432);
nand U1791 (N_1791,N_1288,N_1200);
and U1792 (N_1792,N_1155,N_627);
and U1793 (N_1793,N_1174,N_1373);
and U1794 (N_1794,N_1464,N_900);
nand U1795 (N_1795,N_1176,N_113);
xor U1796 (N_1796,N_897,In_970);
and U1797 (N_1797,N_1375,N_1116);
and U1798 (N_1798,N_1326,In_1812);
nand U1799 (N_1799,N_1337,N_1271);
nand U1800 (N_1800,N_1293,N_924);
nand U1801 (N_1801,N_1344,N_1317);
xor U1802 (N_1802,In_1578,N_1361);
xnor U1803 (N_1803,In_903,N_962);
nor U1804 (N_1804,N_1189,N_1196);
nor U1805 (N_1805,N_1324,N_692);
nand U1806 (N_1806,N_1021,In_39);
xnor U1807 (N_1807,N_1173,In_2097);
and U1808 (N_1808,N_1099,In_1160);
and U1809 (N_1809,N_258,N_1303);
and U1810 (N_1810,N_149,In_640);
nand U1811 (N_1811,N_706,N_889);
and U1812 (N_1812,N_1440,N_1218);
and U1813 (N_1813,N_1291,In_1123);
and U1814 (N_1814,In_518,N_1489);
and U1815 (N_1815,In_171,In_1127);
nor U1816 (N_1816,In_165,In_2493);
or U1817 (N_1817,N_583,N_1429);
xnor U1818 (N_1818,N_1068,N_1198);
and U1819 (N_1819,N_1414,N_1081);
or U1820 (N_1820,N_219,In_2229);
nor U1821 (N_1821,N_1378,N_621);
nand U1822 (N_1822,N_1092,N_1311);
nand U1823 (N_1823,N_1100,N_29);
and U1824 (N_1824,N_1039,N_213);
nand U1825 (N_1825,N_1254,In_1766);
nand U1826 (N_1826,N_1299,In_864);
nand U1827 (N_1827,N_555,N_1069);
or U1828 (N_1828,N_1267,In_1087);
or U1829 (N_1829,N_963,In_287);
nor U1830 (N_1830,In_1606,N_1146);
or U1831 (N_1831,N_751,N_1246);
nand U1832 (N_1832,N_1436,N_1304);
nand U1833 (N_1833,N_1446,N_1457);
xnor U1834 (N_1834,In_1416,N_1130);
nor U1835 (N_1835,N_1472,In_1388);
or U1836 (N_1836,In_2092,N_893);
or U1837 (N_1837,In_2306,In_1163);
nor U1838 (N_1838,N_780,N_1181);
and U1839 (N_1839,N_1272,In_1456);
xnor U1840 (N_1840,N_55,In_447);
or U1841 (N_1841,N_1057,In_2070);
xor U1842 (N_1842,N_1407,N_1406);
xnor U1843 (N_1843,N_1292,In_2471);
and U1844 (N_1844,N_1395,N_1389);
nand U1845 (N_1845,N_293,N_1171);
nand U1846 (N_1846,N_1140,N_911);
nand U1847 (N_1847,N_563,N_504);
nor U1848 (N_1848,N_1011,N_1220);
and U1849 (N_1849,N_1019,In_268);
xnor U1850 (N_1850,N_1463,N_1093);
and U1851 (N_1851,N_1473,N_943);
nor U1852 (N_1852,N_1320,N_1251);
and U1853 (N_1853,In_1049,N_1404);
or U1854 (N_1854,N_1437,N_1410);
xnor U1855 (N_1855,N_1128,N_1479);
nand U1856 (N_1856,N_1461,N_572);
xnor U1857 (N_1857,N_218,N_739);
and U1858 (N_1858,N_589,N_1362);
nor U1859 (N_1859,In_2454,N_1298);
or U1860 (N_1860,N_872,N_505);
xnor U1861 (N_1861,N_1043,N_1280);
or U1862 (N_1862,In_2209,In_1393);
nand U1863 (N_1863,In_1978,In_1555);
nor U1864 (N_1864,N_1386,N_178);
xnor U1865 (N_1865,N_1245,N_1452);
nor U1866 (N_1866,In_386,N_867);
xnor U1867 (N_1867,In_1361,In_11);
and U1868 (N_1868,N_1121,In_559);
xnor U1869 (N_1869,N_1477,In_1169);
xnor U1870 (N_1870,N_1294,In_2112);
or U1871 (N_1871,N_654,N_1308);
or U1872 (N_1872,In_313,N_1309);
or U1873 (N_1873,N_1004,N_582);
nand U1874 (N_1874,N_1289,In_2125);
nand U1875 (N_1875,N_1341,N_1054);
nor U1876 (N_1876,N_1065,N_1061);
xnor U1877 (N_1877,In_1502,N_926);
nand U1878 (N_1878,N_1476,In_552);
xnor U1879 (N_1879,N_1154,N_1157);
nand U1880 (N_1880,In_759,N_1451);
xor U1881 (N_1881,N_1498,N_1101);
xnor U1882 (N_1882,In_1525,In_547);
and U1883 (N_1883,N_839,N_1269);
or U1884 (N_1884,N_795,N_1290);
nor U1885 (N_1885,In_2111,N_242);
and U1886 (N_1886,N_402,In_1485);
and U1887 (N_1887,In_1924,N_1467);
and U1888 (N_1888,N_1072,N_1026);
xnor U1889 (N_1889,N_349,N_881);
nand U1890 (N_1890,N_842,N_593);
or U1891 (N_1891,N_909,In_500);
or U1892 (N_1892,N_1455,N_833);
nand U1893 (N_1893,N_1221,N_1067);
or U1894 (N_1894,N_21,N_1492);
nor U1895 (N_1895,N_1020,N_567);
or U1896 (N_1896,N_1296,N_1003);
nor U1897 (N_1897,In_2008,N_1357);
xor U1898 (N_1898,N_1346,In_1229);
or U1899 (N_1899,N_1287,N_716);
nor U1900 (N_1900,In_2462,In_1045);
nand U1901 (N_1901,N_676,N_1158);
and U1902 (N_1902,N_1111,In_1260);
nor U1903 (N_1903,N_1145,N_1430);
nor U1904 (N_1904,N_1229,N_1106);
xor U1905 (N_1905,In_210,N_1421);
or U1906 (N_1906,N_1441,N_602);
nand U1907 (N_1907,N_1080,N_1073);
nand U1908 (N_1908,N_501,N_1165);
and U1909 (N_1909,N_1445,In_307);
xor U1910 (N_1910,N_1336,N_1000);
xnor U1911 (N_1911,N_1307,In_243);
or U1912 (N_1912,N_552,N_1209);
or U1913 (N_1913,In_1649,N_1051);
nand U1914 (N_1914,In_614,N_1405);
and U1915 (N_1915,N_1098,N_1147);
nand U1916 (N_1916,In_1663,N_1197);
and U1917 (N_1917,N_1338,In_806);
nand U1918 (N_1918,In_2169,In_350);
or U1919 (N_1919,N_1367,N_1325);
xor U1920 (N_1920,N_1233,N_1321);
nor U1921 (N_1921,N_101,In_1154);
nor U1922 (N_1922,N_1259,N_799);
or U1923 (N_1923,N_1052,N_1422);
nor U1924 (N_1924,N_255,N_632);
nand U1925 (N_1925,N_1153,N_1235);
nor U1926 (N_1926,In_692,In_1876);
nor U1927 (N_1927,In_2349,N_1444);
nor U1928 (N_1928,In_821,N_1495);
nand U1929 (N_1929,N_729,In_234);
nor U1930 (N_1930,N_1244,N_374);
xor U1931 (N_1931,N_1193,N_1060);
and U1932 (N_1932,N_1347,In_921);
nor U1933 (N_1933,N_1087,In_2110);
nor U1934 (N_1934,In_2436,N_172);
nand U1935 (N_1935,N_1103,N_1032);
nor U1936 (N_1936,In_2286,N_1258);
or U1937 (N_1937,N_1465,N_451);
xor U1938 (N_1938,N_1348,N_1475);
or U1939 (N_1939,N_1417,N_1487);
and U1940 (N_1940,N_1108,N_958);
nand U1941 (N_1941,N_704,N_546);
nand U1942 (N_1942,N_1001,In_1658);
and U1943 (N_1943,N_810,N_929);
and U1944 (N_1944,N_396,N_1339);
xor U1945 (N_1945,N_946,In_383);
xor U1946 (N_1946,N_1374,In_308);
nand U1947 (N_1947,N_545,N_1049);
and U1948 (N_1948,In_522,N_870);
xor U1949 (N_1949,N_1050,N_1355);
nand U1950 (N_1950,N_1432,N_523);
nor U1951 (N_1951,In_2458,In_0);
nor U1952 (N_1952,N_1075,N_431);
or U1953 (N_1953,N_1186,N_1401);
or U1954 (N_1954,In_975,N_701);
nor U1955 (N_1955,N_1448,N_1110);
nor U1956 (N_1956,N_81,N_1105);
nand U1957 (N_1957,N_1359,N_967);
and U1958 (N_1958,In_403,N_1143);
nor U1959 (N_1959,N_168,N_417);
xor U1960 (N_1960,N_40,N_1199);
nor U1961 (N_1961,In_1860,N_1424);
nor U1962 (N_1962,N_1074,In_193);
and U1963 (N_1963,N_1273,N_1028);
nor U1964 (N_1964,N_1179,In_1151);
nor U1965 (N_1965,In_109,N_571);
or U1966 (N_1966,N_1231,In_812);
and U1967 (N_1967,In_1591,N_1387);
and U1968 (N_1968,N_761,In_535);
or U1969 (N_1969,In_423,In_1599);
and U1970 (N_1970,In_1059,N_516);
xor U1971 (N_1971,In_779,N_1333);
or U1972 (N_1972,N_1332,N_923);
nor U1973 (N_1973,N_1230,N_2);
xor U1974 (N_1974,N_570,N_1172);
nor U1975 (N_1975,In_1757,N_975);
and U1976 (N_1976,N_1211,In_1214);
nor U1977 (N_1977,N_1127,N_1133);
or U1978 (N_1978,N_1194,N_1342);
nand U1979 (N_1979,N_1478,N_344);
nand U1980 (N_1980,N_470,N_1480);
and U1981 (N_1981,N_1059,N_683);
nand U1982 (N_1982,N_144,N_1490);
and U1983 (N_1983,N_382,N_1400);
or U1984 (N_1984,N_119,N_380);
nand U1985 (N_1985,In_172,N_1247);
nor U1986 (N_1986,In_695,N_1202);
nand U1987 (N_1987,N_32,N_1391);
and U1988 (N_1988,N_1469,N_1466);
nand U1989 (N_1989,N_1459,N_1082);
and U1990 (N_1990,N_1409,N_1351);
nor U1991 (N_1991,N_755,In_1367);
xor U1992 (N_1992,N_445,N_340);
xor U1993 (N_1993,N_1094,N_1482);
xnor U1994 (N_1994,In_2198,N_1160);
or U1995 (N_1995,N_1261,In_1849);
nor U1996 (N_1996,N_1219,N_1070);
nor U1997 (N_1997,In_218,N_1460);
xnor U1998 (N_1998,N_1411,N_1449);
and U1999 (N_1999,In_1579,N_1177);
and U2000 (N_2000,N_1547,N_1914);
nand U2001 (N_2001,N_1654,N_1562);
nand U2002 (N_2002,N_1906,N_1863);
nor U2003 (N_2003,N_1725,N_1577);
and U2004 (N_2004,N_1593,N_1613);
nand U2005 (N_2005,N_1698,N_1803);
or U2006 (N_2006,N_1596,N_1890);
xor U2007 (N_2007,N_1757,N_1607);
nor U2008 (N_2008,N_1537,N_1804);
nor U2009 (N_2009,N_1553,N_1550);
and U2010 (N_2010,N_1773,N_1840);
or U2011 (N_2011,N_1776,N_1866);
nand U2012 (N_2012,N_1966,N_1516);
xnor U2013 (N_2013,N_1641,N_1646);
nand U2014 (N_2014,N_1629,N_1627);
or U2015 (N_2015,N_1623,N_1844);
or U2016 (N_2016,N_1879,N_1558);
xor U2017 (N_2017,N_1766,N_1691);
or U2018 (N_2018,N_1928,N_1505);
nand U2019 (N_2019,N_1874,N_1990);
nor U2020 (N_2020,N_1856,N_1848);
and U2021 (N_2021,N_1819,N_1522);
nor U2022 (N_2022,N_1794,N_1769);
xnor U2023 (N_2023,N_1709,N_1650);
nor U2024 (N_2024,N_1560,N_1687);
and U2025 (N_2025,N_1688,N_1947);
or U2026 (N_2026,N_1739,N_1817);
nor U2027 (N_2027,N_1614,N_1587);
nor U2028 (N_2028,N_1948,N_1765);
nor U2029 (N_2029,N_1957,N_1857);
xnor U2030 (N_2030,N_1588,N_1876);
nand U2031 (N_2031,N_1832,N_1865);
xnor U2032 (N_2032,N_1750,N_1677);
and U2033 (N_2033,N_1660,N_1770);
or U2034 (N_2034,N_1667,N_1535);
xnor U2035 (N_2035,N_1884,N_1970);
nand U2036 (N_2036,N_1918,N_1644);
or U2037 (N_2037,N_1532,N_1919);
nor U2038 (N_2038,N_1518,N_1506);
nand U2039 (N_2039,N_1965,N_1942);
and U2040 (N_2040,N_1967,N_1836);
and U2041 (N_2041,N_1612,N_1873);
and U2042 (N_2042,N_1726,N_1599);
xor U2043 (N_2043,N_1665,N_1830);
or U2044 (N_2044,N_1806,N_1915);
nor U2045 (N_2045,N_1943,N_1674);
nor U2046 (N_2046,N_1534,N_1800);
and U2047 (N_2047,N_1802,N_1852);
and U2048 (N_2048,N_1720,N_1713);
xnor U2049 (N_2049,N_1727,N_1814);
or U2050 (N_2050,N_1512,N_1582);
and U2051 (N_2051,N_1741,N_1860);
nor U2052 (N_2052,N_1872,N_1655);
or U2053 (N_2053,N_1785,N_1634);
nor U2054 (N_2054,N_1903,N_1759);
or U2055 (N_2055,N_1944,N_1600);
nand U2056 (N_2056,N_1754,N_1810);
nand U2057 (N_2057,N_1916,N_1690);
and U2058 (N_2058,N_1912,N_1565);
nand U2059 (N_2059,N_1880,N_1743);
nor U2060 (N_2060,N_1870,N_1790);
nand U2061 (N_2061,N_1503,N_1902);
or U2062 (N_2062,N_1778,N_1673);
xnor U2063 (N_2063,N_1526,N_1531);
xor U2064 (N_2064,N_1995,N_1823);
and U2065 (N_2065,N_1847,N_1571);
nand U2066 (N_2066,N_1543,N_1923);
nand U2067 (N_2067,N_1881,N_1556);
and U2068 (N_2068,N_1827,N_1972);
nand U2069 (N_2069,N_1753,N_1930);
xnor U2070 (N_2070,N_1584,N_1793);
or U2071 (N_2071,N_1501,N_1575);
nor U2072 (N_2072,N_1632,N_1960);
or U2073 (N_2073,N_1878,N_1982);
and U2074 (N_2074,N_1816,N_1837);
and U2075 (N_2075,N_1731,N_1714);
xor U2076 (N_2076,N_1764,N_1594);
nor U2077 (N_2077,N_1564,N_1781);
nand U2078 (N_2078,N_1668,N_1786);
nand U2079 (N_2079,N_1898,N_1981);
nand U2080 (N_2080,N_1638,N_1932);
xor U2081 (N_2081,N_1875,N_1984);
nor U2082 (N_2082,N_1729,N_1831);
nor U2083 (N_2083,N_1843,N_1573);
nand U2084 (N_2084,N_1996,N_1973);
or U2085 (N_2085,N_1885,N_1715);
and U2086 (N_2086,N_1894,N_1805);
or U2087 (N_2087,N_1509,N_1969);
nor U2088 (N_2088,N_1985,N_1514);
or U2089 (N_2089,N_1855,N_1620);
nor U2090 (N_2090,N_1771,N_1777);
and U2091 (N_2091,N_1642,N_1988);
or U2092 (N_2092,N_1700,N_1772);
and U2093 (N_2093,N_1854,N_1801);
xor U2094 (N_2094,N_1675,N_1950);
xnor U2095 (N_2095,N_1626,N_1569);
and U2096 (N_2096,N_1616,N_1887);
or U2097 (N_2097,N_1661,N_1929);
nand U2098 (N_2098,N_1630,N_1711);
nor U2099 (N_2099,N_1706,N_1822);
nand U2100 (N_2100,N_1748,N_1845);
nand U2101 (N_2101,N_1888,N_1954);
xnor U2102 (N_2102,N_1751,N_1937);
or U2103 (N_2103,N_1552,N_1774);
or U2104 (N_2104,N_1920,N_1945);
or U2105 (N_2105,N_1733,N_1693);
and U2106 (N_2106,N_1581,N_1633);
xnor U2107 (N_2107,N_1761,N_1762);
and U2108 (N_2108,N_1975,N_1580);
xnor U2109 (N_2109,N_1882,N_1842);
and U2110 (N_2110,N_1609,N_1767);
and U2111 (N_2111,N_1758,N_1656);
or U2112 (N_2112,N_1585,N_1508);
or U2113 (N_2113,N_1997,N_1540);
or U2114 (N_2114,N_1601,N_1940);
or U2115 (N_2115,N_1546,N_1869);
xnor U2116 (N_2116,N_1962,N_1530);
and U2117 (N_2117,N_1597,N_1811);
nand U2118 (N_2118,N_1788,N_1521);
xor U2119 (N_2119,N_1548,N_1527);
xnor U2120 (N_2120,N_1908,N_1680);
nand U2121 (N_2121,N_1724,N_1834);
nor U2122 (N_2122,N_1862,N_1807);
nor U2123 (N_2123,N_1611,N_1998);
xor U2124 (N_2124,N_1694,N_1542);
xor U2125 (N_2125,N_1946,N_1651);
or U2126 (N_2126,N_1555,N_1746);
nor U2127 (N_2127,N_1625,N_1798);
nor U2128 (N_2128,N_1977,N_1523);
nor U2129 (N_2129,N_1853,N_1818);
nand U2130 (N_2130,N_1895,N_1554);
nand U2131 (N_2131,N_1578,N_1663);
xor U2132 (N_2132,N_1708,N_1647);
nor U2133 (N_2133,N_1897,N_1672);
and U2134 (N_2134,N_1636,N_1779);
and U2135 (N_2135,N_1799,N_1605);
nand U2136 (N_2136,N_1952,N_1809);
nand U2137 (N_2137,N_1999,N_1701);
or U2138 (N_2138,N_1783,N_1949);
nand U2139 (N_2139,N_1824,N_1511);
nor U2140 (N_2140,N_1603,N_1592);
xor U2141 (N_2141,N_1519,N_1653);
xor U2142 (N_2142,N_1529,N_1507);
nor U2143 (N_2143,N_1828,N_1924);
xnor U2144 (N_2144,N_1905,N_1576);
nand U2145 (N_2145,N_1787,N_1963);
nor U2146 (N_2146,N_1961,N_1839);
or U2147 (N_2147,N_1846,N_1971);
nor U2148 (N_2148,N_1678,N_1510);
nand U2149 (N_2149,N_1795,N_1652);
or U2150 (N_2150,N_1868,N_1676);
or U2151 (N_2151,N_1864,N_1861);
and U2152 (N_2152,N_1958,N_1911);
nor U2153 (N_2153,N_1728,N_1815);
xnor U2154 (N_2154,N_1978,N_1528);
nand U2155 (N_2155,N_1586,N_1934);
and U2156 (N_2156,N_1956,N_1891);
or U2157 (N_2157,N_1841,N_1721);
nand U2158 (N_2158,N_1504,N_1662);
or U2159 (N_2159,N_1541,N_1719);
or U2160 (N_2160,N_1520,N_1570);
xnor U2161 (N_2161,N_1763,N_1859);
or U2162 (N_2162,N_1533,N_1722);
nor U2163 (N_2163,N_1964,N_1900);
nor U2164 (N_2164,N_1936,N_1849);
and U2165 (N_2165,N_1621,N_1610);
xnor U2166 (N_2166,N_1833,N_1645);
or U2167 (N_2167,N_1567,N_1755);
and U2168 (N_2168,N_1736,N_1659);
or U2169 (N_2169,N_1951,N_1631);
and U2170 (N_2170,N_1976,N_1959);
xor U2171 (N_2171,N_1886,N_1699);
or U2172 (N_2172,N_1838,N_1657);
or U2173 (N_2173,N_1987,N_1517);
nor U2174 (N_2174,N_1835,N_1760);
xnor U2175 (N_2175,N_1695,N_1545);
or U2176 (N_2176,N_1617,N_1723);
nor U2177 (N_2177,N_1538,N_1782);
xor U2178 (N_2178,N_1513,N_1913);
or U2179 (N_2179,N_1789,N_1712);
nand U2180 (N_2180,N_1574,N_1829);
xor U2181 (N_2181,N_1953,N_1705);
or U2182 (N_2182,N_1775,N_1539);
or U2183 (N_2183,N_1608,N_1738);
and U2184 (N_2184,N_1983,N_1525);
or U2185 (N_2185,N_1756,N_1619);
and U2186 (N_2186,N_1635,N_1867);
and U2187 (N_2187,N_1666,N_1780);
nor U2188 (N_2188,N_1909,N_1679);
nor U2189 (N_2189,N_1986,N_1877);
nand U2190 (N_2190,N_1639,N_1544);
nand U2191 (N_2191,N_1640,N_1572);
nor U2192 (N_2192,N_1649,N_1938);
xor U2193 (N_2193,N_1692,N_1922);
or U2194 (N_2194,N_1702,N_1536);
xor U2195 (N_2195,N_1579,N_1910);
and U2196 (N_2196,N_1850,N_1745);
nor U2197 (N_2197,N_1598,N_1551);
nor U2198 (N_2198,N_1648,N_1925);
nor U2199 (N_2199,N_1559,N_1883);
xnor U2200 (N_2200,N_1892,N_1615);
xor U2201 (N_2201,N_1858,N_1591);
and U2202 (N_2202,N_1955,N_1734);
and U2203 (N_2203,N_1606,N_1670);
or U2204 (N_2204,N_1669,N_1685);
nand U2205 (N_2205,N_1622,N_1566);
nand U2206 (N_2206,N_1618,N_1730);
xor U2207 (N_2207,N_1933,N_1931);
nand U2208 (N_2208,N_1941,N_1664);
or U2209 (N_2209,N_1524,N_1899);
and U2210 (N_2210,N_1602,N_1821);
xor U2211 (N_2211,N_1500,N_1684);
and U2212 (N_2212,N_1812,N_1561);
nor U2213 (N_2213,N_1643,N_1502);
xor U2214 (N_2214,N_1683,N_1921);
nor U2215 (N_2215,N_1992,N_1797);
and U2216 (N_2216,N_1628,N_1604);
or U2217 (N_2217,N_1735,N_1991);
nand U2218 (N_2218,N_1682,N_1624);
or U2219 (N_2219,N_1974,N_1686);
and U2220 (N_2220,N_1901,N_1979);
or U2221 (N_2221,N_1896,N_1826);
nor U2222 (N_2222,N_1583,N_1893);
nor U2223 (N_2223,N_1926,N_1825);
xnor U2224 (N_2224,N_1689,N_1968);
and U2225 (N_2225,N_1557,N_1768);
and U2226 (N_2226,N_1590,N_1747);
nand U2227 (N_2227,N_1595,N_1808);
nor U2228 (N_2228,N_1752,N_1904);
nand U2229 (N_2229,N_1589,N_1907);
and U2230 (N_2230,N_1749,N_1742);
xor U2231 (N_2231,N_1980,N_1993);
nand U2232 (N_2232,N_1989,N_1820);
nor U2233 (N_2233,N_1994,N_1637);
nand U2234 (N_2234,N_1737,N_1851);
or U2235 (N_2235,N_1744,N_1697);
or U2236 (N_2236,N_1927,N_1784);
nand U2237 (N_2237,N_1658,N_1707);
and U2238 (N_2238,N_1710,N_1935);
xor U2239 (N_2239,N_1813,N_1704);
nand U2240 (N_2240,N_1568,N_1515);
and U2241 (N_2241,N_1796,N_1671);
or U2242 (N_2242,N_1716,N_1792);
xnor U2243 (N_2243,N_1718,N_1696);
nand U2244 (N_2244,N_1917,N_1871);
nand U2245 (N_2245,N_1791,N_1681);
nand U2246 (N_2246,N_1732,N_1740);
nand U2247 (N_2247,N_1717,N_1703);
or U2248 (N_2248,N_1549,N_1889);
and U2249 (N_2249,N_1563,N_1939);
nor U2250 (N_2250,N_1817,N_1631);
nand U2251 (N_2251,N_1832,N_1887);
or U2252 (N_2252,N_1978,N_1644);
and U2253 (N_2253,N_1537,N_1639);
or U2254 (N_2254,N_1878,N_1970);
xnor U2255 (N_2255,N_1950,N_1782);
nor U2256 (N_2256,N_1639,N_1704);
nor U2257 (N_2257,N_1879,N_1717);
nand U2258 (N_2258,N_1927,N_1718);
or U2259 (N_2259,N_1933,N_1661);
and U2260 (N_2260,N_1813,N_1603);
nor U2261 (N_2261,N_1903,N_1978);
nor U2262 (N_2262,N_1702,N_1529);
or U2263 (N_2263,N_1681,N_1604);
nor U2264 (N_2264,N_1781,N_1647);
and U2265 (N_2265,N_1713,N_1993);
xnor U2266 (N_2266,N_1706,N_1804);
or U2267 (N_2267,N_1713,N_1502);
nand U2268 (N_2268,N_1705,N_1892);
xnor U2269 (N_2269,N_1683,N_1591);
or U2270 (N_2270,N_1624,N_1933);
or U2271 (N_2271,N_1963,N_1782);
or U2272 (N_2272,N_1914,N_1527);
or U2273 (N_2273,N_1902,N_1509);
and U2274 (N_2274,N_1779,N_1680);
xnor U2275 (N_2275,N_1887,N_1838);
or U2276 (N_2276,N_1501,N_1886);
nand U2277 (N_2277,N_1685,N_1673);
nand U2278 (N_2278,N_1727,N_1539);
and U2279 (N_2279,N_1989,N_1935);
xor U2280 (N_2280,N_1789,N_1666);
nand U2281 (N_2281,N_1737,N_1675);
xnor U2282 (N_2282,N_1615,N_1595);
nand U2283 (N_2283,N_1761,N_1595);
or U2284 (N_2284,N_1530,N_1638);
nand U2285 (N_2285,N_1594,N_1695);
xor U2286 (N_2286,N_1755,N_1937);
xor U2287 (N_2287,N_1689,N_1871);
or U2288 (N_2288,N_1907,N_1842);
and U2289 (N_2289,N_1511,N_1552);
and U2290 (N_2290,N_1553,N_1857);
xnor U2291 (N_2291,N_1888,N_1560);
nand U2292 (N_2292,N_1754,N_1619);
nor U2293 (N_2293,N_1866,N_1936);
or U2294 (N_2294,N_1976,N_1603);
xor U2295 (N_2295,N_1546,N_1538);
xnor U2296 (N_2296,N_1625,N_1569);
nor U2297 (N_2297,N_1758,N_1545);
xor U2298 (N_2298,N_1749,N_1785);
nand U2299 (N_2299,N_1592,N_1570);
nand U2300 (N_2300,N_1870,N_1584);
nand U2301 (N_2301,N_1679,N_1761);
xnor U2302 (N_2302,N_1796,N_1784);
xor U2303 (N_2303,N_1510,N_1536);
or U2304 (N_2304,N_1950,N_1887);
nor U2305 (N_2305,N_1847,N_1545);
nor U2306 (N_2306,N_1897,N_1665);
nand U2307 (N_2307,N_1751,N_1736);
nand U2308 (N_2308,N_1645,N_1886);
xnor U2309 (N_2309,N_1875,N_1811);
and U2310 (N_2310,N_1518,N_1924);
xor U2311 (N_2311,N_1721,N_1769);
nor U2312 (N_2312,N_1992,N_1737);
and U2313 (N_2313,N_1874,N_1664);
nor U2314 (N_2314,N_1588,N_1728);
nor U2315 (N_2315,N_1560,N_1862);
and U2316 (N_2316,N_1795,N_1914);
nand U2317 (N_2317,N_1635,N_1743);
and U2318 (N_2318,N_1674,N_1853);
xor U2319 (N_2319,N_1695,N_1570);
xnor U2320 (N_2320,N_1564,N_1679);
and U2321 (N_2321,N_1704,N_1735);
nor U2322 (N_2322,N_1767,N_1889);
and U2323 (N_2323,N_1866,N_1710);
nor U2324 (N_2324,N_1621,N_1550);
or U2325 (N_2325,N_1686,N_1726);
nor U2326 (N_2326,N_1917,N_1541);
or U2327 (N_2327,N_1713,N_1730);
and U2328 (N_2328,N_1702,N_1535);
or U2329 (N_2329,N_1511,N_1784);
and U2330 (N_2330,N_1818,N_1978);
or U2331 (N_2331,N_1744,N_1812);
xnor U2332 (N_2332,N_1585,N_1963);
nand U2333 (N_2333,N_1696,N_1651);
or U2334 (N_2334,N_1797,N_1606);
nand U2335 (N_2335,N_1758,N_1751);
nand U2336 (N_2336,N_1625,N_1663);
and U2337 (N_2337,N_1537,N_1904);
xor U2338 (N_2338,N_1635,N_1585);
or U2339 (N_2339,N_1616,N_1960);
nor U2340 (N_2340,N_1943,N_1816);
and U2341 (N_2341,N_1513,N_1999);
nor U2342 (N_2342,N_1612,N_1854);
and U2343 (N_2343,N_1873,N_1558);
nand U2344 (N_2344,N_1520,N_1564);
xnor U2345 (N_2345,N_1549,N_1937);
nor U2346 (N_2346,N_1979,N_1800);
xnor U2347 (N_2347,N_1678,N_1938);
xor U2348 (N_2348,N_1928,N_1787);
xnor U2349 (N_2349,N_1811,N_1634);
or U2350 (N_2350,N_1685,N_1542);
xnor U2351 (N_2351,N_1760,N_1638);
or U2352 (N_2352,N_1870,N_1594);
nand U2353 (N_2353,N_1681,N_1943);
nor U2354 (N_2354,N_1570,N_1887);
xor U2355 (N_2355,N_1504,N_1977);
and U2356 (N_2356,N_1693,N_1829);
xnor U2357 (N_2357,N_1695,N_1678);
nor U2358 (N_2358,N_1546,N_1770);
xor U2359 (N_2359,N_1783,N_1750);
or U2360 (N_2360,N_1701,N_1865);
nor U2361 (N_2361,N_1575,N_1785);
or U2362 (N_2362,N_1822,N_1986);
and U2363 (N_2363,N_1777,N_1600);
xnor U2364 (N_2364,N_1825,N_1868);
and U2365 (N_2365,N_1908,N_1823);
or U2366 (N_2366,N_1762,N_1541);
or U2367 (N_2367,N_1724,N_1573);
or U2368 (N_2368,N_1938,N_1775);
and U2369 (N_2369,N_1573,N_1749);
or U2370 (N_2370,N_1912,N_1754);
nor U2371 (N_2371,N_1978,N_1691);
nand U2372 (N_2372,N_1597,N_1900);
xnor U2373 (N_2373,N_1805,N_1992);
nand U2374 (N_2374,N_1581,N_1852);
nor U2375 (N_2375,N_1627,N_1924);
nor U2376 (N_2376,N_1777,N_1841);
nand U2377 (N_2377,N_1512,N_1699);
and U2378 (N_2378,N_1686,N_1960);
nor U2379 (N_2379,N_1717,N_1817);
and U2380 (N_2380,N_1571,N_1591);
and U2381 (N_2381,N_1854,N_1909);
xnor U2382 (N_2382,N_1897,N_1776);
or U2383 (N_2383,N_1660,N_1986);
nand U2384 (N_2384,N_1598,N_1653);
nor U2385 (N_2385,N_1569,N_1789);
xor U2386 (N_2386,N_1798,N_1634);
xor U2387 (N_2387,N_1628,N_1696);
and U2388 (N_2388,N_1753,N_1684);
and U2389 (N_2389,N_1973,N_1919);
nand U2390 (N_2390,N_1913,N_1637);
nor U2391 (N_2391,N_1763,N_1882);
and U2392 (N_2392,N_1835,N_1949);
nor U2393 (N_2393,N_1692,N_1571);
xor U2394 (N_2394,N_1590,N_1929);
and U2395 (N_2395,N_1729,N_1803);
nor U2396 (N_2396,N_1726,N_1528);
nor U2397 (N_2397,N_1619,N_1952);
and U2398 (N_2398,N_1526,N_1996);
or U2399 (N_2399,N_1657,N_1539);
nand U2400 (N_2400,N_1964,N_1845);
or U2401 (N_2401,N_1996,N_1612);
or U2402 (N_2402,N_1562,N_1681);
or U2403 (N_2403,N_1551,N_1994);
xnor U2404 (N_2404,N_1747,N_1766);
or U2405 (N_2405,N_1851,N_1820);
xor U2406 (N_2406,N_1543,N_1685);
and U2407 (N_2407,N_1680,N_1520);
nor U2408 (N_2408,N_1999,N_1536);
nand U2409 (N_2409,N_1944,N_1697);
xnor U2410 (N_2410,N_1871,N_1673);
and U2411 (N_2411,N_1978,N_1758);
nor U2412 (N_2412,N_1981,N_1694);
nand U2413 (N_2413,N_1578,N_1619);
nor U2414 (N_2414,N_1569,N_1506);
or U2415 (N_2415,N_1808,N_1566);
nor U2416 (N_2416,N_1872,N_1573);
xor U2417 (N_2417,N_1690,N_1898);
and U2418 (N_2418,N_1979,N_1688);
and U2419 (N_2419,N_1527,N_1851);
and U2420 (N_2420,N_1503,N_1991);
xor U2421 (N_2421,N_1858,N_1559);
nand U2422 (N_2422,N_1832,N_1761);
xor U2423 (N_2423,N_1874,N_1906);
xor U2424 (N_2424,N_1819,N_1998);
xnor U2425 (N_2425,N_1855,N_1591);
and U2426 (N_2426,N_1739,N_1785);
and U2427 (N_2427,N_1548,N_1688);
and U2428 (N_2428,N_1576,N_1704);
xor U2429 (N_2429,N_1870,N_1957);
and U2430 (N_2430,N_1650,N_1772);
xnor U2431 (N_2431,N_1778,N_1641);
and U2432 (N_2432,N_1547,N_1704);
nor U2433 (N_2433,N_1778,N_1672);
nand U2434 (N_2434,N_1746,N_1511);
nor U2435 (N_2435,N_1962,N_1948);
xor U2436 (N_2436,N_1682,N_1663);
or U2437 (N_2437,N_1695,N_1883);
xnor U2438 (N_2438,N_1946,N_1934);
nand U2439 (N_2439,N_1809,N_1576);
xnor U2440 (N_2440,N_1671,N_1722);
nor U2441 (N_2441,N_1656,N_1720);
or U2442 (N_2442,N_1883,N_1531);
nand U2443 (N_2443,N_1741,N_1678);
xor U2444 (N_2444,N_1839,N_1527);
xor U2445 (N_2445,N_1712,N_1732);
nand U2446 (N_2446,N_1714,N_1824);
and U2447 (N_2447,N_1807,N_1881);
and U2448 (N_2448,N_1844,N_1877);
nand U2449 (N_2449,N_1758,N_1886);
and U2450 (N_2450,N_1543,N_1993);
or U2451 (N_2451,N_1949,N_1967);
and U2452 (N_2452,N_1863,N_1630);
nand U2453 (N_2453,N_1593,N_1816);
or U2454 (N_2454,N_1848,N_1557);
or U2455 (N_2455,N_1575,N_1648);
xnor U2456 (N_2456,N_1799,N_1778);
or U2457 (N_2457,N_1810,N_1876);
xnor U2458 (N_2458,N_1507,N_1517);
and U2459 (N_2459,N_1882,N_1747);
and U2460 (N_2460,N_1962,N_1503);
and U2461 (N_2461,N_1871,N_1512);
nor U2462 (N_2462,N_1828,N_1962);
xnor U2463 (N_2463,N_1650,N_1927);
and U2464 (N_2464,N_1932,N_1750);
or U2465 (N_2465,N_1716,N_1584);
nand U2466 (N_2466,N_1624,N_1647);
xnor U2467 (N_2467,N_1775,N_1818);
or U2468 (N_2468,N_1688,N_1848);
xor U2469 (N_2469,N_1811,N_1669);
nand U2470 (N_2470,N_1590,N_1506);
or U2471 (N_2471,N_1900,N_1638);
xor U2472 (N_2472,N_1715,N_1919);
or U2473 (N_2473,N_1838,N_1673);
xnor U2474 (N_2474,N_1868,N_1607);
xor U2475 (N_2475,N_1942,N_1929);
or U2476 (N_2476,N_1547,N_1688);
and U2477 (N_2477,N_1731,N_1506);
nor U2478 (N_2478,N_1926,N_1602);
nand U2479 (N_2479,N_1788,N_1715);
nor U2480 (N_2480,N_1640,N_1648);
xnor U2481 (N_2481,N_1948,N_1589);
nor U2482 (N_2482,N_1879,N_1991);
nand U2483 (N_2483,N_1816,N_1591);
nor U2484 (N_2484,N_1568,N_1636);
and U2485 (N_2485,N_1711,N_1500);
nand U2486 (N_2486,N_1851,N_1977);
nand U2487 (N_2487,N_1732,N_1834);
xnor U2488 (N_2488,N_1810,N_1526);
xor U2489 (N_2489,N_1533,N_1669);
or U2490 (N_2490,N_1796,N_1594);
xor U2491 (N_2491,N_1651,N_1859);
nand U2492 (N_2492,N_1627,N_1526);
nor U2493 (N_2493,N_1558,N_1505);
or U2494 (N_2494,N_1992,N_1935);
xnor U2495 (N_2495,N_1964,N_1682);
and U2496 (N_2496,N_1691,N_1755);
or U2497 (N_2497,N_1951,N_1765);
xnor U2498 (N_2498,N_1535,N_1605);
nor U2499 (N_2499,N_1559,N_1539);
nor U2500 (N_2500,N_2224,N_2231);
or U2501 (N_2501,N_2285,N_2486);
nand U2502 (N_2502,N_2089,N_2357);
nor U2503 (N_2503,N_2120,N_2018);
nand U2504 (N_2504,N_2211,N_2162);
nand U2505 (N_2505,N_2087,N_2293);
or U2506 (N_2506,N_2134,N_2151);
nor U2507 (N_2507,N_2455,N_2277);
nand U2508 (N_2508,N_2114,N_2288);
and U2509 (N_2509,N_2341,N_2164);
nor U2510 (N_2510,N_2079,N_2335);
nor U2511 (N_2511,N_2470,N_2045);
or U2512 (N_2512,N_2083,N_2323);
nor U2513 (N_2513,N_2491,N_2414);
nor U2514 (N_2514,N_2415,N_2013);
and U2515 (N_2515,N_2241,N_2093);
nand U2516 (N_2516,N_2152,N_2050);
xor U2517 (N_2517,N_2354,N_2185);
or U2518 (N_2518,N_2340,N_2249);
nand U2519 (N_2519,N_2084,N_2167);
xor U2520 (N_2520,N_2128,N_2396);
or U2521 (N_2521,N_2266,N_2220);
and U2522 (N_2522,N_2010,N_2142);
or U2523 (N_2523,N_2399,N_2240);
nand U2524 (N_2524,N_2379,N_2011);
or U2525 (N_2525,N_2064,N_2250);
xnor U2526 (N_2526,N_2336,N_2094);
nand U2527 (N_2527,N_2383,N_2177);
nor U2528 (N_2528,N_2187,N_2365);
or U2529 (N_2529,N_2475,N_2276);
nand U2530 (N_2530,N_2061,N_2186);
nand U2531 (N_2531,N_2239,N_2359);
nand U2532 (N_2532,N_2484,N_2074);
nor U2533 (N_2533,N_2313,N_2404);
and U2534 (N_2534,N_2304,N_2222);
and U2535 (N_2535,N_2482,N_2001);
xnor U2536 (N_2536,N_2065,N_2447);
and U2537 (N_2537,N_2438,N_2267);
nand U2538 (N_2538,N_2299,N_2168);
xor U2539 (N_2539,N_2110,N_2219);
nand U2540 (N_2540,N_2442,N_2238);
or U2541 (N_2541,N_2138,N_2048);
and U2542 (N_2542,N_2300,N_2403);
nor U2543 (N_2543,N_2283,N_2075);
xor U2544 (N_2544,N_2003,N_2144);
xnor U2545 (N_2545,N_2189,N_2203);
and U2546 (N_2546,N_2433,N_2392);
nor U2547 (N_2547,N_2369,N_2377);
nand U2548 (N_2548,N_2424,N_2361);
xnor U2549 (N_2549,N_2243,N_2235);
xor U2550 (N_2550,N_2097,N_2319);
xor U2551 (N_2551,N_2312,N_2446);
or U2552 (N_2552,N_2023,N_2479);
or U2553 (N_2553,N_2122,N_2386);
nor U2554 (N_2554,N_2281,N_2096);
xnor U2555 (N_2555,N_2217,N_2124);
nand U2556 (N_2556,N_2019,N_2441);
xor U2557 (N_2557,N_2309,N_2436);
and U2558 (N_2558,N_2161,N_2179);
nor U2559 (N_2559,N_2307,N_2395);
nor U2560 (N_2560,N_2201,N_2368);
or U2561 (N_2561,N_2454,N_2017);
nor U2562 (N_2562,N_2421,N_2090);
nand U2563 (N_2563,N_2067,N_2072);
nor U2564 (N_2564,N_2070,N_2471);
xnor U2565 (N_2565,N_2125,N_2314);
nand U2566 (N_2566,N_2461,N_2228);
xnor U2567 (N_2567,N_2102,N_2492);
nand U2568 (N_2568,N_2043,N_2363);
or U2569 (N_2569,N_2112,N_2247);
and U2570 (N_2570,N_2391,N_2171);
nand U2571 (N_2571,N_2047,N_2024);
nand U2572 (N_2572,N_2119,N_2158);
or U2573 (N_2573,N_2409,N_2420);
or U2574 (N_2574,N_2184,N_2428);
nor U2575 (N_2575,N_2166,N_2347);
nor U2576 (N_2576,N_2477,N_2389);
xor U2577 (N_2577,N_2485,N_2481);
or U2578 (N_2578,N_2209,N_2182);
nand U2579 (N_2579,N_2488,N_2127);
xor U2580 (N_2580,N_2287,N_2205);
nand U2581 (N_2581,N_2212,N_2196);
or U2582 (N_2582,N_2229,N_2371);
or U2583 (N_2583,N_2129,N_2294);
xor U2584 (N_2584,N_2145,N_2257);
and U2585 (N_2585,N_2180,N_2202);
and U2586 (N_2586,N_2155,N_2216);
xnor U2587 (N_2587,N_2413,N_2109);
nor U2588 (N_2588,N_2311,N_2374);
nor U2589 (N_2589,N_2326,N_2040);
nand U2590 (N_2590,N_2355,N_2059);
nand U2591 (N_2591,N_2463,N_2016);
nor U2592 (N_2592,N_2435,N_2159);
or U2593 (N_2593,N_2041,N_2337);
xor U2594 (N_2594,N_2289,N_2262);
nor U2595 (N_2595,N_2260,N_2376);
xor U2596 (N_2596,N_2264,N_2029);
nand U2597 (N_2597,N_2286,N_2092);
xor U2598 (N_2598,N_2057,N_2160);
and U2599 (N_2599,N_2098,N_2136);
nor U2600 (N_2600,N_2246,N_2370);
nor U2601 (N_2601,N_2137,N_2271);
nor U2602 (N_2602,N_2278,N_2150);
xor U2603 (N_2603,N_2223,N_2412);
or U2604 (N_2604,N_2265,N_2086);
xor U2605 (N_2605,N_2373,N_2402);
or U2606 (N_2606,N_2366,N_2418);
nand U2607 (N_2607,N_2440,N_2251);
and U2608 (N_2608,N_2226,N_2444);
nor U2609 (N_2609,N_2105,N_2176);
xnor U2610 (N_2610,N_2234,N_2147);
nand U2611 (N_2611,N_2302,N_2156);
nand U2612 (N_2612,N_2268,N_2324);
xnor U2613 (N_2613,N_2237,N_2430);
nor U2614 (N_2614,N_2106,N_2297);
xnor U2615 (N_2615,N_2437,N_2175);
or U2616 (N_2616,N_2188,N_2101);
and U2617 (N_2617,N_2351,N_2116);
nand U2618 (N_2618,N_2282,N_2480);
and U2619 (N_2619,N_2245,N_2410);
nor U2620 (N_2620,N_2107,N_2375);
or U2621 (N_2621,N_2362,N_2031);
nor U2622 (N_2622,N_2360,N_2450);
or U2623 (N_2623,N_2218,N_2460);
and U2624 (N_2624,N_2473,N_2406);
and U2625 (N_2625,N_2364,N_2465);
nand U2626 (N_2626,N_2056,N_2068);
xnor U2627 (N_2627,N_2398,N_2232);
nor U2628 (N_2628,N_2458,N_2080);
nand U2629 (N_2629,N_2174,N_2382);
xor U2630 (N_2630,N_2385,N_2078);
xor U2631 (N_2631,N_2191,N_2353);
nand U2632 (N_2632,N_2451,N_2133);
nor U2633 (N_2633,N_2103,N_2135);
and U2634 (N_2634,N_2295,N_2493);
or U2635 (N_2635,N_2483,N_2063);
xor U2636 (N_2636,N_2197,N_2328);
and U2637 (N_2637,N_2208,N_2387);
or U2638 (N_2638,N_2380,N_2349);
or U2639 (N_2639,N_2467,N_2496);
nor U2640 (N_2640,N_2457,N_2000);
nand U2641 (N_2641,N_2111,N_2478);
and U2642 (N_2642,N_2405,N_2149);
nand U2643 (N_2643,N_2014,N_2292);
nor U2644 (N_2644,N_2027,N_2419);
nor U2645 (N_2645,N_2334,N_2163);
and U2646 (N_2646,N_2062,N_2123);
nor U2647 (N_2647,N_2181,N_2248);
xnor U2648 (N_2648,N_2178,N_2195);
and U2649 (N_2649,N_2066,N_2055);
xnor U2650 (N_2650,N_2499,N_2258);
nand U2651 (N_2651,N_2397,N_2416);
and U2652 (N_2652,N_2453,N_2192);
nand U2653 (N_2653,N_2275,N_2269);
and U2654 (N_2654,N_2053,N_2172);
nand U2655 (N_2655,N_2306,N_2308);
nand U2656 (N_2656,N_2058,N_2154);
xnor U2657 (N_2657,N_2252,N_2054);
nor U2658 (N_2658,N_2104,N_2099);
or U2659 (N_2659,N_2204,N_2459);
xor U2660 (N_2660,N_2034,N_2207);
or U2661 (N_2661,N_2130,N_2236);
xnor U2662 (N_2662,N_2310,N_2474);
and U2663 (N_2663,N_2032,N_2346);
nand U2664 (N_2664,N_2489,N_2468);
xor U2665 (N_2665,N_2330,N_2329);
xor U2666 (N_2666,N_2298,N_2356);
and U2667 (N_2667,N_2401,N_2321);
or U2668 (N_2668,N_2254,N_2193);
or U2669 (N_2669,N_2487,N_2394);
or U2670 (N_2670,N_2022,N_2456);
xor U2671 (N_2671,N_2206,N_2049);
and U2672 (N_2672,N_2448,N_2315);
xor U2673 (N_2673,N_2439,N_2280);
xnor U2674 (N_2674,N_2263,N_2073);
xnor U2675 (N_2675,N_2253,N_2146);
nor U2676 (N_2676,N_2213,N_2035);
or U2677 (N_2677,N_2350,N_2117);
or U2678 (N_2678,N_2113,N_2227);
nand U2679 (N_2679,N_2331,N_2215);
nor U2680 (N_2680,N_2427,N_2210);
or U2681 (N_2681,N_2118,N_2332);
or U2682 (N_2682,N_2036,N_2230);
xnor U2683 (N_2683,N_2198,N_2352);
xor U2684 (N_2684,N_2449,N_2242);
xnor U2685 (N_2685,N_2452,N_2008);
xor U2686 (N_2686,N_2320,N_2233);
nand U2687 (N_2687,N_2325,N_2132);
xnor U2688 (N_2688,N_2121,N_2490);
and U2689 (N_2689,N_2327,N_2417);
or U2690 (N_2690,N_2339,N_2434);
or U2691 (N_2691,N_2190,N_2051);
and U2692 (N_2692,N_2494,N_2173);
nand U2693 (N_2693,N_2025,N_2274);
nand U2694 (N_2694,N_2153,N_2221);
xor U2695 (N_2695,N_2345,N_2148);
nand U2696 (N_2696,N_2378,N_2046);
or U2697 (N_2697,N_2200,N_2429);
and U2698 (N_2698,N_2466,N_2303);
or U2699 (N_2699,N_2425,N_2199);
nor U2700 (N_2700,N_2462,N_2426);
xor U2701 (N_2701,N_2290,N_2445);
xnor U2702 (N_2702,N_2464,N_2495);
and U2703 (N_2703,N_2021,N_2407);
or U2704 (N_2704,N_2358,N_2039);
xnor U2705 (N_2705,N_2348,N_2076);
nor U2706 (N_2706,N_2038,N_2273);
or U2707 (N_2707,N_2225,N_2020);
nand U2708 (N_2708,N_2390,N_2259);
nand U2709 (N_2709,N_2052,N_2498);
or U2710 (N_2710,N_2244,N_2316);
nand U2711 (N_2711,N_2126,N_2042);
or U2712 (N_2712,N_2169,N_2317);
nand U2713 (N_2713,N_2044,N_2469);
nand U2714 (N_2714,N_2384,N_2443);
nand U2715 (N_2715,N_2422,N_2165);
or U2716 (N_2716,N_2261,N_2408);
nor U2717 (N_2717,N_2108,N_2183);
or U2718 (N_2718,N_2472,N_2431);
xor U2719 (N_2719,N_2476,N_2004);
nor U2720 (N_2720,N_2296,N_2342);
and U2721 (N_2721,N_2400,N_2139);
xnor U2722 (N_2722,N_2214,N_2140);
xnor U2723 (N_2723,N_2131,N_2388);
xnor U2724 (N_2724,N_2081,N_2272);
xnor U2725 (N_2725,N_2060,N_2100);
xor U2726 (N_2726,N_2256,N_2255);
or U2727 (N_2727,N_2082,N_2005);
nor U2728 (N_2728,N_2006,N_2305);
or U2729 (N_2729,N_2279,N_2143);
xor U2730 (N_2730,N_2071,N_2037);
nor U2731 (N_2731,N_2026,N_2381);
or U2732 (N_2732,N_2423,N_2077);
nand U2733 (N_2733,N_2007,N_2301);
nor U2734 (N_2734,N_2338,N_2009);
nand U2735 (N_2735,N_2194,N_2432);
nand U2736 (N_2736,N_2497,N_2270);
or U2737 (N_2737,N_2002,N_2170);
nand U2738 (N_2738,N_2033,N_2318);
or U2739 (N_2739,N_2095,N_2284);
xor U2740 (N_2740,N_2141,N_2030);
xor U2741 (N_2741,N_2343,N_2069);
and U2742 (N_2742,N_2015,N_2322);
or U2743 (N_2743,N_2291,N_2012);
nand U2744 (N_2744,N_2157,N_2091);
xor U2745 (N_2745,N_2115,N_2411);
xnor U2746 (N_2746,N_2333,N_2085);
or U2747 (N_2747,N_2344,N_2088);
xnor U2748 (N_2748,N_2393,N_2367);
or U2749 (N_2749,N_2372,N_2028);
and U2750 (N_2750,N_2244,N_2131);
or U2751 (N_2751,N_2421,N_2436);
xnor U2752 (N_2752,N_2209,N_2423);
and U2753 (N_2753,N_2401,N_2347);
xor U2754 (N_2754,N_2391,N_2173);
nand U2755 (N_2755,N_2025,N_2267);
xnor U2756 (N_2756,N_2004,N_2073);
or U2757 (N_2757,N_2387,N_2416);
or U2758 (N_2758,N_2310,N_2026);
nand U2759 (N_2759,N_2061,N_2143);
and U2760 (N_2760,N_2225,N_2266);
and U2761 (N_2761,N_2443,N_2224);
or U2762 (N_2762,N_2425,N_2130);
nor U2763 (N_2763,N_2479,N_2098);
and U2764 (N_2764,N_2303,N_2406);
xnor U2765 (N_2765,N_2179,N_2005);
nor U2766 (N_2766,N_2455,N_2279);
or U2767 (N_2767,N_2133,N_2236);
and U2768 (N_2768,N_2130,N_2300);
nand U2769 (N_2769,N_2062,N_2435);
nor U2770 (N_2770,N_2305,N_2010);
nand U2771 (N_2771,N_2043,N_2384);
and U2772 (N_2772,N_2370,N_2223);
and U2773 (N_2773,N_2429,N_2357);
or U2774 (N_2774,N_2448,N_2499);
xnor U2775 (N_2775,N_2025,N_2436);
nand U2776 (N_2776,N_2389,N_2395);
or U2777 (N_2777,N_2373,N_2216);
and U2778 (N_2778,N_2368,N_2056);
xor U2779 (N_2779,N_2488,N_2315);
nor U2780 (N_2780,N_2226,N_2381);
nand U2781 (N_2781,N_2139,N_2080);
xnor U2782 (N_2782,N_2458,N_2283);
and U2783 (N_2783,N_2423,N_2210);
xnor U2784 (N_2784,N_2378,N_2431);
and U2785 (N_2785,N_2074,N_2195);
xor U2786 (N_2786,N_2173,N_2338);
or U2787 (N_2787,N_2398,N_2123);
nor U2788 (N_2788,N_2254,N_2024);
nand U2789 (N_2789,N_2220,N_2348);
and U2790 (N_2790,N_2195,N_2101);
and U2791 (N_2791,N_2405,N_2435);
or U2792 (N_2792,N_2018,N_2416);
or U2793 (N_2793,N_2032,N_2209);
nand U2794 (N_2794,N_2113,N_2304);
nor U2795 (N_2795,N_2354,N_2325);
nor U2796 (N_2796,N_2245,N_2156);
nand U2797 (N_2797,N_2143,N_2465);
or U2798 (N_2798,N_2338,N_2070);
nand U2799 (N_2799,N_2404,N_2377);
nor U2800 (N_2800,N_2432,N_2255);
nor U2801 (N_2801,N_2338,N_2006);
xnor U2802 (N_2802,N_2329,N_2112);
nand U2803 (N_2803,N_2273,N_2055);
and U2804 (N_2804,N_2358,N_2157);
nand U2805 (N_2805,N_2034,N_2347);
nor U2806 (N_2806,N_2272,N_2279);
or U2807 (N_2807,N_2226,N_2423);
and U2808 (N_2808,N_2446,N_2496);
xnor U2809 (N_2809,N_2470,N_2277);
or U2810 (N_2810,N_2141,N_2001);
nor U2811 (N_2811,N_2158,N_2429);
or U2812 (N_2812,N_2050,N_2070);
or U2813 (N_2813,N_2263,N_2448);
xor U2814 (N_2814,N_2163,N_2065);
or U2815 (N_2815,N_2145,N_2114);
and U2816 (N_2816,N_2150,N_2492);
or U2817 (N_2817,N_2037,N_2005);
nor U2818 (N_2818,N_2458,N_2484);
nor U2819 (N_2819,N_2170,N_2159);
nor U2820 (N_2820,N_2062,N_2208);
or U2821 (N_2821,N_2027,N_2127);
or U2822 (N_2822,N_2303,N_2311);
and U2823 (N_2823,N_2296,N_2346);
xnor U2824 (N_2824,N_2249,N_2415);
and U2825 (N_2825,N_2341,N_2401);
xnor U2826 (N_2826,N_2137,N_2494);
nor U2827 (N_2827,N_2149,N_2496);
and U2828 (N_2828,N_2454,N_2292);
or U2829 (N_2829,N_2090,N_2244);
nand U2830 (N_2830,N_2240,N_2105);
xnor U2831 (N_2831,N_2355,N_2438);
xor U2832 (N_2832,N_2117,N_2385);
or U2833 (N_2833,N_2195,N_2034);
nor U2834 (N_2834,N_2174,N_2368);
and U2835 (N_2835,N_2220,N_2137);
or U2836 (N_2836,N_2044,N_2265);
nor U2837 (N_2837,N_2346,N_2311);
or U2838 (N_2838,N_2038,N_2419);
or U2839 (N_2839,N_2224,N_2422);
and U2840 (N_2840,N_2100,N_2406);
xor U2841 (N_2841,N_2448,N_2131);
nand U2842 (N_2842,N_2091,N_2035);
nand U2843 (N_2843,N_2449,N_2312);
and U2844 (N_2844,N_2363,N_2230);
xor U2845 (N_2845,N_2347,N_2018);
nor U2846 (N_2846,N_2471,N_2279);
xnor U2847 (N_2847,N_2413,N_2395);
xnor U2848 (N_2848,N_2062,N_2092);
nand U2849 (N_2849,N_2437,N_2336);
xnor U2850 (N_2850,N_2354,N_2261);
nor U2851 (N_2851,N_2198,N_2039);
xnor U2852 (N_2852,N_2070,N_2370);
nand U2853 (N_2853,N_2413,N_2008);
nand U2854 (N_2854,N_2110,N_2039);
nor U2855 (N_2855,N_2493,N_2410);
or U2856 (N_2856,N_2432,N_2382);
nor U2857 (N_2857,N_2354,N_2174);
xor U2858 (N_2858,N_2481,N_2297);
or U2859 (N_2859,N_2296,N_2091);
or U2860 (N_2860,N_2189,N_2472);
xor U2861 (N_2861,N_2263,N_2205);
xnor U2862 (N_2862,N_2299,N_2138);
nor U2863 (N_2863,N_2421,N_2358);
and U2864 (N_2864,N_2405,N_2404);
xnor U2865 (N_2865,N_2359,N_2040);
nor U2866 (N_2866,N_2377,N_2422);
and U2867 (N_2867,N_2484,N_2126);
nor U2868 (N_2868,N_2450,N_2335);
and U2869 (N_2869,N_2410,N_2475);
nand U2870 (N_2870,N_2096,N_2049);
xor U2871 (N_2871,N_2066,N_2266);
xnor U2872 (N_2872,N_2368,N_2164);
xnor U2873 (N_2873,N_2372,N_2090);
xnor U2874 (N_2874,N_2081,N_2091);
xor U2875 (N_2875,N_2030,N_2477);
xnor U2876 (N_2876,N_2212,N_2408);
and U2877 (N_2877,N_2343,N_2333);
and U2878 (N_2878,N_2413,N_2083);
and U2879 (N_2879,N_2099,N_2403);
xnor U2880 (N_2880,N_2417,N_2242);
nand U2881 (N_2881,N_2224,N_2088);
or U2882 (N_2882,N_2270,N_2230);
or U2883 (N_2883,N_2386,N_2004);
and U2884 (N_2884,N_2053,N_2163);
or U2885 (N_2885,N_2459,N_2239);
nor U2886 (N_2886,N_2478,N_2335);
xnor U2887 (N_2887,N_2070,N_2186);
nand U2888 (N_2888,N_2185,N_2468);
or U2889 (N_2889,N_2467,N_2143);
nor U2890 (N_2890,N_2263,N_2143);
and U2891 (N_2891,N_2190,N_2418);
or U2892 (N_2892,N_2345,N_2383);
and U2893 (N_2893,N_2322,N_2098);
or U2894 (N_2894,N_2341,N_2106);
or U2895 (N_2895,N_2142,N_2277);
or U2896 (N_2896,N_2262,N_2388);
or U2897 (N_2897,N_2037,N_2294);
xor U2898 (N_2898,N_2007,N_2098);
and U2899 (N_2899,N_2126,N_2068);
or U2900 (N_2900,N_2181,N_2342);
and U2901 (N_2901,N_2174,N_2225);
nand U2902 (N_2902,N_2332,N_2436);
and U2903 (N_2903,N_2448,N_2447);
or U2904 (N_2904,N_2382,N_2056);
or U2905 (N_2905,N_2021,N_2023);
nor U2906 (N_2906,N_2206,N_2378);
nand U2907 (N_2907,N_2024,N_2236);
nor U2908 (N_2908,N_2062,N_2490);
nand U2909 (N_2909,N_2249,N_2281);
or U2910 (N_2910,N_2186,N_2167);
nand U2911 (N_2911,N_2335,N_2193);
or U2912 (N_2912,N_2117,N_2360);
nand U2913 (N_2913,N_2004,N_2392);
or U2914 (N_2914,N_2323,N_2392);
nor U2915 (N_2915,N_2453,N_2126);
nand U2916 (N_2916,N_2244,N_2496);
and U2917 (N_2917,N_2270,N_2070);
and U2918 (N_2918,N_2363,N_2247);
and U2919 (N_2919,N_2339,N_2035);
xnor U2920 (N_2920,N_2197,N_2239);
xor U2921 (N_2921,N_2140,N_2126);
xor U2922 (N_2922,N_2486,N_2332);
xnor U2923 (N_2923,N_2019,N_2072);
nor U2924 (N_2924,N_2000,N_2331);
and U2925 (N_2925,N_2204,N_2256);
nand U2926 (N_2926,N_2261,N_2303);
nor U2927 (N_2927,N_2423,N_2041);
xnor U2928 (N_2928,N_2269,N_2278);
and U2929 (N_2929,N_2109,N_2149);
and U2930 (N_2930,N_2022,N_2029);
xor U2931 (N_2931,N_2414,N_2436);
and U2932 (N_2932,N_2436,N_2446);
nor U2933 (N_2933,N_2183,N_2362);
xor U2934 (N_2934,N_2011,N_2188);
nor U2935 (N_2935,N_2469,N_2133);
or U2936 (N_2936,N_2112,N_2446);
and U2937 (N_2937,N_2219,N_2166);
or U2938 (N_2938,N_2414,N_2354);
nor U2939 (N_2939,N_2009,N_2115);
nor U2940 (N_2940,N_2082,N_2183);
and U2941 (N_2941,N_2468,N_2141);
xor U2942 (N_2942,N_2289,N_2251);
xnor U2943 (N_2943,N_2149,N_2231);
or U2944 (N_2944,N_2416,N_2056);
and U2945 (N_2945,N_2466,N_2379);
and U2946 (N_2946,N_2375,N_2222);
and U2947 (N_2947,N_2242,N_2451);
nor U2948 (N_2948,N_2214,N_2262);
xnor U2949 (N_2949,N_2141,N_2022);
nor U2950 (N_2950,N_2420,N_2422);
or U2951 (N_2951,N_2126,N_2351);
or U2952 (N_2952,N_2120,N_2012);
nor U2953 (N_2953,N_2267,N_2235);
and U2954 (N_2954,N_2220,N_2457);
nand U2955 (N_2955,N_2108,N_2345);
or U2956 (N_2956,N_2470,N_2092);
xor U2957 (N_2957,N_2059,N_2073);
and U2958 (N_2958,N_2461,N_2335);
or U2959 (N_2959,N_2144,N_2186);
nand U2960 (N_2960,N_2220,N_2070);
and U2961 (N_2961,N_2438,N_2450);
and U2962 (N_2962,N_2436,N_2046);
nand U2963 (N_2963,N_2333,N_2490);
and U2964 (N_2964,N_2449,N_2164);
nor U2965 (N_2965,N_2371,N_2083);
xor U2966 (N_2966,N_2487,N_2418);
or U2967 (N_2967,N_2090,N_2360);
or U2968 (N_2968,N_2213,N_2443);
xnor U2969 (N_2969,N_2227,N_2332);
nand U2970 (N_2970,N_2221,N_2452);
nor U2971 (N_2971,N_2352,N_2205);
or U2972 (N_2972,N_2142,N_2086);
xor U2973 (N_2973,N_2289,N_2234);
nor U2974 (N_2974,N_2108,N_2142);
xnor U2975 (N_2975,N_2147,N_2453);
or U2976 (N_2976,N_2448,N_2126);
and U2977 (N_2977,N_2173,N_2419);
xor U2978 (N_2978,N_2259,N_2458);
nor U2979 (N_2979,N_2014,N_2188);
nand U2980 (N_2980,N_2142,N_2152);
or U2981 (N_2981,N_2190,N_2318);
or U2982 (N_2982,N_2255,N_2225);
and U2983 (N_2983,N_2019,N_2423);
or U2984 (N_2984,N_2498,N_2016);
xor U2985 (N_2985,N_2484,N_2428);
xor U2986 (N_2986,N_2470,N_2121);
and U2987 (N_2987,N_2034,N_2217);
xnor U2988 (N_2988,N_2444,N_2495);
and U2989 (N_2989,N_2168,N_2443);
and U2990 (N_2990,N_2130,N_2340);
nor U2991 (N_2991,N_2337,N_2336);
xnor U2992 (N_2992,N_2117,N_2447);
nand U2993 (N_2993,N_2403,N_2143);
or U2994 (N_2994,N_2314,N_2018);
and U2995 (N_2995,N_2273,N_2202);
and U2996 (N_2996,N_2076,N_2452);
nand U2997 (N_2997,N_2374,N_2166);
or U2998 (N_2998,N_2403,N_2376);
or U2999 (N_2999,N_2107,N_2309);
and U3000 (N_3000,N_2902,N_2963);
or U3001 (N_3001,N_2819,N_2727);
or U3002 (N_3002,N_2805,N_2940);
nor U3003 (N_3003,N_2845,N_2979);
nor U3004 (N_3004,N_2740,N_2705);
nor U3005 (N_3005,N_2753,N_2726);
nor U3006 (N_3006,N_2767,N_2711);
nand U3007 (N_3007,N_2646,N_2776);
xnor U3008 (N_3008,N_2633,N_2997);
xor U3009 (N_3009,N_2783,N_2590);
xnor U3010 (N_3010,N_2565,N_2680);
nor U3011 (N_3011,N_2862,N_2866);
or U3012 (N_3012,N_2534,N_2771);
and U3013 (N_3013,N_2630,N_2786);
nor U3014 (N_3014,N_2548,N_2739);
and U3015 (N_3015,N_2540,N_2906);
or U3016 (N_3016,N_2977,N_2609);
or U3017 (N_3017,N_2752,N_2974);
nand U3018 (N_3018,N_2794,N_2958);
or U3019 (N_3019,N_2774,N_2584);
and U3020 (N_3020,N_2651,N_2856);
nor U3021 (N_3021,N_2511,N_2538);
nor U3022 (N_3022,N_2735,N_2885);
and U3023 (N_3023,N_2702,N_2564);
nor U3024 (N_3024,N_2524,N_2725);
nor U3025 (N_3025,N_2861,N_2718);
nand U3026 (N_3026,N_2982,N_2615);
nor U3027 (N_3027,N_2852,N_2684);
nor U3028 (N_3028,N_2549,N_2972);
xor U3029 (N_3029,N_2579,N_2695);
or U3030 (N_3030,N_2729,N_2841);
and U3031 (N_3031,N_2879,N_2987);
nand U3032 (N_3032,N_2994,N_2766);
nor U3033 (N_3033,N_2883,N_2928);
xnor U3034 (N_3034,N_2556,N_2535);
and U3035 (N_3035,N_2793,N_2693);
nand U3036 (N_3036,N_2872,N_2723);
xor U3037 (N_3037,N_2569,N_2658);
or U3038 (N_3038,N_2789,N_2728);
and U3039 (N_3039,N_2521,N_2580);
nand U3040 (N_3040,N_2865,N_2890);
and U3041 (N_3041,N_2675,N_2650);
nand U3042 (N_3042,N_2961,N_2973);
or U3043 (N_3043,N_2561,N_2593);
or U3044 (N_3044,N_2810,N_2777);
nand U3045 (N_3045,N_2661,N_2606);
xor U3046 (N_3046,N_2578,N_2500);
nand U3047 (N_3047,N_2859,N_2560);
nor U3048 (N_3048,N_2934,N_2536);
xor U3049 (N_3049,N_2826,N_2738);
xnor U3050 (N_3050,N_2712,N_2623);
or U3051 (N_3051,N_2932,N_2635);
nor U3052 (N_3052,N_2597,N_2998);
nor U3053 (N_3053,N_2751,N_2848);
and U3054 (N_3054,N_2806,N_2992);
and U3055 (N_3055,N_2889,N_2835);
nand U3056 (N_3056,N_2969,N_2531);
nor U3057 (N_3057,N_2795,N_2652);
or U3058 (N_3058,N_2860,N_2923);
nor U3059 (N_3059,N_2917,N_2807);
nor U3060 (N_3060,N_2891,N_2991);
and U3061 (N_3061,N_2857,N_2601);
nand U3062 (N_3062,N_2950,N_2980);
or U3063 (N_3063,N_2863,N_2689);
xnor U3064 (N_3064,N_2539,N_2914);
xnor U3065 (N_3065,N_2975,N_2545);
and U3066 (N_3066,N_2612,N_2758);
and U3067 (N_3067,N_2634,N_2804);
or U3068 (N_3068,N_2710,N_2756);
nor U3069 (N_3069,N_2638,N_2873);
or U3070 (N_3070,N_2583,N_2530);
xor U3071 (N_3071,N_2813,N_2567);
and U3072 (N_3072,N_2822,N_2724);
nand U3073 (N_3073,N_2659,N_2853);
xnor U3074 (N_3074,N_2760,N_2614);
nand U3075 (N_3075,N_2617,N_2830);
xor U3076 (N_3076,N_2818,N_2855);
nor U3077 (N_3077,N_2965,N_2745);
nor U3078 (N_3078,N_2611,N_2666);
nor U3079 (N_3079,N_2796,N_2690);
xnor U3080 (N_3080,N_2838,N_2527);
and U3081 (N_3081,N_2839,N_2893);
and U3082 (N_3082,N_2546,N_2772);
nand U3083 (N_3083,N_2894,N_2836);
nor U3084 (N_3084,N_2631,N_2517);
nor U3085 (N_3085,N_2909,N_2912);
xor U3086 (N_3086,N_2533,N_2506);
or U3087 (N_3087,N_2574,N_2828);
nand U3088 (N_3088,N_2968,N_2798);
or U3089 (N_3089,N_2757,N_2938);
or U3090 (N_3090,N_2592,N_2955);
and U3091 (N_3091,N_2790,N_2800);
xnor U3092 (N_3092,N_2878,N_2781);
and U3093 (N_3093,N_2624,N_2936);
nand U3094 (N_3094,N_2526,N_2755);
nor U3095 (N_3095,N_2887,N_2605);
nor U3096 (N_3096,N_2553,N_2637);
xnor U3097 (N_3097,N_2692,N_2874);
and U3098 (N_3098,N_2736,N_2985);
nand U3099 (N_3099,N_2532,N_2515);
nor U3100 (N_3100,N_2763,N_2586);
or U3101 (N_3101,N_2898,N_2983);
nand U3102 (N_3102,N_2881,N_2507);
nor U3103 (N_3103,N_2596,N_2904);
and U3104 (N_3104,N_2743,N_2884);
nor U3105 (N_3105,N_2984,N_2730);
nor U3106 (N_3106,N_2844,N_2832);
nor U3107 (N_3107,N_2951,N_2552);
nor U3108 (N_3108,N_2981,N_2669);
nand U3109 (N_3109,N_2570,N_2922);
nand U3110 (N_3110,N_2620,N_2698);
and U3111 (N_3111,N_2817,N_2952);
nor U3112 (N_3112,N_2875,N_2707);
nand U3113 (N_3113,N_2670,N_2554);
xnor U3114 (N_3114,N_2673,N_2559);
or U3115 (N_3115,N_2709,N_2843);
or U3116 (N_3116,N_2820,N_2908);
or U3117 (N_3117,N_2996,N_2930);
nand U3118 (N_3118,N_2880,N_2660);
nand U3119 (N_3119,N_2557,N_2713);
xnor U3120 (N_3120,N_2665,N_2607);
nor U3121 (N_3121,N_2537,N_2871);
nor U3122 (N_3122,N_2582,N_2516);
nor U3123 (N_3123,N_2957,N_2999);
nor U3124 (N_3124,N_2575,N_2558);
nand U3125 (N_3125,N_2555,N_2916);
nor U3126 (N_3126,N_2761,N_2608);
xor U3127 (N_3127,N_2791,N_2945);
and U3128 (N_3128,N_2667,N_2664);
nand U3129 (N_3129,N_2870,N_2547);
xor U3130 (N_3130,N_2905,N_2748);
nand U3131 (N_3131,N_2773,N_2716);
or U3132 (N_3132,N_2787,N_2851);
xor U3133 (N_3133,N_2769,N_2788);
xor U3134 (N_3134,N_2683,N_2747);
nor U3135 (N_3135,N_2837,N_2868);
and U3136 (N_3136,N_2779,N_2986);
and U3137 (N_3137,N_2503,N_2943);
or U3138 (N_3138,N_2602,N_2812);
and U3139 (N_3139,N_2926,N_2944);
nor U3140 (N_3140,N_2573,N_2882);
nand U3141 (N_3141,N_2677,N_2920);
nand U3142 (N_3142,N_2610,N_2719);
nand U3143 (N_3143,N_2825,N_2672);
nand U3144 (N_3144,N_2967,N_2799);
xnor U3145 (N_3145,N_2588,N_2896);
nor U3146 (N_3146,N_2703,N_2656);
nand U3147 (N_3147,N_2948,N_2746);
nand U3148 (N_3148,N_2892,N_2662);
nor U3149 (N_3149,N_2708,N_2613);
nand U3150 (N_3150,N_2840,N_2847);
or U3151 (N_3151,N_2543,N_2505);
xor U3152 (N_3152,N_2643,N_2595);
nand U3153 (N_3153,N_2768,N_2571);
and U3154 (N_3154,N_2642,N_2947);
and U3155 (N_3155,N_2551,N_2519);
and U3156 (N_3156,N_2589,N_2903);
or U3157 (N_3157,N_2598,N_2850);
or U3158 (N_3158,N_2895,N_2834);
and U3159 (N_3159,N_2886,N_2603);
nor U3160 (N_3160,N_2685,N_2577);
and U3161 (N_3161,N_2962,N_2681);
nand U3162 (N_3162,N_2949,N_2541);
xnor U3163 (N_3163,N_2585,N_2854);
nor U3164 (N_3164,N_2566,N_2528);
or U3165 (N_3165,N_2915,N_2792);
xnor U3166 (N_3166,N_2918,N_2864);
or U3167 (N_3167,N_2842,N_2679);
xnor U3168 (N_3168,N_2935,N_2504);
nor U3169 (N_3169,N_2959,N_2544);
or U3170 (N_3170,N_2648,N_2741);
nand U3171 (N_3171,N_2563,N_2737);
nor U3172 (N_3172,N_2816,N_2626);
and U3173 (N_3173,N_2686,N_2636);
nand U3174 (N_3174,N_2645,N_2901);
or U3175 (N_3175,N_2510,N_2801);
nand U3176 (N_3176,N_2688,N_2668);
or U3177 (N_3177,N_2629,N_2775);
and U3178 (N_3178,N_2988,N_2699);
nor U3179 (N_3179,N_2576,N_2717);
or U3180 (N_3180,N_2942,N_2911);
or U3181 (N_3181,N_2802,N_2604);
or U3182 (N_3182,N_2900,N_2759);
xor U3183 (N_3183,N_2764,N_2946);
nand U3184 (N_3184,N_2846,N_2572);
nand U3185 (N_3185,N_2867,N_2618);
xnor U3186 (N_3186,N_2811,N_2663);
nand U3187 (N_3187,N_2933,N_2704);
nand U3188 (N_3188,N_2523,N_2765);
and U3189 (N_3189,N_2518,N_2821);
xnor U3190 (N_3190,N_2976,N_2966);
nand U3191 (N_3191,N_2931,N_2954);
or U3192 (N_3192,N_2734,N_2815);
or U3193 (N_3193,N_2941,N_2720);
nand U3194 (N_3194,N_2639,N_2622);
xnor U3195 (N_3195,N_2899,N_2628);
nand U3196 (N_3196,N_2823,N_2919);
nor U3197 (N_3197,N_2621,N_2619);
nor U3198 (N_3198,N_2877,N_2785);
nand U3199 (N_3199,N_2897,N_2581);
nor U3200 (N_3200,N_2653,N_2525);
and U3201 (N_3201,N_2625,N_2964);
or U3202 (N_3202,N_2676,N_2989);
and U3203 (N_3203,N_2888,N_2978);
xor U3204 (N_3204,N_2956,N_2647);
and U3205 (N_3205,N_2778,N_2522);
nand U3206 (N_3206,N_2501,N_2754);
or U3207 (N_3207,N_2696,N_2782);
or U3208 (N_3208,N_2514,N_2678);
nand U3209 (N_3209,N_2587,N_2568);
nor U3210 (N_3210,N_2706,N_2762);
xor U3211 (N_3211,N_2562,N_2700);
xnor U3212 (N_3212,N_2814,N_2824);
xor U3213 (N_3213,N_2520,N_2869);
xor U3214 (N_3214,N_2970,N_2694);
xor U3215 (N_3215,N_2849,N_2937);
and U3216 (N_3216,N_2701,N_2594);
nand U3217 (N_3217,N_2714,N_2591);
and U3218 (N_3218,N_2509,N_2732);
nor U3219 (N_3219,N_2927,N_2829);
xnor U3220 (N_3220,N_2913,N_2657);
xnor U3221 (N_3221,N_2939,N_2742);
and U3222 (N_3222,N_2627,N_2827);
xor U3223 (N_3223,N_2808,N_2731);
xor U3224 (N_3224,N_2502,N_2924);
and U3225 (N_3225,N_2921,N_2655);
nand U3226 (N_3226,N_2671,N_2833);
nor U3227 (N_3227,N_2995,N_2876);
or U3228 (N_3228,N_2797,N_2644);
nor U3229 (N_3229,N_2925,N_2529);
nor U3230 (N_3230,N_2929,N_2780);
or U3231 (N_3231,N_2691,N_2858);
and U3232 (N_3232,N_2960,N_2831);
and U3233 (N_3233,N_2971,N_2907);
xor U3234 (N_3234,N_2993,N_2512);
xnor U3235 (N_3235,N_2508,N_2697);
or U3236 (N_3236,N_2674,N_2809);
or U3237 (N_3237,N_2542,N_2513);
and U3238 (N_3238,N_2744,N_2715);
and U3239 (N_3239,N_2953,N_2640);
nor U3240 (N_3240,N_2600,N_2616);
nand U3241 (N_3241,N_2722,N_2687);
or U3242 (N_3242,N_2632,N_2682);
nand U3243 (N_3243,N_2750,N_2770);
and U3244 (N_3244,N_2784,N_2721);
nand U3245 (N_3245,N_2910,N_2990);
xnor U3246 (N_3246,N_2550,N_2641);
and U3247 (N_3247,N_2649,N_2654);
and U3248 (N_3248,N_2749,N_2803);
or U3249 (N_3249,N_2599,N_2733);
and U3250 (N_3250,N_2535,N_2614);
xor U3251 (N_3251,N_2700,N_2504);
xnor U3252 (N_3252,N_2549,N_2615);
nor U3253 (N_3253,N_2589,N_2823);
xnor U3254 (N_3254,N_2545,N_2652);
and U3255 (N_3255,N_2683,N_2642);
or U3256 (N_3256,N_2813,N_2738);
or U3257 (N_3257,N_2710,N_2780);
or U3258 (N_3258,N_2700,N_2658);
xnor U3259 (N_3259,N_2746,N_2696);
and U3260 (N_3260,N_2797,N_2617);
xor U3261 (N_3261,N_2595,N_2789);
or U3262 (N_3262,N_2905,N_2783);
and U3263 (N_3263,N_2677,N_2684);
or U3264 (N_3264,N_2526,N_2564);
or U3265 (N_3265,N_2766,N_2733);
or U3266 (N_3266,N_2549,N_2800);
nand U3267 (N_3267,N_2923,N_2922);
or U3268 (N_3268,N_2671,N_2508);
and U3269 (N_3269,N_2857,N_2573);
or U3270 (N_3270,N_2775,N_2696);
nor U3271 (N_3271,N_2730,N_2890);
xor U3272 (N_3272,N_2992,N_2922);
nor U3273 (N_3273,N_2761,N_2600);
and U3274 (N_3274,N_2772,N_2647);
and U3275 (N_3275,N_2504,N_2839);
and U3276 (N_3276,N_2867,N_2696);
or U3277 (N_3277,N_2866,N_2787);
xor U3278 (N_3278,N_2949,N_2974);
or U3279 (N_3279,N_2931,N_2727);
nor U3280 (N_3280,N_2752,N_2837);
xnor U3281 (N_3281,N_2518,N_2938);
nand U3282 (N_3282,N_2592,N_2544);
and U3283 (N_3283,N_2703,N_2943);
nand U3284 (N_3284,N_2622,N_2508);
and U3285 (N_3285,N_2527,N_2824);
nand U3286 (N_3286,N_2641,N_2847);
nand U3287 (N_3287,N_2517,N_2681);
or U3288 (N_3288,N_2974,N_2610);
or U3289 (N_3289,N_2678,N_2568);
or U3290 (N_3290,N_2993,N_2795);
and U3291 (N_3291,N_2875,N_2767);
xnor U3292 (N_3292,N_2797,N_2895);
and U3293 (N_3293,N_2986,N_2879);
xnor U3294 (N_3294,N_2915,N_2511);
xor U3295 (N_3295,N_2849,N_2879);
nor U3296 (N_3296,N_2613,N_2991);
nand U3297 (N_3297,N_2870,N_2846);
nor U3298 (N_3298,N_2907,N_2678);
xnor U3299 (N_3299,N_2941,N_2815);
nor U3300 (N_3300,N_2900,N_2983);
or U3301 (N_3301,N_2849,N_2896);
xnor U3302 (N_3302,N_2916,N_2541);
and U3303 (N_3303,N_2576,N_2632);
nor U3304 (N_3304,N_2613,N_2916);
or U3305 (N_3305,N_2828,N_2630);
nand U3306 (N_3306,N_2738,N_2814);
nand U3307 (N_3307,N_2970,N_2640);
and U3308 (N_3308,N_2935,N_2925);
and U3309 (N_3309,N_2778,N_2886);
nand U3310 (N_3310,N_2811,N_2986);
or U3311 (N_3311,N_2817,N_2593);
nand U3312 (N_3312,N_2742,N_2965);
and U3313 (N_3313,N_2741,N_2561);
and U3314 (N_3314,N_2789,N_2815);
nand U3315 (N_3315,N_2631,N_2661);
nor U3316 (N_3316,N_2829,N_2860);
nor U3317 (N_3317,N_2604,N_2544);
or U3318 (N_3318,N_2904,N_2566);
or U3319 (N_3319,N_2853,N_2869);
xor U3320 (N_3320,N_2572,N_2765);
nor U3321 (N_3321,N_2606,N_2926);
nand U3322 (N_3322,N_2929,N_2955);
nor U3323 (N_3323,N_2948,N_2856);
and U3324 (N_3324,N_2585,N_2883);
nand U3325 (N_3325,N_2763,N_2571);
or U3326 (N_3326,N_2903,N_2766);
nand U3327 (N_3327,N_2527,N_2615);
and U3328 (N_3328,N_2851,N_2640);
and U3329 (N_3329,N_2749,N_2961);
or U3330 (N_3330,N_2715,N_2594);
or U3331 (N_3331,N_2707,N_2801);
or U3332 (N_3332,N_2958,N_2802);
and U3333 (N_3333,N_2868,N_2622);
and U3334 (N_3334,N_2655,N_2878);
or U3335 (N_3335,N_2819,N_2918);
nand U3336 (N_3336,N_2815,N_2802);
xor U3337 (N_3337,N_2797,N_2782);
nor U3338 (N_3338,N_2997,N_2917);
nand U3339 (N_3339,N_2941,N_2748);
or U3340 (N_3340,N_2757,N_2740);
nor U3341 (N_3341,N_2615,N_2727);
nor U3342 (N_3342,N_2879,N_2665);
xor U3343 (N_3343,N_2959,N_2548);
xnor U3344 (N_3344,N_2899,N_2730);
and U3345 (N_3345,N_2824,N_2719);
and U3346 (N_3346,N_2985,N_2621);
nand U3347 (N_3347,N_2659,N_2593);
or U3348 (N_3348,N_2547,N_2567);
nor U3349 (N_3349,N_2834,N_2827);
or U3350 (N_3350,N_2724,N_2777);
nand U3351 (N_3351,N_2684,N_2671);
xor U3352 (N_3352,N_2848,N_2999);
nand U3353 (N_3353,N_2956,N_2662);
nor U3354 (N_3354,N_2986,N_2891);
xor U3355 (N_3355,N_2924,N_2660);
or U3356 (N_3356,N_2794,N_2608);
and U3357 (N_3357,N_2630,N_2838);
nand U3358 (N_3358,N_2943,N_2850);
nand U3359 (N_3359,N_2660,N_2935);
and U3360 (N_3360,N_2549,N_2757);
nor U3361 (N_3361,N_2806,N_2757);
and U3362 (N_3362,N_2610,N_2538);
or U3363 (N_3363,N_2574,N_2851);
nor U3364 (N_3364,N_2726,N_2938);
xnor U3365 (N_3365,N_2679,N_2806);
nor U3366 (N_3366,N_2691,N_2835);
xnor U3367 (N_3367,N_2888,N_2615);
and U3368 (N_3368,N_2520,N_2533);
or U3369 (N_3369,N_2627,N_2570);
nand U3370 (N_3370,N_2534,N_2826);
nand U3371 (N_3371,N_2941,N_2733);
or U3372 (N_3372,N_2618,N_2558);
nand U3373 (N_3373,N_2823,N_2755);
xnor U3374 (N_3374,N_2836,N_2993);
or U3375 (N_3375,N_2998,N_2934);
and U3376 (N_3376,N_2567,N_2852);
nor U3377 (N_3377,N_2514,N_2552);
xor U3378 (N_3378,N_2869,N_2672);
and U3379 (N_3379,N_2606,N_2674);
nor U3380 (N_3380,N_2650,N_2545);
xor U3381 (N_3381,N_2776,N_2893);
nor U3382 (N_3382,N_2822,N_2626);
nor U3383 (N_3383,N_2550,N_2697);
or U3384 (N_3384,N_2936,N_2886);
or U3385 (N_3385,N_2637,N_2687);
or U3386 (N_3386,N_2671,N_2549);
nand U3387 (N_3387,N_2732,N_2686);
xor U3388 (N_3388,N_2831,N_2689);
nor U3389 (N_3389,N_2834,N_2503);
xor U3390 (N_3390,N_2910,N_2500);
xor U3391 (N_3391,N_2547,N_2786);
xnor U3392 (N_3392,N_2851,N_2540);
nor U3393 (N_3393,N_2993,N_2539);
nand U3394 (N_3394,N_2636,N_2708);
and U3395 (N_3395,N_2605,N_2886);
nand U3396 (N_3396,N_2736,N_2759);
nor U3397 (N_3397,N_2597,N_2527);
or U3398 (N_3398,N_2870,N_2903);
nand U3399 (N_3399,N_2981,N_2846);
and U3400 (N_3400,N_2603,N_2717);
or U3401 (N_3401,N_2582,N_2715);
and U3402 (N_3402,N_2595,N_2711);
and U3403 (N_3403,N_2538,N_2622);
nor U3404 (N_3404,N_2549,N_2811);
or U3405 (N_3405,N_2736,N_2975);
and U3406 (N_3406,N_2710,N_2993);
or U3407 (N_3407,N_2788,N_2599);
or U3408 (N_3408,N_2529,N_2777);
xnor U3409 (N_3409,N_2650,N_2519);
and U3410 (N_3410,N_2613,N_2753);
or U3411 (N_3411,N_2873,N_2613);
nand U3412 (N_3412,N_2721,N_2889);
nand U3413 (N_3413,N_2628,N_2932);
or U3414 (N_3414,N_2872,N_2911);
nand U3415 (N_3415,N_2565,N_2751);
nor U3416 (N_3416,N_2759,N_2801);
and U3417 (N_3417,N_2761,N_2616);
nor U3418 (N_3418,N_2680,N_2678);
nand U3419 (N_3419,N_2823,N_2757);
nor U3420 (N_3420,N_2750,N_2848);
xnor U3421 (N_3421,N_2607,N_2739);
nor U3422 (N_3422,N_2763,N_2949);
nand U3423 (N_3423,N_2850,N_2724);
xor U3424 (N_3424,N_2776,N_2918);
or U3425 (N_3425,N_2914,N_2617);
nor U3426 (N_3426,N_2812,N_2777);
nand U3427 (N_3427,N_2745,N_2514);
and U3428 (N_3428,N_2714,N_2770);
or U3429 (N_3429,N_2723,N_2612);
nand U3430 (N_3430,N_2943,N_2531);
and U3431 (N_3431,N_2934,N_2776);
and U3432 (N_3432,N_2796,N_2773);
or U3433 (N_3433,N_2586,N_2908);
and U3434 (N_3434,N_2513,N_2819);
nand U3435 (N_3435,N_2539,N_2562);
nand U3436 (N_3436,N_2725,N_2665);
nor U3437 (N_3437,N_2936,N_2769);
nand U3438 (N_3438,N_2860,N_2928);
or U3439 (N_3439,N_2870,N_2676);
xor U3440 (N_3440,N_2541,N_2745);
and U3441 (N_3441,N_2555,N_2949);
xor U3442 (N_3442,N_2949,N_2729);
xor U3443 (N_3443,N_2539,N_2822);
nor U3444 (N_3444,N_2861,N_2583);
xor U3445 (N_3445,N_2638,N_2796);
or U3446 (N_3446,N_2872,N_2856);
or U3447 (N_3447,N_2765,N_2702);
xor U3448 (N_3448,N_2898,N_2730);
or U3449 (N_3449,N_2776,N_2552);
and U3450 (N_3450,N_2614,N_2910);
or U3451 (N_3451,N_2619,N_2939);
nand U3452 (N_3452,N_2531,N_2538);
nor U3453 (N_3453,N_2882,N_2528);
and U3454 (N_3454,N_2672,N_2854);
and U3455 (N_3455,N_2737,N_2627);
nor U3456 (N_3456,N_2510,N_2796);
nor U3457 (N_3457,N_2755,N_2751);
nand U3458 (N_3458,N_2980,N_2780);
nor U3459 (N_3459,N_2548,N_2993);
nand U3460 (N_3460,N_2561,N_2719);
nand U3461 (N_3461,N_2696,N_2592);
nand U3462 (N_3462,N_2720,N_2725);
and U3463 (N_3463,N_2933,N_2615);
or U3464 (N_3464,N_2962,N_2628);
nand U3465 (N_3465,N_2901,N_2985);
nand U3466 (N_3466,N_2925,N_2874);
xor U3467 (N_3467,N_2552,N_2731);
xor U3468 (N_3468,N_2768,N_2932);
nor U3469 (N_3469,N_2716,N_2740);
xnor U3470 (N_3470,N_2960,N_2699);
or U3471 (N_3471,N_2954,N_2994);
nand U3472 (N_3472,N_2623,N_2889);
xor U3473 (N_3473,N_2647,N_2991);
or U3474 (N_3474,N_2992,N_2730);
nand U3475 (N_3475,N_2792,N_2564);
nand U3476 (N_3476,N_2623,N_2983);
and U3477 (N_3477,N_2825,N_2578);
xnor U3478 (N_3478,N_2795,N_2845);
and U3479 (N_3479,N_2844,N_2946);
xor U3480 (N_3480,N_2939,N_2673);
nor U3481 (N_3481,N_2625,N_2722);
and U3482 (N_3482,N_2903,N_2718);
nand U3483 (N_3483,N_2949,N_2688);
nor U3484 (N_3484,N_2501,N_2800);
nor U3485 (N_3485,N_2872,N_2608);
nand U3486 (N_3486,N_2791,N_2640);
or U3487 (N_3487,N_2884,N_2835);
nor U3488 (N_3488,N_2721,N_2765);
xnor U3489 (N_3489,N_2839,N_2698);
or U3490 (N_3490,N_2575,N_2552);
nor U3491 (N_3491,N_2878,N_2701);
and U3492 (N_3492,N_2934,N_2640);
xor U3493 (N_3493,N_2900,N_2640);
xor U3494 (N_3494,N_2710,N_2817);
xnor U3495 (N_3495,N_2682,N_2961);
xor U3496 (N_3496,N_2627,N_2890);
xnor U3497 (N_3497,N_2642,N_2946);
xor U3498 (N_3498,N_2613,N_2510);
and U3499 (N_3499,N_2534,N_2917);
nand U3500 (N_3500,N_3287,N_3152);
or U3501 (N_3501,N_3151,N_3265);
xor U3502 (N_3502,N_3492,N_3069);
and U3503 (N_3503,N_3298,N_3293);
and U3504 (N_3504,N_3436,N_3462);
nor U3505 (N_3505,N_3381,N_3208);
xor U3506 (N_3506,N_3183,N_3187);
or U3507 (N_3507,N_3249,N_3203);
nand U3508 (N_3508,N_3380,N_3311);
or U3509 (N_3509,N_3474,N_3005);
nand U3510 (N_3510,N_3410,N_3202);
nand U3511 (N_3511,N_3021,N_3269);
or U3512 (N_3512,N_3169,N_3391);
nor U3513 (N_3513,N_3161,N_3285);
or U3514 (N_3514,N_3344,N_3351);
or U3515 (N_3515,N_3482,N_3240);
or U3516 (N_3516,N_3128,N_3211);
nand U3517 (N_3517,N_3075,N_3115);
and U3518 (N_3518,N_3369,N_3233);
nand U3519 (N_3519,N_3071,N_3460);
nor U3520 (N_3520,N_3363,N_3100);
or U3521 (N_3521,N_3254,N_3135);
nor U3522 (N_3522,N_3372,N_3461);
xnor U3523 (N_3523,N_3347,N_3076);
xnor U3524 (N_3524,N_3070,N_3330);
xnor U3525 (N_3525,N_3230,N_3166);
xnor U3526 (N_3526,N_3379,N_3019);
xnor U3527 (N_3527,N_3471,N_3095);
nand U3528 (N_3528,N_3270,N_3283);
xor U3529 (N_3529,N_3332,N_3335);
nor U3530 (N_3530,N_3341,N_3091);
xnor U3531 (N_3531,N_3286,N_3360);
xnor U3532 (N_3532,N_3093,N_3246);
and U3533 (N_3533,N_3419,N_3013);
nand U3534 (N_3534,N_3188,N_3025);
or U3535 (N_3535,N_3088,N_3168);
or U3536 (N_3536,N_3144,N_3141);
and U3537 (N_3537,N_3412,N_3239);
xnor U3538 (N_3538,N_3043,N_3241);
and U3539 (N_3539,N_3484,N_3117);
xnor U3540 (N_3540,N_3264,N_3138);
nand U3541 (N_3541,N_3464,N_3159);
nand U3542 (N_3542,N_3050,N_3487);
nor U3543 (N_3543,N_3328,N_3001);
or U3544 (N_3544,N_3319,N_3062);
and U3545 (N_3545,N_3139,N_3416);
nand U3546 (N_3546,N_3178,N_3185);
or U3547 (N_3547,N_3219,N_3366);
nor U3548 (N_3548,N_3370,N_3180);
and U3549 (N_3549,N_3130,N_3408);
or U3550 (N_3550,N_3457,N_3313);
nor U3551 (N_3551,N_3488,N_3068);
nand U3552 (N_3552,N_3358,N_3172);
xnor U3553 (N_3553,N_3498,N_3384);
or U3554 (N_3554,N_3491,N_3237);
or U3555 (N_3555,N_3432,N_3429);
or U3556 (N_3556,N_3404,N_3063);
and U3557 (N_3557,N_3163,N_3158);
nor U3558 (N_3558,N_3496,N_3060);
and U3559 (N_3559,N_3026,N_3442);
nand U3560 (N_3560,N_3094,N_3009);
xnor U3561 (N_3561,N_3251,N_3247);
or U3562 (N_3562,N_3443,N_3170);
nor U3563 (N_3563,N_3295,N_3108);
or U3564 (N_3564,N_3036,N_3015);
nand U3565 (N_3565,N_3260,N_3463);
nand U3566 (N_3566,N_3055,N_3216);
or U3567 (N_3567,N_3282,N_3389);
or U3568 (N_3568,N_3343,N_3054);
and U3569 (N_3569,N_3092,N_3024);
nand U3570 (N_3570,N_3248,N_3387);
and U3571 (N_3571,N_3477,N_3478);
or U3572 (N_3572,N_3084,N_3284);
xor U3573 (N_3573,N_3255,N_3263);
and U3574 (N_3574,N_3048,N_3225);
nor U3575 (N_3575,N_3258,N_3367);
nor U3576 (N_3576,N_3215,N_3278);
and U3577 (N_3577,N_3401,N_3197);
nor U3578 (N_3578,N_3354,N_3087);
nand U3579 (N_3579,N_3164,N_3348);
and U3580 (N_3580,N_3171,N_3276);
and U3581 (N_3581,N_3101,N_3450);
or U3582 (N_3582,N_3281,N_3148);
or U3583 (N_3583,N_3065,N_3362);
nand U3584 (N_3584,N_3377,N_3274);
and U3585 (N_3585,N_3074,N_3103);
nand U3586 (N_3586,N_3038,N_3323);
or U3587 (N_3587,N_3481,N_3018);
or U3588 (N_3588,N_3205,N_3275);
nand U3589 (N_3589,N_3453,N_3376);
and U3590 (N_3590,N_3353,N_3226);
or U3591 (N_3591,N_3468,N_3245);
xnor U3592 (N_3592,N_3058,N_3427);
or U3593 (N_3593,N_3433,N_3217);
nor U3594 (N_3594,N_3243,N_3256);
nor U3595 (N_3595,N_3489,N_3388);
nand U3596 (N_3596,N_3244,N_3032);
nand U3597 (N_3597,N_3181,N_3102);
nand U3598 (N_3598,N_3470,N_3198);
xor U3599 (N_3599,N_3459,N_3368);
and U3600 (N_3600,N_3097,N_3434);
and U3601 (N_3601,N_3324,N_3157);
nand U3602 (N_3602,N_3339,N_3131);
nor U3603 (N_3603,N_3266,N_3016);
xnor U3604 (N_3604,N_3320,N_3020);
xor U3605 (N_3605,N_3277,N_3235);
xor U3606 (N_3606,N_3194,N_3415);
nor U3607 (N_3607,N_3373,N_3007);
xnor U3608 (N_3608,N_3112,N_3150);
nand U3609 (N_3609,N_3064,N_3073);
xnor U3610 (N_3610,N_3398,N_3333);
and U3611 (N_3611,N_3458,N_3405);
or U3612 (N_3612,N_3124,N_3214);
or U3613 (N_3613,N_3155,N_3302);
nand U3614 (N_3614,N_3116,N_3307);
or U3615 (N_3615,N_3126,N_3114);
or U3616 (N_3616,N_3083,N_3191);
xnor U3617 (N_3617,N_3306,N_3223);
or U3618 (N_3618,N_3394,N_3209);
xnor U3619 (N_3619,N_3140,N_3454);
nor U3620 (N_3620,N_3082,N_3123);
and U3621 (N_3621,N_3400,N_3292);
xnor U3622 (N_3622,N_3467,N_3029);
and U3623 (N_3623,N_3494,N_3099);
xor U3624 (N_3624,N_3035,N_3145);
xor U3625 (N_3625,N_3407,N_3109);
or U3626 (N_3626,N_3193,N_3111);
or U3627 (N_3627,N_3120,N_3200);
nand U3628 (N_3628,N_3066,N_3056);
xor U3629 (N_3629,N_3149,N_3315);
or U3630 (N_3630,N_3497,N_3395);
xor U3631 (N_3631,N_3196,N_3228);
nor U3632 (N_3632,N_3049,N_3080);
xnor U3633 (N_3633,N_3231,N_3397);
and U3634 (N_3634,N_3238,N_3143);
or U3635 (N_3635,N_3014,N_3051);
or U3636 (N_3636,N_3137,N_3349);
or U3637 (N_3637,N_3411,N_3096);
and U3638 (N_3638,N_3224,N_3352);
xor U3639 (N_3639,N_3012,N_3086);
xnor U3640 (N_3640,N_3418,N_3406);
nor U3641 (N_3641,N_3437,N_3428);
nand U3642 (N_3642,N_3227,N_3345);
nor U3643 (N_3643,N_3420,N_3299);
and U3644 (N_3644,N_3493,N_3179);
nand U3645 (N_3645,N_3375,N_3318);
nand U3646 (N_3646,N_3220,N_3340);
and U3647 (N_3647,N_3403,N_3210);
or U3648 (N_3648,N_3393,N_3356);
nor U3649 (N_3649,N_3153,N_3317);
nor U3650 (N_3650,N_3221,N_3003);
nand U3651 (N_3651,N_3177,N_3127);
xor U3652 (N_3652,N_3142,N_3472);
nor U3653 (N_3653,N_3473,N_3113);
nand U3654 (N_3654,N_3034,N_3273);
xor U3655 (N_3655,N_3422,N_3378);
or U3656 (N_3656,N_3479,N_3184);
xor U3657 (N_3657,N_3288,N_3175);
nand U3658 (N_3658,N_3030,N_3077);
and U3659 (N_3659,N_3465,N_3390);
nand U3660 (N_3660,N_3441,N_3399);
and U3661 (N_3661,N_3485,N_3119);
and U3662 (N_3662,N_3371,N_3483);
nand U3663 (N_3663,N_3106,N_3162);
and U3664 (N_3664,N_3435,N_3259);
nand U3665 (N_3665,N_3331,N_3440);
xnor U3666 (N_3666,N_3052,N_3027);
nand U3667 (N_3667,N_3334,N_3006);
xnor U3668 (N_3668,N_3300,N_3361);
or U3669 (N_3669,N_3438,N_3396);
nor U3670 (N_3670,N_3122,N_3059);
nor U3671 (N_3671,N_3325,N_3469);
or U3672 (N_3672,N_3312,N_3046);
or U3673 (N_3673,N_3409,N_3426);
and U3674 (N_3674,N_3207,N_3303);
nand U3675 (N_3675,N_3451,N_3297);
or U3676 (N_3676,N_3425,N_3495);
and U3677 (N_3677,N_3133,N_3037);
nand U3678 (N_3678,N_3189,N_3430);
nor U3679 (N_3679,N_3304,N_3008);
and U3680 (N_3680,N_3085,N_3147);
nand U3681 (N_3681,N_3456,N_3121);
and U3682 (N_3682,N_3039,N_3364);
and U3683 (N_3683,N_3212,N_3421);
nand U3684 (N_3684,N_3042,N_3402);
xnor U3685 (N_3685,N_3031,N_3480);
xnor U3686 (N_3686,N_3218,N_3466);
xor U3687 (N_3687,N_3053,N_3195);
xor U3688 (N_3688,N_3268,N_3250);
xor U3689 (N_3689,N_3475,N_3321);
or U3690 (N_3690,N_3261,N_3444);
or U3691 (N_3691,N_3308,N_3327);
and U3692 (N_3692,N_3182,N_3383);
and U3693 (N_3693,N_3253,N_3090);
nor U3694 (N_3694,N_3301,N_3252);
and U3695 (N_3695,N_3271,N_3448);
xnor U3696 (N_3696,N_3222,N_3173);
nor U3697 (N_3697,N_3431,N_3232);
or U3698 (N_3698,N_3004,N_3326);
nor U3699 (N_3699,N_3417,N_3079);
or U3700 (N_3700,N_3040,N_3022);
xor U3701 (N_3701,N_3165,N_3010);
nand U3702 (N_3702,N_3146,N_3002);
nand U3703 (N_3703,N_3374,N_3045);
nand U3704 (N_3704,N_3176,N_3229);
xor U3705 (N_3705,N_3309,N_3291);
nand U3706 (N_3706,N_3098,N_3033);
and U3707 (N_3707,N_3338,N_3105);
nor U3708 (N_3708,N_3199,N_3129);
nor U3709 (N_3709,N_3186,N_3204);
nand U3710 (N_3710,N_3242,N_3439);
xor U3711 (N_3711,N_3452,N_3365);
xor U3712 (N_3712,N_3447,N_3322);
and U3713 (N_3713,N_3446,N_3310);
nor U3714 (N_3714,N_3262,N_3167);
xor U3715 (N_3715,N_3044,N_3089);
and U3716 (N_3716,N_3067,N_3078);
xnor U3717 (N_3717,N_3386,N_3449);
and U3718 (N_3718,N_3424,N_3294);
xor U3719 (N_3719,N_3414,N_3041);
xnor U3720 (N_3720,N_3190,N_3160);
nor U3721 (N_3721,N_3455,N_3342);
or U3722 (N_3722,N_3104,N_3423);
or U3723 (N_3723,N_3234,N_3017);
nor U3724 (N_3724,N_3192,N_3314);
xor U3725 (N_3725,N_3476,N_3201);
and U3726 (N_3726,N_3280,N_3305);
nor U3727 (N_3727,N_3499,N_3000);
and U3728 (N_3728,N_3174,N_3486);
nand U3729 (N_3729,N_3107,N_3490);
and U3730 (N_3730,N_3154,N_3257);
nor U3731 (N_3731,N_3385,N_3357);
nor U3732 (N_3732,N_3296,N_3359);
and U3733 (N_3733,N_3011,N_3057);
and U3734 (N_3734,N_3156,N_3445);
or U3735 (N_3735,N_3350,N_3329);
xnor U3736 (N_3736,N_3316,N_3213);
or U3737 (N_3737,N_3337,N_3336);
nand U3738 (N_3738,N_3125,N_3118);
nand U3739 (N_3739,N_3081,N_3132);
or U3740 (N_3740,N_3028,N_3047);
nor U3741 (N_3741,N_3289,N_3272);
nand U3742 (N_3742,N_3061,N_3206);
nand U3743 (N_3743,N_3413,N_3236);
and U3744 (N_3744,N_3023,N_3136);
or U3745 (N_3745,N_3072,N_3290);
and U3746 (N_3746,N_3382,N_3346);
xor U3747 (N_3747,N_3134,N_3279);
nand U3748 (N_3748,N_3267,N_3392);
nand U3749 (N_3749,N_3110,N_3355);
xnor U3750 (N_3750,N_3415,N_3417);
xnor U3751 (N_3751,N_3044,N_3425);
xor U3752 (N_3752,N_3473,N_3367);
xnor U3753 (N_3753,N_3403,N_3481);
nor U3754 (N_3754,N_3442,N_3189);
nand U3755 (N_3755,N_3167,N_3131);
and U3756 (N_3756,N_3232,N_3334);
nor U3757 (N_3757,N_3073,N_3198);
and U3758 (N_3758,N_3132,N_3431);
xnor U3759 (N_3759,N_3275,N_3181);
xor U3760 (N_3760,N_3386,N_3049);
xnor U3761 (N_3761,N_3482,N_3239);
or U3762 (N_3762,N_3315,N_3037);
nand U3763 (N_3763,N_3342,N_3196);
or U3764 (N_3764,N_3033,N_3339);
nand U3765 (N_3765,N_3155,N_3339);
nor U3766 (N_3766,N_3273,N_3195);
nand U3767 (N_3767,N_3291,N_3176);
nor U3768 (N_3768,N_3370,N_3468);
nand U3769 (N_3769,N_3095,N_3419);
or U3770 (N_3770,N_3209,N_3492);
or U3771 (N_3771,N_3369,N_3381);
xor U3772 (N_3772,N_3468,N_3312);
nor U3773 (N_3773,N_3315,N_3064);
nand U3774 (N_3774,N_3275,N_3062);
or U3775 (N_3775,N_3291,N_3184);
or U3776 (N_3776,N_3099,N_3419);
nor U3777 (N_3777,N_3417,N_3264);
xnor U3778 (N_3778,N_3019,N_3332);
or U3779 (N_3779,N_3338,N_3083);
and U3780 (N_3780,N_3270,N_3252);
xor U3781 (N_3781,N_3038,N_3041);
xor U3782 (N_3782,N_3015,N_3491);
and U3783 (N_3783,N_3273,N_3456);
xnor U3784 (N_3784,N_3372,N_3122);
xor U3785 (N_3785,N_3398,N_3026);
or U3786 (N_3786,N_3462,N_3207);
or U3787 (N_3787,N_3092,N_3103);
or U3788 (N_3788,N_3125,N_3202);
nand U3789 (N_3789,N_3460,N_3022);
xnor U3790 (N_3790,N_3470,N_3407);
nand U3791 (N_3791,N_3025,N_3424);
nor U3792 (N_3792,N_3115,N_3256);
nand U3793 (N_3793,N_3001,N_3342);
nand U3794 (N_3794,N_3279,N_3357);
nor U3795 (N_3795,N_3342,N_3144);
or U3796 (N_3796,N_3315,N_3226);
nor U3797 (N_3797,N_3432,N_3161);
nor U3798 (N_3798,N_3300,N_3014);
nand U3799 (N_3799,N_3428,N_3031);
nand U3800 (N_3800,N_3348,N_3481);
nand U3801 (N_3801,N_3098,N_3144);
nor U3802 (N_3802,N_3152,N_3253);
and U3803 (N_3803,N_3354,N_3031);
nand U3804 (N_3804,N_3330,N_3363);
nor U3805 (N_3805,N_3344,N_3011);
and U3806 (N_3806,N_3474,N_3322);
xor U3807 (N_3807,N_3057,N_3459);
or U3808 (N_3808,N_3104,N_3469);
nor U3809 (N_3809,N_3470,N_3403);
xnor U3810 (N_3810,N_3355,N_3303);
or U3811 (N_3811,N_3485,N_3339);
nor U3812 (N_3812,N_3210,N_3320);
and U3813 (N_3813,N_3297,N_3487);
xnor U3814 (N_3814,N_3363,N_3021);
nor U3815 (N_3815,N_3047,N_3434);
and U3816 (N_3816,N_3251,N_3406);
or U3817 (N_3817,N_3087,N_3162);
nor U3818 (N_3818,N_3121,N_3087);
nand U3819 (N_3819,N_3345,N_3146);
nor U3820 (N_3820,N_3443,N_3039);
or U3821 (N_3821,N_3062,N_3130);
xor U3822 (N_3822,N_3359,N_3334);
xnor U3823 (N_3823,N_3305,N_3177);
nor U3824 (N_3824,N_3000,N_3318);
xor U3825 (N_3825,N_3330,N_3045);
or U3826 (N_3826,N_3385,N_3325);
xor U3827 (N_3827,N_3461,N_3381);
nor U3828 (N_3828,N_3199,N_3013);
and U3829 (N_3829,N_3208,N_3274);
nor U3830 (N_3830,N_3297,N_3357);
and U3831 (N_3831,N_3150,N_3016);
or U3832 (N_3832,N_3280,N_3479);
and U3833 (N_3833,N_3413,N_3374);
and U3834 (N_3834,N_3365,N_3297);
nand U3835 (N_3835,N_3245,N_3177);
xor U3836 (N_3836,N_3119,N_3064);
nand U3837 (N_3837,N_3058,N_3118);
or U3838 (N_3838,N_3086,N_3050);
xor U3839 (N_3839,N_3087,N_3019);
nand U3840 (N_3840,N_3290,N_3241);
nor U3841 (N_3841,N_3309,N_3076);
or U3842 (N_3842,N_3350,N_3464);
or U3843 (N_3843,N_3209,N_3002);
nand U3844 (N_3844,N_3091,N_3271);
xnor U3845 (N_3845,N_3164,N_3156);
nand U3846 (N_3846,N_3007,N_3487);
and U3847 (N_3847,N_3397,N_3235);
xor U3848 (N_3848,N_3083,N_3072);
nor U3849 (N_3849,N_3176,N_3352);
nor U3850 (N_3850,N_3155,N_3321);
and U3851 (N_3851,N_3055,N_3488);
xor U3852 (N_3852,N_3179,N_3337);
xor U3853 (N_3853,N_3419,N_3077);
xnor U3854 (N_3854,N_3452,N_3329);
or U3855 (N_3855,N_3459,N_3378);
xor U3856 (N_3856,N_3083,N_3412);
xnor U3857 (N_3857,N_3148,N_3267);
xnor U3858 (N_3858,N_3299,N_3163);
or U3859 (N_3859,N_3062,N_3041);
xnor U3860 (N_3860,N_3095,N_3149);
xor U3861 (N_3861,N_3408,N_3412);
or U3862 (N_3862,N_3280,N_3255);
or U3863 (N_3863,N_3398,N_3148);
nor U3864 (N_3864,N_3423,N_3122);
or U3865 (N_3865,N_3443,N_3333);
or U3866 (N_3866,N_3180,N_3462);
and U3867 (N_3867,N_3411,N_3331);
xnor U3868 (N_3868,N_3215,N_3369);
xor U3869 (N_3869,N_3278,N_3393);
nand U3870 (N_3870,N_3428,N_3438);
nand U3871 (N_3871,N_3188,N_3349);
nand U3872 (N_3872,N_3491,N_3330);
or U3873 (N_3873,N_3457,N_3352);
nor U3874 (N_3874,N_3379,N_3432);
or U3875 (N_3875,N_3172,N_3035);
nor U3876 (N_3876,N_3020,N_3037);
and U3877 (N_3877,N_3400,N_3020);
nand U3878 (N_3878,N_3065,N_3462);
nor U3879 (N_3879,N_3119,N_3284);
and U3880 (N_3880,N_3368,N_3341);
and U3881 (N_3881,N_3180,N_3393);
xnor U3882 (N_3882,N_3212,N_3487);
nand U3883 (N_3883,N_3289,N_3265);
nand U3884 (N_3884,N_3334,N_3466);
or U3885 (N_3885,N_3223,N_3355);
and U3886 (N_3886,N_3474,N_3313);
nor U3887 (N_3887,N_3281,N_3405);
xor U3888 (N_3888,N_3285,N_3496);
nand U3889 (N_3889,N_3139,N_3037);
or U3890 (N_3890,N_3202,N_3071);
xnor U3891 (N_3891,N_3471,N_3339);
xnor U3892 (N_3892,N_3259,N_3222);
and U3893 (N_3893,N_3315,N_3488);
or U3894 (N_3894,N_3021,N_3156);
or U3895 (N_3895,N_3218,N_3140);
and U3896 (N_3896,N_3272,N_3227);
xor U3897 (N_3897,N_3030,N_3333);
nor U3898 (N_3898,N_3176,N_3202);
and U3899 (N_3899,N_3046,N_3497);
or U3900 (N_3900,N_3230,N_3168);
xnor U3901 (N_3901,N_3007,N_3315);
nor U3902 (N_3902,N_3311,N_3206);
or U3903 (N_3903,N_3427,N_3339);
and U3904 (N_3904,N_3048,N_3435);
nor U3905 (N_3905,N_3145,N_3459);
nand U3906 (N_3906,N_3273,N_3431);
and U3907 (N_3907,N_3048,N_3208);
nand U3908 (N_3908,N_3409,N_3342);
and U3909 (N_3909,N_3063,N_3384);
xnor U3910 (N_3910,N_3380,N_3301);
and U3911 (N_3911,N_3022,N_3443);
and U3912 (N_3912,N_3254,N_3113);
xor U3913 (N_3913,N_3274,N_3218);
nand U3914 (N_3914,N_3051,N_3497);
xnor U3915 (N_3915,N_3113,N_3325);
nand U3916 (N_3916,N_3333,N_3272);
nor U3917 (N_3917,N_3146,N_3261);
or U3918 (N_3918,N_3301,N_3098);
xnor U3919 (N_3919,N_3231,N_3002);
nand U3920 (N_3920,N_3467,N_3435);
nor U3921 (N_3921,N_3090,N_3429);
and U3922 (N_3922,N_3499,N_3058);
nor U3923 (N_3923,N_3280,N_3090);
or U3924 (N_3924,N_3020,N_3496);
or U3925 (N_3925,N_3250,N_3328);
xnor U3926 (N_3926,N_3364,N_3144);
or U3927 (N_3927,N_3259,N_3138);
xor U3928 (N_3928,N_3319,N_3418);
or U3929 (N_3929,N_3435,N_3104);
nand U3930 (N_3930,N_3350,N_3398);
nand U3931 (N_3931,N_3302,N_3499);
or U3932 (N_3932,N_3218,N_3077);
and U3933 (N_3933,N_3276,N_3485);
nand U3934 (N_3934,N_3157,N_3044);
xor U3935 (N_3935,N_3022,N_3234);
xor U3936 (N_3936,N_3042,N_3380);
or U3937 (N_3937,N_3308,N_3110);
and U3938 (N_3938,N_3140,N_3000);
or U3939 (N_3939,N_3124,N_3332);
nor U3940 (N_3940,N_3488,N_3129);
nor U3941 (N_3941,N_3099,N_3340);
xor U3942 (N_3942,N_3481,N_3276);
xor U3943 (N_3943,N_3365,N_3417);
xor U3944 (N_3944,N_3074,N_3118);
or U3945 (N_3945,N_3446,N_3118);
and U3946 (N_3946,N_3107,N_3221);
or U3947 (N_3947,N_3018,N_3085);
or U3948 (N_3948,N_3069,N_3237);
or U3949 (N_3949,N_3474,N_3470);
or U3950 (N_3950,N_3346,N_3138);
nand U3951 (N_3951,N_3180,N_3040);
nand U3952 (N_3952,N_3289,N_3105);
and U3953 (N_3953,N_3239,N_3410);
nand U3954 (N_3954,N_3320,N_3060);
nor U3955 (N_3955,N_3278,N_3106);
or U3956 (N_3956,N_3486,N_3050);
and U3957 (N_3957,N_3394,N_3139);
and U3958 (N_3958,N_3301,N_3034);
nand U3959 (N_3959,N_3448,N_3256);
xor U3960 (N_3960,N_3385,N_3333);
xnor U3961 (N_3961,N_3143,N_3424);
or U3962 (N_3962,N_3104,N_3498);
nand U3963 (N_3963,N_3340,N_3079);
nor U3964 (N_3964,N_3280,N_3339);
or U3965 (N_3965,N_3384,N_3094);
and U3966 (N_3966,N_3050,N_3064);
nand U3967 (N_3967,N_3389,N_3472);
and U3968 (N_3968,N_3235,N_3091);
xor U3969 (N_3969,N_3446,N_3479);
nor U3970 (N_3970,N_3258,N_3123);
and U3971 (N_3971,N_3391,N_3492);
nor U3972 (N_3972,N_3446,N_3121);
xor U3973 (N_3973,N_3191,N_3445);
nand U3974 (N_3974,N_3453,N_3207);
nor U3975 (N_3975,N_3289,N_3071);
or U3976 (N_3976,N_3058,N_3350);
xnor U3977 (N_3977,N_3395,N_3417);
nand U3978 (N_3978,N_3190,N_3221);
and U3979 (N_3979,N_3136,N_3421);
or U3980 (N_3980,N_3153,N_3265);
nand U3981 (N_3981,N_3254,N_3474);
or U3982 (N_3982,N_3108,N_3315);
and U3983 (N_3983,N_3123,N_3233);
xor U3984 (N_3984,N_3350,N_3308);
or U3985 (N_3985,N_3390,N_3023);
and U3986 (N_3986,N_3227,N_3329);
xor U3987 (N_3987,N_3495,N_3203);
nor U3988 (N_3988,N_3399,N_3114);
nor U3989 (N_3989,N_3451,N_3021);
xor U3990 (N_3990,N_3111,N_3226);
and U3991 (N_3991,N_3227,N_3261);
nand U3992 (N_3992,N_3358,N_3028);
or U3993 (N_3993,N_3170,N_3395);
nor U3994 (N_3994,N_3219,N_3194);
xnor U3995 (N_3995,N_3300,N_3488);
nor U3996 (N_3996,N_3375,N_3431);
xnor U3997 (N_3997,N_3472,N_3088);
and U3998 (N_3998,N_3363,N_3135);
or U3999 (N_3999,N_3174,N_3293);
xor U4000 (N_4000,N_3589,N_3896);
xnor U4001 (N_4001,N_3904,N_3549);
or U4002 (N_4002,N_3895,N_3544);
xor U4003 (N_4003,N_3835,N_3829);
and U4004 (N_4004,N_3581,N_3543);
nor U4005 (N_4005,N_3652,N_3721);
or U4006 (N_4006,N_3719,N_3909);
nand U4007 (N_4007,N_3618,N_3849);
xnor U4008 (N_4008,N_3729,N_3922);
xor U4009 (N_4009,N_3881,N_3833);
or U4010 (N_4010,N_3750,N_3523);
xnor U4011 (N_4011,N_3999,N_3793);
and U4012 (N_4012,N_3805,N_3850);
nor U4013 (N_4013,N_3848,N_3605);
and U4014 (N_4014,N_3563,N_3948);
nand U4015 (N_4015,N_3715,N_3570);
nand U4016 (N_4016,N_3816,N_3866);
nor U4017 (N_4017,N_3954,N_3545);
nor U4018 (N_4018,N_3770,N_3837);
xor U4019 (N_4019,N_3513,N_3594);
nand U4020 (N_4020,N_3892,N_3553);
nor U4021 (N_4021,N_3635,N_3655);
or U4022 (N_4022,N_3644,N_3834);
xnor U4023 (N_4023,N_3539,N_3855);
xor U4024 (N_4024,N_3813,N_3661);
nand U4025 (N_4025,N_3502,N_3871);
xor U4026 (N_4026,N_3706,N_3559);
and U4027 (N_4027,N_3615,N_3981);
nand U4028 (N_4028,N_3970,N_3908);
xnor U4029 (N_4029,N_3645,N_3976);
xor U4030 (N_4030,N_3572,N_3932);
and U4031 (N_4031,N_3510,N_3529);
xnor U4032 (N_4032,N_3936,N_3868);
or U4033 (N_4033,N_3537,N_3643);
or U4034 (N_4034,N_3769,N_3694);
xor U4035 (N_4035,N_3962,N_3957);
and U4036 (N_4036,N_3608,N_3956);
xnor U4037 (N_4037,N_3836,N_3761);
nor U4038 (N_4038,N_3940,N_3565);
or U4039 (N_4039,N_3937,N_3610);
and U4040 (N_4040,N_3910,N_3822);
nor U4041 (N_4041,N_3964,N_3617);
xnor U4042 (N_4042,N_3671,N_3782);
xor U4043 (N_4043,N_3784,N_3975);
or U4044 (N_4044,N_3906,N_3742);
or U4045 (N_4045,N_3744,N_3709);
and U4046 (N_4046,N_3753,N_3585);
xnor U4047 (N_4047,N_3823,N_3710);
nand U4048 (N_4048,N_3607,N_3959);
nand U4049 (N_4049,N_3503,N_3686);
or U4050 (N_4050,N_3552,N_3548);
and U4051 (N_4051,N_3984,N_3526);
and U4052 (N_4052,N_3820,N_3575);
or U4053 (N_4053,N_3878,N_3807);
xnor U4054 (N_4054,N_3724,N_3638);
xnor U4055 (N_4055,N_3772,N_3560);
or U4056 (N_4056,N_3893,N_3625);
xor U4057 (N_4057,N_3576,N_3612);
and U4058 (N_4058,N_3691,N_3872);
nor U4059 (N_4059,N_3704,N_3765);
xnor U4060 (N_4060,N_3851,N_3831);
nand U4061 (N_4061,N_3662,N_3762);
or U4062 (N_4062,N_3681,N_3799);
nand U4063 (N_4063,N_3883,N_3597);
nor U4064 (N_4064,N_3989,N_3876);
nor U4065 (N_4065,N_3860,N_3651);
nor U4066 (N_4066,N_3916,N_3749);
nand U4067 (N_4067,N_3887,N_3619);
xor U4068 (N_4068,N_3740,N_3828);
nand U4069 (N_4069,N_3821,N_3663);
nand U4070 (N_4070,N_3569,N_3856);
nand U4071 (N_4071,N_3726,N_3693);
xnor U4072 (N_4072,N_3930,N_3787);
xor U4073 (N_4073,N_3789,N_3527);
and U4074 (N_4074,N_3616,N_3689);
or U4075 (N_4075,N_3889,N_3777);
nand U4076 (N_4076,N_3997,N_3556);
and U4077 (N_4077,N_3773,N_3683);
and U4078 (N_4078,N_3796,N_3631);
nor U4079 (N_4079,N_3657,N_3621);
nor U4080 (N_4080,N_3938,N_3590);
nand U4081 (N_4081,N_3842,N_3562);
xnor U4082 (N_4082,N_3682,N_3911);
or U4083 (N_4083,N_3953,N_3500);
or U4084 (N_4084,N_3532,N_3687);
nor U4085 (N_4085,N_3546,N_3806);
nor U4086 (N_4086,N_3763,N_3571);
xor U4087 (N_4087,N_3656,N_3741);
xnor U4088 (N_4088,N_3788,N_3604);
xor U4089 (N_4089,N_3992,N_3944);
nand U4090 (N_4090,N_3733,N_3776);
and U4091 (N_4091,N_3918,N_3901);
xor U4092 (N_4092,N_3504,N_3880);
and U4093 (N_4093,N_3598,N_3913);
or U4094 (N_4094,N_3809,N_3637);
nor U4095 (N_4095,N_3923,N_3915);
and U4096 (N_4096,N_3790,N_3942);
nand U4097 (N_4097,N_3819,N_3648);
nand U4098 (N_4098,N_3963,N_3949);
nor U4099 (N_4099,N_3755,N_3952);
xnor U4100 (N_4100,N_3567,N_3622);
or U4101 (N_4101,N_3812,N_3522);
nor U4102 (N_4102,N_3903,N_3982);
or U4103 (N_4103,N_3700,N_3533);
nor U4104 (N_4104,N_3641,N_3929);
or U4105 (N_4105,N_3875,N_3584);
or U4106 (N_4106,N_3863,N_3670);
or U4107 (N_4107,N_3877,N_3905);
or U4108 (N_4108,N_3558,N_3582);
or U4109 (N_4109,N_3639,N_3826);
and U4110 (N_4110,N_3852,N_3780);
and U4111 (N_4111,N_3583,N_3841);
and U4112 (N_4112,N_3939,N_3974);
xor U4113 (N_4113,N_3623,N_3511);
nor U4114 (N_4114,N_3536,N_3707);
and U4115 (N_4115,N_3606,N_3611);
or U4116 (N_4116,N_3557,N_3517);
and U4117 (N_4117,N_3705,N_3534);
nand U4118 (N_4118,N_3767,N_3673);
nor U4119 (N_4119,N_3547,N_3731);
nand U4120 (N_4120,N_3718,N_3794);
and U4121 (N_4121,N_3737,N_3966);
xnor U4122 (N_4122,N_3603,N_3775);
or U4123 (N_4123,N_3506,N_3814);
or U4124 (N_4124,N_3679,N_3847);
xor U4125 (N_4125,N_3926,N_3843);
xor U4126 (N_4126,N_3587,N_3519);
or U4127 (N_4127,N_3745,N_3697);
nor U4128 (N_4128,N_3924,N_3508);
nor U4129 (N_4129,N_3858,N_3988);
and U4130 (N_4130,N_3665,N_3595);
nand U4131 (N_4131,N_3902,N_3779);
nand U4132 (N_4132,N_3853,N_3596);
nand U4133 (N_4133,N_3830,N_3946);
xnor U4134 (N_4134,N_3566,N_3739);
nand U4135 (N_4135,N_3531,N_3521);
nor U4136 (N_4136,N_3890,N_3907);
nand U4137 (N_4137,N_3934,N_3840);
nor U4138 (N_4138,N_3732,N_3771);
xor U4139 (N_4139,N_3817,N_3630);
or U4140 (N_4140,N_3685,N_3698);
and U4141 (N_4141,N_3525,N_3757);
xor U4142 (N_4142,N_3854,N_3586);
xor U4143 (N_4143,N_3978,N_3973);
nor U4144 (N_4144,N_3735,N_3738);
and U4145 (N_4145,N_3632,N_3714);
or U4146 (N_4146,N_3925,N_3897);
xnor U4147 (N_4147,N_3542,N_3520);
nand U4148 (N_4148,N_3554,N_3713);
nand U4149 (N_4149,N_3752,N_3985);
nor U4150 (N_4150,N_3561,N_3620);
nand U4151 (N_4151,N_3869,N_3690);
nand U4152 (N_4152,N_3550,N_3990);
xor U4153 (N_4153,N_3825,N_3873);
nand U4154 (N_4154,N_3882,N_3800);
xnor U4155 (N_4155,N_3688,N_3748);
and U4156 (N_4156,N_3518,N_3955);
or U4157 (N_4157,N_3960,N_3991);
and U4158 (N_4158,N_3803,N_3899);
or U4159 (N_4159,N_3845,N_3633);
or U4160 (N_4160,N_3658,N_3797);
nor U4161 (N_4161,N_3951,N_3666);
or U4162 (N_4162,N_3993,N_3592);
xnor U4163 (N_4163,N_3920,N_3599);
and U4164 (N_4164,N_3839,N_3676);
xor U4165 (N_4165,N_3678,N_3950);
and U4166 (N_4166,N_3514,N_3540);
nand U4167 (N_4167,N_3660,N_3675);
and U4168 (N_4168,N_3535,N_3695);
and U4169 (N_4169,N_3811,N_3818);
or U4170 (N_4170,N_3986,N_3600);
nor U4171 (N_4171,N_3696,N_3580);
nor U4172 (N_4172,N_3931,N_3838);
and U4173 (N_4173,N_3867,N_3998);
and U4174 (N_4174,N_3588,N_3528);
nor U4175 (N_4175,N_3703,N_3568);
nor U4176 (N_4176,N_3827,N_3798);
nand U4177 (N_4177,N_3774,N_3968);
or U4178 (N_4178,N_3751,N_3971);
xor U4179 (N_4179,N_3958,N_3538);
or U4180 (N_4180,N_3870,N_3824);
nand U4181 (N_4181,N_3720,N_3626);
and U4182 (N_4182,N_3781,N_3579);
nor U4183 (N_4183,N_3783,N_3601);
nand U4184 (N_4184,N_3564,N_3636);
and U4185 (N_4185,N_3702,N_3524);
xor U4186 (N_4186,N_3766,N_3578);
xnor U4187 (N_4187,N_3791,N_3802);
nand U4188 (N_4188,N_3865,N_3634);
nand U4189 (N_4189,N_3515,N_3972);
nor U4190 (N_4190,N_3627,N_3747);
and U4191 (N_4191,N_3602,N_3743);
or U4192 (N_4192,N_3888,N_3857);
or U4193 (N_4193,N_3995,N_3754);
nand U4194 (N_4194,N_3609,N_3987);
xnor U4195 (N_4195,N_3591,N_3967);
nand U4196 (N_4196,N_3912,N_3680);
nand U4197 (N_4197,N_3507,N_3624);
xnor U4198 (N_4198,N_3884,N_3760);
nand U4199 (N_4199,N_3674,N_3629);
xnor U4200 (N_4200,N_3501,N_3891);
and U4201 (N_4201,N_3977,N_3917);
and U4202 (N_4202,N_3722,N_3677);
and U4203 (N_4203,N_3961,N_3933);
xor U4204 (N_4204,N_3921,N_3699);
nand U4205 (N_4205,N_3654,N_3672);
xnor U4206 (N_4206,N_3900,N_3832);
or U4207 (N_4207,N_3684,N_3945);
and U4208 (N_4208,N_3885,N_3725);
or U4209 (N_4209,N_3659,N_3530);
and U4210 (N_4210,N_3717,N_3759);
nand U4211 (N_4211,N_3555,N_3758);
xor U4212 (N_4212,N_3516,N_3914);
xnor U4213 (N_4213,N_3943,N_3716);
xnor U4214 (N_4214,N_3574,N_3804);
xor U4215 (N_4215,N_3736,N_3711);
xnor U4216 (N_4216,N_3509,N_3669);
and U4217 (N_4217,N_3996,N_3668);
nand U4218 (N_4218,N_3746,N_3730);
xor U4219 (N_4219,N_3894,N_3667);
xor U4220 (N_4220,N_3898,N_3756);
and U4221 (N_4221,N_3768,N_3649);
or U4222 (N_4222,N_3573,N_3593);
or U4223 (N_4223,N_3815,N_3701);
nand U4224 (N_4224,N_3708,N_3614);
and U4225 (N_4225,N_3613,N_3935);
xor U4226 (N_4226,N_3640,N_3664);
xnor U4227 (N_4227,N_3928,N_3505);
or U4228 (N_4228,N_3653,N_3941);
xnor U4229 (N_4229,N_3778,N_3846);
nand U4230 (N_4230,N_3808,N_3785);
or U4231 (N_4231,N_3650,N_3795);
nand U4232 (N_4232,N_3927,N_3628);
and U4233 (N_4233,N_3879,N_3994);
or U4234 (N_4234,N_3844,N_3727);
nor U4235 (N_4235,N_3692,N_3786);
nand U4236 (N_4236,N_3764,N_3712);
xor U4237 (N_4237,N_3969,N_3647);
nor U4238 (N_4238,N_3980,N_3577);
nand U4239 (N_4239,N_3979,N_3541);
xnor U4240 (N_4240,N_3792,N_3919);
nor U4241 (N_4241,N_3728,N_3864);
or U4242 (N_4242,N_3965,N_3512);
and U4243 (N_4243,N_3859,N_3551);
or U4244 (N_4244,N_3886,N_3723);
nor U4245 (N_4245,N_3642,N_3861);
xnor U4246 (N_4246,N_3801,N_3983);
xnor U4247 (N_4247,N_3862,N_3874);
nand U4248 (N_4248,N_3734,N_3646);
xor U4249 (N_4249,N_3947,N_3810);
xnor U4250 (N_4250,N_3940,N_3694);
nor U4251 (N_4251,N_3730,N_3781);
and U4252 (N_4252,N_3622,N_3764);
nand U4253 (N_4253,N_3643,N_3585);
and U4254 (N_4254,N_3609,N_3957);
or U4255 (N_4255,N_3950,N_3713);
nor U4256 (N_4256,N_3795,N_3615);
nor U4257 (N_4257,N_3584,N_3890);
nor U4258 (N_4258,N_3998,N_3762);
or U4259 (N_4259,N_3757,N_3651);
nand U4260 (N_4260,N_3936,N_3844);
or U4261 (N_4261,N_3991,N_3506);
or U4262 (N_4262,N_3590,N_3879);
nor U4263 (N_4263,N_3747,N_3956);
or U4264 (N_4264,N_3758,N_3878);
xnor U4265 (N_4265,N_3631,N_3936);
and U4266 (N_4266,N_3954,N_3919);
xnor U4267 (N_4267,N_3785,N_3893);
or U4268 (N_4268,N_3811,N_3950);
xnor U4269 (N_4269,N_3653,N_3936);
nand U4270 (N_4270,N_3765,N_3777);
xor U4271 (N_4271,N_3865,N_3522);
and U4272 (N_4272,N_3644,N_3645);
nand U4273 (N_4273,N_3797,N_3694);
and U4274 (N_4274,N_3742,N_3640);
nand U4275 (N_4275,N_3983,N_3500);
nor U4276 (N_4276,N_3569,N_3869);
nor U4277 (N_4277,N_3580,N_3721);
nor U4278 (N_4278,N_3661,N_3725);
and U4279 (N_4279,N_3641,N_3508);
nand U4280 (N_4280,N_3974,N_3828);
or U4281 (N_4281,N_3887,N_3967);
xor U4282 (N_4282,N_3746,N_3786);
nand U4283 (N_4283,N_3549,N_3930);
nor U4284 (N_4284,N_3926,N_3704);
and U4285 (N_4285,N_3862,N_3532);
xor U4286 (N_4286,N_3609,N_3820);
nor U4287 (N_4287,N_3718,N_3614);
nor U4288 (N_4288,N_3591,N_3787);
nor U4289 (N_4289,N_3526,N_3811);
nor U4290 (N_4290,N_3944,N_3695);
nand U4291 (N_4291,N_3589,N_3772);
nand U4292 (N_4292,N_3884,N_3952);
nor U4293 (N_4293,N_3698,N_3560);
nand U4294 (N_4294,N_3705,N_3686);
xor U4295 (N_4295,N_3898,N_3572);
nand U4296 (N_4296,N_3873,N_3723);
nor U4297 (N_4297,N_3956,N_3819);
nand U4298 (N_4298,N_3837,N_3561);
nor U4299 (N_4299,N_3932,N_3770);
or U4300 (N_4300,N_3926,N_3959);
or U4301 (N_4301,N_3992,N_3993);
and U4302 (N_4302,N_3519,N_3612);
xnor U4303 (N_4303,N_3697,N_3721);
or U4304 (N_4304,N_3972,N_3956);
nor U4305 (N_4305,N_3542,N_3740);
and U4306 (N_4306,N_3620,N_3717);
nor U4307 (N_4307,N_3584,N_3752);
nand U4308 (N_4308,N_3849,N_3807);
xnor U4309 (N_4309,N_3567,N_3692);
nor U4310 (N_4310,N_3963,N_3673);
and U4311 (N_4311,N_3824,N_3641);
nand U4312 (N_4312,N_3547,N_3884);
and U4313 (N_4313,N_3677,N_3746);
xnor U4314 (N_4314,N_3934,N_3534);
nor U4315 (N_4315,N_3984,N_3986);
nand U4316 (N_4316,N_3619,N_3545);
xnor U4317 (N_4317,N_3946,N_3810);
and U4318 (N_4318,N_3699,N_3817);
or U4319 (N_4319,N_3708,N_3730);
xor U4320 (N_4320,N_3989,N_3705);
or U4321 (N_4321,N_3529,N_3655);
nand U4322 (N_4322,N_3858,N_3688);
or U4323 (N_4323,N_3669,N_3684);
or U4324 (N_4324,N_3713,N_3758);
nor U4325 (N_4325,N_3802,N_3970);
and U4326 (N_4326,N_3602,N_3519);
or U4327 (N_4327,N_3794,N_3590);
or U4328 (N_4328,N_3759,N_3501);
nand U4329 (N_4329,N_3545,N_3961);
nand U4330 (N_4330,N_3977,N_3957);
nand U4331 (N_4331,N_3711,N_3943);
and U4332 (N_4332,N_3598,N_3989);
nor U4333 (N_4333,N_3541,N_3893);
or U4334 (N_4334,N_3857,N_3965);
and U4335 (N_4335,N_3657,N_3762);
nor U4336 (N_4336,N_3515,N_3505);
nor U4337 (N_4337,N_3695,N_3890);
and U4338 (N_4338,N_3560,N_3845);
xor U4339 (N_4339,N_3600,N_3910);
nand U4340 (N_4340,N_3600,N_3837);
or U4341 (N_4341,N_3627,N_3830);
and U4342 (N_4342,N_3539,N_3700);
xor U4343 (N_4343,N_3514,N_3774);
or U4344 (N_4344,N_3926,N_3875);
and U4345 (N_4345,N_3826,N_3646);
and U4346 (N_4346,N_3677,N_3619);
xnor U4347 (N_4347,N_3852,N_3980);
or U4348 (N_4348,N_3767,N_3895);
nand U4349 (N_4349,N_3935,N_3948);
or U4350 (N_4350,N_3573,N_3982);
xnor U4351 (N_4351,N_3796,N_3581);
nor U4352 (N_4352,N_3741,N_3546);
xnor U4353 (N_4353,N_3998,N_3975);
and U4354 (N_4354,N_3730,N_3920);
xor U4355 (N_4355,N_3546,N_3654);
or U4356 (N_4356,N_3905,N_3741);
and U4357 (N_4357,N_3853,N_3844);
nand U4358 (N_4358,N_3864,N_3909);
xnor U4359 (N_4359,N_3686,N_3567);
xnor U4360 (N_4360,N_3512,N_3945);
and U4361 (N_4361,N_3902,N_3805);
or U4362 (N_4362,N_3628,N_3891);
or U4363 (N_4363,N_3799,N_3914);
nand U4364 (N_4364,N_3988,N_3996);
and U4365 (N_4365,N_3629,N_3583);
nand U4366 (N_4366,N_3941,N_3750);
and U4367 (N_4367,N_3520,N_3867);
or U4368 (N_4368,N_3588,N_3999);
nor U4369 (N_4369,N_3866,N_3771);
nand U4370 (N_4370,N_3995,N_3607);
nand U4371 (N_4371,N_3649,N_3949);
and U4372 (N_4372,N_3729,N_3844);
xnor U4373 (N_4373,N_3819,N_3774);
nand U4374 (N_4374,N_3901,N_3919);
xnor U4375 (N_4375,N_3938,N_3935);
xor U4376 (N_4376,N_3873,N_3881);
nor U4377 (N_4377,N_3789,N_3635);
or U4378 (N_4378,N_3986,N_3913);
nand U4379 (N_4379,N_3885,N_3950);
xnor U4380 (N_4380,N_3774,N_3734);
and U4381 (N_4381,N_3539,N_3839);
nand U4382 (N_4382,N_3861,N_3796);
or U4383 (N_4383,N_3540,N_3813);
and U4384 (N_4384,N_3568,N_3550);
xnor U4385 (N_4385,N_3533,N_3841);
nor U4386 (N_4386,N_3836,N_3941);
nor U4387 (N_4387,N_3664,N_3794);
or U4388 (N_4388,N_3630,N_3739);
nand U4389 (N_4389,N_3542,N_3585);
and U4390 (N_4390,N_3781,N_3793);
nand U4391 (N_4391,N_3959,N_3800);
nor U4392 (N_4392,N_3852,N_3609);
xor U4393 (N_4393,N_3807,N_3520);
nor U4394 (N_4394,N_3752,N_3891);
nand U4395 (N_4395,N_3979,N_3921);
or U4396 (N_4396,N_3801,N_3607);
nand U4397 (N_4397,N_3886,N_3969);
nor U4398 (N_4398,N_3714,N_3666);
xnor U4399 (N_4399,N_3888,N_3739);
and U4400 (N_4400,N_3711,N_3740);
or U4401 (N_4401,N_3578,N_3521);
and U4402 (N_4402,N_3845,N_3867);
nor U4403 (N_4403,N_3717,N_3909);
xnor U4404 (N_4404,N_3944,N_3805);
and U4405 (N_4405,N_3794,N_3957);
xor U4406 (N_4406,N_3693,N_3959);
nand U4407 (N_4407,N_3535,N_3942);
nand U4408 (N_4408,N_3572,N_3778);
and U4409 (N_4409,N_3955,N_3570);
nand U4410 (N_4410,N_3501,N_3794);
nor U4411 (N_4411,N_3723,N_3934);
or U4412 (N_4412,N_3579,N_3651);
nand U4413 (N_4413,N_3545,N_3802);
or U4414 (N_4414,N_3839,N_3583);
xnor U4415 (N_4415,N_3560,N_3525);
nand U4416 (N_4416,N_3648,N_3634);
nor U4417 (N_4417,N_3571,N_3560);
nand U4418 (N_4418,N_3928,N_3758);
xor U4419 (N_4419,N_3904,N_3836);
xor U4420 (N_4420,N_3909,N_3722);
and U4421 (N_4421,N_3752,N_3707);
nor U4422 (N_4422,N_3710,N_3754);
nand U4423 (N_4423,N_3533,N_3966);
or U4424 (N_4424,N_3814,N_3787);
nor U4425 (N_4425,N_3995,N_3832);
nand U4426 (N_4426,N_3952,N_3730);
or U4427 (N_4427,N_3510,N_3741);
xnor U4428 (N_4428,N_3749,N_3847);
or U4429 (N_4429,N_3971,N_3848);
xnor U4430 (N_4430,N_3866,N_3994);
and U4431 (N_4431,N_3950,N_3810);
xnor U4432 (N_4432,N_3958,N_3793);
and U4433 (N_4433,N_3653,N_3761);
and U4434 (N_4434,N_3868,N_3850);
and U4435 (N_4435,N_3923,N_3605);
nand U4436 (N_4436,N_3804,N_3952);
and U4437 (N_4437,N_3558,N_3943);
xor U4438 (N_4438,N_3520,N_3577);
xnor U4439 (N_4439,N_3925,N_3772);
nor U4440 (N_4440,N_3857,N_3619);
xor U4441 (N_4441,N_3993,N_3916);
nor U4442 (N_4442,N_3771,N_3673);
nand U4443 (N_4443,N_3763,N_3981);
or U4444 (N_4444,N_3633,N_3809);
and U4445 (N_4445,N_3817,N_3860);
nor U4446 (N_4446,N_3564,N_3701);
and U4447 (N_4447,N_3515,N_3944);
nand U4448 (N_4448,N_3825,N_3608);
nand U4449 (N_4449,N_3634,N_3782);
nor U4450 (N_4450,N_3567,N_3587);
xor U4451 (N_4451,N_3742,N_3589);
nor U4452 (N_4452,N_3947,N_3613);
nor U4453 (N_4453,N_3816,N_3749);
nor U4454 (N_4454,N_3800,N_3593);
nand U4455 (N_4455,N_3591,N_3814);
nand U4456 (N_4456,N_3890,N_3744);
xor U4457 (N_4457,N_3843,N_3708);
xor U4458 (N_4458,N_3753,N_3846);
nor U4459 (N_4459,N_3553,N_3956);
or U4460 (N_4460,N_3998,N_3950);
nand U4461 (N_4461,N_3766,N_3721);
xor U4462 (N_4462,N_3911,N_3686);
nor U4463 (N_4463,N_3624,N_3709);
xnor U4464 (N_4464,N_3797,N_3944);
nor U4465 (N_4465,N_3815,N_3956);
xor U4466 (N_4466,N_3923,N_3924);
nand U4467 (N_4467,N_3852,N_3506);
or U4468 (N_4468,N_3691,N_3844);
nand U4469 (N_4469,N_3971,N_3792);
nor U4470 (N_4470,N_3938,N_3623);
or U4471 (N_4471,N_3637,N_3613);
xor U4472 (N_4472,N_3519,N_3938);
nand U4473 (N_4473,N_3732,N_3533);
xor U4474 (N_4474,N_3750,N_3774);
xnor U4475 (N_4475,N_3786,N_3616);
or U4476 (N_4476,N_3871,N_3731);
or U4477 (N_4477,N_3524,N_3595);
nor U4478 (N_4478,N_3791,N_3671);
and U4479 (N_4479,N_3535,N_3950);
and U4480 (N_4480,N_3844,N_3705);
nand U4481 (N_4481,N_3956,N_3706);
xor U4482 (N_4482,N_3834,N_3699);
nand U4483 (N_4483,N_3857,N_3735);
nand U4484 (N_4484,N_3640,N_3617);
nor U4485 (N_4485,N_3544,N_3660);
nor U4486 (N_4486,N_3867,N_3815);
or U4487 (N_4487,N_3541,N_3845);
or U4488 (N_4488,N_3996,N_3631);
xnor U4489 (N_4489,N_3934,N_3814);
nor U4490 (N_4490,N_3590,N_3993);
nor U4491 (N_4491,N_3657,N_3797);
nor U4492 (N_4492,N_3704,N_3965);
and U4493 (N_4493,N_3882,N_3728);
or U4494 (N_4494,N_3594,N_3613);
or U4495 (N_4495,N_3844,N_3745);
or U4496 (N_4496,N_3946,N_3985);
and U4497 (N_4497,N_3847,N_3825);
xnor U4498 (N_4498,N_3643,N_3851);
nor U4499 (N_4499,N_3540,N_3561);
or U4500 (N_4500,N_4040,N_4436);
and U4501 (N_4501,N_4478,N_4056);
nor U4502 (N_4502,N_4295,N_4074);
nor U4503 (N_4503,N_4270,N_4389);
and U4504 (N_4504,N_4324,N_4087);
nor U4505 (N_4505,N_4227,N_4150);
or U4506 (N_4506,N_4058,N_4396);
xor U4507 (N_4507,N_4197,N_4151);
and U4508 (N_4508,N_4114,N_4276);
or U4509 (N_4509,N_4112,N_4440);
nor U4510 (N_4510,N_4143,N_4242);
or U4511 (N_4511,N_4362,N_4264);
and U4512 (N_4512,N_4186,N_4119);
or U4513 (N_4513,N_4002,N_4431);
or U4514 (N_4514,N_4003,N_4130);
or U4515 (N_4515,N_4022,N_4366);
nand U4516 (N_4516,N_4424,N_4020);
or U4517 (N_4517,N_4164,N_4344);
xor U4518 (N_4518,N_4419,N_4069);
xnor U4519 (N_4519,N_4350,N_4443);
xor U4520 (N_4520,N_4499,N_4065);
and U4521 (N_4521,N_4116,N_4356);
xor U4522 (N_4522,N_4289,N_4059);
and U4523 (N_4523,N_4086,N_4325);
nor U4524 (N_4524,N_4391,N_4206);
or U4525 (N_4525,N_4024,N_4070);
nor U4526 (N_4526,N_4146,N_4081);
nand U4527 (N_4527,N_4266,N_4472);
nand U4528 (N_4528,N_4029,N_4100);
xnor U4529 (N_4529,N_4294,N_4099);
nand U4530 (N_4530,N_4042,N_4037);
nand U4531 (N_4531,N_4192,N_4371);
nand U4532 (N_4532,N_4488,N_4032);
or U4533 (N_4533,N_4133,N_4171);
nor U4534 (N_4534,N_4177,N_4101);
xnor U4535 (N_4535,N_4298,N_4082);
nor U4536 (N_4536,N_4135,N_4202);
or U4537 (N_4537,N_4327,N_4441);
nand U4538 (N_4538,N_4148,N_4169);
nand U4539 (N_4539,N_4231,N_4317);
nor U4540 (N_4540,N_4288,N_4492);
xnor U4541 (N_4541,N_4010,N_4140);
and U4542 (N_4542,N_4398,N_4246);
nor U4543 (N_4543,N_4115,N_4016);
nand U4544 (N_4544,N_4291,N_4428);
xnor U4545 (N_4545,N_4092,N_4282);
nand U4546 (N_4546,N_4374,N_4085);
or U4547 (N_4547,N_4057,N_4489);
and U4548 (N_4548,N_4377,N_4018);
xor U4549 (N_4549,N_4027,N_4342);
xnor U4550 (N_4550,N_4222,N_4215);
xnor U4551 (N_4551,N_4256,N_4267);
or U4552 (N_4552,N_4038,N_4439);
or U4553 (N_4553,N_4455,N_4471);
nor U4554 (N_4554,N_4111,N_4296);
nor U4555 (N_4555,N_4201,N_4425);
or U4556 (N_4556,N_4286,N_4163);
xor U4557 (N_4557,N_4254,N_4383);
nor U4558 (N_4558,N_4360,N_4370);
nor U4559 (N_4559,N_4262,N_4249);
nor U4560 (N_4560,N_4292,N_4039);
nor U4561 (N_4561,N_4104,N_4494);
or U4562 (N_4562,N_4071,N_4308);
and U4563 (N_4563,N_4060,N_4180);
and U4564 (N_4564,N_4109,N_4329);
xnor U4565 (N_4565,N_4273,N_4028);
nor U4566 (N_4566,N_4481,N_4390);
or U4567 (N_4567,N_4218,N_4339);
xnor U4568 (N_4568,N_4012,N_4280);
and U4569 (N_4569,N_4093,N_4077);
nand U4570 (N_4570,N_4462,N_4330);
nand U4571 (N_4571,N_4051,N_4278);
and U4572 (N_4572,N_4106,N_4036);
and U4573 (N_4573,N_4458,N_4275);
or U4574 (N_4574,N_4126,N_4376);
xnor U4575 (N_4575,N_4001,N_4220);
nor U4576 (N_4576,N_4303,N_4486);
or U4577 (N_4577,N_4435,N_4427);
or U4578 (N_4578,N_4351,N_4041);
and U4579 (N_4579,N_4411,N_4026);
nand U4580 (N_4580,N_4234,N_4166);
and U4581 (N_4581,N_4083,N_4252);
or U4582 (N_4582,N_4145,N_4283);
xor U4583 (N_4583,N_4449,N_4117);
xnor U4584 (N_4584,N_4284,N_4346);
and U4585 (N_4585,N_4238,N_4033);
or U4586 (N_4586,N_4442,N_4023);
nand U4587 (N_4587,N_4347,N_4451);
or U4588 (N_4588,N_4399,N_4408);
nand U4589 (N_4589,N_4352,N_4341);
and U4590 (N_4590,N_4009,N_4415);
or U4591 (N_4591,N_4063,N_4345);
and U4592 (N_4592,N_4405,N_4088);
or U4593 (N_4593,N_4107,N_4250);
nand U4594 (N_4594,N_4476,N_4105);
nor U4595 (N_4595,N_4331,N_4263);
nand U4596 (N_4596,N_4230,N_4307);
or U4597 (N_4597,N_4300,N_4365);
and U4598 (N_4598,N_4168,N_4233);
xor U4599 (N_4599,N_4011,N_4387);
nor U4600 (N_4600,N_4248,N_4096);
or U4601 (N_4601,N_4224,N_4239);
and U4602 (N_4602,N_4064,N_4310);
or U4603 (N_4603,N_4272,N_4416);
or U4604 (N_4604,N_4091,N_4279);
and U4605 (N_4605,N_4301,N_4102);
nand U4606 (N_4606,N_4223,N_4355);
or U4607 (N_4607,N_4311,N_4477);
xor U4608 (N_4608,N_4373,N_4050);
xnor U4609 (N_4609,N_4113,N_4174);
nand U4610 (N_4610,N_4067,N_4313);
or U4611 (N_4611,N_4004,N_4209);
xor U4612 (N_4612,N_4090,N_4097);
or U4613 (N_4613,N_4053,N_4395);
and U4614 (N_4614,N_4255,N_4228);
nand U4615 (N_4615,N_4274,N_4429);
nor U4616 (N_4616,N_4221,N_4400);
nand U4617 (N_4617,N_4258,N_4229);
nand U4618 (N_4618,N_4332,N_4123);
or U4619 (N_4619,N_4485,N_4170);
nand U4620 (N_4620,N_4072,N_4196);
xor U4621 (N_4621,N_4384,N_4375);
nand U4622 (N_4622,N_4464,N_4453);
nand U4623 (N_4623,N_4232,N_4179);
or U4624 (N_4624,N_4075,N_4021);
and U4625 (N_4625,N_4066,N_4208);
nand U4626 (N_4626,N_4259,N_4401);
and U4627 (N_4627,N_4412,N_4445);
or U4628 (N_4628,N_4446,N_4349);
nand U4629 (N_4629,N_4095,N_4277);
or U4630 (N_4630,N_4413,N_4461);
nor U4631 (N_4631,N_4434,N_4318);
and U4632 (N_4632,N_4369,N_4414);
and U4633 (N_4633,N_4194,N_4203);
nor U4634 (N_4634,N_4118,N_4237);
xor U4635 (N_4635,N_4245,N_4156);
xor U4636 (N_4636,N_4185,N_4198);
nor U4637 (N_4637,N_4199,N_4493);
or U4638 (N_4638,N_4079,N_4271);
or U4639 (N_4639,N_4187,N_4147);
nor U4640 (N_4640,N_4315,N_4423);
nor U4641 (N_4641,N_4265,N_4212);
and U4642 (N_4642,N_4404,N_4172);
or U4643 (N_4643,N_4139,N_4162);
xnor U4644 (N_4644,N_4410,N_4188);
nor U4645 (N_4645,N_4189,N_4054);
nand U4646 (N_4646,N_4025,N_4035);
nand U4647 (N_4647,N_4055,N_4382);
and U4648 (N_4648,N_4154,N_4491);
or U4649 (N_4649,N_4498,N_4019);
or U4650 (N_4650,N_4062,N_4463);
and U4651 (N_4651,N_4049,N_4497);
nor U4652 (N_4652,N_4293,N_4084);
xnor U4653 (N_4653,N_4098,N_4184);
nor U4654 (N_4654,N_4321,N_4142);
or U4655 (N_4655,N_4269,N_4473);
xor U4656 (N_4656,N_4363,N_4468);
nand U4657 (N_4657,N_4261,N_4122);
or U4658 (N_4658,N_4178,N_4046);
nand U4659 (N_4659,N_4422,N_4030);
nor U4660 (N_4660,N_4433,N_4299);
xnor U4661 (N_4661,N_4323,N_4125);
and U4662 (N_4662,N_4474,N_4452);
nand U4663 (N_4663,N_4225,N_4044);
and U4664 (N_4664,N_4136,N_4240);
nand U4665 (N_4665,N_4287,N_4159);
nand U4666 (N_4666,N_4052,N_4448);
xor U4667 (N_4667,N_4161,N_4421);
and U4668 (N_4668,N_4467,N_4333);
nor U4669 (N_4669,N_4454,N_4359);
and U4670 (N_4670,N_4204,N_4361);
xnor U4671 (N_4671,N_4379,N_4432);
xor U4672 (N_4672,N_4348,N_4137);
nor U4673 (N_4673,N_4153,N_4381);
and U4674 (N_4674,N_4406,N_4495);
xnor U4675 (N_4675,N_4110,N_4320);
and U4676 (N_4676,N_4173,N_4155);
nand U4677 (N_4677,N_4141,N_4068);
and U4678 (N_4678,N_4005,N_4243);
nand U4679 (N_4679,N_4484,N_4129);
or U4680 (N_4680,N_4437,N_4205);
nand U4681 (N_4681,N_4089,N_4364);
and U4682 (N_4682,N_4182,N_4380);
xnor U4683 (N_4683,N_4285,N_4268);
nor U4684 (N_4684,N_4014,N_4236);
nor U4685 (N_4685,N_4482,N_4103);
or U4686 (N_4686,N_4034,N_4131);
and U4687 (N_4687,N_4343,N_4195);
nor U4688 (N_4688,N_4127,N_4334);
or U4689 (N_4689,N_4388,N_4403);
or U4690 (N_4690,N_4251,N_4470);
nand U4691 (N_4691,N_4466,N_4183);
nor U4692 (N_4692,N_4017,N_4043);
and U4693 (N_4693,N_4314,N_4358);
and U4694 (N_4694,N_4418,N_4080);
xor U4695 (N_4695,N_4336,N_4340);
nand U4696 (N_4696,N_4322,N_4337);
and U4697 (N_4697,N_4121,N_4487);
nor U4698 (N_4698,N_4152,N_4480);
nor U4699 (N_4699,N_4447,N_4312);
nor U4700 (N_4700,N_4465,N_4392);
and U4701 (N_4701,N_4409,N_4305);
nand U4702 (N_4702,N_4354,N_4216);
or U4703 (N_4703,N_4357,N_4213);
and U4704 (N_4704,N_4200,N_4438);
nor U4705 (N_4705,N_4149,N_4257);
and U4706 (N_4706,N_4469,N_4385);
nor U4707 (N_4707,N_4045,N_4290);
and U4708 (N_4708,N_4031,N_4047);
and U4709 (N_4709,N_4247,N_4302);
nor U4710 (N_4710,N_4253,N_4326);
xnor U4711 (N_4711,N_4160,N_4015);
xor U4712 (N_4712,N_4475,N_4158);
or U4713 (N_4713,N_4444,N_4426);
and U4714 (N_4714,N_4479,N_4217);
and U4715 (N_4715,N_4193,N_4260);
and U4716 (N_4716,N_4459,N_4165);
and U4717 (N_4717,N_4191,N_4378);
nor U4718 (N_4718,N_4397,N_4190);
and U4719 (N_4719,N_4367,N_4214);
xor U4720 (N_4720,N_4394,N_4061);
nor U4721 (N_4721,N_4496,N_4013);
xor U4722 (N_4722,N_4006,N_4128);
nand U4723 (N_4723,N_4297,N_4456);
and U4724 (N_4724,N_4450,N_4306);
xor U4725 (N_4725,N_4393,N_4417);
or U4726 (N_4726,N_4210,N_4008);
nor U4727 (N_4727,N_4134,N_4244);
nor U4728 (N_4728,N_4007,N_4144);
or U4729 (N_4729,N_4167,N_4407);
and U4730 (N_4730,N_4460,N_4207);
or U4731 (N_4731,N_4157,N_4386);
xnor U4732 (N_4732,N_4132,N_4335);
and U4733 (N_4733,N_4120,N_4176);
nor U4734 (N_4734,N_4353,N_4368);
nand U4735 (N_4735,N_4000,N_4235);
xnor U4736 (N_4736,N_4219,N_4490);
nor U4737 (N_4737,N_4175,N_4241);
and U4738 (N_4738,N_4338,N_4094);
nand U4739 (N_4739,N_4076,N_4181);
xor U4740 (N_4740,N_4226,N_4078);
xnor U4741 (N_4741,N_4048,N_4211);
xnor U4742 (N_4742,N_4124,N_4328);
and U4743 (N_4743,N_4309,N_4138);
nand U4744 (N_4744,N_4483,N_4319);
and U4745 (N_4745,N_4372,N_4108);
nand U4746 (N_4746,N_4420,N_4316);
and U4747 (N_4747,N_4457,N_4402);
and U4748 (N_4748,N_4073,N_4430);
nand U4749 (N_4749,N_4281,N_4304);
nand U4750 (N_4750,N_4159,N_4280);
nor U4751 (N_4751,N_4301,N_4225);
nor U4752 (N_4752,N_4241,N_4481);
or U4753 (N_4753,N_4061,N_4014);
and U4754 (N_4754,N_4498,N_4074);
or U4755 (N_4755,N_4381,N_4116);
and U4756 (N_4756,N_4297,N_4061);
or U4757 (N_4757,N_4097,N_4441);
nand U4758 (N_4758,N_4263,N_4458);
nor U4759 (N_4759,N_4362,N_4304);
or U4760 (N_4760,N_4356,N_4084);
nor U4761 (N_4761,N_4116,N_4450);
xnor U4762 (N_4762,N_4044,N_4458);
nor U4763 (N_4763,N_4058,N_4263);
nand U4764 (N_4764,N_4326,N_4413);
xor U4765 (N_4765,N_4026,N_4071);
nor U4766 (N_4766,N_4472,N_4441);
or U4767 (N_4767,N_4052,N_4083);
xnor U4768 (N_4768,N_4049,N_4346);
or U4769 (N_4769,N_4267,N_4244);
or U4770 (N_4770,N_4267,N_4417);
nand U4771 (N_4771,N_4098,N_4278);
and U4772 (N_4772,N_4204,N_4453);
xnor U4773 (N_4773,N_4105,N_4200);
or U4774 (N_4774,N_4435,N_4022);
nand U4775 (N_4775,N_4381,N_4076);
and U4776 (N_4776,N_4201,N_4232);
nand U4777 (N_4777,N_4236,N_4351);
nor U4778 (N_4778,N_4135,N_4320);
nor U4779 (N_4779,N_4224,N_4430);
or U4780 (N_4780,N_4032,N_4146);
xor U4781 (N_4781,N_4456,N_4271);
or U4782 (N_4782,N_4326,N_4435);
and U4783 (N_4783,N_4418,N_4336);
nor U4784 (N_4784,N_4166,N_4047);
nand U4785 (N_4785,N_4139,N_4020);
xnor U4786 (N_4786,N_4463,N_4298);
or U4787 (N_4787,N_4457,N_4044);
nor U4788 (N_4788,N_4257,N_4148);
xor U4789 (N_4789,N_4461,N_4152);
nand U4790 (N_4790,N_4167,N_4065);
nand U4791 (N_4791,N_4061,N_4155);
and U4792 (N_4792,N_4487,N_4065);
nor U4793 (N_4793,N_4082,N_4278);
and U4794 (N_4794,N_4067,N_4483);
and U4795 (N_4795,N_4355,N_4115);
or U4796 (N_4796,N_4064,N_4366);
and U4797 (N_4797,N_4297,N_4358);
xor U4798 (N_4798,N_4327,N_4495);
nand U4799 (N_4799,N_4187,N_4351);
nand U4800 (N_4800,N_4365,N_4422);
or U4801 (N_4801,N_4125,N_4247);
nand U4802 (N_4802,N_4163,N_4425);
xor U4803 (N_4803,N_4324,N_4185);
nand U4804 (N_4804,N_4355,N_4305);
and U4805 (N_4805,N_4383,N_4007);
or U4806 (N_4806,N_4113,N_4098);
and U4807 (N_4807,N_4105,N_4001);
xor U4808 (N_4808,N_4044,N_4357);
nand U4809 (N_4809,N_4069,N_4447);
nand U4810 (N_4810,N_4001,N_4201);
nand U4811 (N_4811,N_4407,N_4347);
xor U4812 (N_4812,N_4362,N_4059);
nand U4813 (N_4813,N_4354,N_4027);
nand U4814 (N_4814,N_4302,N_4469);
or U4815 (N_4815,N_4038,N_4426);
nor U4816 (N_4816,N_4073,N_4359);
xnor U4817 (N_4817,N_4437,N_4186);
xor U4818 (N_4818,N_4414,N_4277);
xor U4819 (N_4819,N_4139,N_4119);
xnor U4820 (N_4820,N_4499,N_4226);
nor U4821 (N_4821,N_4470,N_4482);
or U4822 (N_4822,N_4010,N_4098);
and U4823 (N_4823,N_4195,N_4015);
and U4824 (N_4824,N_4429,N_4120);
and U4825 (N_4825,N_4096,N_4356);
xnor U4826 (N_4826,N_4150,N_4405);
or U4827 (N_4827,N_4407,N_4361);
and U4828 (N_4828,N_4372,N_4367);
and U4829 (N_4829,N_4205,N_4335);
nor U4830 (N_4830,N_4152,N_4044);
xor U4831 (N_4831,N_4389,N_4118);
nand U4832 (N_4832,N_4330,N_4435);
and U4833 (N_4833,N_4405,N_4201);
nor U4834 (N_4834,N_4007,N_4358);
nand U4835 (N_4835,N_4351,N_4313);
or U4836 (N_4836,N_4299,N_4321);
and U4837 (N_4837,N_4296,N_4223);
xnor U4838 (N_4838,N_4460,N_4068);
nand U4839 (N_4839,N_4041,N_4225);
nor U4840 (N_4840,N_4263,N_4403);
nor U4841 (N_4841,N_4414,N_4386);
xor U4842 (N_4842,N_4198,N_4458);
nand U4843 (N_4843,N_4183,N_4275);
xnor U4844 (N_4844,N_4481,N_4228);
and U4845 (N_4845,N_4392,N_4277);
xor U4846 (N_4846,N_4494,N_4161);
nor U4847 (N_4847,N_4476,N_4076);
or U4848 (N_4848,N_4046,N_4341);
xor U4849 (N_4849,N_4114,N_4349);
and U4850 (N_4850,N_4483,N_4078);
nor U4851 (N_4851,N_4151,N_4445);
nor U4852 (N_4852,N_4207,N_4011);
nor U4853 (N_4853,N_4095,N_4141);
or U4854 (N_4854,N_4458,N_4290);
nand U4855 (N_4855,N_4260,N_4000);
or U4856 (N_4856,N_4261,N_4110);
nand U4857 (N_4857,N_4354,N_4098);
and U4858 (N_4858,N_4023,N_4096);
and U4859 (N_4859,N_4043,N_4395);
nor U4860 (N_4860,N_4034,N_4283);
nor U4861 (N_4861,N_4492,N_4297);
or U4862 (N_4862,N_4479,N_4116);
xnor U4863 (N_4863,N_4321,N_4399);
xor U4864 (N_4864,N_4003,N_4298);
nor U4865 (N_4865,N_4354,N_4453);
or U4866 (N_4866,N_4199,N_4474);
and U4867 (N_4867,N_4322,N_4015);
xnor U4868 (N_4868,N_4379,N_4136);
xor U4869 (N_4869,N_4014,N_4464);
or U4870 (N_4870,N_4294,N_4379);
and U4871 (N_4871,N_4108,N_4050);
and U4872 (N_4872,N_4356,N_4292);
nand U4873 (N_4873,N_4022,N_4027);
or U4874 (N_4874,N_4375,N_4003);
or U4875 (N_4875,N_4248,N_4339);
and U4876 (N_4876,N_4079,N_4317);
and U4877 (N_4877,N_4085,N_4465);
or U4878 (N_4878,N_4196,N_4261);
and U4879 (N_4879,N_4195,N_4421);
or U4880 (N_4880,N_4228,N_4017);
and U4881 (N_4881,N_4364,N_4241);
and U4882 (N_4882,N_4196,N_4182);
nor U4883 (N_4883,N_4022,N_4033);
xor U4884 (N_4884,N_4310,N_4289);
nor U4885 (N_4885,N_4384,N_4387);
and U4886 (N_4886,N_4266,N_4458);
nor U4887 (N_4887,N_4075,N_4354);
or U4888 (N_4888,N_4074,N_4215);
or U4889 (N_4889,N_4138,N_4110);
xnor U4890 (N_4890,N_4204,N_4247);
and U4891 (N_4891,N_4373,N_4023);
xnor U4892 (N_4892,N_4044,N_4226);
and U4893 (N_4893,N_4069,N_4044);
and U4894 (N_4894,N_4106,N_4287);
or U4895 (N_4895,N_4320,N_4109);
and U4896 (N_4896,N_4430,N_4160);
or U4897 (N_4897,N_4158,N_4387);
or U4898 (N_4898,N_4218,N_4323);
and U4899 (N_4899,N_4369,N_4116);
and U4900 (N_4900,N_4396,N_4197);
and U4901 (N_4901,N_4074,N_4384);
nand U4902 (N_4902,N_4295,N_4118);
and U4903 (N_4903,N_4455,N_4385);
nand U4904 (N_4904,N_4499,N_4326);
nand U4905 (N_4905,N_4378,N_4401);
or U4906 (N_4906,N_4155,N_4146);
or U4907 (N_4907,N_4311,N_4483);
or U4908 (N_4908,N_4140,N_4098);
xor U4909 (N_4909,N_4292,N_4499);
and U4910 (N_4910,N_4313,N_4025);
nand U4911 (N_4911,N_4464,N_4183);
nor U4912 (N_4912,N_4431,N_4343);
xnor U4913 (N_4913,N_4141,N_4114);
nand U4914 (N_4914,N_4061,N_4424);
xnor U4915 (N_4915,N_4438,N_4318);
or U4916 (N_4916,N_4459,N_4315);
or U4917 (N_4917,N_4176,N_4260);
or U4918 (N_4918,N_4410,N_4233);
or U4919 (N_4919,N_4371,N_4255);
nor U4920 (N_4920,N_4191,N_4190);
and U4921 (N_4921,N_4354,N_4466);
nand U4922 (N_4922,N_4433,N_4061);
or U4923 (N_4923,N_4458,N_4406);
nor U4924 (N_4924,N_4108,N_4325);
nand U4925 (N_4925,N_4322,N_4467);
nand U4926 (N_4926,N_4045,N_4429);
nor U4927 (N_4927,N_4453,N_4240);
nor U4928 (N_4928,N_4028,N_4185);
xor U4929 (N_4929,N_4247,N_4382);
nand U4930 (N_4930,N_4161,N_4284);
xnor U4931 (N_4931,N_4314,N_4113);
xnor U4932 (N_4932,N_4129,N_4051);
nand U4933 (N_4933,N_4227,N_4348);
and U4934 (N_4934,N_4019,N_4131);
nand U4935 (N_4935,N_4222,N_4340);
xor U4936 (N_4936,N_4342,N_4241);
and U4937 (N_4937,N_4195,N_4030);
or U4938 (N_4938,N_4042,N_4346);
nor U4939 (N_4939,N_4464,N_4448);
xnor U4940 (N_4940,N_4065,N_4257);
or U4941 (N_4941,N_4062,N_4474);
nand U4942 (N_4942,N_4248,N_4457);
nand U4943 (N_4943,N_4043,N_4214);
or U4944 (N_4944,N_4051,N_4411);
or U4945 (N_4945,N_4367,N_4061);
xnor U4946 (N_4946,N_4027,N_4435);
and U4947 (N_4947,N_4032,N_4319);
and U4948 (N_4948,N_4489,N_4229);
nand U4949 (N_4949,N_4104,N_4240);
and U4950 (N_4950,N_4000,N_4343);
or U4951 (N_4951,N_4394,N_4434);
nor U4952 (N_4952,N_4281,N_4301);
nand U4953 (N_4953,N_4153,N_4452);
nor U4954 (N_4954,N_4446,N_4325);
or U4955 (N_4955,N_4063,N_4469);
and U4956 (N_4956,N_4350,N_4298);
or U4957 (N_4957,N_4398,N_4467);
nor U4958 (N_4958,N_4331,N_4031);
and U4959 (N_4959,N_4494,N_4026);
or U4960 (N_4960,N_4137,N_4149);
or U4961 (N_4961,N_4286,N_4245);
xnor U4962 (N_4962,N_4002,N_4172);
or U4963 (N_4963,N_4207,N_4231);
xnor U4964 (N_4964,N_4212,N_4456);
and U4965 (N_4965,N_4125,N_4210);
nor U4966 (N_4966,N_4480,N_4034);
nand U4967 (N_4967,N_4295,N_4190);
or U4968 (N_4968,N_4071,N_4265);
and U4969 (N_4969,N_4238,N_4080);
xor U4970 (N_4970,N_4458,N_4211);
nor U4971 (N_4971,N_4278,N_4348);
and U4972 (N_4972,N_4303,N_4168);
nand U4973 (N_4973,N_4149,N_4007);
or U4974 (N_4974,N_4130,N_4334);
nor U4975 (N_4975,N_4414,N_4377);
or U4976 (N_4976,N_4038,N_4454);
nand U4977 (N_4977,N_4249,N_4390);
nand U4978 (N_4978,N_4025,N_4261);
or U4979 (N_4979,N_4308,N_4155);
nand U4980 (N_4980,N_4477,N_4040);
or U4981 (N_4981,N_4223,N_4133);
or U4982 (N_4982,N_4372,N_4420);
and U4983 (N_4983,N_4423,N_4220);
nor U4984 (N_4984,N_4007,N_4018);
nand U4985 (N_4985,N_4284,N_4208);
or U4986 (N_4986,N_4397,N_4131);
xor U4987 (N_4987,N_4122,N_4392);
xnor U4988 (N_4988,N_4467,N_4377);
nand U4989 (N_4989,N_4324,N_4437);
and U4990 (N_4990,N_4009,N_4351);
nand U4991 (N_4991,N_4499,N_4420);
xor U4992 (N_4992,N_4396,N_4262);
and U4993 (N_4993,N_4347,N_4467);
xor U4994 (N_4994,N_4230,N_4203);
xor U4995 (N_4995,N_4226,N_4393);
nor U4996 (N_4996,N_4158,N_4030);
or U4997 (N_4997,N_4031,N_4225);
nor U4998 (N_4998,N_4421,N_4329);
xor U4999 (N_4999,N_4134,N_4162);
and U5000 (N_5000,N_4532,N_4744);
nand U5001 (N_5001,N_4993,N_4746);
xor U5002 (N_5002,N_4907,N_4726);
and U5003 (N_5003,N_4972,N_4650);
xnor U5004 (N_5004,N_4736,N_4863);
nand U5005 (N_5005,N_4600,N_4692);
nand U5006 (N_5006,N_4775,N_4823);
or U5007 (N_5007,N_4740,N_4541);
xnor U5008 (N_5008,N_4612,N_4534);
xnor U5009 (N_5009,N_4565,N_4614);
and U5010 (N_5010,N_4618,N_4872);
xor U5011 (N_5011,N_4952,N_4771);
and U5012 (N_5012,N_4531,N_4737);
xnor U5013 (N_5013,N_4877,N_4825);
nor U5014 (N_5014,N_4566,N_4797);
or U5015 (N_5015,N_4851,N_4954);
xor U5016 (N_5016,N_4686,N_4873);
nor U5017 (N_5017,N_4820,N_4828);
nor U5018 (N_5018,N_4789,N_4561);
or U5019 (N_5019,N_4968,N_4783);
xnor U5020 (N_5020,N_4764,N_4850);
xnor U5021 (N_5021,N_4538,N_4948);
nor U5022 (N_5022,N_4504,N_4845);
xor U5023 (N_5023,N_4846,N_4832);
or U5024 (N_5024,N_4928,N_4556);
xnor U5025 (N_5025,N_4507,N_4675);
xnor U5026 (N_5026,N_4676,N_4944);
nand U5027 (N_5027,N_4610,N_4943);
xor U5028 (N_5028,N_4754,N_4909);
xor U5029 (N_5029,N_4712,N_4557);
and U5030 (N_5030,N_4788,N_4896);
or U5031 (N_5031,N_4906,N_4970);
or U5032 (N_5032,N_4628,N_4812);
or U5033 (N_5033,N_4790,N_4839);
nand U5034 (N_5034,N_4515,N_4503);
nor U5035 (N_5035,N_4843,N_4743);
xnor U5036 (N_5036,N_4625,N_4999);
nand U5037 (N_5037,N_4732,N_4886);
xor U5038 (N_5038,N_4632,N_4997);
nor U5039 (N_5039,N_4959,N_4669);
nor U5040 (N_5040,N_4947,N_4802);
nand U5041 (N_5041,N_4753,N_4777);
xnor U5042 (N_5042,N_4933,N_4693);
nor U5043 (N_5043,N_4995,N_4941);
xor U5044 (N_5044,N_4567,N_4587);
or U5045 (N_5045,N_4553,N_4808);
and U5046 (N_5046,N_4640,N_4853);
nor U5047 (N_5047,N_4898,N_4711);
or U5048 (N_5048,N_4539,N_4511);
and U5049 (N_5049,N_4800,N_4509);
or U5050 (N_5050,N_4582,N_4656);
nor U5051 (N_5051,N_4537,N_4918);
nand U5052 (N_5052,N_4831,N_4763);
nor U5053 (N_5053,N_4857,N_4938);
or U5054 (N_5054,N_4706,N_4755);
xnor U5055 (N_5055,N_4624,N_4888);
or U5056 (N_5056,N_4665,N_4864);
nor U5057 (N_5057,N_4689,N_4822);
or U5058 (N_5058,N_4894,N_4757);
xnor U5059 (N_5059,N_4935,N_4786);
nor U5060 (N_5060,N_4987,N_4801);
or U5061 (N_5061,N_4583,N_4639);
and U5062 (N_5062,N_4733,N_4805);
nand U5063 (N_5063,N_4663,N_4964);
and U5064 (N_5064,N_4714,N_4929);
and U5065 (N_5065,N_4871,N_4700);
xnor U5066 (N_5066,N_4593,N_4579);
or U5067 (N_5067,N_4885,N_4932);
nand U5068 (N_5068,N_4721,N_4591);
nand U5069 (N_5069,N_4976,N_4841);
and U5070 (N_5070,N_4983,N_4694);
nand U5071 (N_5071,N_4814,N_4984);
or U5072 (N_5072,N_4701,N_4629);
nand U5073 (N_5073,N_4770,N_4602);
and U5074 (N_5074,N_4926,N_4868);
or U5075 (N_5075,N_4697,N_4974);
or U5076 (N_5076,N_4978,N_4601);
or U5077 (N_5077,N_4953,N_4578);
nand U5078 (N_5078,N_4728,N_4646);
or U5079 (N_5079,N_4560,N_4980);
nor U5080 (N_5080,N_4680,N_4750);
and U5081 (N_5081,N_4641,N_4513);
or U5082 (N_5082,N_4804,N_4965);
nor U5083 (N_5083,N_4768,N_4549);
nor U5084 (N_5084,N_4588,N_4621);
xnor U5085 (N_5085,N_4793,N_4779);
nand U5086 (N_5086,N_4862,N_4861);
or U5087 (N_5087,N_4875,N_4869);
xor U5088 (N_5088,N_4573,N_4631);
xnor U5089 (N_5089,N_4668,N_4923);
nand U5090 (N_5090,N_4530,N_4544);
xor U5091 (N_5091,N_4759,N_4774);
nor U5092 (N_5092,N_4838,N_4604);
nor U5093 (N_5093,N_4930,N_4795);
or U5094 (N_5094,N_4596,N_4727);
or U5095 (N_5095,N_4854,N_4682);
and U5096 (N_5096,N_4595,N_4899);
or U5097 (N_5097,N_4807,N_4897);
xnor U5098 (N_5098,N_4992,N_4985);
or U5099 (N_5099,N_4571,N_4844);
nand U5100 (N_5100,N_4829,N_4905);
nor U5101 (N_5101,N_4558,N_4772);
nor U5102 (N_5102,N_4562,N_4773);
and U5103 (N_5103,N_4921,N_4840);
nand U5104 (N_5104,N_4834,N_4816);
nor U5105 (N_5105,N_4528,N_4842);
nor U5106 (N_5106,N_4900,N_4989);
nor U5107 (N_5107,N_4506,N_4688);
xnor U5108 (N_5108,N_4599,N_4502);
nand U5109 (N_5109,N_4551,N_4908);
nor U5110 (N_5110,N_4778,N_4501);
nor U5111 (N_5111,N_4780,N_4613);
xnor U5112 (N_5112,N_4542,N_4644);
or U5113 (N_5113,N_4514,N_4769);
and U5114 (N_5114,N_4852,N_4643);
nor U5115 (N_5115,N_4880,N_4517);
nand U5116 (N_5116,N_4914,N_4705);
nor U5117 (N_5117,N_4710,N_4633);
nor U5118 (N_5118,N_4891,N_4991);
nand U5119 (N_5119,N_4796,N_4611);
and U5120 (N_5120,N_4917,N_4603);
and U5121 (N_5121,N_4522,N_4903);
or U5122 (N_5122,N_4520,N_4654);
nor U5123 (N_5123,N_4742,N_4901);
xnor U5124 (N_5124,N_4961,N_4671);
xor U5125 (N_5125,N_4887,N_4708);
nand U5126 (N_5126,N_4568,N_4655);
xor U5127 (N_5127,N_4510,N_4855);
nand U5128 (N_5128,N_4882,N_4735);
and U5129 (N_5129,N_4902,N_4904);
and U5130 (N_5130,N_4787,N_4837);
xor U5131 (N_5131,N_4749,N_4791);
and U5132 (N_5132,N_4616,N_4766);
nand U5133 (N_5133,N_4859,N_4696);
or U5134 (N_5134,N_4518,N_4924);
nand U5135 (N_5135,N_4519,N_4758);
and U5136 (N_5136,N_4821,N_4684);
or U5137 (N_5137,N_4653,N_4934);
xnor U5138 (N_5138,N_4533,N_4971);
and U5139 (N_5139,N_4713,N_4678);
xnor U5140 (N_5140,N_4605,N_4945);
nor U5141 (N_5141,N_4927,N_4949);
nand U5142 (N_5142,N_4942,N_4833);
or U5143 (N_5143,N_4826,N_4883);
or U5144 (N_5144,N_4637,N_4725);
xnor U5145 (N_5145,N_4648,N_4659);
and U5146 (N_5146,N_4792,N_4670);
xor U5147 (N_5147,N_4627,N_4642);
nand U5148 (N_5148,N_4581,N_4724);
nor U5149 (N_5149,N_4940,N_4765);
and U5150 (N_5150,N_4647,N_4516);
xnor U5151 (N_5151,N_4580,N_4535);
and U5152 (N_5152,N_4752,N_4973);
xor U5153 (N_5153,N_4683,N_4982);
nand U5154 (N_5154,N_4572,N_4794);
and U5155 (N_5155,N_4975,N_4806);
nor U5156 (N_5156,N_4652,N_4738);
xor U5157 (N_5157,N_4681,N_4785);
and U5158 (N_5158,N_4608,N_4525);
or U5159 (N_5159,N_4748,N_4527);
and U5160 (N_5160,N_4811,N_4607);
and U5161 (N_5161,N_4956,N_4847);
xnor U5162 (N_5162,N_4919,N_4979);
nor U5163 (N_5163,N_4889,N_4815);
and U5164 (N_5164,N_4672,N_4895);
nor U5165 (N_5165,N_4619,N_4922);
xnor U5166 (N_5166,N_4597,N_4951);
xnor U5167 (N_5167,N_4645,N_4634);
nor U5168 (N_5168,N_4704,N_4819);
and U5169 (N_5169,N_4575,N_4879);
or U5170 (N_5170,N_4760,N_4723);
or U5171 (N_5171,N_4555,N_4691);
nand U5172 (N_5172,N_4667,N_4529);
or U5173 (N_5173,N_4782,N_4761);
and U5174 (N_5174,N_4911,N_4835);
or U5175 (N_5175,N_4803,N_4626);
or U5176 (N_5176,N_4698,N_4589);
xnor U5177 (N_5177,N_4849,N_4685);
nor U5178 (N_5178,N_4776,N_4666);
and U5179 (N_5179,N_4699,N_4981);
xor U5180 (N_5180,N_4827,N_4677);
nand U5181 (N_5181,N_4717,N_4623);
nor U5182 (N_5182,N_4598,N_4617);
nand U5183 (N_5183,N_4878,N_4876);
nand U5184 (N_5184,N_4563,N_4865);
or U5185 (N_5185,N_4939,N_4848);
nand U5186 (N_5186,N_4756,N_4931);
and U5187 (N_5187,N_4962,N_4925);
and U5188 (N_5188,N_4884,N_4998);
xor U5189 (N_5189,N_4813,N_4818);
nor U5190 (N_5190,N_4784,N_4798);
xnor U5191 (N_5191,N_4523,N_4867);
xnor U5192 (N_5192,N_4977,N_4936);
xor U5193 (N_5193,N_4649,N_4660);
nand U5194 (N_5194,N_4702,N_4540);
and U5195 (N_5195,N_4661,N_4767);
nand U5196 (N_5196,N_4963,N_4548);
xnor U5197 (N_5197,N_4635,N_4543);
nand U5198 (N_5198,N_4590,N_4734);
and U5199 (N_5199,N_4521,N_4662);
nor U5200 (N_5200,N_4550,N_4615);
or U5201 (N_5201,N_4609,N_4651);
or U5202 (N_5202,N_4703,N_4709);
and U5203 (N_5203,N_4547,N_4569);
nor U5204 (N_5204,N_4584,N_4592);
nand U5205 (N_5205,N_4564,N_4690);
and U5206 (N_5206,N_4870,N_4524);
or U5207 (N_5207,N_4966,N_4718);
or U5208 (N_5208,N_4799,N_4817);
and U5209 (N_5209,N_4687,N_4574);
and U5210 (N_5210,N_4585,N_4741);
xor U5211 (N_5211,N_4950,N_4673);
xor U5212 (N_5212,N_4570,N_4781);
nand U5213 (N_5213,N_4967,N_4722);
nor U5214 (N_5214,N_4960,N_4500);
nor U5215 (N_5215,N_4664,N_4715);
nand U5216 (N_5216,N_4638,N_4657);
nand U5217 (N_5217,N_4536,N_4739);
nand U5218 (N_5218,N_4874,N_4505);
nand U5219 (N_5219,N_4915,N_4719);
and U5220 (N_5220,N_4594,N_4679);
xnor U5221 (N_5221,N_4747,N_4892);
nor U5222 (N_5222,N_4916,N_4858);
or U5223 (N_5223,N_4912,N_4695);
xnor U5224 (N_5224,N_4762,N_4920);
nand U5225 (N_5225,N_4658,N_4881);
nor U5226 (N_5226,N_4910,N_4824);
nor U5227 (N_5227,N_4957,N_4830);
nor U5228 (N_5228,N_4577,N_4707);
or U5229 (N_5229,N_4512,N_4893);
xnor U5230 (N_5230,N_4674,N_4586);
and U5231 (N_5231,N_4620,N_4836);
and U5232 (N_5232,N_4994,N_4545);
nand U5233 (N_5233,N_4729,N_4526);
nand U5234 (N_5234,N_4554,N_4810);
nand U5235 (N_5235,N_4606,N_4630);
xnor U5236 (N_5236,N_4946,N_4860);
xnor U5237 (N_5237,N_4730,N_4955);
or U5238 (N_5238,N_4751,N_4716);
xnor U5239 (N_5239,N_4636,N_4988);
nor U5240 (N_5240,N_4559,N_4731);
and U5241 (N_5241,N_4622,N_4937);
or U5242 (N_5242,N_4890,N_4856);
and U5243 (N_5243,N_4809,N_4969);
nor U5244 (N_5244,N_4745,N_4866);
or U5245 (N_5245,N_4986,N_4913);
nand U5246 (N_5246,N_4508,N_4576);
nor U5247 (N_5247,N_4990,N_4552);
or U5248 (N_5248,N_4720,N_4958);
nor U5249 (N_5249,N_4996,N_4546);
xnor U5250 (N_5250,N_4977,N_4640);
and U5251 (N_5251,N_4581,N_4772);
nor U5252 (N_5252,N_4968,N_4510);
nand U5253 (N_5253,N_4747,N_4745);
xor U5254 (N_5254,N_4581,N_4661);
nor U5255 (N_5255,N_4656,N_4681);
or U5256 (N_5256,N_4861,N_4584);
xnor U5257 (N_5257,N_4717,N_4613);
nand U5258 (N_5258,N_4561,N_4681);
nor U5259 (N_5259,N_4672,N_4734);
nand U5260 (N_5260,N_4708,N_4528);
nor U5261 (N_5261,N_4991,N_4545);
xnor U5262 (N_5262,N_4689,N_4540);
nor U5263 (N_5263,N_4924,N_4556);
xor U5264 (N_5264,N_4668,N_4595);
or U5265 (N_5265,N_4513,N_4819);
nor U5266 (N_5266,N_4763,N_4609);
and U5267 (N_5267,N_4924,N_4678);
and U5268 (N_5268,N_4589,N_4826);
and U5269 (N_5269,N_4549,N_4795);
nand U5270 (N_5270,N_4738,N_4681);
and U5271 (N_5271,N_4708,N_4604);
and U5272 (N_5272,N_4672,N_4642);
nor U5273 (N_5273,N_4747,N_4674);
and U5274 (N_5274,N_4711,N_4678);
nor U5275 (N_5275,N_4927,N_4502);
nor U5276 (N_5276,N_4787,N_4651);
or U5277 (N_5277,N_4817,N_4507);
nor U5278 (N_5278,N_4857,N_4722);
nand U5279 (N_5279,N_4777,N_4937);
nor U5280 (N_5280,N_4717,N_4737);
or U5281 (N_5281,N_4701,N_4900);
and U5282 (N_5282,N_4660,N_4874);
and U5283 (N_5283,N_4662,N_4678);
or U5284 (N_5284,N_4620,N_4706);
and U5285 (N_5285,N_4900,N_4916);
xnor U5286 (N_5286,N_4583,N_4753);
nor U5287 (N_5287,N_4848,N_4863);
and U5288 (N_5288,N_4814,N_4722);
and U5289 (N_5289,N_4668,N_4985);
and U5290 (N_5290,N_4563,N_4949);
nand U5291 (N_5291,N_4875,N_4833);
or U5292 (N_5292,N_4557,N_4927);
nand U5293 (N_5293,N_4741,N_4924);
or U5294 (N_5294,N_4790,N_4979);
and U5295 (N_5295,N_4814,N_4832);
nor U5296 (N_5296,N_4588,N_4907);
nor U5297 (N_5297,N_4793,N_4588);
nor U5298 (N_5298,N_4596,N_4531);
nor U5299 (N_5299,N_4702,N_4550);
nand U5300 (N_5300,N_4928,N_4995);
nor U5301 (N_5301,N_4943,N_4969);
and U5302 (N_5302,N_4706,N_4851);
or U5303 (N_5303,N_4996,N_4685);
or U5304 (N_5304,N_4824,N_4674);
nand U5305 (N_5305,N_4884,N_4573);
and U5306 (N_5306,N_4913,N_4861);
and U5307 (N_5307,N_4757,N_4658);
and U5308 (N_5308,N_4904,N_4887);
or U5309 (N_5309,N_4588,N_4669);
and U5310 (N_5310,N_4673,N_4695);
nor U5311 (N_5311,N_4755,N_4506);
or U5312 (N_5312,N_4847,N_4964);
nand U5313 (N_5313,N_4807,N_4633);
nor U5314 (N_5314,N_4659,N_4816);
and U5315 (N_5315,N_4822,N_4740);
nand U5316 (N_5316,N_4815,N_4710);
and U5317 (N_5317,N_4521,N_4635);
xor U5318 (N_5318,N_4870,N_4703);
nor U5319 (N_5319,N_4821,N_4780);
nand U5320 (N_5320,N_4802,N_4940);
or U5321 (N_5321,N_4524,N_4612);
or U5322 (N_5322,N_4558,N_4566);
nand U5323 (N_5323,N_4761,N_4762);
nand U5324 (N_5324,N_4603,N_4867);
and U5325 (N_5325,N_4795,N_4852);
or U5326 (N_5326,N_4732,N_4512);
or U5327 (N_5327,N_4535,N_4837);
xor U5328 (N_5328,N_4914,N_4980);
or U5329 (N_5329,N_4761,N_4962);
xor U5330 (N_5330,N_4762,N_4740);
or U5331 (N_5331,N_4958,N_4707);
xnor U5332 (N_5332,N_4867,N_4589);
xor U5333 (N_5333,N_4575,N_4872);
or U5334 (N_5334,N_4759,N_4640);
and U5335 (N_5335,N_4998,N_4563);
or U5336 (N_5336,N_4618,N_4652);
nand U5337 (N_5337,N_4712,N_4881);
and U5338 (N_5338,N_4683,N_4992);
xnor U5339 (N_5339,N_4812,N_4538);
or U5340 (N_5340,N_4790,N_4966);
nor U5341 (N_5341,N_4910,N_4563);
xnor U5342 (N_5342,N_4528,N_4652);
nand U5343 (N_5343,N_4589,N_4998);
nand U5344 (N_5344,N_4975,N_4677);
xnor U5345 (N_5345,N_4958,N_4886);
nor U5346 (N_5346,N_4606,N_4847);
or U5347 (N_5347,N_4572,N_4903);
nor U5348 (N_5348,N_4599,N_4973);
nand U5349 (N_5349,N_4790,N_4572);
and U5350 (N_5350,N_4722,N_4773);
or U5351 (N_5351,N_4836,N_4932);
nand U5352 (N_5352,N_4706,N_4651);
nor U5353 (N_5353,N_4773,N_4973);
xnor U5354 (N_5354,N_4672,N_4984);
nor U5355 (N_5355,N_4946,N_4826);
or U5356 (N_5356,N_4847,N_4677);
xnor U5357 (N_5357,N_4774,N_4755);
nor U5358 (N_5358,N_4778,N_4537);
or U5359 (N_5359,N_4857,N_4544);
nor U5360 (N_5360,N_4647,N_4845);
nor U5361 (N_5361,N_4705,N_4747);
nand U5362 (N_5362,N_4886,N_4635);
nand U5363 (N_5363,N_4668,N_4583);
nor U5364 (N_5364,N_4626,N_4511);
nand U5365 (N_5365,N_4908,N_4627);
or U5366 (N_5366,N_4818,N_4945);
or U5367 (N_5367,N_4760,N_4918);
nor U5368 (N_5368,N_4609,N_4848);
and U5369 (N_5369,N_4858,N_4657);
and U5370 (N_5370,N_4985,N_4511);
xor U5371 (N_5371,N_4773,N_4755);
nor U5372 (N_5372,N_4959,N_4554);
or U5373 (N_5373,N_4931,N_4684);
nand U5374 (N_5374,N_4640,N_4770);
xnor U5375 (N_5375,N_4764,N_4548);
xnor U5376 (N_5376,N_4973,N_4992);
nor U5377 (N_5377,N_4802,N_4913);
xnor U5378 (N_5378,N_4850,N_4822);
nand U5379 (N_5379,N_4743,N_4607);
nand U5380 (N_5380,N_4863,N_4841);
and U5381 (N_5381,N_4613,N_4690);
or U5382 (N_5382,N_4861,N_4511);
xor U5383 (N_5383,N_4704,N_4571);
xnor U5384 (N_5384,N_4712,N_4880);
or U5385 (N_5385,N_4934,N_4871);
xnor U5386 (N_5386,N_4792,N_4981);
and U5387 (N_5387,N_4539,N_4990);
nor U5388 (N_5388,N_4520,N_4580);
and U5389 (N_5389,N_4668,N_4673);
nor U5390 (N_5390,N_4884,N_4880);
xnor U5391 (N_5391,N_4996,N_4740);
and U5392 (N_5392,N_4755,N_4705);
or U5393 (N_5393,N_4838,N_4691);
nand U5394 (N_5394,N_4966,N_4780);
and U5395 (N_5395,N_4865,N_4999);
xnor U5396 (N_5396,N_4894,N_4819);
xnor U5397 (N_5397,N_4634,N_4560);
nor U5398 (N_5398,N_4910,N_4626);
nor U5399 (N_5399,N_4587,N_4559);
xnor U5400 (N_5400,N_4798,N_4856);
xor U5401 (N_5401,N_4564,N_4583);
nor U5402 (N_5402,N_4605,N_4930);
nand U5403 (N_5403,N_4864,N_4742);
xnor U5404 (N_5404,N_4872,N_4663);
nor U5405 (N_5405,N_4754,N_4801);
or U5406 (N_5406,N_4860,N_4606);
xor U5407 (N_5407,N_4612,N_4512);
or U5408 (N_5408,N_4817,N_4908);
and U5409 (N_5409,N_4894,N_4943);
or U5410 (N_5410,N_4975,N_4907);
or U5411 (N_5411,N_4968,N_4883);
nor U5412 (N_5412,N_4512,N_4998);
or U5413 (N_5413,N_4834,N_4569);
or U5414 (N_5414,N_4650,N_4945);
and U5415 (N_5415,N_4693,N_4710);
or U5416 (N_5416,N_4866,N_4627);
or U5417 (N_5417,N_4628,N_4782);
and U5418 (N_5418,N_4732,N_4849);
nor U5419 (N_5419,N_4663,N_4978);
xnor U5420 (N_5420,N_4823,N_4554);
nor U5421 (N_5421,N_4558,N_4669);
xnor U5422 (N_5422,N_4740,N_4631);
or U5423 (N_5423,N_4873,N_4905);
or U5424 (N_5424,N_4686,N_4956);
nor U5425 (N_5425,N_4586,N_4997);
xor U5426 (N_5426,N_4637,N_4818);
nor U5427 (N_5427,N_4957,N_4842);
nand U5428 (N_5428,N_4995,N_4902);
nor U5429 (N_5429,N_4908,N_4935);
and U5430 (N_5430,N_4944,N_4741);
nor U5431 (N_5431,N_4611,N_4835);
xnor U5432 (N_5432,N_4686,N_4634);
nor U5433 (N_5433,N_4754,N_4535);
and U5434 (N_5434,N_4997,N_4726);
nor U5435 (N_5435,N_4514,N_4980);
or U5436 (N_5436,N_4517,N_4668);
xor U5437 (N_5437,N_4507,N_4646);
xnor U5438 (N_5438,N_4689,N_4900);
nand U5439 (N_5439,N_4874,N_4651);
nor U5440 (N_5440,N_4778,N_4787);
or U5441 (N_5441,N_4547,N_4815);
or U5442 (N_5442,N_4749,N_4909);
or U5443 (N_5443,N_4761,N_4517);
nor U5444 (N_5444,N_4994,N_4960);
and U5445 (N_5445,N_4605,N_4990);
or U5446 (N_5446,N_4586,N_4718);
and U5447 (N_5447,N_4616,N_4946);
nor U5448 (N_5448,N_4780,N_4527);
nor U5449 (N_5449,N_4815,N_4741);
xnor U5450 (N_5450,N_4564,N_4608);
or U5451 (N_5451,N_4869,N_4890);
nand U5452 (N_5452,N_4773,N_4810);
and U5453 (N_5453,N_4711,N_4773);
nor U5454 (N_5454,N_4948,N_4851);
or U5455 (N_5455,N_4509,N_4888);
xor U5456 (N_5456,N_4690,N_4761);
and U5457 (N_5457,N_4715,N_4771);
and U5458 (N_5458,N_4701,N_4644);
xnor U5459 (N_5459,N_4889,N_4877);
or U5460 (N_5460,N_4981,N_4574);
and U5461 (N_5461,N_4845,N_4836);
nand U5462 (N_5462,N_4740,N_4928);
and U5463 (N_5463,N_4967,N_4587);
and U5464 (N_5464,N_4872,N_4580);
nor U5465 (N_5465,N_4622,N_4956);
nor U5466 (N_5466,N_4564,N_4716);
xnor U5467 (N_5467,N_4636,N_4688);
and U5468 (N_5468,N_4683,N_4657);
or U5469 (N_5469,N_4905,N_4824);
nor U5470 (N_5470,N_4744,N_4712);
and U5471 (N_5471,N_4882,N_4661);
and U5472 (N_5472,N_4733,N_4616);
nand U5473 (N_5473,N_4578,N_4634);
nor U5474 (N_5474,N_4791,N_4684);
xor U5475 (N_5475,N_4851,N_4511);
nand U5476 (N_5476,N_4610,N_4727);
nor U5477 (N_5477,N_4676,N_4673);
xnor U5478 (N_5478,N_4886,N_4950);
or U5479 (N_5479,N_4927,N_4644);
nor U5480 (N_5480,N_4819,N_4902);
nand U5481 (N_5481,N_4853,N_4694);
nand U5482 (N_5482,N_4976,N_4910);
and U5483 (N_5483,N_4589,N_4594);
nand U5484 (N_5484,N_4693,N_4879);
or U5485 (N_5485,N_4526,N_4549);
and U5486 (N_5486,N_4508,N_4960);
xnor U5487 (N_5487,N_4781,N_4617);
or U5488 (N_5488,N_4753,N_4715);
xnor U5489 (N_5489,N_4846,N_4947);
or U5490 (N_5490,N_4826,N_4634);
nor U5491 (N_5491,N_4718,N_4574);
and U5492 (N_5492,N_4654,N_4978);
nor U5493 (N_5493,N_4850,N_4718);
nand U5494 (N_5494,N_4900,N_4936);
or U5495 (N_5495,N_4658,N_4538);
nor U5496 (N_5496,N_4635,N_4848);
or U5497 (N_5497,N_4546,N_4823);
nor U5498 (N_5498,N_4772,N_4928);
xnor U5499 (N_5499,N_4812,N_4570);
and U5500 (N_5500,N_5258,N_5080);
xor U5501 (N_5501,N_5338,N_5234);
and U5502 (N_5502,N_5054,N_5144);
nor U5503 (N_5503,N_5344,N_5077);
and U5504 (N_5504,N_5262,N_5064);
xor U5505 (N_5505,N_5098,N_5298);
and U5506 (N_5506,N_5277,N_5390);
nand U5507 (N_5507,N_5255,N_5000);
and U5508 (N_5508,N_5470,N_5044);
or U5509 (N_5509,N_5206,N_5129);
and U5510 (N_5510,N_5100,N_5304);
nand U5511 (N_5511,N_5491,N_5463);
or U5512 (N_5512,N_5221,N_5349);
xor U5513 (N_5513,N_5251,N_5430);
and U5514 (N_5514,N_5253,N_5417);
or U5515 (N_5515,N_5185,N_5365);
and U5516 (N_5516,N_5090,N_5075);
nor U5517 (N_5517,N_5330,N_5172);
and U5518 (N_5518,N_5056,N_5293);
nor U5519 (N_5519,N_5362,N_5252);
xnor U5520 (N_5520,N_5379,N_5266);
xor U5521 (N_5521,N_5455,N_5243);
xor U5522 (N_5522,N_5345,N_5209);
xnor U5523 (N_5523,N_5245,N_5196);
nor U5524 (N_5524,N_5194,N_5211);
nand U5525 (N_5525,N_5024,N_5416);
nor U5526 (N_5526,N_5326,N_5040);
or U5527 (N_5527,N_5411,N_5178);
nor U5528 (N_5528,N_5469,N_5367);
or U5529 (N_5529,N_5110,N_5399);
or U5530 (N_5530,N_5495,N_5219);
xor U5531 (N_5531,N_5460,N_5393);
xor U5532 (N_5532,N_5214,N_5383);
nor U5533 (N_5533,N_5215,N_5055);
nand U5534 (N_5534,N_5318,N_5193);
nor U5535 (N_5535,N_5394,N_5320);
or U5536 (N_5536,N_5296,N_5352);
and U5537 (N_5537,N_5078,N_5012);
nand U5538 (N_5538,N_5138,N_5335);
and U5539 (N_5539,N_5357,N_5405);
nor U5540 (N_5540,N_5333,N_5380);
xor U5541 (N_5541,N_5042,N_5006);
or U5542 (N_5542,N_5364,N_5294);
nor U5543 (N_5543,N_5385,N_5179);
nor U5544 (N_5544,N_5081,N_5249);
xnor U5545 (N_5545,N_5324,N_5124);
or U5546 (N_5546,N_5112,N_5093);
xnor U5547 (N_5547,N_5143,N_5225);
or U5548 (N_5548,N_5133,N_5311);
xnor U5549 (N_5549,N_5322,N_5480);
or U5550 (N_5550,N_5408,N_5232);
xnor U5551 (N_5551,N_5014,N_5286);
nand U5552 (N_5552,N_5271,N_5037);
nor U5553 (N_5553,N_5210,N_5229);
xnor U5554 (N_5554,N_5290,N_5069);
nand U5555 (N_5555,N_5097,N_5487);
nor U5556 (N_5556,N_5459,N_5461);
or U5557 (N_5557,N_5072,N_5376);
xnor U5558 (N_5558,N_5045,N_5414);
or U5559 (N_5559,N_5388,N_5472);
nand U5560 (N_5560,N_5424,N_5287);
nand U5561 (N_5561,N_5354,N_5264);
nor U5562 (N_5562,N_5198,N_5273);
xor U5563 (N_5563,N_5351,N_5094);
and U5564 (N_5564,N_5403,N_5401);
nand U5565 (N_5565,N_5114,N_5451);
or U5566 (N_5566,N_5125,N_5233);
nor U5567 (N_5567,N_5076,N_5246);
nor U5568 (N_5568,N_5442,N_5306);
or U5569 (N_5569,N_5420,N_5065);
nor U5570 (N_5570,N_5453,N_5171);
and U5571 (N_5571,N_5268,N_5305);
or U5572 (N_5572,N_5189,N_5329);
nor U5573 (N_5573,N_5265,N_5492);
or U5574 (N_5574,N_5248,N_5190);
or U5575 (N_5575,N_5360,N_5025);
xnor U5576 (N_5576,N_5377,N_5140);
or U5577 (N_5577,N_5008,N_5468);
xnor U5578 (N_5578,N_5106,N_5422);
and U5579 (N_5579,N_5395,N_5205);
or U5580 (N_5580,N_5220,N_5496);
nand U5581 (N_5581,N_5195,N_5498);
xor U5582 (N_5582,N_5426,N_5485);
and U5583 (N_5583,N_5348,N_5481);
nand U5584 (N_5584,N_5434,N_5446);
or U5585 (N_5585,N_5458,N_5026);
xnor U5586 (N_5586,N_5123,N_5325);
or U5587 (N_5587,N_5062,N_5166);
xnor U5588 (N_5588,N_5115,N_5427);
or U5589 (N_5589,N_5309,N_5016);
and U5590 (N_5590,N_5315,N_5436);
nand U5591 (N_5591,N_5327,N_5439);
and U5592 (N_5592,N_5235,N_5337);
and U5593 (N_5593,N_5095,N_5445);
nand U5594 (N_5594,N_5060,N_5247);
xor U5595 (N_5595,N_5130,N_5373);
nand U5596 (N_5596,N_5378,N_5161);
nor U5597 (N_5597,N_5188,N_5389);
nor U5598 (N_5598,N_5339,N_5152);
xor U5599 (N_5599,N_5162,N_5228);
xor U5600 (N_5600,N_5341,N_5475);
xnor U5601 (N_5601,N_5462,N_5023);
or U5602 (N_5602,N_5218,N_5011);
or U5603 (N_5603,N_5250,N_5203);
nor U5604 (N_5604,N_5347,N_5031);
or U5605 (N_5605,N_5432,N_5361);
or U5606 (N_5606,N_5331,N_5200);
nand U5607 (N_5607,N_5402,N_5392);
nor U5608 (N_5608,N_5300,N_5053);
or U5609 (N_5609,N_5254,N_5438);
xnor U5610 (N_5610,N_5494,N_5127);
xor U5611 (N_5611,N_5034,N_5085);
or U5612 (N_5612,N_5413,N_5267);
xor U5613 (N_5613,N_5073,N_5175);
nor U5614 (N_5614,N_5021,N_5039);
nor U5615 (N_5615,N_5099,N_5036);
nor U5616 (N_5616,N_5299,N_5103);
nand U5617 (N_5617,N_5108,N_5168);
and U5618 (N_5618,N_5313,N_5227);
nor U5619 (N_5619,N_5412,N_5375);
nor U5620 (N_5620,N_5409,N_5048);
nand U5621 (N_5621,N_5415,N_5447);
xor U5622 (N_5622,N_5479,N_5371);
or U5623 (N_5623,N_5181,N_5467);
and U5624 (N_5624,N_5259,N_5288);
and U5625 (N_5625,N_5067,N_5289);
and U5626 (N_5626,N_5120,N_5167);
xnor U5627 (N_5627,N_5109,N_5473);
nand U5628 (N_5628,N_5239,N_5033);
or U5629 (N_5629,N_5102,N_5160);
xnor U5630 (N_5630,N_5433,N_5117);
nand U5631 (N_5631,N_5435,N_5010);
xor U5632 (N_5632,N_5483,N_5041);
nand U5633 (N_5633,N_5141,N_5116);
nor U5634 (N_5634,N_5493,N_5238);
or U5635 (N_5635,N_5270,N_5242);
nand U5636 (N_5636,N_5312,N_5499);
nand U5637 (N_5637,N_5136,N_5015);
xnor U5638 (N_5638,N_5122,N_5066);
nor U5639 (N_5639,N_5437,N_5118);
and U5640 (N_5640,N_5132,N_5230);
nand U5641 (N_5641,N_5135,N_5274);
or U5642 (N_5642,N_5059,N_5396);
xnor U5643 (N_5643,N_5423,N_5374);
and U5644 (N_5644,N_5187,N_5223);
xnor U5645 (N_5645,N_5151,N_5088);
and U5646 (N_5646,N_5017,N_5263);
nand U5647 (N_5647,N_5372,N_5256);
nand U5648 (N_5648,N_5028,N_5278);
or U5649 (N_5649,N_5005,N_5450);
xor U5650 (N_5650,N_5369,N_5295);
nand U5651 (N_5651,N_5244,N_5201);
or U5652 (N_5652,N_5001,N_5192);
nor U5653 (N_5653,N_5004,N_5350);
xor U5654 (N_5654,N_5334,N_5465);
or U5655 (N_5655,N_5444,N_5176);
or U5656 (N_5656,N_5150,N_5174);
nand U5657 (N_5657,N_5043,N_5029);
and U5658 (N_5658,N_5302,N_5292);
nor U5659 (N_5659,N_5443,N_5049);
nor U5660 (N_5660,N_5191,N_5038);
nand U5661 (N_5661,N_5355,N_5119);
or U5662 (N_5662,N_5237,N_5082);
or U5663 (N_5663,N_5303,N_5449);
xor U5664 (N_5664,N_5022,N_5419);
xor U5665 (N_5665,N_5317,N_5113);
xor U5666 (N_5666,N_5323,N_5207);
nor U5667 (N_5667,N_5052,N_5007);
and U5668 (N_5668,N_5079,N_5276);
and U5669 (N_5669,N_5063,N_5368);
or U5670 (N_5670,N_5019,N_5440);
or U5671 (N_5671,N_5370,N_5083);
nand U5672 (N_5672,N_5226,N_5386);
xnor U5673 (N_5673,N_5020,N_5184);
and U5674 (N_5674,N_5421,N_5398);
nand U5675 (N_5675,N_5158,N_5061);
nand U5676 (N_5676,N_5404,N_5328);
nor U5677 (N_5677,N_5157,N_5476);
nor U5678 (N_5678,N_5428,N_5202);
and U5679 (N_5679,N_5240,N_5222);
and U5680 (N_5680,N_5154,N_5297);
xnor U5681 (N_5681,N_5173,N_5418);
and U5682 (N_5682,N_5101,N_5260);
or U5683 (N_5683,N_5321,N_5477);
and U5684 (N_5684,N_5261,N_5310);
or U5685 (N_5685,N_5387,N_5197);
xnor U5686 (N_5686,N_5382,N_5177);
xnor U5687 (N_5687,N_5486,N_5018);
or U5688 (N_5688,N_5488,N_5105);
nand U5689 (N_5689,N_5163,N_5165);
nand U5690 (N_5690,N_5003,N_5308);
and U5691 (N_5691,N_5283,N_5087);
nand U5692 (N_5692,N_5231,N_5159);
xnor U5693 (N_5693,N_5126,N_5280);
or U5694 (N_5694,N_5121,N_5457);
nor U5695 (N_5695,N_5156,N_5363);
and U5696 (N_5696,N_5282,N_5204);
and U5697 (N_5697,N_5285,N_5346);
or U5698 (N_5698,N_5236,N_5149);
xor U5699 (N_5699,N_5111,N_5448);
or U5700 (N_5700,N_5180,N_5284);
nor U5701 (N_5701,N_5316,N_5107);
nand U5702 (N_5702,N_5058,N_5381);
nor U5703 (N_5703,N_5410,N_5484);
nor U5704 (N_5704,N_5452,N_5137);
nor U5705 (N_5705,N_5314,N_5057);
nor U5706 (N_5706,N_5291,N_5425);
xnor U5707 (N_5707,N_5092,N_5406);
or U5708 (N_5708,N_5147,N_5343);
xnor U5709 (N_5709,N_5279,N_5340);
or U5710 (N_5710,N_5047,N_5489);
nand U5711 (N_5711,N_5359,N_5397);
nor U5712 (N_5712,N_5241,N_5301);
or U5713 (N_5713,N_5155,N_5074);
and U5714 (N_5714,N_5471,N_5086);
nor U5715 (N_5715,N_5153,N_5128);
nor U5716 (N_5716,N_5068,N_5213);
nor U5717 (N_5717,N_5032,N_5035);
nand U5718 (N_5718,N_5089,N_5070);
nand U5719 (N_5719,N_5186,N_5164);
nand U5720 (N_5720,N_5217,N_5046);
xnor U5721 (N_5721,N_5071,N_5009);
or U5722 (N_5722,N_5490,N_5169);
nand U5723 (N_5723,N_5454,N_5429);
and U5724 (N_5724,N_5139,N_5170);
nor U5725 (N_5725,N_5224,N_5482);
or U5726 (N_5726,N_5366,N_5391);
and U5727 (N_5727,N_5030,N_5051);
and U5728 (N_5728,N_5384,N_5281);
xnor U5729 (N_5729,N_5407,N_5146);
nand U5730 (N_5730,N_5319,N_5208);
xnor U5731 (N_5731,N_5332,N_5131);
or U5732 (N_5732,N_5134,N_5182);
nand U5733 (N_5733,N_5272,N_5142);
and U5734 (N_5734,N_5441,N_5353);
nand U5735 (N_5735,N_5199,N_5466);
xor U5736 (N_5736,N_5013,N_5478);
and U5737 (N_5737,N_5216,N_5104);
and U5738 (N_5738,N_5183,N_5336);
nand U5739 (N_5739,N_5358,N_5027);
nand U5740 (N_5740,N_5356,N_5091);
nor U5741 (N_5741,N_5212,N_5474);
nand U5742 (N_5742,N_5084,N_5145);
nand U5743 (N_5743,N_5307,N_5002);
nand U5744 (N_5744,N_5050,N_5148);
nor U5745 (N_5745,N_5431,N_5096);
and U5746 (N_5746,N_5456,N_5275);
or U5747 (N_5747,N_5464,N_5257);
nor U5748 (N_5748,N_5400,N_5497);
xor U5749 (N_5749,N_5269,N_5342);
or U5750 (N_5750,N_5272,N_5293);
or U5751 (N_5751,N_5174,N_5454);
and U5752 (N_5752,N_5059,N_5298);
nor U5753 (N_5753,N_5179,N_5288);
nor U5754 (N_5754,N_5239,N_5089);
nand U5755 (N_5755,N_5023,N_5475);
nor U5756 (N_5756,N_5364,N_5460);
and U5757 (N_5757,N_5059,N_5256);
nor U5758 (N_5758,N_5185,N_5286);
or U5759 (N_5759,N_5017,N_5086);
xnor U5760 (N_5760,N_5008,N_5415);
nor U5761 (N_5761,N_5110,N_5360);
or U5762 (N_5762,N_5110,N_5430);
nor U5763 (N_5763,N_5206,N_5229);
or U5764 (N_5764,N_5051,N_5032);
and U5765 (N_5765,N_5467,N_5193);
nor U5766 (N_5766,N_5045,N_5050);
and U5767 (N_5767,N_5071,N_5257);
and U5768 (N_5768,N_5226,N_5180);
xnor U5769 (N_5769,N_5405,N_5491);
nand U5770 (N_5770,N_5285,N_5221);
and U5771 (N_5771,N_5062,N_5165);
xor U5772 (N_5772,N_5195,N_5497);
nand U5773 (N_5773,N_5197,N_5493);
and U5774 (N_5774,N_5100,N_5233);
nand U5775 (N_5775,N_5036,N_5392);
nor U5776 (N_5776,N_5257,N_5190);
and U5777 (N_5777,N_5047,N_5210);
or U5778 (N_5778,N_5445,N_5470);
nand U5779 (N_5779,N_5361,N_5393);
and U5780 (N_5780,N_5449,N_5034);
nor U5781 (N_5781,N_5122,N_5423);
nor U5782 (N_5782,N_5382,N_5481);
xor U5783 (N_5783,N_5289,N_5346);
nand U5784 (N_5784,N_5328,N_5443);
nand U5785 (N_5785,N_5016,N_5049);
xnor U5786 (N_5786,N_5498,N_5486);
or U5787 (N_5787,N_5060,N_5140);
and U5788 (N_5788,N_5431,N_5235);
nor U5789 (N_5789,N_5484,N_5198);
nor U5790 (N_5790,N_5212,N_5211);
nand U5791 (N_5791,N_5167,N_5094);
nand U5792 (N_5792,N_5458,N_5181);
xor U5793 (N_5793,N_5362,N_5165);
nand U5794 (N_5794,N_5344,N_5225);
nand U5795 (N_5795,N_5020,N_5083);
and U5796 (N_5796,N_5010,N_5162);
nand U5797 (N_5797,N_5444,N_5089);
and U5798 (N_5798,N_5167,N_5022);
nand U5799 (N_5799,N_5205,N_5050);
and U5800 (N_5800,N_5109,N_5086);
or U5801 (N_5801,N_5322,N_5142);
or U5802 (N_5802,N_5090,N_5150);
nor U5803 (N_5803,N_5433,N_5457);
and U5804 (N_5804,N_5274,N_5210);
xor U5805 (N_5805,N_5409,N_5041);
nand U5806 (N_5806,N_5258,N_5485);
nor U5807 (N_5807,N_5226,N_5081);
and U5808 (N_5808,N_5048,N_5336);
nor U5809 (N_5809,N_5070,N_5170);
xor U5810 (N_5810,N_5411,N_5441);
nor U5811 (N_5811,N_5204,N_5484);
or U5812 (N_5812,N_5276,N_5494);
or U5813 (N_5813,N_5240,N_5109);
xnor U5814 (N_5814,N_5343,N_5179);
nand U5815 (N_5815,N_5082,N_5327);
or U5816 (N_5816,N_5308,N_5422);
nor U5817 (N_5817,N_5407,N_5289);
nor U5818 (N_5818,N_5205,N_5165);
and U5819 (N_5819,N_5497,N_5267);
nand U5820 (N_5820,N_5214,N_5335);
xnor U5821 (N_5821,N_5006,N_5131);
nor U5822 (N_5822,N_5367,N_5333);
xor U5823 (N_5823,N_5053,N_5137);
nand U5824 (N_5824,N_5247,N_5475);
xnor U5825 (N_5825,N_5419,N_5471);
and U5826 (N_5826,N_5069,N_5487);
nand U5827 (N_5827,N_5488,N_5368);
or U5828 (N_5828,N_5111,N_5112);
or U5829 (N_5829,N_5222,N_5119);
nand U5830 (N_5830,N_5134,N_5492);
or U5831 (N_5831,N_5131,N_5335);
nand U5832 (N_5832,N_5054,N_5348);
nand U5833 (N_5833,N_5033,N_5045);
xnor U5834 (N_5834,N_5321,N_5287);
xor U5835 (N_5835,N_5130,N_5371);
nand U5836 (N_5836,N_5244,N_5163);
and U5837 (N_5837,N_5337,N_5326);
or U5838 (N_5838,N_5273,N_5137);
xnor U5839 (N_5839,N_5199,N_5239);
or U5840 (N_5840,N_5033,N_5030);
and U5841 (N_5841,N_5297,N_5030);
xor U5842 (N_5842,N_5316,N_5013);
nor U5843 (N_5843,N_5147,N_5322);
or U5844 (N_5844,N_5150,N_5274);
nand U5845 (N_5845,N_5321,N_5498);
xnor U5846 (N_5846,N_5379,N_5004);
and U5847 (N_5847,N_5380,N_5214);
xnor U5848 (N_5848,N_5481,N_5205);
xor U5849 (N_5849,N_5446,N_5166);
or U5850 (N_5850,N_5248,N_5108);
and U5851 (N_5851,N_5069,N_5309);
xnor U5852 (N_5852,N_5287,N_5044);
and U5853 (N_5853,N_5144,N_5046);
nor U5854 (N_5854,N_5456,N_5440);
or U5855 (N_5855,N_5050,N_5017);
or U5856 (N_5856,N_5122,N_5100);
and U5857 (N_5857,N_5282,N_5192);
and U5858 (N_5858,N_5478,N_5011);
nand U5859 (N_5859,N_5427,N_5423);
nor U5860 (N_5860,N_5024,N_5357);
and U5861 (N_5861,N_5433,N_5266);
nand U5862 (N_5862,N_5388,N_5024);
nand U5863 (N_5863,N_5189,N_5072);
nand U5864 (N_5864,N_5198,N_5309);
nor U5865 (N_5865,N_5394,N_5260);
or U5866 (N_5866,N_5178,N_5410);
xnor U5867 (N_5867,N_5416,N_5184);
nor U5868 (N_5868,N_5282,N_5001);
nand U5869 (N_5869,N_5302,N_5471);
or U5870 (N_5870,N_5275,N_5234);
xor U5871 (N_5871,N_5078,N_5123);
nor U5872 (N_5872,N_5340,N_5225);
nand U5873 (N_5873,N_5230,N_5306);
xor U5874 (N_5874,N_5202,N_5096);
xor U5875 (N_5875,N_5124,N_5171);
and U5876 (N_5876,N_5398,N_5089);
xnor U5877 (N_5877,N_5102,N_5123);
nand U5878 (N_5878,N_5347,N_5165);
or U5879 (N_5879,N_5346,N_5272);
xnor U5880 (N_5880,N_5120,N_5268);
nand U5881 (N_5881,N_5375,N_5253);
or U5882 (N_5882,N_5140,N_5444);
and U5883 (N_5883,N_5459,N_5435);
xor U5884 (N_5884,N_5374,N_5307);
nor U5885 (N_5885,N_5466,N_5001);
or U5886 (N_5886,N_5215,N_5201);
nand U5887 (N_5887,N_5067,N_5017);
and U5888 (N_5888,N_5336,N_5017);
nand U5889 (N_5889,N_5407,N_5360);
nand U5890 (N_5890,N_5377,N_5416);
or U5891 (N_5891,N_5216,N_5089);
nand U5892 (N_5892,N_5141,N_5464);
or U5893 (N_5893,N_5138,N_5028);
nand U5894 (N_5894,N_5055,N_5323);
xor U5895 (N_5895,N_5310,N_5204);
xor U5896 (N_5896,N_5271,N_5279);
or U5897 (N_5897,N_5092,N_5442);
nand U5898 (N_5898,N_5247,N_5010);
or U5899 (N_5899,N_5346,N_5476);
xor U5900 (N_5900,N_5414,N_5066);
nand U5901 (N_5901,N_5169,N_5380);
nand U5902 (N_5902,N_5306,N_5493);
or U5903 (N_5903,N_5201,N_5060);
nor U5904 (N_5904,N_5097,N_5365);
nand U5905 (N_5905,N_5346,N_5074);
nor U5906 (N_5906,N_5048,N_5097);
xnor U5907 (N_5907,N_5256,N_5203);
xnor U5908 (N_5908,N_5221,N_5279);
or U5909 (N_5909,N_5303,N_5483);
nor U5910 (N_5910,N_5176,N_5226);
xnor U5911 (N_5911,N_5256,N_5130);
xnor U5912 (N_5912,N_5084,N_5344);
xnor U5913 (N_5913,N_5258,N_5162);
nor U5914 (N_5914,N_5060,N_5332);
nor U5915 (N_5915,N_5438,N_5199);
and U5916 (N_5916,N_5303,N_5055);
xor U5917 (N_5917,N_5046,N_5030);
and U5918 (N_5918,N_5437,N_5334);
or U5919 (N_5919,N_5493,N_5153);
and U5920 (N_5920,N_5118,N_5488);
nand U5921 (N_5921,N_5142,N_5168);
nor U5922 (N_5922,N_5227,N_5199);
or U5923 (N_5923,N_5047,N_5369);
nand U5924 (N_5924,N_5401,N_5234);
nand U5925 (N_5925,N_5052,N_5269);
nand U5926 (N_5926,N_5460,N_5271);
and U5927 (N_5927,N_5249,N_5140);
xnor U5928 (N_5928,N_5449,N_5347);
nand U5929 (N_5929,N_5110,N_5478);
nand U5930 (N_5930,N_5021,N_5202);
nand U5931 (N_5931,N_5189,N_5146);
xnor U5932 (N_5932,N_5341,N_5116);
or U5933 (N_5933,N_5150,N_5306);
nand U5934 (N_5934,N_5309,N_5289);
or U5935 (N_5935,N_5104,N_5156);
and U5936 (N_5936,N_5040,N_5077);
or U5937 (N_5937,N_5018,N_5211);
nand U5938 (N_5938,N_5357,N_5181);
or U5939 (N_5939,N_5352,N_5160);
or U5940 (N_5940,N_5188,N_5372);
nand U5941 (N_5941,N_5438,N_5018);
and U5942 (N_5942,N_5368,N_5445);
nor U5943 (N_5943,N_5182,N_5098);
nand U5944 (N_5944,N_5278,N_5069);
nor U5945 (N_5945,N_5215,N_5371);
xnor U5946 (N_5946,N_5315,N_5048);
and U5947 (N_5947,N_5109,N_5420);
nand U5948 (N_5948,N_5194,N_5426);
and U5949 (N_5949,N_5025,N_5054);
xnor U5950 (N_5950,N_5361,N_5191);
nor U5951 (N_5951,N_5056,N_5086);
xnor U5952 (N_5952,N_5147,N_5377);
nor U5953 (N_5953,N_5328,N_5020);
xnor U5954 (N_5954,N_5219,N_5181);
or U5955 (N_5955,N_5038,N_5358);
and U5956 (N_5956,N_5233,N_5278);
or U5957 (N_5957,N_5036,N_5096);
and U5958 (N_5958,N_5376,N_5094);
nor U5959 (N_5959,N_5114,N_5463);
xnor U5960 (N_5960,N_5365,N_5276);
nand U5961 (N_5961,N_5235,N_5294);
nor U5962 (N_5962,N_5346,N_5308);
and U5963 (N_5963,N_5357,N_5410);
and U5964 (N_5964,N_5085,N_5427);
and U5965 (N_5965,N_5196,N_5334);
nor U5966 (N_5966,N_5446,N_5157);
or U5967 (N_5967,N_5208,N_5305);
nand U5968 (N_5968,N_5054,N_5499);
xor U5969 (N_5969,N_5017,N_5192);
nand U5970 (N_5970,N_5414,N_5436);
nand U5971 (N_5971,N_5071,N_5190);
nor U5972 (N_5972,N_5031,N_5218);
xnor U5973 (N_5973,N_5005,N_5006);
or U5974 (N_5974,N_5190,N_5306);
and U5975 (N_5975,N_5062,N_5099);
xor U5976 (N_5976,N_5298,N_5442);
or U5977 (N_5977,N_5407,N_5023);
nor U5978 (N_5978,N_5271,N_5244);
xor U5979 (N_5979,N_5301,N_5117);
nand U5980 (N_5980,N_5418,N_5378);
xnor U5981 (N_5981,N_5051,N_5485);
xor U5982 (N_5982,N_5022,N_5401);
and U5983 (N_5983,N_5228,N_5296);
or U5984 (N_5984,N_5495,N_5336);
nor U5985 (N_5985,N_5297,N_5402);
xnor U5986 (N_5986,N_5257,N_5302);
or U5987 (N_5987,N_5118,N_5009);
nor U5988 (N_5988,N_5475,N_5310);
and U5989 (N_5989,N_5414,N_5018);
nor U5990 (N_5990,N_5194,N_5256);
nand U5991 (N_5991,N_5366,N_5027);
and U5992 (N_5992,N_5447,N_5143);
or U5993 (N_5993,N_5342,N_5364);
or U5994 (N_5994,N_5091,N_5228);
nand U5995 (N_5995,N_5135,N_5088);
xor U5996 (N_5996,N_5418,N_5410);
xor U5997 (N_5997,N_5008,N_5326);
and U5998 (N_5998,N_5202,N_5152);
xnor U5999 (N_5999,N_5225,N_5331);
nand U6000 (N_6000,N_5937,N_5806);
or U6001 (N_6001,N_5925,N_5655);
or U6002 (N_6002,N_5871,N_5886);
xor U6003 (N_6003,N_5973,N_5972);
nand U6004 (N_6004,N_5620,N_5847);
and U6005 (N_6005,N_5903,N_5965);
xnor U6006 (N_6006,N_5692,N_5898);
nor U6007 (N_6007,N_5833,N_5667);
or U6008 (N_6008,N_5567,N_5990);
and U6009 (N_6009,N_5911,N_5938);
or U6010 (N_6010,N_5525,N_5701);
xnor U6011 (N_6011,N_5890,N_5555);
nand U6012 (N_6012,N_5939,N_5538);
or U6013 (N_6013,N_5659,N_5974);
nor U6014 (N_6014,N_5604,N_5571);
nor U6015 (N_6015,N_5829,N_5810);
nor U6016 (N_6016,N_5896,N_5794);
xor U6017 (N_6017,N_5653,N_5980);
nand U6018 (N_6018,N_5891,N_5504);
and U6019 (N_6019,N_5500,N_5636);
xnor U6020 (N_6020,N_5707,N_5734);
and U6021 (N_6021,N_5987,N_5675);
or U6022 (N_6022,N_5738,N_5543);
nand U6023 (N_6023,N_5897,N_5637);
xnor U6024 (N_6024,N_5730,N_5857);
or U6025 (N_6025,N_5695,N_5761);
nand U6026 (N_6026,N_5874,N_5901);
or U6027 (N_6027,N_5600,N_5688);
or U6028 (N_6028,N_5586,N_5536);
xor U6029 (N_6029,N_5762,N_5619);
or U6030 (N_6030,N_5617,N_5670);
xnor U6031 (N_6031,N_5785,N_5817);
nand U6032 (N_6032,N_5658,N_5927);
or U6033 (N_6033,N_5855,N_5912);
nand U6034 (N_6034,N_5867,N_5507);
and U6035 (N_6035,N_5608,N_5698);
nand U6036 (N_6036,N_5622,N_5852);
nand U6037 (N_6037,N_5501,N_5862);
nand U6038 (N_6038,N_5728,N_5663);
or U6039 (N_6039,N_5529,N_5958);
nand U6040 (N_6040,N_5657,N_5624);
xor U6041 (N_6041,N_5917,N_5724);
and U6042 (N_6042,N_5683,N_5934);
xnor U6043 (N_6043,N_5775,N_5589);
nand U6044 (N_6044,N_5506,N_5892);
or U6045 (N_6045,N_5685,N_5566);
nor U6046 (N_6046,N_5941,N_5635);
or U6047 (N_6047,N_5792,N_5848);
or U6048 (N_6048,N_5825,N_5537);
and U6049 (N_6049,N_5557,N_5588);
nor U6050 (N_6050,N_5929,N_5665);
xor U6051 (N_6051,N_5978,N_5598);
and U6052 (N_6052,N_5573,N_5826);
or U6053 (N_6053,N_5520,N_5765);
or U6054 (N_6054,N_5832,N_5576);
nor U6055 (N_6055,N_5603,N_5596);
nor U6056 (N_6056,N_5554,N_5986);
xor U6057 (N_6057,N_5781,N_5584);
xnor U6058 (N_6058,N_5725,N_5764);
or U6059 (N_6059,N_5805,N_5813);
and U6060 (N_6060,N_5945,N_5577);
and U6061 (N_6061,N_5766,N_5668);
nand U6062 (N_6062,N_5514,N_5900);
or U6063 (N_6063,N_5613,N_5689);
nor U6064 (N_6064,N_5642,N_5732);
and U6065 (N_6065,N_5513,N_5627);
or U6066 (N_6066,N_5932,N_5643);
and U6067 (N_6067,N_5672,N_5928);
or U6068 (N_6068,N_5835,N_5870);
nor U6069 (N_6069,N_5691,N_5943);
or U6070 (N_6070,N_5547,N_5797);
nor U6071 (N_6071,N_5541,N_5854);
or U6072 (N_6072,N_5906,N_5998);
nand U6073 (N_6073,N_5646,N_5976);
and U6074 (N_6074,N_5840,N_5907);
nor U6075 (N_6075,N_5649,N_5522);
nand U6076 (N_6076,N_5539,N_5790);
nor U6077 (N_6077,N_5581,N_5988);
nand U6078 (N_6078,N_5585,N_5739);
or U6079 (N_6079,N_5666,N_5760);
or U6080 (N_6080,N_5621,N_5632);
nand U6081 (N_6081,N_5851,N_5748);
nand U6082 (N_6082,N_5517,N_5592);
nand U6083 (N_6083,N_5737,N_5673);
or U6084 (N_6084,N_5580,N_5952);
xor U6085 (N_6085,N_5863,N_5532);
and U6086 (N_6086,N_5908,N_5800);
nor U6087 (N_6087,N_5887,N_5570);
and U6088 (N_6088,N_5503,N_5718);
or U6089 (N_6089,N_5744,N_5936);
or U6090 (N_6090,N_5818,N_5526);
or U6091 (N_6091,N_5989,N_5772);
or U6092 (N_6092,N_5644,N_5796);
and U6093 (N_6093,N_5582,N_5742);
xnor U6094 (N_6094,N_5966,N_5647);
xnor U6095 (N_6095,N_5696,N_5860);
or U6096 (N_6096,N_5815,N_5572);
or U6097 (N_6097,N_5599,N_5700);
nand U6098 (N_6098,N_5618,N_5814);
xor U6099 (N_6099,N_5930,N_5823);
nand U6100 (N_6100,N_5713,N_5678);
and U6101 (N_6101,N_5793,N_5975);
xor U6102 (N_6102,N_5578,N_5949);
xor U6103 (N_6103,N_5662,N_5575);
or U6104 (N_6104,N_5704,N_5940);
or U6105 (N_6105,N_5615,N_5866);
nand U6106 (N_6106,N_5770,N_5864);
or U6107 (N_6107,N_5579,N_5991);
and U6108 (N_6108,N_5716,N_5697);
or U6109 (N_6109,N_5933,N_5816);
or U6110 (N_6110,N_5953,N_5558);
xor U6111 (N_6111,N_5623,N_5527);
or U6112 (N_6112,N_5523,N_5992);
nand U6113 (N_6113,N_5856,N_5768);
nand U6114 (N_6114,N_5758,N_5902);
nor U6115 (N_6115,N_5755,N_5609);
nand U6116 (N_6116,N_5594,N_5510);
and U6117 (N_6117,N_5719,N_5798);
or U6118 (N_6118,N_5751,N_5509);
nand U6119 (N_6119,N_5920,N_5648);
xnor U6120 (N_6120,N_5574,N_5569);
nand U6121 (N_6121,N_5703,N_5954);
nor U6122 (N_6122,N_5551,N_5721);
nor U6123 (N_6123,N_5838,N_5802);
or U6124 (N_6124,N_5553,N_5693);
and U6125 (N_6125,N_5819,N_5605);
nand U6126 (N_6126,N_5947,N_5904);
xor U6127 (N_6127,N_5512,N_5858);
or U6128 (N_6128,N_5893,N_5740);
or U6129 (N_6129,N_5749,N_5656);
and U6130 (N_6130,N_5562,N_5565);
nand U6131 (N_6131,N_5834,N_5951);
or U6132 (N_6132,N_5787,N_5593);
xor U6133 (N_6133,N_5731,N_5950);
or U6134 (N_6134,N_5528,N_5752);
and U6135 (N_6135,N_5877,N_5982);
nand U6136 (N_6136,N_5804,N_5922);
and U6137 (N_6137,N_5779,N_5881);
or U6138 (N_6138,N_5616,N_5850);
nand U6139 (N_6139,N_5763,N_5519);
and U6140 (N_6140,N_5607,N_5597);
nand U6141 (N_6141,N_5601,N_5963);
or U6142 (N_6142,N_5694,N_5780);
and U6143 (N_6143,N_5924,N_5531);
and U6144 (N_6144,N_5511,N_5849);
nor U6145 (N_6145,N_5610,N_5914);
and U6146 (N_6146,N_5722,N_5777);
xnor U6147 (N_6147,N_5630,N_5747);
nor U6148 (N_6148,N_5899,N_5710);
and U6149 (N_6149,N_5996,N_5652);
and U6150 (N_6150,N_5782,N_5709);
or U6151 (N_6151,N_5638,N_5746);
xnor U6152 (N_6152,N_5669,N_5743);
or U6153 (N_6153,N_5705,N_5960);
xnor U6154 (N_6154,N_5808,N_5828);
nor U6155 (N_6155,N_5803,N_5677);
nor U6156 (N_6156,N_5639,N_5880);
xor U6157 (N_6157,N_5961,N_5641);
or U6158 (N_6158,N_5591,N_5985);
nand U6159 (N_6159,N_5625,N_5645);
nor U6160 (N_6160,N_5769,N_5865);
xor U6161 (N_6161,N_5905,N_5587);
xnor U6162 (N_6162,N_5708,N_5595);
or U6163 (N_6163,N_5773,N_5611);
and U6164 (N_6164,N_5799,N_5970);
nand U6165 (N_6165,N_5962,N_5699);
xor U6166 (N_6166,N_5712,N_5729);
nand U6167 (N_6167,N_5508,N_5983);
or U6168 (N_6168,N_5872,N_5869);
or U6169 (N_6169,N_5836,N_5923);
or U6170 (N_6170,N_5629,N_5502);
xnor U6171 (N_6171,N_5842,N_5868);
nor U6172 (N_6172,N_5521,N_5711);
nor U6173 (N_6173,N_5757,N_5778);
xnor U6174 (N_6174,N_5861,N_5631);
nor U6175 (N_6175,N_5956,N_5843);
or U6176 (N_6176,N_5984,N_5682);
nor U6177 (N_6177,N_5795,N_5686);
or U6178 (N_6178,N_5767,N_5942);
and U6179 (N_6179,N_5759,N_5735);
or U6180 (N_6180,N_5919,N_5727);
nor U6181 (N_6181,N_5981,N_5745);
xor U6182 (N_6182,N_5690,N_5967);
nor U6183 (N_6183,N_5791,N_5602);
xor U6184 (N_6184,N_5968,N_5807);
nor U6185 (N_6185,N_5918,N_5559);
nor U6186 (N_6186,N_5926,N_5831);
nand U6187 (N_6187,N_5606,N_5651);
or U6188 (N_6188,N_5921,N_5590);
nor U6189 (N_6189,N_5946,N_5754);
nor U6190 (N_6190,N_5977,N_5999);
xnor U6191 (N_6191,N_5664,N_5997);
and U6192 (N_6192,N_5715,N_5812);
nand U6193 (N_6193,N_5530,N_5549);
and U6194 (N_6194,N_5811,N_5534);
and U6195 (N_6195,N_5994,N_5830);
or U6196 (N_6196,N_5957,N_5827);
nor U6197 (N_6197,N_5895,N_5505);
nor U6198 (N_6198,N_5614,N_5995);
or U6199 (N_6199,N_5824,N_5518);
nand U6200 (N_6200,N_5839,N_5809);
or U6201 (N_6201,N_5959,N_5654);
nor U6202 (N_6202,N_5674,N_5640);
xor U6203 (N_6203,N_5671,N_5633);
xnor U6204 (N_6204,N_5550,N_5789);
nand U6205 (N_6205,N_5756,N_5971);
or U6206 (N_6206,N_5913,N_5948);
nand U6207 (N_6207,N_5786,N_5944);
nor U6208 (N_6208,N_5841,N_5822);
nand U6209 (N_6209,N_5563,N_5516);
xor U6210 (N_6210,N_5628,N_5568);
or U6211 (N_6211,N_5533,N_5684);
xnor U6212 (N_6212,N_5821,N_5626);
xor U6213 (N_6213,N_5964,N_5878);
nor U6214 (N_6214,N_5583,N_5717);
nand U6215 (N_6215,N_5879,N_5969);
and U6216 (N_6216,N_5801,N_5845);
nand U6217 (N_6217,N_5535,N_5883);
nand U6218 (N_6218,N_5931,N_5788);
nand U6219 (N_6219,N_5820,N_5771);
or U6220 (N_6220,N_5916,N_5650);
nand U6221 (N_6221,N_5844,N_5979);
xnor U6222 (N_6222,N_5774,N_5873);
nand U6223 (N_6223,N_5540,N_5876);
and U6224 (N_6224,N_5723,N_5889);
xor U6225 (N_6225,N_5676,N_5783);
or U6226 (N_6226,N_5955,N_5634);
and U6227 (N_6227,N_5884,N_5679);
and U6228 (N_6228,N_5859,N_5875);
nand U6229 (N_6229,N_5776,N_5935);
nand U6230 (N_6230,N_5993,N_5885);
and U6231 (N_6231,N_5733,N_5687);
nand U6232 (N_6232,N_5544,N_5560);
or U6233 (N_6233,N_5888,N_5612);
nand U6234 (N_6234,N_5545,N_5915);
and U6235 (N_6235,N_5894,N_5546);
xnor U6236 (N_6236,N_5515,N_5702);
nand U6237 (N_6237,N_5661,N_5846);
and U6238 (N_6238,N_5542,N_5882);
nand U6239 (N_6239,N_5741,N_5853);
nand U6240 (N_6240,N_5784,N_5524);
nand U6241 (N_6241,N_5736,N_5910);
or U6242 (N_6242,N_5564,N_5909);
nand U6243 (N_6243,N_5680,N_5660);
nand U6244 (N_6244,N_5726,N_5753);
nand U6245 (N_6245,N_5720,N_5561);
nor U6246 (N_6246,N_5706,N_5681);
xnor U6247 (N_6247,N_5750,N_5714);
or U6248 (N_6248,N_5837,N_5548);
and U6249 (N_6249,N_5556,N_5552);
nand U6250 (N_6250,N_5607,N_5781);
xnor U6251 (N_6251,N_5547,N_5940);
or U6252 (N_6252,N_5513,N_5823);
xor U6253 (N_6253,N_5694,N_5865);
nor U6254 (N_6254,N_5882,N_5516);
and U6255 (N_6255,N_5984,N_5670);
or U6256 (N_6256,N_5696,N_5800);
nand U6257 (N_6257,N_5632,N_5821);
nor U6258 (N_6258,N_5831,N_5698);
or U6259 (N_6259,N_5803,N_5755);
nand U6260 (N_6260,N_5801,N_5713);
or U6261 (N_6261,N_5653,N_5750);
nor U6262 (N_6262,N_5711,N_5930);
or U6263 (N_6263,N_5985,N_5944);
nand U6264 (N_6264,N_5831,N_5565);
or U6265 (N_6265,N_5504,N_5952);
nand U6266 (N_6266,N_5762,N_5838);
or U6267 (N_6267,N_5708,N_5732);
xnor U6268 (N_6268,N_5709,N_5523);
xor U6269 (N_6269,N_5846,N_5759);
and U6270 (N_6270,N_5837,N_5865);
xor U6271 (N_6271,N_5964,N_5620);
and U6272 (N_6272,N_5984,N_5748);
xor U6273 (N_6273,N_5507,N_5862);
nand U6274 (N_6274,N_5620,N_5797);
nand U6275 (N_6275,N_5853,N_5755);
or U6276 (N_6276,N_5728,N_5527);
nand U6277 (N_6277,N_5792,N_5878);
or U6278 (N_6278,N_5629,N_5907);
nor U6279 (N_6279,N_5794,N_5565);
or U6280 (N_6280,N_5898,N_5810);
nor U6281 (N_6281,N_5681,N_5878);
or U6282 (N_6282,N_5613,N_5621);
nor U6283 (N_6283,N_5825,N_5714);
nand U6284 (N_6284,N_5889,N_5565);
nor U6285 (N_6285,N_5520,N_5552);
nand U6286 (N_6286,N_5812,N_5925);
nand U6287 (N_6287,N_5982,N_5770);
nor U6288 (N_6288,N_5695,N_5691);
nand U6289 (N_6289,N_5860,N_5893);
xor U6290 (N_6290,N_5663,N_5617);
xnor U6291 (N_6291,N_5913,N_5783);
nor U6292 (N_6292,N_5932,N_5601);
xnor U6293 (N_6293,N_5765,N_5826);
xnor U6294 (N_6294,N_5884,N_5962);
or U6295 (N_6295,N_5851,N_5904);
xor U6296 (N_6296,N_5532,N_5742);
xnor U6297 (N_6297,N_5739,N_5842);
nand U6298 (N_6298,N_5943,N_5611);
xnor U6299 (N_6299,N_5876,N_5574);
xor U6300 (N_6300,N_5505,N_5792);
xnor U6301 (N_6301,N_5682,N_5766);
or U6302 (N_6302,N_5791,N_5649);
xor U6303 (N_6303,N_5856,N_5802);
and U6304 (N_6304,N_5890,N_5887);
and U6305 (N_6305,N_5923,N_5678);
and U6306 (N_6306,N_5589,N_5676);
xnor U6307 (N_6307,N_5700,N_5721);
or U6308 (N_6308,N_5769,N_5651);
and U6309 (N_6309,N_5978,N_5914);
nor U6310 (N_6310,N_5848,N_5582);
nand U6311 (N_6311,N_5912,N_5944);
xnor U6312 (N_6312,N_5614,N_5875);
xnor U6313 (N_6313,N_5977,N_5952);
and U6314 (N_6314,N_5612,N_5760);
xnor U6315 (N_6315,N_5833,N_5611);
or U6316 (N_6316,N_5646,N_5998);
nor U6317 (N_6317,N_5677,N_5518);
nor U6318 (N_6318,N_5726,N_5508);
xor U6319 (N_6319,N_5883,N_5699);
nor U6320 (N_6320,N_5854,N_5928);
xnor U6321 (N_6321,N_5704,N_5515);
and U6322 (N_6322,N_5805,N_5527);
nand U6323 (N_6323,N_5547,N_5620);
xor U6324 (N_6324,N_5574,N_5674);
xnor U6325 (N_6325,N_5630,N_5960);
and U6326 (N_6326,N_5561,N_5678);
nor U6327 (N_6327,N_5529,N_5564);
and U6328 (N_6328,N_5938,N_5742);
or U6329 (N_6329,N_5617,N_5863);
nor U6330 (N_6330,N_5578,N_5956);
nor U6331 (N_6331,N_5820,N_5985);
and U6332 (N_6332,N_5886,N_5601);
and U6333 (N_6333,N_5639,N_5848);
nor U6334 (N_6334,N_5958,N_5760);
nand U6335 (N_6335,N_5581,N_5647);
nand U6336 (N_6336,N_5581,N_5864);
and U6337 (N_6337,N_5586,N_5769);
or U6338 (N_6338,N_5507,N_5511);
or U6339 (N_6339,N_5592,N_5716);
nor U6340 (N_6340,N_5894,N_5656);
or U6341 (N_6341,N_5606,N_5796);
nand U6342 (N_6342,N_5885,N_5738);
and U6343 (N_6343,N_5926,N_5868);
xnor U6344 (N_6344,N_5919,N_5760);
or U6345 (N_6345,N_5522,N_5697);
or U6346 (N_6346,N_5613,N_5675);
xor U6347 (N_6347,N_5995,N_5887);
and U6348 (N_6348,N_5900,N_5907);
nand U6349 (N_6349,N_5912,N_5572);
xor U6350 (N_6350,N_5554,N_5720);
or U6351 (N_6351,N_5698,N_5940);
nand U6352 (N_6352,N_5586,N_5821);
nand U6353 (N_6353,N_5881,N_5559);
and U6354 (N_6354,N_5839,N_5916);
xor U6355 (N_6355,N_5699,N_5715);
or U6356 (N_6356,N_5759,N_5987);
or U6357 (N_6357,N_5867,N_5992);
nand U6358 (N_6358,N_5750,N_5828);
or U6359 (N_6359,N_5994,N_5863);
or U6360 (N_6360,N_5556,N_5721);
nand U6361 (N_6361,N_5501,N_5984);
and U6362 (N_6362,N_5705,N_5613);
or U6363 (N_6363,N_5834,N_5509);
nor U6364 (N_6364,N_5691,N_5597);
or U6365 (N_6365,N_5948,N_5551);
nor U6366 (N_6366,N_5694,N_5822);
xnor U6367 (N_6367,N_5952,N_5805);
and U6368 (N_6368,N_5881,N_5891);
nor U6369 (N_6369,N_5699,N_5979);
nor U6370 (N_6370,N_5842,N_5534);
xnor U6371 (N_6371,N_5602,N_5706);
nand U6372 (N_6372,N_5622,N_5806);
nor U6373 (N_6373,N_5638,N_5910);
xor U6374 (N_6374,N_5688,N_5604);
nor U6375 (N_6375,N_5519,N_5657);
xor U6376 (N_6376,N_5523,N_5796);
nand U6377 (N_6377,N_5954,N_5878);
xor U6378 (N_6378,N_5616,N_5514);
and U6379 (N_6379,N_5585,N_5795);
or U6380 (N_6380,N_5703,N_5811);
and U6381 (N_6381,N_5991,N_5573);
xor U6382 (N_6382,N_5877,N_5936);
xnor U6383 (N_6383,N_5783,N_5777);
xor U6384 (N_6384,N_5924,N_5948);
and U6385 (N_6385,N_5570,N_5504);
and U6386 (N_6386,N_5654,N_5572);
and U6387 (N_6387,N_5903,N_5692);
or U6388 (N_6388,N_5665,N_5982);
nor U6389 (N_6389,N_5849,N_5620);
xnor U6390 (N_6390,N_5957,N_5971);
nor U6391 (N_6391,N_5672,N_5729);
nor U6392 (N_6392,N_5715,N_5543);
or U6393 (N_6393,N_5864,N_5758);
nand U6394 (N_6394,N_5572,N_5792);
or U6395 (N_6395,N_5609,N_5687);
nor U6396 (N_6396,N_5754,N_5686);
xor U6397 (N_6397,N_5956,N_5911);
nor U6398 (N_6398,N_5779,N_5752);
xnor U6399 (N_6399,N_5915,N_5708);
nand U6400 (N_6400,N_5589,N_5507);
nand U6401 (N_6401,N_5691,N_5517);
and U6402 (N_6402,N_5717,N_5829);
or U6403 (N_6403,N_5740,N_5987);
xor U6404 (N_6404,N_5658,N_5629);
and U6405 (N_6405,N_5602,N_5622);
and U6406 (N_6406,N_5584,N_5849);
and U6407 (N_6407,N_5983,N_5942);
and U6408 (N_6408,N_5944,N_5799);
nor U6409 (N_6409,N_5948,N_5753);
xnor U6410 (N_6410,N_5815,N_5888);
nand U6411 (N_6411,N_5605,N_5644);
xnor U6412 (N_6412,N_5950,N_5546);
or U6413 (N_6413,N_5755,N_5665);
xnor U6414 (N_6414,N_5770,N_5830);
nor U6415 (N_6415,N_5513,N_5710);
nand U6416 (N_6416,N_5609,N_5971);
xnor U6417 (N_6417,N_5819,N_5718);
nor U6418 (N_6418,N_5817,N_5660);
nand U6419 (N_6419,N_5905,N_5537);
nor U6420 (N_6420,N_5503,N_5754);
xnor U6421 (N_6421,N_5951,N_5712);
xnor U6422 (N_6422,N_5530,N_5976);
nand U6423 (N_6423,N_5969,N_5755);
or U6424 (N_6424,N_5591,N_5868);
nand U6425 (N_6425,N_5571,N_5547);
and U6426 (N_6426,N_5940,N_5718);
xnor U6427 (N_6427,N_5832,N_5543);
and U6428 (N_6428,N_5568,N_5610);
or U6429 (N_6429,N_5741,N_5672);
nor U6430 (N_6430,N_5871,N_5774);
xor U6431 (N_6431,N_5721,N_5550);
or U6432 (N_6432,N_5781,N_5633);
or U6433 (N_6433,N_5629,N_5630);
and U6434 (N_6434,N_5501,N_5957);
or U6435 (N_6435,N_5880,N_5686);
and U6436 (N_6436,N_5706,N_5857);
nor U6437 (N_6437,N_5974,N_5715);
xnor U6438 (N_6438,N_5779,N_5727);
or U6439 (N_6439,N_5698,N_5951);
or U6440 (N_6440,N_5905,N_5562);
nor U6441 (N_6441,N_5963,N_5636);
or U6442 (N_6442,N_5796,N_5989);
nand U6443 (N_6443,N_5548,N_5604);
nand U6444 (N_6444,N_5725,N_5844);
nor U6445 (N_6445,N_5903,N_5835);
nand U6446 (N_6446,N_5642,N_5988);
nor U6447 (N_6447,N_5515,N_5684);
or U6448 (N_6448,N_5508,N_5795);
and U6449 (N_6449,N_5743,N_5961);
and U6450 (N_6450,N_5542,N_5856);
xor U6451 (N_6451,N_5728,N_5986);
and U6452 (N_6452,N_5779,N_5940);
nand U6453 (N_6453,N_5674,N_5940);
and U6454 (N_6454,N_5798,N_5608);
nor U6455 (N_6455,N_5698,N_5948);
and U6456 (N_6456,N_5648,N_5834);
and U6457 (N_6457,N_5675,N_5925);
xnor U6458 (N_6458,N_5967,N_5503);
or U6459 (N_6459,N_5976,N_5504);
and U6460 (N_6460,N_5912,N_5804);
and U6461 (N_6461,N_5753,N_5679);
or U6462 (N_6462,N_5781,N_5729);
or U6463 (N_6463,N_5689,N_5535);
nand U6464 (N_6464,N_5790,N_5620);
nand U6465 (N_6465,N_5960,N_5957);
or U6466 (N_6466,N_5960,N_5578);
or U6467 (N_6467,N_5823,N_5797);
nand U6468 (N_6468,N_5673,N_5626);
or U6469 (N_6469,N_5818,N_5503);
nor U6470 (N_6470,N_5744,N_5750);
or U6471 (N_6471,N_5925,N_5778);
xor U6472 (N_6472,N_5667,N_5613);
or U6473 (N_6473,N_5976,N_5569);
nor U6474 (N_6474,N_5844,N_5512);
and U6475 (N_6475,N_5614,N_5770);
or U6476 (N_6476,N_5823,N_5830);
or U6477 (N_6477,N_5896,N_5890);
or U6478 (N_6478,N_5980,N_5866);
nand U6479 (N_6479,N_5741,N_5841);
nor U6480 (N_6480,N_5780,N_5815);
nor U6481 (N_6481,N_5986,N_5975);
and U6482 (N_6482,N_5897,N_5627);
nor U6483 (N_6483,N_5809,N_5961);
and U6484 (N_6484,N_5821,N_5818);
nand U6485 (N_6485,N_5527,N_5778);
nand U6486 (N_6486,N_5697,N_5565);
nor U6487 (N_6487,N_5875,N_5507);
nand U6488 (N_6488,N_5513,N_5779);
nand U6489 (N_6489,N_5714,N_5564);
nand U6490 (N_6490,N_5708,N_5676);
xnor U6491 (N_6491,N_5514,N_5777);
nor U6492 (N_6492,N_5710,N_5860);
nand U6493 (N_6493,N_5923,N_5958);
and U6494 (N_6494,N_5876,N_5751);
xor U6495 (N_6495,N_5790,N_5826);
or U6496 (N_6496,N_5534,N_5949);
nand U6497 (N_6497,N_5672,N_5593);
nand U6498 (N_6498,N_5740,N_5849);
xnor U6499 (N_6499,N_5693,N_5608);
xor U6500 (N_6500,N_6143,N_6185);
xor U6501 (N_6501,N_6047,N_6235);
nor U6502 (N_6502,N_6425,N_6126);
xor U6503 (N_6503,N_6370,N_6402);
xnor U6504 (N_6504,N_6065,N_6009);
or U6505 (N_6505,N_6321,N_6341);
and U6506 (N_6506,N_6265,N_6045);
nor U6507 (N_6507,N_6162,N_6286);
xnor U6508 (N_6508,N_6444,N_6429);
nand U6509 (N_6509,N_6069,N_6024);
nor U6510 (N_6510,N_6379,N_6033);
xnor U6511 (N_6511,N_6175,N_6147);
xor U6512 (N_6512,N_6249,N_6075);
xnor U6513 (N_6513,N_6308,N_6112);
nand U6514 (N_6514,N_6316,N_6405);
and U6515 (N_6515,N_6046,N_6263);
xor U6516 (N_6516,N_6407,N_6160);
nor U6517 (N_6517,N_6246,N_6456);
nor U6518 (N_6518,N_6424,N_6153);
nor U6519 (N_6519,N_6278,N_6351);
or U6520 (N_6520,N_6353,N_6027);
xor U6521 (N_6521,N_6105,N_6292);
and U6522 (N_6522,N_6417,N_6089);
or U6523 (N_6523,N_6161,N_6117);
nor U6524 (N_6524,N_6433,N_6347);
nand U6525 (N_6525,N_6349,N_6420);
nand U6526 (N_6526,N_6334,N_6496);
nor U6527 (N_6527,N_6206,N_6123);
nand U6528 (N_6528,N_6179,N_6101);
and U6529 (N_6529,N_6216,N_6019);
and U6530 (N_6530,N_6231,N_6422);
or U6531 (N_6531,N_6129,N_6189);
nand U6532 (N_6532,N_6188,N_6088);
and U6533 (N_6533,N_6016,N_6022);
and U6534 (N_6534,N_6310,N_6282);
and U6535 (N_6535,N_6136,N_6066);
or U6536 (N_6536,N_6004,N_6079);
xnor U6537 (N_6537,N_6168,N_6494);
xor U6538 (N_6538,N_6318,N_6234);
xnor U6539 (N_6539,N_6176,N_6335);
nand U6540 (N_6540,N_6319,N_6317);
or U6541 (N_6541,N_6103,N_6244);
xnor U6542 (N_6542,N_6002,N_6118);
or U6543 (N_6543,N_6108,N_6042);
or U6544 (N_6544,N_6166,N_6084);
xor U6545 (N_6545,N_6455,N_6256);
nor U6546 (N_6546,N_6119,N_6459);
and U6547 (N_6547,N_6437,N_6314);
xor U6548 (N_6548,N_6289,N_6039);
xnor U6549 (N_6549,N_6177,N_6356);
xnor U6550 (N_6550,N_6350,N_6387);
xor U6551 (N_6551,N_6329,N_6109);
nor U6552 (N_6552,N_6304,N_6025);
and U6553 (N_6553,N_6354,N_6200);
or U6554 (N_6554,N_6100,N_6472);
and U6555 (N_6555,N_6184,N_6201);
and U6556 (N_6556,N_6450,N_6110);
or U6557 (N_6557,N_6464,N_6158);
or U6558 (N_6558,N_6380,N_6048);
xor U6559 (N_6559,N_6301,N_6213);
or U6560 (N_6560,N_6011,N_6017);
nand U6561 (N_6561,N_6217,N_6489);
and U6562 (N_6562,N_6107,N_6478);
nor U6563 (N_6563,N_6378,N_6159);
xor U6564 (N_6564,N_6102,N_6006);
or U6565 (N_6565,N_6373,N_6428);
nand U6566 (N_6566,N_6280,N_6365);
xnor U6567 (N_6567,N_6151,N_6195);
nand U6568 (N_6568,N_6245,N_6055);
nand U6569 (N_6569,N_6233,N_6077);
xor U6570 (N_6570,N_6348,N_6115);
and U6571 (N_6571,N_6204,N_6196);
nand U6572 (N_6572,N_6072,N_6388);
nand U6573 (N_6573,N_6332,N_6255);
and U6574 (N_6574,N_6013,N_6061);
and U6575 (N_6575,N_6164,N_6477);
nor U6576 (N_6576,N_6141,N_6412);
nor U6577 (N_6577,N_6127,N_6431);
nor U6578 (N_6578,N_6259,N_6410);
or U6579 (N_6579,N_6355,N_6393);
or U6580 (N_6580,N_6202,N_6497);
or U6581 (N_6581,N_6254,N_6165);
xnor U6582 (N_6582,N_6174,N_6030);
or U6583 (N_6583,N_6044,N_6469);
and U6584 (N_6584,N_6148,N_6205);
xnor U6585 (N_6585,N_6253,N_6029);
xor U6586 (N_6586,N_6181,N_6416);
nor U6587 (N_6587,N_6395,N_6443);
nor U6588 (N_6588,N_6376,N_6389);
xor U6589 (N_6589,N_6083,N_6482);
nand U6590 (N_6590,N_6113,N_6293);
and U6591 (N_6591,N_6071,N_6135);
and U6592 (N_6592,N_6149,N_6237);
nand U6593 (N_6593,N_6021,N_6481);
nor U6594 (N_6594,N_6359,N_6390);
and U6595 (N_6595,N_6312,N_6284);
xnor U6596 (N_6596,N_6453,N_6190);
nor U6597 (N_6597,N_6418,N_6173);
nor U6598 (N_6598,N_6197,N_6493);
nor U6599 (N_6599,N_6228,N_6054);
xnor U6600 (N_6600,N_6441,N_6068);
nand U6601 (N_6601,N_6210,N_6404);
xor U6602 (N_6602,N_6330,N_6276);
and U6603 (N_6603,N_6480,N_6302);
or U6604 (N_6604,N_6183,N_6303);
nor U6605 (N_6605,N_6252,N_6260);
nand U6606 (N_6606,N_6266,N_6096);
nor U6607 (N_6607,N_6250,N_6134);
nand U6608 (N_6608,N_6460,N_6451);
and U6609 (N_6609,N_6313,N_6471);
and U6610 (N_6610,N_6005,N_6169);
and U6611 (N_6611,N_6426,N_6050);
xnor U6612 (N_6612,N_6095,N_6081);
nor U6613 (N_6613,N_6311,N_6458);
nor U6614 (N_6614,N_6466,N_6020);
nor U6615 (N_6615,N_6251,N_6218);
and U6616 (N_6616,N_6333,N_6297);
nor U6617 (N_6617,N_6399,N_6093);
xnor U6618 (N_6618,N_6036,N_6034);
xnor U6619 (N_6619,N_6120,N_6327);
nor U6620 (N_6620,N_6128,N_6492);
or U6621 (N_6621,N_6080,N_6230);
nand U6622 (N_6622,N_6275,N_6248);
or U6623 (N_6623,N_6085,N_6012);
or U6624 (N_6624,N_6461,N_6099);
nor U6625 (N_6625,N_6485,N_6475);
nand U6626 (N_6626,N_6074,N_6130);
and U6627 (N_6627,N_6104,N_6467);
and U6628 (N_6628,N_6242,N_6106);
nand U6629 (N_6629,N_6452,N_6375);
xnor U6630 (N_6630,N_6357,N_6053);
xnor U6631 (N_6631,N_6076,N_6434);
and U6632 (N_6632,N_6091,N_6421);
nor U6633 (N_6633,N_6191,N_6155);
or U6634 (N_6634,N_6374,N_6232);
nor U6635 (N_6635,N_6163,N_6447);
xor U6636 (N_6636,N_6137,N_6215);
or U6637 (N_6637,N_6057,N_6345);
and U6638 (N_6638,N_6052,N_6131);
nor U6639 (N_6639,N_6346,N_6331);
nor U6640 (N_6640,N_6470,N_6037);
and U6641 (N_6641,N_6290,N_6269);
or U6642 (N_6642,N_6325,N_6145);
nand U6643 (N_6643,N_6299,N_6384);
nor U6644 (N_6644,N_6491,N_6396);
or U6645 (N_6645,N_6032,N_6221);
nor U6646 (N_6646,N_6010,N_6398);
nand U6647 (N_6647,N_6454,N_6211);
xor U6648 (N_6648,N_6473,N_6000);
or U6649 (N_6649,N_6171,N_6440);
xnor U6650 (N_6650,N_6257,N_6474);
nor U6651 (N_6651,N_6003,N_6015);
nor U6652 (N_6652,N_6360,N_6060);
nand U6653 (N_6653,N_6063,N_6427);
nor U6654 (N_6654,N_6328,N_6111);
or U6655 (N_6655,N_6187,N_6008);
xnor U6656 (N_6656,N_6490,N_6320);
or U6657 (N_6657,N_6182,N_6144);
nand U6658 (N_6658,N_6170,N_6307);
or U6659 (N_6659,N_6476,N_6340);
xor U6660 (N_6660,N_6116,N_6309);
xor U6661 (N_6661,N_6086,N_6371);
xor U6662 (N_6662,N_6457,N_6383);
and U6663 (N_6663,N_6018,N_6436);
nand U6664 (N_6664,N_6062,N_6058);
or U6665 (N_6665,N_6367,N_6363);
nand U6666 (N_6666,N_6400,N_6180);
and U6667 (N_6667,N_6090,N_6368);
and U6668 (N_6668,N_6358,N_6059);
nand U6669 (N_6669,N_6121,N_6445);
or U6670 (N_6670,N_6446,N_6487);
nand U6671 (N_6671,N_6392,N_6300);
or U6672 (N_6672,N_6031,N_6465);
and U6673 (N_6673,N_6291,N_6337);
and U6674 (N_6674,N_6463,N_6192);
and U6675 (N_6675,N_6157,N_6040);
xnor U6676 (N_6676,N_6122,N_6271);
nand U6677 (N_6677,N_6222,N_6391);
and U6678 (N_6678,N_6414,N_6369);
nand U6679 (N_6679,N_6468,N_6070);
and U6680 (N_6680,N_6236,N_6268);
nor U6681 (N_6681,N_6067,N_6411);
or U6682 (N_6682,N_6423,N_6140);
and U6683 (N_6683,N_6274,N_6406);
or U6684 (N_6684,N_6295,N_6339);
and U6685 (N_6685,N_6324,N_6486);
xnor U6686 (N_6686,N_6078,N_6167);
and U6687 (N_6687,N_6056,N_6064);
nand U6688 (N_6688,N_6285,N_6092);
and U6689 (N_6689,N_6362,N_6098);
or U6690 (N_6690,N_6133,N_6483);
nor U6691 (N_6691,N_6156,N_6146);
nand U6692 (N_6692,N_6343,N_6223);
xor U6693 (N_6693,N_6366,N_6270);
or U6694 (N_6694,N_6209,N_6364);
xor U6695 (N_6695,N_6142,N_6479);
nor U6696 (N_6696,N_6124,N_6051);
or U6697 (N_6697,N_6279,N_6336);
xnor U6698 (N_6698,N_6305,N_6227);
and U6699 (N_6699,N_6306,N_6262);
or U6700 (N_6700,N_6342,N_6198);
or U6701 (N_6701,N_6413,N_6240);
nor U6702 (N_6702,N_6484,N_6462);
or U6703 (N_6703,N_6401,N_6041);
nand U6704 (N_6704,N_6283,N_6220);
nor U6705 (N_6705,N_6243,N_6229);
nand U6706 (N_6706,N_6043,N_6322);
nor U6707 (N_6707,N_6132,N_6495);
xnor U6708 (N_6708,N_6023,N_6372);
nand U6709 (N_6709,N_6326,N_6225);
nor U6710 (N_6710,N_6439,N_6403);
or U6711 (N_6711,N_6415,N_6087);
and U6712 (N_6712,N_6224,N_6408);
and U6713 (N_6713,N_6203,N_6386);
nand U6714 (N_6714,N_6381,N_6498);
nor U6715 (N_6715,N_6296,N_6352);
and U6716 (N_6716,N_6172,N_6409);
or U6717 (N_6717,N_6035,N_6344);
and U6718 (N_6718,N_6448,N_6219);
nor U6719 (N_6719,N_6226,N_6432);
and U6720 (N_6720,N_6264,N_6287);
or U6721 (N_6721,N_6323,N_6014);
nor U6722 (N_6722,N_6488,N_6247);
xnor U6723 (N_6723,N_6267,N_6338);
and U6724 (N_6724,N_6208,N_6207);
nor U6725 (N_6725,N_6212,N_6150);
xor U6726 (N_6726,N_6007,N_6385);
and U6727 (N_6727,N_6097,N_6154);
nand U6728 (N_6728,N_6214,N_6001);
nand U6729 (N_6729,N_6435,N_6186);
nand U6730 (N_6730,N_6377,N_6049);
nor U6731 (N_6731,N_6382,N_6294);
nor U6732 (N_6732,N_6193,N_6438);
xnor U6733 (N_6733,N_6449,N_6194);
xor U6734 (N_6734,N_6125,N_6397);
nand U6735 (N_6735,N_6239,N_6238);
or U6736 (N_6736,N_6419,N_6288);
or U6737 (N_6737,N_6273,N_6298);
nor U6738 (N_6738,N_6026,N_6199);
nor U6739 (N_6739,N_6442,N_6082);
or U6740 (N_6740,N_6094,N_6178);
nor U6741 (N_6741,N_6361,N_6114);
nor U6742 (N_6742,N_6138,N_6499);
and U6743 (N_6743,N_6430,N_6315);
or U6744 (N_6744,N_6272,N_6139);
and U6745 (N_6745,N_6038,N_6152);
nor U6746 (N_6746,N_6241,N_6073);
xnor U6747 (N_6747,N_6277,N_6258);
or U6748 (N_6748,N_6281,N_6394);
nor U6749 (N_6749,N_6261,N_6028);
or U6750 (N_6750,N_6090,N_6466);
nor U6751 (N_6751,N_6438,N_6437);
or U6752 (N_6752,N_6291,N_6260);
nor U6753 (N_6753,N_6192,N_6362);
nor U6754 (N_6754,N_6348,N_6036);
and U6755 (N_6755,N_6443,N_6422);
and U6756 (N_6756,N_6216,N_6249);
xor U6757 (N_6757,N_6075,N_6032);
nand U6758 (N_6758,N_6093,N_6173);
and U6759 (N_6759,N_6490,N_6499);
xor U6760 (N_6760,N_6224,N_6498);
nand U6761 (N_6761,N_6216,N_6115);
xnor U6762 (N_6762,N_6353,N_6382);
or U6763 (N_6763,N_6008,N_6359);
and U6764 (N_6764,N_6160,N_6040);
and U6765 (N_6765,N_6434,N_6373);
nand U6766 (N_6766,N_6137,N_6020);
nand U6767 (N_6767,N_6435,N_6437);
xnor U6768 (N_6768,N_6025,N_6133);
or U6769 (N_6769,N_6042,N_6073);
and U6770 (N_6770,N_6244,N_6442);
nor U6771 (N_6771,N_6295,N_6358);
xor U6772 (N_6772,N_6233,N_6146);
xor U6773 (N_6773,N_6066,N_6196);
nor U6774 (N_6774,N_6110,N_6093);
nand U6775 (N_6775,N_6079,N_6116);
xor U6776 (N_6776,N_6196,N_6389);
nand U6777 (N_6777,N_6299,N_6469);
nor U6778 (N_6778,N_6322,N_6479);
or U6779 (N_6779,N_6036,N_6309);
and U6780 (N_6780,N_6279,N_6120);
or U6781 (N_6781,N_6209,N_6010);
xnor U6782 (N_6782,N_6274,N_6122);
nand U6783 (N_6783,N_6142,N_6259);
or U6784 (N_6784,N_6359,N_6469);
or U6785 (N_6785,N_6368,N_6013);
and U6786 (N_6786,N_6071,N_6173);
xor U6787 (N_6787,N_6050,N_6171);
or U6788 (N_6788,N_6246,N_6425);
or U6789 (N_6789,N_6214,N_6120);
nor U6790 (N_6790,N_6113,N_6407);
xnor U6791 (N_6791,N_6474,N_6060);
xnor U6792 (N_6792,N_6138,N_6127);
xor U6793 (N_6793,N_6469,N_6342);
xor U6794 (N_6794,N_6324,N_6069);
and U6795 (N_6795,N_6257,N_6100);
nand U6796 (N_6796,N_6092,N_6416);
nand U6797 (N_6797,N_6220,N_6030);
nand U6798 (N_6798,N_6274,N_6232);
or U6799 (N_6799,N_6333,N_6437);
and U6800 (N_6800,N_6468,N_6339);
xnor U6801 (N_6801,N_6106,N_6415);
xor U6802 (N_6802,N_6145,N_6258);
nand U6803 (N_6803,N_6063,N_6470);
and U6804 (N_6804,N_6406,N_6059);
nand U6805 (N_6805,N_6344,N_6374);
nand U6806 (N_6806,N_6456,N_6431);
nor U6807 (N_6807,N_6054,N_6289);
xnor U6808 (N_6808,N_6304,N_6409);
or U6809 (N_6809,N_6212,N_6077);
nand U6810 (N_6810,N_6168,N_6039);
nand U6811 (N_6811,N_6080,N_6414);
and U6812 (N_6812,N_6141,N_6088);
xnor U6813 (N_6813,N_6389,N_6343);
or U6814 (N_6814,N_6255,N_6046);
nor U6815 (N_6815,N_6359,N_6143);
or U6816 (N_6816,N_6164,N_6064);
and U6817 (N_6817,N_6080,N_6077);
xnor U6818 (N_6818,N_6254,N_6072);
or U6819 (N_6819,N_6169,N_6237);
xor U6820 (N_6820,N_6128,N_6424);
and U6821 (N_6821,N_6124,N_6214);
xor U6822 (N_6822,N_6054,N_6306);
nor U6823 (N_6823,N_6054,N_6127);
nand U6824 (N_6824,N_6472,N_6300);
or U6825 (N_6825,N_6347,N_6081);
nor U6826 (N_6826,N_6295,N_6269);
nand U6827 (N_6827,N_6266,N_6360);
nor U6828 (N_6828,N_6125,N_6020);
and U6829 (N_6829,N_6108,N_6278);
nor U6830 (N_6830,N_6443,N_6446);
xor U6831 (N_6831,N_6091,N_6349);
nor U6832 (N_6832,N_6384,N_6050);
xor U6833 (N_6833,N_6439,N_6384);
nand U6834 (N_6834,N_6423,N_6125);
or U6835 (N_6835,N_6073,N_6499);
nand U6836 (N_6836,N_6294,N_6283);
and U6837 (N_6837,N_6337,N_6219);
or U6838 (N_6838,N_6250,N_6329);
or U6839 (N_6839,N_6175,N_6067);
and U6840 (N_6840,N_6181,N_6115);
xor U6841 (N_6841,N_6323,N_6210);
nor U6842 (N_6842,N_6225,N_6204);
xnor U6843 (N_6843,N_6418,N_6402);
xnor U6844 (N_6844,N_6197,N_6464);
xor U6845 (N_6845,N_6209,N_6121);
xnor U6846 (N_6846,N_6089,N_6266);
nand U6847 (N_6847,N_6157,N_6150);
xnor U6848 (N_6848,N_6123,N_6467);
and U6849 (N_6849,N_6362,N_6443);
xnor U6850 (N_6850,N_6266,N_6441);
nand U6851 (N_6851,N_6085,N_6402);
and U6852 (N_6852,N_6207,N_6292);
or U6853 (N_6853,N_6111,N_6082);
nand U6854 (N_6854,N_6391,N_6408);
xor U6855 (N_6855,N_6256,N_6236);
nand U6856 (N_6856,N_6238,N_6138);
nand U6857 (N_6857,N_6372,N_6274);
or U6858 (N_6858,N_6058,N_6007);
or U6859 (N_6859,N_6023,N_6435);
nor U6860 (N_6860,N_6150,N_6092);
or U6861 (N_6861,N_6351,N_6465);
nor U6862 (N_6862,N_6495,N_6464);
nor U6863 (N_6863,N_6112,N_6492);
or U6864 (N_6864,N_6195,N_6074);
nand U6865 (N_6865,N_6444,N_6155);
or U6866 (N_6866,N_6069,N_6385);
nand U6867 (N_6867,N_6058,N_6173);
and U6868 (N_6868,N_6094,N_6228);
or U6869 (N_6869,N_6158,N_6304);
nand U6870 (N_6870,N_6321,N_6473);
nor U6871 (N_6871,N_6353,N_6030);
xor U6872 (N_6872,N_6120,N_6243);
nand U6873 (N_6873,N_6204,N_6442);
and U6874 (N_6874,N_6198,N_6137);
and U6875 (N_6875,N_6294,N_6481);
nand U6876 (N_6876,N_6223,N_6095);
and U6877 (N_6877,N_6382,N_6213);
and U6878 (N_6878,N_6274,N_6082);
nor U6879 (N_6879,N_6028,N_6181);
and U6880 (N_6880,N_6338,N_6039);
xnor U6881 (N_6881,N_6086,N_6497);
or U6882 (N_6882,N_6244,N_6092);
nand U6883 (N_6883,N_6400,N_6402);
nor U6884 (N_6884,N_6018,N_6151);
and U6885 (N_6885,N_6262,N_6071);
nor U6886 (N_6886,N_6250,N_6083);
or U6887 (N_6887,N_6021,N_6043);
or U6888 (N_6888,N_6291,N_6107);
nand U6889 (N_6889,N_6320,N_6204);
nand U6890 (N_6890,N_6474,N_6092);
or U6891 (N_6891,N_6405,N_6452);
and U6892 (N_6892,N_6192,N_6290);
xnor U6893 (N_6893,N_6291,N_6497);
and U6894 (N_6894,N_6056,N_6347);
and U6895 (N_6895,N_6027,N_6101);
and U6896 (N_6896,N_6247,N_6177);
nor U6897 (N_6897,N_6168,N_6024);
or U6898 (N_6898,N_6025,N_6212);
and U6899 (N_6899,N_6493,N_6105);
nand U6900 (N_6900,N_6278,N_6223);
or U6901 (N_6901,N_6189,N_6073);
nor U6902 (N_6902,N_6415,N_6025);
and U6903 (N_6903,N_6263,N_6217);
nand U6904 (N_6904,N_6369,N_6372);
and U6905 (N_6905,N_6211,N_6448);
or U6906 (N_6906,N_6336,N_6226);
nor U6907 (N_6907,N_6065,N_6043);
xnor U6908 (N_6908,N_6265,N_6247);
xnor U6909 (N_6909,N_6479,N_6260);
nand U6910 (N_6910,N_6484,N_6387);
or U6911 (N_6911,N_6325,N_6388);
xnor U6912 (N_6912,N_6154,N_6063);
nand U6913 (N_6913,N_6416,N_6378);
and U6914 (N_6914,N_6254,N_6060);
nor U6915 (N_6915,N_6492,N_6324);
or U6916 (N_6916,N_6326,N_6157);
nand U6917 (N_6917,N_6488,N_6400);
nor U6918 (N_6918,N_6418,N_6082);
and U6919 (N_6919,N_6486,N_6297);
nor U6920 (N_6920,N_6240,N_6070);
nor U6921 (N_6921,N_6057,N_6389);
xnor U6922 (N_6922,N_6332,N_6442);
and U6923 (N_6923,N_6495,N_6126);
xor U6924 (N_6924,N_6064,N_6068);
nor U6925 (N_6925,N_6402,N_6432);
xor U6926 (N_6926,N_6160,N_6438);
xor U6927 (N_6927,N_6421,N_6061);
and U6928 (N_6928,N_6489,N_6248);
xnor U6929 (N_6929,N_6054,N_6245);
xnor U6930 (N_6930,N_6238,N_6333);
and U6931 (N_6931,N_6266,N_6477);
and U6932 (N_6932,N_6117,N_6095);
xnor U6933 (N_6933,N_6386,N_6146);
nand U6934 (N_6934,N_6144,N_6068);
nand U6935 (N_6935,N_6092,N_6403);
nor U6936 (N_6936,N_6346,N_6315);
xor U6937 (N_6937,N_6457,N_6191);
and U6938 (N_6938,N_6252,N_6483);
nor U6939 (N_6939,N_6104,N_6431);
or U6940 (N_6940,N_6082,N_6499);
nor U6941 (N_6941,N_6171,N_6405);
and U6942 (N_6942,N_6276,N_6386);
nor U6943 (N_6943,N_6023,N_6262);
nor U6944 (N_6944,N_6240,N_6407);
nand U6945 (N_6945,N_6092,N_6007);
nand U6946 (N_6946,N_6016,N_6212);
and U6947 (N_6947,N_6308,N_6472);
nand U6948 (N_6948,N_6003,N_6005);
xor U6949 (N_6949,N_6467,N_6000);
or U6950 (N_6950,N_6463,N_6065);
nand U6951 (N_6951,N_6220,N_6451);
nor U6952 (N_6952,N_6296,N_6414);
nor U6953 (N_6953,N_6160,N_6228);
and U6954 (N_6954,N_6028,N_6468);
and U6955 (N_6955,N_6488,N_6187);
xor U6956 (N_6956,N_6053,N_6268);
nor U6957 (N_6957,N_6446,N_6058);
nor U6958 (N_6958,N_6205,N_6197);
nand U6959 (N_6959,N_6379,N_6167);
nand U6960 (N_6960,N_6435,N_6045);
xnor U6961 (N_6961,N_6059,N_6335);
or U6962 (N_6962,N_6033,N_6266);
nand U6963 (N_6963,N_6432,N_6388);
nand U6964 (N_6964,N_6387,N_6278);
nand U6965 (N_6965,N_6292,N_6342);
nor U6966 (N_6966,N_6437,N_6421);
and U6967 (N_6967,N_6273,N_6093);
xnor U6968 (N_6968,N_6252,N_6111);
and U6969 (N_6969,N_6113,N_6415);
nor U6970 (N_6970,N_6329,N_6309);
and U6971 (N_6971,N_6493,N_6470);
nand U6972 (N_6972,N_6393,N_6378);
xor U6973 (N_6973,N_6134,N_6494);
or U6974 (N_6974,N_6095,N_6004);
and U6975 (N_6975,N_6462,N_6089);
xnor U6976 (N_6976,N_6164,N_6342);
nand U6977 (N_6977,N_6367,N_6143);
nor U6978 (N_6978,N_6342,N_6485);
and U6979 (N_6979,N_6253,N_6116);
xnor U6980 (N_6980,N_6409,N_6040);
nor U6981 (N_6981,N_6462,N_6239);
nand U6982 (N_6982,N_6478,N_6032);
xor U6983 (N_6983,N_6143,N_6235);
or U6984 (N_6984,N_6278,N_6397);
nand U6985 (N_6985,N_6476,N_6101);
or U6986 (N_6986,N_6271,N_6408);
xnor U6987 (N_6987,N_6386,N_6234);
or U6988 (N_6988,N_6402,N_6094);
and U6989 (N_6989,N_6410,N_6217);
or U6990 (N_6990,N_6268,N_6492);
and U6991 (N_6991,N_6296,N_6496);
and U6992 (N_6992,N_6164,N_6321);
and U6993 (N_6993,N_6488,N_6418);
and U6994 (N_6994,N_6036,N_6149);
and U6995 (N_6995,N_6441,N_6418);
or U6996 (N_6996,N_6463,N_6284);
or U6997 (N_6997,N_6428,N_6322);
xnor U6998 (N_6998,N_6026,N_6044);
nor U6999 (N_6999,N_6461,N_6396);
and U7000 (N_7000,N_6937,N_6595);
and U7001 (N_7001,N_6500,N_6577);
and U7002 (N_7002,N_6603,N_6985);
nand U7003 (N_7003,N_6829,N_6510);
and U7004 (N_7004,N_6888,N_6569);
and U7005 (N_7005,N_6855,N_6667);
and U7006 (N_7006,N_6934,N_6687);
xor U7007 (N_7007,N_6781,N_6601);
and U7008 (N_7008,N_6862,N_6796);
nor U7009 (N_7009,N_6597,N_6815);
nand U7010 (N_7010,N_6795,N_6693);
xor U7011 (N_7011,N_6915,N_6988);
xor U7012 (N_7012,N_6555,N_6733);
xnor U7013 (N_7013,N_6546,N_6877);
xnor U7014 (N_7014,N_6843,N_6907);
and U7015 (N_7015,N_6557,N_6686);
and U7016 (N_7016,N_6953,N_6997);
nor U7017 (N_7017,N_6732,N_6870);
nor U7018 (N_7018,N_6755,N_6673);
and U7019 (N_7019,N_6926,N_6731);
and U7020 (N_7020,N_6632,N_6730);
or U7021 (N_7021,N_6824,N_6628);
or U7022 (N_7022,N_6668,N_6900);
xnor U7023 (N_7023,N_6548,N_6854);
or U7024 (N_7024,N_6952,N_6778);
nand U7025 (N_7025,N_6891,N_6702);
and U7026 (N_7026,N_6852,N_6990);
xnor U7027 (N_7027,N_6684,N_6503);
and U7028 (N_7028,N_6991,N_6951);
or U7029 (N_7029,N_6660,N_6764);
nand U7030 (N_7030,N_6680,N_6513);
xor U7031 (N_7031,N_6580,N_6901);
nor U7032 (N_7032,N_6780,N_6699);
or U7033 (N_7033,N_6771,N_6588);
and U7034 (N_7034,N_6689,N_6960);
nor U7035 (N_7035,N_6909,N_6665);
nand U7036 (N_7036,N_6656,N_6972);
nor U7037 (N_7037,N_6512,N_6837);
nor U7038 (N_7038,N_6842,N_6627);
and U7039 (N_7039,N_6658,N_6703);
and U7040 (N_7040,N_6614,N_6986);
and U7041 (N_7041,N_6899,N_6898);
xnor U7042 (N_7042,N_6941,N_6695);
and U7043 (N_7043,N_6596,N_6633);
nand U7044 (N_7044,N_6841,N_6762);
and U7045 (N_7045,N_6599,N_6681);
and U7046 (N_7046,N_6607,N_6685);
or U7047 (N_7047,N_6549,N_6919);
and U7048 (N_7048,N_6757,N_6938);
xor U7049 (N_7049,N_6650,N_6920);
nor U7050 (N_7050,N_6818,N_6825);
nand U7051 (N_7051,N_6823,N_6609);
xor U7052 (N_7052,N_6790,N_6871);
nand U7053 (N_7053,N_6657,N_6638);
and U7054 (N_7054,N_6677,N_6947);
nand U7055 (N_7055,N_6690,N_6783);
nor U7056 (N_7056,N_6949,N_6616);
nand U7057 (N_7057,N_6749,N_6848);
nor U7058 (N_7058,N_6501,N_6956);
nand U7059 (N_7059,N_6563,N_6922);
nand U7060 (N_7060,N_6845,N_6706);
xnor U7061 (N_7061,N_6648,N_6736);
or U7062 (N_7062,N_6530,N_6725);
or U7063 (N_7063,N_6674,N_6911);
or U7064 (N_7064,N_6808,N_6866);
and U7065 (N_7065,N_6525,N_6805);
nand U7066 (N_7066,N_6821,N_6679);
or U7067 (N_7067,N_6968,N_6923);
nand U7068 (N_7068,N_6618,N_6751);
and U7069 (N_7069,N_6675,N_6758);
or U7070 (N_7070,N_6741,N_6789);
nand U7071 (N_7071,N_6539,N_6662);
nand U7072 (N_7072,N_6545,N_6881);
xnor U7073 (N_7073,N_6728,N_6630);
nand U7074 (N_7074,N_6720,N_6570);
nor U7075 (N_7075,N_6582,N_6860);
nor U7076 (N_7076,N_6943,N_6816);
nand U7077 (N_7077,N_6586,N_6645);
or U7078 (N_7078,N_6567,N_6715);
nor U7079 (N_7079,N_6777,N_6939);
xor U7080 (N_7080,N_6566,N_6772);
xnor U7081 (N_7081,N_6664,N_6998);
xor U7082 (N_7082,N_6869,N_6791);
nor U7083 (N_7083,N_6520,N_6640);
and U7084 (N_7084,N_6857,N_6587);
xor U7085 (N_7085,N_6739,N_6814);
nand U7086 (N_7086,N_6526,N_6559);
or U7087 (N_7087,N_6773,N_6834);
and U7088 (N_7088,N_6697,N_6621);
nor U7089 (N_7089,N_6910,N_6813);
xor U7090 (N_7090,N_6999,N_6885);
or U7091 (N_7091,N_6593,N_6889);
and U7092 (N_7092,N_6971,N_6615);
nand U7093 (N_7093,N_6847,N_6692);
nor U7094 (N_7094,N_6827,N_6917);
and U7095 (N_7095,N_6625,N_6647);
or U7096 (N_7096,N_6722,N_6637);
xnor U7097 (N_7097,N_6565,N_6529);
xor U7098 (N_7098,N_6552,N_6895);
or U7099 (N_7099,N_6718,N_6806);
nand U7100 (N_7100,N_6849,N_6760);
nor U7101 (N_7101,N_6636,N_6822);
and U7102 (N_7102,N_6994,N_6613);
or U7103 (N_7103,N_6708,N_6654);
and U7104 (N_7104,N_6634,N_6787);
and U7105 (N_7105,N_6989,N_6942);
nand U7106 (N_7106,N_6519,N_6832);
or U7107 (N_7107,N_6554,N_6629);
and U7108 (N_7108,N_6876,N_6502);
or U7109 (N_7109,N_6584,N_6624);
nand U7110 (N_7110,N_6717,N_6756);
or U7111 (N_7111,N_6768,N_6535);
and U7112 (N_7112,N_6882,N_6556);
and U7113 (N_7113,N_6913,N_6562);
nor U7114 (N_7114,N_6663,N_6819);
or U7115 (N_7115,N_6826,N_6518);
nor U7116 (N_7116,N_6831,N_6779);
nor U7117 (N_7117,N_6817,N_6746);
xnor U7118 (N_7118,N_6859,N_6537);
nor U7119 (N_7119,N_6868,N_6788);
or U7120 (N_7120,N_6969,N_6880);
nand U7121 (N_7121,N_6523,N_6966);
xor U7122 (N_7122,N_6924,N_6948);
or U7123 (N_7123,N_6564,N_6793);
nor U7124 (N_7124,N_6710,N_6765);
or U7125 (N_7125,N_6521,N_6631);
and U7126 (N_7126,N_6867,N_6887);
and U7127 (N_7127,N_6622,N_6669);
nor U7128 (N_7128,N_6700,N_6950);
nand U7129 (N_7129,N_6786,N_6661);
xor U7130 (N_7130,N_6916,N_6602);
xnor U7131 (N_7131,N_6527,N_6550);
or U7132 (N_7132,N_6861,N_6707);
nand U7133 (N_7133,N_6716,N_6612);
nor U7134 (N_7134,N_6863,N_6709);
and U7135 (N_7135,N_6833,N_6811);
nand U7136 (N_7136,N_6522,N_6610);
nor U7137 (N_7137,N_6646,N_6740);
nor U7138 (N_7138,N_6914,N_6879);
and U7139 (N_7139,N_6865,N_6704);
nand U7140 (N_7140,N_6711,N_6802);
nor U7141 (N_7141,N_6551,N_6835);
xor U7142 (N_7142,N_6878,N_6642);
and U7143 (N_7143,N_6921,N_6698);
or U7144 (N_7144,N_6723,N_6608);
nand U7145 (N_7145,N_6536,N_6678);
or U7146 (N_7146,N_6846,N_6604);
nor U7147 (N_7147,N_6970,N_6932);
or U7148 (N_7148,N_6931,N_6828);
nor U7149 (N_7149,N_6524,N_6744);
xor U7150 (N_7150,N_6830,N_6903);
nand U7151 (N_7151,N_6944,N_6724);
nand U7152 (N_7152,N_6683,N_6605);
nand U7153 (N_7153,N_6585,N_6694);
and U7154 (N_7154,N_6886,N_6511);
nand U7155 (N_7155,N_6558,N_6649);
or U7156 (N_7156,N_6544,N_6721);
and U7157 (N_7157,N_6590,N_6547);
and U7158 (N_7158,N_6873,N_6505);
xor U7159 (N_7159,N_6714,N_6935);
nor U7160 (N_7160,N_6965,N_6560);
nand U7161 (N_7161,N_6600,N_6753);
or U7162 (N_7162,N_6531,N_6574);
and U7163 (N_7163,N_6961,N_6517);
or U7164 (N_7164,N_6713,N_6639);
or U7165 (N_7165,N_6872,N_6810);
xnor U7166 (N_7166,N_6928,N_6927);
or U7167 (N_7167,N_6620,N_6853);
or U7168 (N_7168,N_6712,N_6532);
nor U7169 (N_7169,N_6743,N_6807);
and U7170 (N_7170,N_6992,N_6884);
xnor U7171 (N_7171,N_6874,N_6946);
nand U7172 (N_7172,N_6973,N_6809);
and U7173 (N_7173,N_6995,N_6775);
and U7174 (N_7174,N_6666,N_6509);
nand U7175 (N_7175,N_6897,N_6643);
and U7176 (N_7176,N_6672,N_6984);
xnor U7177 (N_7177,N_6504,N_6906);
nor U7178 (N_7178,N_6575,N_6987);
xnor U7179 (N_7179,N_6726,N_6967);
or U7180 (N_7180,N_6528,N_6896);
xnor U7181 (N_7181,N_6737,N_6974);
nor U7182 (N_7182,N_6800,N_6976);
nor U7183 (N_7183,N_6594,N_6626);
or U7184 (N_7184,N_6571,N_6515);
xnor U7185 (N_7185,N_6635,N_6671);
nand U7186 (N_7186,N_6576,N_6676);
and U7187 (N_7187,N_6641,N_6890);
or U7188 (N_7188,N_6670,N_6553);
xor U7189 (N_7189,N_6804,N_6691);
xnor U7190 (N_7190,N_6836,N_6918);
or U7191 (N_7191,N_6975,N_6514);
nand U7192 (N_7192,N_6792,N_6623);
or U7193 (N_7193,N_6581,N_6912);
or U7194 (N_7194,N_6981,N_6840);
nand U7195 (N_7195,N_6682,N_6782);
nand U7196 (N_7196,N_6930,N_6894);
nand U7197 (N_7197,N_6606,N_6902);
or U7198 (N_7198,N_6750,N_6655);
or U7199 (N_7199,N_6534,N_6591);
xnor U7200 (N_7200,N_6747,N_6541);
and U7201 (N_7201,N_6644,N_6839);
xor U7202 (N_7202,N_6738,N_6977);
nor U7203 (N_7203,N_6980,N_6933);
nand U7204 (N_7204,N_6893,N_6929);
nor U7205 (N_7205,N_6763,N_6583);
nor U7206 (N_7206,N_6652,N_6651);
or U7207 (N_7207,N_6617,N_6908);
and U7208 (N_7208,N_6940,N_6957);
xor U7209 (N_7209,N_6838,N_6696);
and U7210 (N_7210,N_6752,N_6543);
xnor U7211 (N_7211,N_6729,N_6759);
or U7212 (N_7212,N_6905,N_6844);
or U7213 (N_7213,N_6785,N_6542);
xnor U7214 (N_7214,N_6979,N_6540);
and U7215 (N_7215,N_6799,N_6801);
xnor U7216 (N_7216,N_6761,N_6561);
and U7217 (N_7217,N_6516,N_6573);
nor U7218 (N_7218,N_6767,N_6572);
xor U7219 (N_7219,N_6996,N_6820);
or U7220 (N_7220,N_6533,N_6892);
or U7221 (N_7221,N_6803,N_6856);
nor U7222 (N_7222,N_6982,N_6945);
nor U7223 (N_7223,N_6579,N_6776);
nor U7224 (N_7224,N_6954,N_6993);
nor U7225 (N_7225,N_6745,N_6904);
and U7226 (N_7226,N_6719,N_6688);
and U7227 (N_7227,N_6592,N_6705);
xnor U7228 (N_7228,N_6589,N_6812);
nor U7229 (N_7229,N_6851,N_6797);
and U7230 (N_7230,N_6766,N_6925);
xnor U7231 (N_7231,N_6794,N_6875);
nand U7232 (N_7232,N_6955,N_6963);
nor U7233 (N_7233,N_6754,N_6735);
xor U7234 (N_7234,N_6883,N_6611);
nor U7235 (N_7235,N_6619,N_6769);
and U7236 (N_7236,N_6727,N_6568);
nand U7237 (N_7237,N_6701,N_6983);
nor U7238 (N_7238,N_6748,N_6506);
xnor U7239 (N_7239,N_6958,N_6962);
or U7240 (N_7240,N_6864,N_6508);
and U7241 (N_7241,N_6798,N_6659);
nor U7242 (N_7242,N_6653,N_6742);
nor U7243 (N_7243,N_6936,N_6774);
or U7244 (N_7244,N_6598,N_6959);
nand U7245 (N_7245,N_6734,N_6964);
xor U7246 (N_7246,N_6858,N_6578);
xor U7247 (N_7247,N_6978,N_6507);
nand U7248 (N_7248,N_6850,N_6538);
nor U7249 (N_7249,N_6784,N_6770);
nor U7250 (N_7250,N_6989,N_6507);
or U7251 (N_7251,N_6926,N_6996);
nor U7252 (N_7252,N_6883,N_6872);
xor U7253 (N_7253,N_6803,N_6698);
nand U7254 (N_7254,N_6775,N_6910);
and U7255 (N_7255,N_6886,N_6866);
nor U7256 (N_7256,N_6955,N_6827);
nand U7257 (N_7257,N_6806,N_6886);
or U7258 (N_7258,N_6554,N_6644);
nand U7259 (N_7259,N_6974,N_6556);
or U7260 (N_7260,N_6536,N_6693);
nand U7261 (N_7261,N_6689,N_6979);
nor U7262 (N_7262,N_6909,N_6574);
or U7263 (N_7263,N_6725,N_6695);
nand U7264 (N_7264,N_6740,N_6828);
and U7265 (N_7265,N_6872,N_6845);
and U7266 (N_7266,N_6682,N_6571);
nand U7267 (N_7267,N_6822,N_6891);
and U7268 (N_7268,N_6519,N_6587);
and U7269 (N_7269,N_6500,N_6835);
xor U7270 (N_7270,N_6927,N_6655);
and U7271 (N_7271,N_6768,N_6620);
xor U7272 (N_7272,N_6745,N_6628);
or U7273 (N_7273,N_6660,N_6819);
and U7274 (N_7274,N_6850,N_6653);
nor U7275 (N_7275,N_6924,N_6940);
or U7276 (N_7276,N_6980,N_6679);
or U7277 (N_7277,N_6650,N_6761);
or U7278 (N_7278,N_6657,N_6958);
or U7279 (N_7279,N_6914,N_6503);
nand U7280 (N_7280,N_6761,N_6604);
or U7281 (N_7281,N_6818,N_6732);
nor U7282 (N_7282,N_6634,N_6949);
or U7283 (N_7283,N_6635,N_6611);
nand U7284 (N_7284,N_6676,N_6786);
nor U7285 (N_7285,N_6697,N_6928);
nand U7286 (N_7286,N_6841,N_6623);
xnor U7287 (N_7287,N_6964,N_6710);
or U7288 (N_7288,N_6506,N_6556);
xnor U7289 (N_7289,N_6620,N_6539);
and U7290 (N_7290,N_6537,N_6781);
nor U7291 (N_7291,N_6798,N_6997);
or U7292 (N_7292,N_6546,N_6651);
or U7293 (N_7293,N_6704,N_6631);
and U7294 (N_7294,N_6842,N_6909);
nand U7295 (N_7295,N_6756,N_6850);
or U7296 (N_7296,N_6936,N_6569);
xor U7297 (N_7297,N_6718,N_6708);
or U7298 (N_7298,N_6636,N_6922);
nor U7299 (N_7299,N_6920,N_6677);
or U7300 (N_7300,N_6900,N_6553);
nand U7301 (N_7301,N_6688,N_6964);
or U7302 (N_7302,N_6515,N_6913);
nand U7303 (N_7303,N_6959,N_6621);
nand U7304 (N_7304,N_6581,N_6672);
nor U7305 (N_7305,N_6989,N_6679);
or U7306 (N_7306,N_6558,N_6786);
nor U7307 (N_7307,N_6645,N_6930);
or U7308 (N_7308,N_6552,N_6604);
and U7309 (N_7309,N_6544,N_6951);
nand U7310 (N_7310,N_6778,N_6567);
xor U7311 (N_7311,N_6915,N_6847);
nand U7312 (N_7312,N_6571,N_6901);
and U7313 (N_7313,N_6654,N_6617);
nand U7314 (N_7314,N_6648,N_6966);
and U7315 (N_7315,N_6783,N_6681);
nand U7316 (N_7316,N_6518,N_6761);
xor U7317 (N_7317,N_6775,N_6667);
nor U7318 (N_7318,N_6974,N_6544);
nand U7319 (N_7319,N_6551,N_6651);
nand U7320 (N_7320,N_6756,N_6831);
nand U7321 (N_7321,N_6730,N_6580);
nand U7322 (N_7322,N_6833,N_6555);
and U7323 (N_7323,N_6906,N_6841);
nand U7324 (N_7324,N_6763,N_6856);
nor U7325 (N_7325,N_6571,N_6668);
nand U7326 (N_7326,N_6838,N_6794);
and U7327 (N_7327,N_6759,N_6951);
xnor U7328 (N_7328,N_6870,N_6512);
nand U7329 (N_7329,N_6886,N_6765);
nand U7330 (N_7330,N_6702,N_6511);
xor U7331 (N_7331,N_6946,N_6608);
nand U7332 (N_7332,N_6938,N_6907);
and U7333 (N_7333,N_6769,N_6593);
xnor U7334 (N_7334,N_6639,N_6796);
xor U7335 (N_7335,N_6675,N_6612);
nand U7336 (N_7336,N_6875,N_6663);
and U7337 (N_7337,N_6504,N_6537);
xnor U7338 (N_7338,N_6680,N_6847);
or U7339 (N_7339,N_6686,N_6834);
or U7340 (N_7340,N_6857,N_6794);
or U7341 (N_7341,N_6841,N_6554);
nand U7342 (N_7342,N_6935,N_6518);
and U7343 (N_7343,N_6920,N_6727);
nor U7344 (N_7344,N_6728,N_6867);
xnor U7345 (N_7345,N_6652,N_6738);
xor U7346 (N_7346,N_6729,N_6632);
xor U7347 (N_7347,N_6866,N_6558);
nor U7348 (N_7348,N_6787,N_6837);
nand U7349 (N_7349,N_6799,N_6842);
and U7350 (N_7350,N_6590,N_6942);
nor U7351 (N_7351,N_6764,N_6690);
or U7352 (N_7352,N_6983,N_6631);
and U7353 (N_7353,N_6677,N_6861);
or U7354 (N_7354,N_6709,N_6627);
or U7355 (N_7355,N_6514,N_6776);
xnor U7356 (N_7356,N_6804,N_6579);
xor U7357 (N_7357,N_6747,N_6717);
and U7358 (N_7358,N_6706,N_6559);
nor U7359 (N_7359,N_6819,N_6750);
nand U7360 (N_7360,N_6973,N_6796);
xnor U7361 (N_7361,N_6977,N_6552);
and U7362 (N_7362,N_6772,N_6714);
nor U7363 (N_7363,N_6690,N_6934);
or U7364 (N_7364,N_6719,N_6761);
and U7365 (N_7365,N_6961,N_6749);
or U7366 (N_7366,N_6572,N_6860);
and U7367 (N_7367,N_6888,N_6912);
and U7368 (N_7368,N_6699,N_6834);
nand U7369 (N_7369,N_6684,N_6645);
nor U7370 (N_7370,N_6857,N_6875);
or U7371 (N_7371,N_6708,N_6864);
nand U7372 (N_7372,N_6744,N_6807);
nand U7373 (N_7373,N_6987,N_6824);
nand U7374 (N_7374,N_6674,N_6766);
nor U7375 (N_7375,N_6890,N_6586);
or U7376 (N_7376,N_6814,N_6645);
nand U7377 (N_7377,N_6835,N_6992);
nor U7378 (N_7378,N_6928,N_6590);
and U7379 (N_7379,N_6560,N_6724);
or U7380 (N_7380,N_6656,N_6721);
nand U7381 (N_7381,N_6906,N_6777);
and U7382 (N_7382,N_6577,N_6773);
or U7383 (N_7383,N_6569,N_6622);
nor U7384 (N_7384,N_6951,N_6955);
or U7385 (N_7385,N_6520,N_6941);
nor U7386 (N_7386,N_6836,N_6899);
nor U7387 (N_7387,N_6528,N_6519);
nor U7388 (N_7388,N_6785,N_6979);
xor U7389 (N_7389,N_6821,N_6622);
and U7390 (N_7390,N_6572,N_6750);
nand U7391 (N_7391,N_6884,N_6827);
or U7392 (N_7392,N_6880,N_6624);
nand U7393 (N_7393,N_6730,N_6933);
nand U7394 (N_7394,N_6811,N_6916);
nor U7395 (N_7395,N_6552,N_6845);
or U7396 (N_7396,N_6757,N_6932);
nor U7397 (N_7397,N_6605,N_6558);
nor U7398 (N_7398,N_6595,N_6596);
xor U7399 (N_7399,N_6616,N_6717);
nand U7400 (N_7400,N_6634,N_6976);
and U7401 (N_7401,N_6990,N_6694);
nor U7402 (N_7402,N_6682,N_6574);
nor U7403 (N_7403,N_6721,N_6886);
nand U7404 (N_7404,N_6621,N_6924);
nor U7405 (N_7405,N_6681,N_6653);
or U7406 (N_7406,N_6909,N_6785);
nor U7407 (N_7407,N_6568,N_6521);
and U7408 (N_7408,N_6698,N_6746);
xnor U7409 (N_7409,N_6532,N_6683);
nor U7410 (N_7410,N_6847,N_6797);
nand U7411 (N_7411,N_6519,N_6708);
xnor U7412 (N_7412,N_6599,N_6796);
nor U7413 (N_7413,N_6644,N_6954);
or U7414 (N_7414,N_6551,N_6562);
xnor U7415 (N_7415,N_6826,N_6601);
and U7416 (N_7416,N_6872,N_6560);
xor U7417 (N_7417,N_6812,N_6533);
nor U7418 (N_7418,N_6518,N_6932);
xnor U7419 (N_7419,N_6709,N_6732);
or U7420 (N_7420,N_6659,N_6537);
xnor U7421 (N_7421,N_6603,N_6774);
nand U7422 (N_7422,N_6843,N_6949);
or U7423 (N_7423,N_6583,N_6639);
xor U7424 (N_7424,N_6941,N_6537);
or U7425 (N_7425,N_6867,N_6848);
xor U7426 (N_7426,N_6949,N_6740);
or U7427 (N_7427,N_6965,N_6765);
nor U7428 (N_7428,N_6858,N_6949);
or U7429 (N_7429,N_6789,N_6621);
nor U7430 (N_7430,N_6530,N_6584);
nand U7431 (N_7431,N_6716,N_6662);
nor U7432 (N_7432,N_6958,N_6800);
xnor U7433 (N_7433,N_6661,N_6741);
or U7434 (N_7434,N_6972,N_6763);
or U7435 (N_7435,N_6549,N_6977);
nor U7436 (N_7436,N_6596,N_6950);
or U7437 (N_7437,N_6817,N_6538);
or U7438 (N_7438,N_6539,N_6757);
or U7439 (N_7439,N_6997,N_6852);
or U7440 (N_7440,N_6876,N_6918);
nor U7441 (N_7441,N_6917,N_6590);
and U7442 (N_7442,N_6923,N_6634);
or U7443 (N_7443,N_6603,N_6523);
nand U7444 (N_7444,N_6956,N_6701);
and U7445 (N_7445,N_6651,N_6860);
and U7446 (N_7446,N_6838,N_6803);
and U7447 (N_7447,N_6642,N_6626);
nand U7448 (N_7448,N_6529,N_6630);
or U7449 (N_7449,N_6955,N_6799);
nor U7450 (N_7450,N_6919,N_6681);
xor U7451 (N_7451,N_6592,N_6702);
and U7452 (N_7452,N_6643,N_6955);
xor U7453 (N_7453,N_6561,N_6873);
xnor U7454 (N_7454,N_6644,N_6964);
xnor U7455 (N_7455,N_6563,N_6999);
xnor U7456 (N_7456,N_6565,N_6634);
nand U7457 (N_7457,N_6513,N_6970);
or U7458 (N_7458,N_6743,N_6902);
or U7459 (N_7459,N_6814,N_6964);
nand U7460 (N_7460,N_6753,N_6698);
nand U7461 (N_7461,N_6894,N_6963);
xnor U7462 (N_7462,N_6611,N_6811);
nor U7463 (N_7463,N_6705,N_6915);
nand U7464 (N_7464,N_6823,N_6804);
nor U7465 (N_7465,N_6577,N_6524);
nor U7466 (N_7466,N_6781,N_6837);
xnor U7467 (N_7467,N_6964,N_6779);
xnor U7468 (N_7468,N_6986,N_6670);
nand U7469 (N_7469,N_6853,N_6904);
xor U7470 (N_7470,N_6761,N_6590);
and U7471 (N_7471,N_6984,N_6813);
nand U7472 (N_7472,N_6926,N_6836);
nand U7473 (N_7473,N_6808,N_6601);
nor U7474 (N_7474,N_6897,N_6545);
and U7475 (N_7475,N_6877,N_6553);
nand U7476 (N_7476,N_6614,N_6516);
and U7477 (N_7477,N_6846,N_6962);
or U7478 (N_7478,N_6962,N_6723);
and U7479 (N_7479,N_6526,N_6712);
and U7480 (N_7480,N_6627,N_6590);
xor U7481 (N_7481,N_6978,N_6722);
or U7482 (N_7482,N_6601,N_6621);
or U7483 (N_7483,N_6815,N_6910);
or U7484 (N_7484,N_6929,N_6961);
or U7485 (N_7485,N_6954,N_6724);
and U7486 (N_7486,N_6515,N_6848);
and U7487 (N_7487,N_6855,N_6987);
nand U7488 (N_7488,N_6813,N_6689);
or U7489 (N_7489,N_6562,N_6849);
xor U7490 (N_7490,N_6622,N_6793);
and U7491 (N_7491,N_6671,N_6535);
nand U7492 (N_7492,N_6554,N_6996);
or U7493 (N_7493,N_6574,N_6614);
and U7494 (N_7494,N_6830,N_6930);
and U7495 (N_7495,N_6703,N_6752);
or U7496 (N_7496,N_6627,N_6701);
or U7497 (N_7497,N_6789,N_6867);
and U7498 (N_7498,N_6975,N_6849);
nand U7499 (N_7499,N_6900,N_6970);
or U7500 (N_7500,N_7441,N_7062);
or U7501 (N_7501,N_7416,N_7382);
nor U7502 (N_7502,N_7443,N_7040);
or U7503 (N_7503,N_7006,N_7207);
and U7504 (N_7504,N_7402,N_7083);
nor U7505 (N_7505,N_7464,N_7347);
nor U7506 (N_7506,N_7194,N_7242);
or U7507 (N_7507,N_7037,N_7051);
and U7508 (N_7508,N_7213,N_7004);
and U7509 (N_7509,N_7081,N_7078);
or U7510 (N_7510,N_7336,N_7294);
xnor U7511 (N_7511,N_7262,N_7179);
nor U7512 (N_7512,N_7011,N_7188);
or U7513 (N_7513,N_7461,N_7360);
nand U7514 (N_7514,N_7344,N_7252);
or U7515 (N_7515,N_7109,N_7233);
or U7516 (N_7516,N_7293,N_7270);
or U7517 (N_7517,N_7150,N_7246);
xor U7518 (N_7518,N_7239,N_7258);
or U7519 (N_7519,N_7259,N_7266);
and U7520 (N_7520,N_7003,N_7395);
xor U7521 (N_7521,N_7303,N_7248);
xnor U7522 (N_7522,N_7495,N_7131);
nor U7523 (N_7523,N_7136,N_7088);
nand U7524 (N_7524,N_7352,N_7404);
or U7525 (N_7525,N_7057,N_7103);
xor U7526 (N_7526,N_7029,N_7177);
or U7527 (N_7527,N_7376,N_7257);
or U7528 (N_7528,N_7363,N_7287);
or U7529 (N_7529,N_7280,N_7216);
xor U7530 (N_7530,N_7403,N_7309);
nor U7531 (N_7531,N_7351,N_7438);
or U7532 (N_7532,N_7412,N_7359);
nor U7533 (N_7533,N_7159,N_7277);
and U7534 (N_7534,N_7086,N_7473);
xnor U7535 (N_7535,N_7429,N_7295);
or U7536 (N_7536,N_7132,N_7275);
nand U7537 (N_7537,N_7299,N_7015);
and U7538 (N_7538,N_7307,N_7151);
and U7539 (N_7539,N_7420,N_7430);
nand U7540 (N_7540,N_7219,N_7191);
and U7541 (N_7541,N_7452,N_7138);
nand U7542 (N_7542,N_7285,N_7223);
and U7543 (N_7543,N_7073,N_7459);
or U7544 (N_7544,N_7397,N_7494);
or U7545 (N_7545,N_7341,N_7311);
and U7546 (N_7546,N_7399,N_7025);
and U7547 (N_7547,N_7163,N_7424);
xnor U7548 (N_7548,N_7445,N_7018);
xnor U7549 (N_7549,N_7212,N_7240);
and U7550 (N_7550,N_7271,N_7053);
nand U7551 (N_7551,N_7471,N_7155);
and U7552 (N_7552,N_7224,N_7465);
and U7553 (N_7553,N_7182,N_7426);
xnor U7554 (N_7554,N_7115,N_7400);
nand U7555 (N_7555,N_7178,N_7306);
and U7556 (N_7556,N_7398,N_7047);
xor U7557 (N_7557,N_7192,N_7470);
or U7558 (N_7558,N_7368,N_7444);
nor U7559 (N_7559,N_7033,N_7002);
xor U7560 (N_7560,N_7048,N_7496);
and U7561 (N_7561,N_7263,N_7268);
or U7562 (N_7562,N_7054,N_7378);
and U7563 (N_7563,N_7091,N_7034);
nor U7564 (N_7564,N_7431,N_7238);
or U7565 (N_7565,N_7020,N_7321);
nor U7566 (N_7566,N_7462,N_7050);
xnor U7567 (N_7567,N_7154,N_7110);
nor U7568 (N_7568,N_7032,N_7437);
nor U7569 (N_7569,N_7408,N_7350);
nand U7570 (N_7570,N_7362,N_7035);
nor U7571 (N_7571,N_7377,N_7128);
nand U7572 (N_7572,N_7147,N_7354);
and U7573 (N_7573,N_7393,N_7189);
and U7574 (N_7574,N_7121,N_7381);
or U7575 (N_7575,N_7292,N_7435);
xor U7576 (N_7576,N_7476,N_7217);
nor U7577 (N_7577,N_7288,N_7272);
nand U7578 (N_7578,N_7406,N_7079);
and U7579 (N_7579,N_7409,N_7319);
or U7580 (N_7580,N_7488,N_7273);
xnor U7581 (N_7581,N_7168,N_7227);
nor U7582 (N_7582,N_7195,N_7332);
nor U7583 (N_7583,N_7475,N_7129);
nand U7584 (N_7584,N_7484,N_7099);
xor U7585 (N_7585,N_7201,N_7281);
or U7586 (N_7586,N_7049,N_7236);
nor U7587 (N_7587,N_7125,N_7463);
xnor U7588 (N_7588,N_7372,N_7481);
and U7589 (N_7589,N_7064,N_7067);
nor U7590 (N_7590,N_7442,N_7228);
nand U7591 (N_7591,N_7282,N_7187);
nor U7592 (N_7592,N_7142,N_7413);
nand U7593 (N_7593,N_7204,N_7071);
nor U7594 (N_7594,N_7490,N_7483);
and U7595 (N_7595,N_7209,N_7183);
nor U7596 (N_7596,N_7491,N_7302);
or U7597 (N_7597,N_7254,N_7021);
nand U7598 (N_7598,N_7096,N_7357);
and U7599 (N_7599,N_7027,N_7371);
nand U7600 (N_7600,N_7127,N_7199);
or U7601 (N_7601,N_7203,N_7405);
or U7602 (N_7602,N_7036,N_7366);
xnor U7603 (N_7603,N_7458,N_7331);
and U7604 (N_7604,N_7065,N_7433);
nor U7605 (N_7605,N_7226,N_7184);
xnor U7606 (N_7606,N_7338,N_7356);
or U7607 (N_7607,N_7022,N_7056);
xnor U7608 (N_7608,N_7094,N_7044);
xnor U7609 (N_7609,N_7104,N_7485);
nor U7610 (N_7610,N_7324,N_7101);
nand U7611 (N_7611,N_7012,N_7063);
or U7612 (N_7612,N_7122,N_7353);
or U7613 (N_7613,N_7333,N_7250);
and U7614 (N_7614,N_7206,N_7396);
nor U7615 (N_7615,N_7215,N_7264);
or U7616 (N_7616,N_7477,N_7369);
or U7617 (N_7617,N_7031,N_7123);
and U7618 (N_7618,N_7421,N_7276);
nand U7619 (N_7619,N_7451,N_7193);
and U7620 (N_7620,N_7211,N_7161);
xor U7621 (N_7621,N_7170,N_7419);
or U7622 (N_7622,N_7326,N_7247);
and U7623 (N_7623,N_7417,N_7074);
or U7624 (N_7624,N_7148,N_7106);
nor U7625 (N_7625,N_7210,N_7385);
or U7626 (N_7626,N_7448,N_7348);
or U7627 (N_7627,N_7283,N_7414);
xnor U7628 (N_7628,N_7434,N_7260);
xnor U7629 (N_7629,N_7315,N_7274);
and U7630 (N_7630,N_7328,N_7139);
or U7631 (N_7631,N_7411,N_7460);
nand U7632 (N_7632,N_7119,N_7384);
or U7633 (N_7633,N_7305,N_7087);
xor U7634 (N_7634,N_7089,N_7410);
xor U7635 (N_7635,N_7007,N_7042);
or U7636 (N_7636,N_7265,N_7137);
or U7637 (N_7637,N_7449,N_7023);
nand U7638 (N_7638,N_7135,N_7279);
nor U7639 (N_7639,N_7166,N_7221);
xor U7640 (N_7640,N_7208,N_7296);
xor U7641 (N_7641,N_7244,N_7092);
xnor U7642 (N_7642,N_7069,N_7316);
and U7643 (N_7643,N_7190,N_7454);
nand U7644 (N_7644,N_7149,N_7145);
or U7645 (N_7645,N_7304,N_7472);
or U7646 (N_7646,N_7167,N_7026);
and U7647 (N_7647,N_7231,N_7017);
or U7648 (N_7648,N_7428,N_7176);
or U7649 (N_7649,N_7261,N_7133);
xnor U7650 (N_7650,N_7152,N_7425);
nand U7651 (N_7651,N_7058,N_7156);
nor U7652 (N_7652,N_7334,N_7269);
nand U7653 (N_7653,N_7180,N_7478);
xnor U7654 (N_7654,N_7346,N_7169);
and U7655 (N_7655,N_7432,N_7016);
or U7656 (N_7656,N_7267,N_7427);
nor U7657 (N_7657,N_7300,N_7340);
and U7658 (N_7658,N_7289,N_7329);
or U7659 (N_7659,N_7019,N_7097);
xor U7660 (N_7660,N_7039,N_7255);
nor U7661 (N_7661,N_7066,N_7114);
and U7662 (N_7662,N_7230,N_7290);
and U7663 (N_7663,N_7418,N_7489);
or U7664 (N_7664,N_7222,N_7243);
xor U7665 (N_7665,N_7301,N_7038);
xnor U7666 (N_7666,N_7415,N_7120);
and U7667 (N_7667,N_7113,N_7325);
nand U7668 (N_7668,N_7095,N_7486);
nor U7669 (N_7669,N_7361,N_7162);
xor U7670 (N_7670,N_7389,N_7380);
nand U7671 (N_7671,N_7140,N_7077);
or U7672 (N_7672,N_7497,N_7010);
nor U7673 (N_7673,N_7084,N_7196);
xnor U7674 (N_7674,N_7253,N_7153);
nor U7675 (N_7675,N_7028,N_7157);
or U7676 (N_7676,N_7480,N_7436);
nor U7677 (N_7677,N_7374,N_7358);
xor U7678 (N_7678,N_7327,N_7466);
xor U7679 (N_7679,N_7030,N_7107);
nand U7680 (N_7680,N_7308,N_7256);
nand U7681 (N_7681,N_7298,N_7278);
nand U7682 (N_7682,N_7116,N_7102);
and U7683 (N_7683,N_7474,N_7364);
or U7684 (N_7684,N_7450,N_7313);
and U7685 (N_7685,N_7317,N_7447);
xor U7686 (N_7686,N_7080,N_7482);
xor U7687 (N_7687,N_7009,N_7072);
or U7688 (N_7688,N_7108,N_7446);
and U7689 (N_7689,N_7312,N_7249);
xor U7690 (N_7690,N_7499,N_7493);
or U7691 (N_7691,N_7008,N_7043);
nand U7692 (N_7692,N_7141,N_7202);
nor U7693 (N_7693,N_7245,N_7082);
nor U7694 (N_7694,N_7185,N_7370);
nand U7695 (N_7695,N_7387,N_7041);
and U7696 (N_7696,N_7342,N_7124);
nand U7697 (N_7697,N_7343,N_7111);
nand U7698 (N_7698,N_7457,N_7117);
nor U7699 (N_7699,N_7479,N_7394);
or U7700 (N_7700,N_7205,N_7158);
nand U7701 (N_7701,N_7144,N_7143);
or U7702 (N_7702,N_7367,N_7234);
or U7703 (N_7703,N_7439,N_7171);
xor U7704 (N_7704,N_7001,N_7455);
nor U7705 (N_7705,N_7229,N_7045);
and U7706 (N_7706,N_7173,N_7061);
nor U7707 (N_7707,N_7105,N_7492);
or U7708 (N_7708,N_7320,N_7024);
and U7709 (N_7709,N_7407,N_7456);
and U7710 (N_7710,N_7068,N_7052);
nand U7711 (N_7711,N_7355,N_7126);
nor U7712 (N_7712,N_7098,N_7375);
nor U7713 (N_7713,N_7453,N_7401);
and U7714 (N_7714,N_7379,N_7422);
xnor U7715 (N_7715,N_7314,N_7232);
nor U7716 (N_7716,N_7165,N_7174);
nor U7717 (N_7717,N_7172,N_7112);
nand U7718 (N_7718,N_7218,N_7323);
nor U7719 (N_7719,N_7487,N_7286);
xor U7720 (N_7720,N_7130,N_7345);
xor U7721 (N_7721,N_7055,N_7337);
or U7722 (N_7722,N_7467,N_7059);
xnor U7723 (N_7723,N_7093,N_7000);
or U7724 (N_7724,N_7085,N_7146);
nor U7725 (N_7725,N_7214,N_7391);
nor U7726 (N_7726,N_7198,N_7498);
or U7727 (N_7727,N_7160,N_7322);
nor U7728 (N_7728,N_7200,N_7392);
xnor U7729 (N_7729,N_7386,N_7164);
or U7730 (N_7730,N_7297,N_7284);
and U7731 (N_7731,N_7076,N_7349);
and U7732 (N_7732,N_7070,N_7335);
xnor U7733 (N_7733,N_7339,N_7318);
or U7734 (N_7734,N_7423,N_7468);
or U7735 (N_7735,N_7291,N_7235);
nor U7736 (N_7736,N_7175,N_7440);
nor U7737 (N_7737,N_7373,N_7090);
xor U7738 (N_7738,N_7005,N_7225);
xor U7739 (N_7739,N_7100,N_7013);
nand U7740 (N_7740,N_7075,N_7469);
xnor U7741 (N_7741,N_7330,N_7186);
nor U7742 (N_7742,N_7383,N_7197);
xor U7743 (N_7743,N_7220,N_7118);
xor U7744 (N_7744,N_7046,N_7365);
nor U7745 (N_7745,N_7134,N_7060);
xnor U7746 (N_7746,N_7390,N_7241);
xor U7747 (N_7747,N_7388,N_7181);
and U7748 (N_7748,N_7237,N_7310);
and U7749 (N_7749,N_7251,N_7014);
xnor U7750 (N_7750,N_7223,N_7039);
nor U7751 (N_7751,N_7240,N_7140);
xor U7752 (N_7752,N_7085,N_7064);
nand U7753 (N_7753,N_7185,N_7229);
nand U7754 (N_7754,N_7298,N_7467);
and U7755 (N_7755,N_7407,N_7167);
or U7756 (N_7756,N_7358,N_7398);
nor U7757 (N_7757,N_7337,N_7345);
nor U7758 (N_7758,N_7025,N_7242);
nand U7759 (N_7759,N_7270,N_7267);
nor U7760 (N_7760,N_7491,N_7397);
and U7761 (N_7761,N_7314,N_7003);
xnor U7762 (N_7762,N_7196,N_7348);
nor U7763 (N_7763,N_7270,N_7279);
and U7764 (N_7764,N_7270,N_7175);
nand U7765 (N_7765,N_7398,N_7390);
and U7766 (N_7766,N_7388,N_7439);
or U7767 (N_7767,N_7196,N_7121);
nand U7768 (N_7768,N_7471,N_7346);
nand U7769 (N_7769,N_7425,N_7283);
nor U7770 (N_7770,N_7304,N_7014);
nand U7771 (N_7771,N_7494,N_7310);
nand U7772 (N_7772,N_7323,N_7024);
and U7773 (N_7773,N_7349,N_7261);
nand U7774 (N_7774,N_7404,N_7327);
and U7775 (N_7775,N_7293,N_7045);
and U7776 (N_7776,N_7158,N_7233);
nor U7777 (N_7777,N_7406,N_7125);
nand U7778 (N_7778,N_7167,N_7203);
or U7779 (N_7779,N_7203,N_7142);
nor U7780 (N_7780,N_7005,N_7033);
nor U7781 (N_7781,N_7134,N_7468);
and U7782 (N_7782,N_7035,N_7247);
or U7783 (N_7783,N_7210,N_7417);
and U7784 (N_7784,N_7086,N_7489);
or U7785 (N_7785,N_7065,N_7288);
and U7786 (N_7786,N_7146,N_7052);
xor U7787 (N_7787,N_7387,N_7193);
or U7788 (N_7788,N_7402,N_7346);
and U7789 (N_7789,N_7152,N_7368);
nor U7790 (N_7790,N_7387,N_7244);
xor U7791 (N_7791,N_7257,N_7407);
nor U7792 (N_7792,N_7038,N_7378);
nand U7793 (N_7793,N_7490,N_7439);
xnor U7794 (N_7794,N_7190,N_7251);
nand U7795 (N_7795,N_7304,N_7248);
and U7796 (N_7796,N_7410,N_7346);
and U7797 (N_7797,N_7292,N_7105);
and U7798 (N_7798,N_7022,N_7434);
or U7799 (N_7799,N_7078,N_7153);
nand U7800 (N_7800,N_7316,N_7207);
or U7801 (N_7801,N_7373,N_7217);
nor U7802 (N_7802,N_7122,N_7201);
xor U7803 (N_7803,N_7259,N_7041);
nand U7804 (N_7804,N_7089,N_7150);
nor U7805 (N_7805,N_7104,N_7102);
and U7806 (N_7806,N_7066,N_7495);
or U7807 (N_7807,N_7043,N_7384);
or U7808 (N_7808,N_7272,N_7369);
or U7809 (N_7809,N_7013,N_7469);
nor U7810 (N_7810,N_7349,N_7429);
or U7811 (N_7811,N_7261,N_7456);
nor U7812 (N_7812,N_7042,N_7108);
xor U7813 (N_7813,N_7084,N_7135);
nand U7814 (N_7814,N_7202,N_7361);
nor U7815 (N_7815,N_7341,N_7097);
or U7816 (N_7816,N_7425,N_7194);
and U7817 (N_7817,N_7354,N_7331);
xnor U7818 (N_7818,N_7265,N_7494);
or U7819 (N_7819,N_7200,N_7109);
nand U7820 (N_7820,N_7251,N_7472);
or U7821 (N_7821,N_7055,N_7282);
nand U7822 (N_7822,N_7391,N_7191);
nand U7823 (N_7823,N_7445,N_7439);
nor U7824 (N_7824,N_7497,N_7498);
or U7825 (N_7825,N_7128,N_7401);
nor U7826 (N_7826,N_7144,N_7233);
xor U7827 (N_7827,N_7456,N_7481);
or U7828 (N_7828,N_7173,N_7016);
xnor U7829 (N_7829,N_7443,N_7225);
xnor U7830 (N_7830,N_7064,N_7447);
and U7831 (N_7831,N_7047,N_7497);
nor U7832 (N_7832,N_7408,N_7393);
nand U7833 (N_7833,N_7441,N_7434);
nand U7834 (N_7834,N_7254,N_7012);
xnor U7835 (N_7835,N_7180,N_7410);
and U7836 (N_7836,N_7409,N_7306);
and U7837 (N_7837,N_7451,N_7085);
or U7838 (N_7838,N_7067,N_7424);
nand U7839 (N_7839,N_7352,N_7231);
nand U7840 (N_7840,N_7283,N_7490);
nand U7841 (N_7841,N_7113,N_7423);
xor U7842 (N_7842,N_7088,N_7286);
nor U7843 (N_7843,N_7459,N_7192);
and U7844 (N_7844,N_7487,N_7355);
xor U7845 (N_7845,N_7432,N_7015);
nor U7846 (N_7846,N_7263,N_7356);
nor U7847 (N_7847,N_7046,N_7430);
nor U7848 (N_7848,N_7036,N_7317);
or U7849 (N_7849,N_7164,N_7374);
and U7850 (N_7850,N_7389,N_7470);
or U7851 (N_7851,N_7237,N_7212);
xor U7852 (N_7852,N_7341,N_7416);
nand U7853 (N_7853,N_7315,N_7413);
and U7854 (N_7854,N_7380,N_7073);
xor U7855 (N_7855,N_7015,N_7161);
nor U7856 (N_7856,N_7407,N_7457);
xor U7857 (N_7857,N_7174,N_7111);
and U7858 (N_7858,N_7373,N_7002);
xnor U7859 (N_7859,N_7274,N_7056);
xor U7860 (N_7860,N_7462,N_7306);
nor U7861 (N_7861,N_7119,N_7288);
xor U7862 (N_7862,N_7231,N_7422);
nor U7863 (N_7863,N_7379,N_7285);
or U7864 (N_7864,N_7353,N_7339);
and U7865 (N_7865,N_7282,N_7362);
nand U7866 (N_7866,N_7156,N_7052);
nand U7867 (N_7867,N_7168,N_7045);
nor U7868 (N_7868,N_7233,N_7167);
and U7869 (N_7869,N_7298,N_7084);
nor U7870 (N_7870,N_7228,N_7429);
nor U7871 (N_7871,N_7128,N_7372);
nor U7872 (N_7872,N_7074,N_7290);
nor U7873 (N_7873,N_7377,N_7302);
and U7874 (N_7874,N_7192,N_7089);
nand U7875 (N_7875,N_7130,N_7478);
and U7876 (N_7876,N_7118,N_7446);
nor U7877 (N_7877,N_7417,N_7253);
xnor U7878 (N_7878,N_7466,N_7066);
xor U7879 (N_7879,N_7082,N_7455);
xor U7880 (N_7880,N_7179,N_7182);
xor U7881 (N_7881,N_7155,N_7413);
nand U7882 (N_7882,N_7306,N_7118);
or U7883 (N_7883,N_7376,N_7248);
and U7884 (N_7884,N_7228,N_7449);
xor U7885 (N_7885,N_7416,N_7380);
nor U7886 (N_7886,N_7149,N_7137);
or U7887 (N_7887,N_7415,N_7285);
xor U7888 (N_7888,N_7433,N_7316);
xnor U7889 (N_7889,N_7203,N_7249);
nand U7890 (N_7890,N_7231,N_7390);
nand U7891 (N_7891,N_7178,N_7403);
nor U7892 (N_7892,N_7252,N_7035);
and U7893 (N_7893,N_7486,N_7498);
xnor U7894 (N_7894,N_7075,N_7434);
xnor U7895 (N_7895,N_7162,N_7427);
xnor U7896 (N_7896,N_7322,N_7394);
or U7897 (N_7897,N_7186,N_7416);
or U7898 (N_7898,N_7457,N_7274);
and U7899 (N_7899,N_7372,N_7386);
or U7900 (N_7900,N_7277,N_7132);
or U7901 (N_7901,N_7311,N_7061);
and U7902 (N_7902,N_7474,N_7437);
nand U7903 (N_7903,N_7045,N_7126);
and U7904 (N_7904,N_7240,N_7432);
nand U7905 (N_7905,N_7281,N_7090);
xor U7906 (N_7906,N_7059,N_7046);
xnor U7907 (N_7907,N_7400,N_7342);
or U7908 (N_7908,N_7144,N_7397);
or U7909 (N_7909,N_7428,N_7208);
or U7910 (N_7910,N_7132,N_7212);
nand U7911 (N_7911,N_7253,N_7009);
or U7912 (N_7912,N_7317,N_7264);
nor U7913 (N_7913,N_7415,N_7239);
and U7914 (N_7914,N_7188,N_7141);
xor U7915 (N_7915,N_7448,N_7181);
and U7916 (N_7916,N_7398,N_7017);
xor U7917 (N_7917,N_7407,N_7486);
and U7918 (N_7918,N_7322,N_7193);
xnor U7919 (N_7919,N_7218,N_7142);
and U7920 (N_7920,N_7110,N_7138);
xnor U7921 (N_7921,N_7478,N_7033);
xnor U7922 (N_7922,N_7159,N_7199);
or U7923 (N_7923,N_7313,N_7219);
nand U7924 (N_7924,N_7248,N_7259);
and U7925 (N_7925,N_7103,N_7474);
nor U7926 (N_7926,N_7436,N_7286);
xor U7927 (N_7927,N_7230,N_7148);
nor U7928 (N_7928,N_7080,N_7146);
nor U7929 (N_7929,N_7090,N_7011);
xor U7930 (N_7930,N_7120,N_7283);
or U7931 (N_7931,N_7374,N_7209);
nand U7932 (N_7932,N_7482,N_7346);
nor U7933 (N_7933,N_7330,N_7275);
nor U7934 (N_7934,N_7117,N_7232);
nor U7935 (N_7935,N_7073,N_7002);
and U7936 (N_7936,N_7008,N_7218);
nor U7937 (N_7937,N_7147,N_7358);
and U7938 (N_7938,N_7045,N_7078);
xor U7939 (N_7939,N_7039,N_7021);
and U7940 (N_7940,N_7160,N_7467);
nand U7941 (N_7941,N_7105,N_7440);
or U7942 (N_7942,N_7104,N_7372);
or U7943 (N_7943,N_7207,N_7152);
or U7944 (N_7944,N_7498,N_7376);
nand U7945 (N_7945,N_7360,N_7009);
or U7946 (N_7946,N_7318,N_7050);
xnor U7947 (N_7947,N_7304,N_7167);
nand U7948 (N_7948,N_7204,N_7490);
or U7949 (N_7949,N_7374,N_7322);
nand U7950 (N_7950,N_7092,N_7475);
nand U7951 (N_7951,N_7192,N_7167);
nand U7952 (N_7952,N_7496,N_7201);
xnor U7953 (N_7953,N_7406,N_7042);
nor U7954 (N_7954,N_7461,N_7019);
nand U7955 (N_7955,N_7158,N_7324);
and U7956 (N_7956,N_7208,N_7305);
xnor U7957 (N_7957,N_7264,N_7428);
or U7958 (N_7958,N_7094,N_7275);
nand U7959 (N_7959,N_7418,N_7465);
nand U7960 (N_7960,N_7386,N_7402);
and U7961 (N_7961,N_7330,N_7295);
nand U7962 (N_7962,N_7413,N_7019);
nor U7963 (N_7963,N_7140,N_7115);
nor U7964 (N_7964,N_7155,N_7345);
xor U7965 (N_7965,N_7473,N_7101);
xnor U7966 (N_7966,N_7151,N_7389);
nand U7967 (N_7967,N_7225,N_7201);
nor U7968 (N_7968,N_7151,N_7088);
or U7969 (N_7969,N_7324,N_7029);
nand U7970 (N_7970,N_7158,N_7144);
xnor U7971 (N_7971,N_7493,N_7240);
nor U7972 (N_7972,N_7489,N_7244);
and U7973 (N_7973,N_7280,N_7115);
nand U7974 (N_7974,N_7337,N_7077);
and U7975 (N_7975,N_7199,N_7327);
xnor U7976 (N_7976,N_7132,N_7371);
nand U7977 (N_7977,N_7115,N_7181);
and U7978 (N_7978,N_7126,N_7316);
and U7979 (N_7979,N_7287,N_7414);
nand U7980 (N_7980,N_7116,N_7284);
nand U7981 (N_7981,N_7346,N_7150);
and U7982 (N_7982,N_7391,N_7245);
xor U7983 (N_7983,N_7363,N_7199);
nor U7984 (N_7984,N_7408,N_7221);
nand U7985 (N_7985,N_7452,N_7292);
nand U7986 (N_7986,N_7260,N_7110);
or U7987 (N_7987,N_7188,N_7255);
and U7988 (N_7988,N_7026,N_7153);
or U7989 (N_7989,N_7252,N_7114);
nand U7990 (N_7990,N_7492,N_7348);
nor U7991 (N_7991,N_7237,N_7292);
nand U7992 (N_7992,N_7192,N_7361);
or U7993 (N_7993,N_7139,N_7204);
and U7994 (N_7994,N_7092,N_7248);
and U7995 (N_7995,N_7044,N_7477);
or U7996 (N_7996,N_7131,N_7329);
and U7997 (N_7997,N_7076,N_7079);
and U7998 (N_7998,N_7377,N_7223);
and U7999 (N_7999,N_7249,N_7488);
nor U8000 (N_8000,N_7794,N_7865);
nor U8001 (N_8001,N_7917,N_7783);
nand U8002 (N_8002,N_7712,N_7887);
nor U8003 (N_8003,N_7749,N_7812);
or U8004 (N_8004,N_7822,N_7759);
and U8005 (N_8005,N_7616,N_7641);
nand U8006 (N_8006,N_7752,N_7744);
or U8007 (N_8007,N_7802,N_7946);
or U8008 (N_8008,N_7986,N_7629);
nand U8009 (N_8009,N_7782,N_7922);
and U8010 (N_8010,N_7524,N_7723);
nand U8011 (N_8011,N_7951,N_7988);
nand U8012 (N_8012,N_7554,N_7726);
nand U8013 (N_8013,N_7732,N_7549);
nand U8014 (N_8014,N_7800,N_7973);
or U8015 (N_8015,N_7608,N_7828);
nand U8016 (N_8016,N_7728,N_7531);
or U8017 (N_8017,N_7792,N_7952);
and U8018 (N_8018,N_7909,N_7716);
nor U8019 (N_8019,N_7795,N_7704);
xnor U8020 (N_8020,N_7850,N_7619);
or U8021 (N_8021,N_7544,N_7501);
or U8022 (N_8022,N_7970,N_7517);
nor U8023 (N_8023,N_7769,N_7523);
nor U8024 (N_8024,N_7817,N_7740);
nand U8025 (N_8025,N_7854,N_7706);
xnor U8026 (N_8026,N_7867,N_7957);
or U8027 (N_8027,N_7572,N_7844);
and U8028 (N_8028,N_7627,N_7881);
nor U8029 (N_8029,N_7760,N_7858);
nand U8030 (N_8030,N_7511,N_7924);
and U8031 (N_8031,N_7969,N_7929);
nand U8032 (N_8032,N_7990,N_7503);
nand U8033 (N_8033,N_7636,N_7600);
xor U8034 (N_8034,N_7985,N_7567);
xnor U8035 (N_8035,N_7787,N_7649);
xor U8036 (N_8036,N_7743,N_7642);
or U8037 (N_8037,N_7918,N_7692);
or U8038 (N_8038,N_7856,N_7886);
xor U8039 (N_8039,N_7774,N_7741);
and U8040 (N_8040,N_7701,N_7606);
xor U8041 (N_8041,N_7984,N_7950);
or U8042 (N_8042,N_7789,N_7597);
and U8043 (N_8043,N_7763,N_7781);
xor U8044 (N_8044,N_7602,N_7633);
and U8045 (N_8045,N_7813,N_7528);
or U8046 (N_8046,N_7579,N_7588);
nand U8047 (N_8047,N_7776,N_7956);
or U8048 (N_8048,N_7637,N_7559);
and U8049 (N_8049,N_7713,N_7804);
nor U8050 (N_8050,N_7902,N_7773);
nand U8051 (N_8051,N_7987,N_7966);
xnor U8052 (N_8052,N_7573,N_7648);
xnor U8053 (N_8053,N_7532,N_7691);
xnor U8054 (N_8054,N_7976,N_7715);
or U8055 (N_8055,N_7672,N_7820);
nand U8056 (N_8056,N_7996,N_7780);
or U8057 (N_8057,N_7786,N_7623);
and U8058 (N_8058,N_7639,N_7937);
xnor U8059 (N_8059,N_7870,N_7831);
nor U8060 (N_8060,N_7862,N_7718);
and U8061 (N_8061,N_7734,N_7905);
xor U8062 (N_8062,N_7832,N_7989);
xnor U8063 (N_8063,N_7992,N_7907);
nor U8064 (N_8064,N_7837,N_7654);
or U8065 (N_8065,N_7555,N_7647);
nor U8066 (N_8066,N_7537,N_7819);
and U8067 (N_8067,N_7615,N_7620);
xor U8068 (N_8068,N_7618,N_7583);
and U8069 (N_8069,N_7689,N_7582);
nor U8070 (N_8070,N_7936,N_7586);
or U8071 (N_8071,N_7888,N_7981);
and U8072 (N_8072,N_7680,N_7851);
or U8073 (N_8073,N_7906,N_7546);
xor U8074 (N_8074,N_7519,N_7975);
nor U8075 (N_8075,N_7810,N_7551);
nor U8076 (N_8076,N_7872,N_7643);
and U8077 (N_8077,N_7940,N_7660);
nor U8078 (N_8078,N_7681,N_7742);
nor U8079 (N_8079,N_7500,N_7694);
or U8080 (N_8080,N_7977,N_7612);
or U8081 (N_8081,N_7892,N_7703);
and U8082 (N_8082,N_7964,N_7864);
nand U8083 (N_8083,N_7558,N_7978);
nor U8084 (N_8084,N_7852,N_7893);
nand U8085 (N_8085,N_7811,N_7842);
nand U8086 (N_8086,N_7841,N_7663);
and U8087 (N_8087,N_7754,N_7825);
xnor U8088 (N_8088,N_7614,N_7891);
and U8089 (N_8089,N_7974,N_7829);
and U8090 (N_8090,N_7836,N_7507);
xnor U8091 (N_8091,N_7980,N_7840);
and U8092 (N_8092,N_7745,N_7729);
nand U8093 (N_8093,N_7834,N_7827);
nand U8094 (N_8094,N_7671,N_7679);
and U8095 (N_8095,N_7958,N_7928);
nor U8096 (N_8096,N_7527,N_7762);
or U8097 (N_8097,N_7576,N_7658);
and U8098 (N_8098,N_7592,N_7653);
xor U8099 (N_8099,N_7839,N_7591);
and U8100 (N_8100,N_7747,N_7538);
and U8101 (N_8101,N_7874,N_7536);
nand U8102 (N_8102,N_7935,N_7962);
and U8103 (N_8103,N_7635,N_7569);
nand U8104 (N_8104,N_7667,N_7912);
and U8105 (N_8105,N_7934,N_7961);
nor U8106 (N_8106,N_7584,N_7542);
nor U8107 (N_8107,N_7847,N_7550);
nand U8108 (N_8108,N_7796,N_7863);
or U8109 (N_8109,N_7798,N_7801);
or U8110 (N_8110,N_7738,N_7580);
xnor U8111 (N_8111,N_7669,N_7705);
nand U8112 (N_8112,N_7943,N_7899);
nor U8113 (N_8113,N_7965,N_7530);
or U8114 (N_8114,N_7512,N_7947);
or U8115 (N_8115,N_7662,N_7901);
nand U8116 (N_8116,N_7739,N_7750);
xor U8117 (N_8117,N_7939,N_7522);
nand U8118 (N_8118,N_7545,N_7577);
nor U8119 (N_8119,N_7562,N_7855);
xnor U8120 (N_8120,N_7815,N_7510);
xor U8121 (N_8121,N_7735,N_7720);
nand U8122 (N_8122,N_7652,N_7682);
or U8123 (N_8123,N_7868,N_7799);
or U8124 (N_8124,N_7697,N_7910);
and U8125 (N_8125,N_7931,N_7757);
nor U8126 (N_8126,N_7727,N_7793);
and U8127 (N_8127,N_7890,N_7574);
nor U8128 (N_8128,N_7625,N_7730);
or U8129 (N_8129,N_7932,N_7993);
and U8130 (N_8130,N_7814,N_7930);
nand U8131 (N_8131,N_7646,N_7661);
nand U8132 (N_8132,N_7553,N_7945);
and U8133 (N_8133,N_7684,N_7609);
or U8134 (N_8134,N_7807,N_7502);
nor U8135 (N_8135,N_7761,N_7748);
or U8136 (N_8136,N_7861,N_7626);
xor U8137 (N_8137,N_7920,N_7768);
or U8138 (N_8138,N_7913,N_7610);
and U8139 (N_8139,N_7674,N_7710);
and U8140 (N_8140,N_7803,N_7896);
nor U8141 (N_8141,N_7736,N_7830);
nor U8142 (N_8142,N_7687,N_7882);
nor U8143 (N_8143,N_7919,N_7566);
xnor U8144 (N_8144,N_7826,N_7999);
nor U8145 (N_8145,N_7504,N_7708);
xnor U8146 (N_8146,N_7560,N_7714);
xnor U8147 (N_8147,N_7790,N_7571);
or U8148 (N_8148,N_7685,N_7645);
nor U8149 (N_8149,N_7529,N_7547);
nand U8150 (N_8150,N_7678,N_7628);
xor U8151 (N_8151,N_7823,N_7657);
xnor U8152 (N_8152,N_7696,N_7894);
or U8153 (N_8153,N_7816,N_7765);
xnor U8154 (N_8154,N_7656,N_7664);
nand U8155 (N_8155,N_7877,N_7771);
nor U8156 (N_8156,N_7556,N_7777);
or U8157 (N_8157,N_7721,N_7944);
or U8158 (N_8158,N_7514,N_7561);
nor U8159 (N_8159,N_7702,N_7630);
or U8160 (N_8160,N_7959,N_7880);
nor U8161 (N_8161,N_7764,N_7770);
and U8162 (N_8162,N_7541,N_7808);
and U8163 (N_8163,N_7543,N_7991);
xnor U8164 (N_8164,N_7960,N_7568);
and U8165 (N_8165,N_7889,N_7857);
nand U8166 (N_8166,N_7766,N_7621);
or U8167 (N_8167,N_7797,N_7695);
and U8168 (N_8168,N_7533,N_7921);
and U8169 (N_8169,N_7673,N_7693);
or U8170 (N_8170,N_7968,N_7904);
nand U8171 (N_8171,N_7785,N_7949);
or U8172 (N_8172,N_7724,N_7897);
xor U8173 (N_8173,N_7665,N_7873);
nor U8174 (N_8174,N_7860,N_7638);
nor U8175 (N_8175,N_7971,N_7589);
or U8176 (N_8176,N_7594,N_7683);
nor U8177 (N_8177,N_7731,N_7942);
nand U8178 (N_8178,N_7737,N_7775);
nand U8179 (N_8179,N_7967,N_7878);
nand U8180 (N_8180,N_7845,N_7599);
nand U8181 (N_8181,N_7846,N_7779);
or U8182 (N_8182,N_7565,N_7911);
xor U8183 (N_8183,N_7613,N_7982);
nand U8184 (N_8184,N_7733,N_7908);
xnor U8185 (N_8185,N_7518,N_7688);
and U8186 (N_8186,N_7895,N_7644);
nand U8187 (N_8187,N_7746,N_7916);
and U8188 (N_8188,N_7884,N_7564);
xnor U8189 (N_8189,N_7915,N_7994);
and U8190 (N_8190,N_7534,N_7900);
nor U8191 (N_8191,N_7651,N_7711);
nand U8192 (N_8192,N_7806,N_7725);
or U8193 (N_8193,N_7707,N_7521);
or U8194 (N_8194,N_7631,N_7938);
nand U8195 (N_8195,N_7535,N_7885);
nor U8196 (N_8196,N_7593,N_7853);
nor U8197 (N_8197,N_7595,N_7575);
nand U8198 (N_8198,N_7650,N_7563);
nand U8199 (N_8199,N_7525,N_7578);
nor U8200 (N_8200,N_7756,N_7607);
nand U8201 (N_8201,N_7859,N_7869);
nor U8202 (N_8202,N_7883,N_7505);
and U8203 (N_8203,N_7605,N_7824);
nor U8204 (N_8204,N_7675,N_7601);
or U8205 (N_8205,N_7767,N_7866);
nor U8206 (N_8206,N_7784,N_7772);
xnor U8207 (N_8207,N_7997,N_7552);
and U8208 (N_8208,N_7581,N_7753);
xor U8209 (N_8209,N_7722,N_7791);
and U8210 (N_8210,N_7963,N_7634);
xor U8211 (N_8211,N_7898,N_7698);
or U8212 (N_8212,N_7818,N_7506);
and U8213 (N_8213,N_7596,N_7876);
xnor U8214 (N_8214,N_7700,N_7998);
or U8215 (N_8215,N_7948,N_7717);
xor U8216 (N_8216,N_7686,N_7875);
xnor U8217 (N_8217,N_7604,N_7871);
or U8218 (N_8218,N_7632,N_7515);
nand U8219 (N_8219,N_7699,N_7690);
and U8220 (N_8220,N_7659,N_7603);
nor U8221 (N_8221,N_7655,N_7622);
nor U8222 (N_8222,N_7955,N_7520);
nand U8223 (N_8223,N_7755,N_7668);
nand U8224 (N_8224,N_7927,N_7983);
or U8225 (N_8225,N_7914,N_7587);
or U8226 (N_8226,N_7548,N_7508);
or U8227 (N_8227,N_7640,N_7821);
and U8228 (N_8228,N_7585,N_7933);
nand U8229 (N_8229,N_7617,N_7879);
or U8230 (N_8230,N_7539,N_7709);
nand U8231 (N_8231,N_7758,N_7833);
and U8232 (N_8232,N_7995,N_7719);
xor U8233 (N_8233,N_7666,N_7835);
or U8234 (N_8234,N_7979,N_7509);
or U8235 (N_8235,N_7923,N_7670);
and U8236 (N_8236,N_7809,N_7751);
xor U8237 (N_8237,N_7941,N_7843);
xor U8238 (N_8238,N_7513,N_7611);
xnor U8239 (N_8239,N_7954,N_7838);
or U8240 (N_8240,N_7953,N_7788);
nand U8241 (N_8241,N_7926,N_7805);
or U8242 (N_8242,N_7676,N_7903);
or U8243 (N_8243,N_7598,N_7516);
or U8244 (N_8244,N_7849,N_7570);
xnor U8245 (N_8245,N_7925,N_7540);
nand U8246 (N_8246,N_7526,N_7972);
or U8247 (N_8247,N_7624,N_7557);
or U8248 (N_8248,N_7590,N_7848);
xor U8249 (N_8249,N_7677,N_7778);
nor U8250 (N_8250,N_7682,N_7610);
nand U8251 (N_8251,N_7869,N_7843);
xor U8252 (N_8252,N_7637,N_7699);
nor U8253 (N_8253,N_7954,N_7590);
or U8254 (N_8254,N_7507,N_7599);
xor U8255 (N_8255,N_7528,N_7567);
or U8256 (N_8256,N_7951,N_7914);
nand U8257 (N_8257,N_7675,N_7812);
nor U8258 (N_8258,N_7647,N_7940);
nor U8259 (N_8259,N_7574,N_7579);
nor U8260 (N_8260,N_7724,N_7609);
nand U8261 (N_8261,N_7753,N_7630);
or U8262 (N_8262,N_7929,N_7699);
and U8263 (N_8263,N_7806,N_7521);
xnor U8264 (N_8264,N_7815,N_7739);
or U8265 (N_8265,N_7654,N_7974);
xor U8266 (N_8266,N_7738,N_7955);
or U8267 (N_8267,N_7985,N_7534);
nor U8268 (N_8268,N_7911,N_7900);
xnor U8269 (N_8269,N_7682,N_7924);
nand U8270 (N_8270,N_7642,N_7756);
and U8271 (N_8271,N_7511,N_7566);
xnor U8272 (N_8272,N_7575,N_7914);
xor U8273 (N_8273,N_7847,N_7575);
xor U8274 (N_8274,N_7768,N_7664);
nor U8275 (N_8275,N_7562,N_7872);
and U8276 (N_8276,N_7507,N_7705);
or U8277 (N_8277,N_7544,N_7560);
nand U8278 (N_8278,N_7782,N_7640);
nor U8279 (N_8279,N_7851,N_7684);
nor U8280 (N_8280,N_7762,N_7568);
xor U8281 (N_8281,N_7872,N_7651);
nor U8282 (N_8282,N_7680,N_7802);
or U8283 (N_8283,N_7812,N_7699);
nor U8284 (N_8284,N_7555,N_7998);
and U8285 (N_8285,N_7733,N_7615);
or U8286 (N_8286,N_7781,N_7746);
nor U8287 (N_8287,N_7549,N_7771);
and U8288 (N_8288,N_7909,N_7809);
or U8289 (N_8289,N_7961,N_7740);
xor U8290 (N_8290,N_7507,N_7718);
nor U8291 (N_8291,N_7512,N_7835);
and U8292 (N_8292,N_7550,N_7692);
nand U8293 (N_8293,N_7545,N_7971);
nor U8294 (N_8294,N_7763,N_7656);
nand U8295 (N_8295,N_7959,N_7576);
nand U8296 (N_8296,N_7520,N_7994);
nand U8297 (N_8297,N_7931,N_7998);
nand U8298 (N_8298,N_7646,N_7584);
xor U8299 (N_8299,N_7763,N_7805);
nand U8300 (N_8300,N_7937,N_7611);
xnor U8301 (N_8301,N_7972,N_7867);
xor U8302 (N_8302,N_7547,N_7908);
nor U8303 (N_8303,N_7695,N_7965);
or U8304 (N_8304,N_7829,N_7843);
or U8305 (N_8305,N_7759,N_7674);
xnor U8306 (N_8306,N_7860,N_7893);
nor U8307 (N_8307,N_7718,N_7931);
xor U8308 (N_8308,N_7604,N_7930);
nor U8309 (N_8309,N_7660,N_7937);
nand U8310 (N_8310,N_7583,N_7810);
nor U8311 (N_8311,N_7777,N_7626);
nand U8312 (N_8312,N_7751,N_7975);
xor U8313 (N_8313,N_7725,N_7501);
nor U8314 (N_8314,N_7978,N_7527);
or U8315 (N_8315,N_7870,N_7948);
or U8316 (N_8316,N_7654,N_7700);
nand U8317 (N_8317,N_7568,N_7961);
and U8318 (N_8318,N_7529,N_7801);
and U8319 (N_8319,N_7541,N_7824);
nor U8320 (N_8320,N_7896,N_7773);
nand U8321 (N_8321,N_7557,N_7573);
xor U8322 (N_8322,N_7752,N_7716);
and U8323 (N_8323,N_7500,N_7622);
and U8324 (N_8324,N_7697,N_7511);
nand U8325 (N_8325,N_7694,N_7771);
nor U8326 (N_8326,N_7888,N_7777);
and U8327 (N_8327,N_7746,N_7714);
and U8328 (N_8328,N_7737,N_7842);
nor U8329 (N_8329,N_7715,N_7949);
nor U8330 (N_8330,N_7785,N_7522);
nand U8331 (N_8331,N_7700,N_7688);
and U8332 (N_8332,N_7541,N_7506);
and U8333 (N_8333,N_7989,N_7781);
xor U8334 (N_8334,N_7818,N_7978);
nand U8335 (N_8335,N_7716,N_7508);
or U8336 (N_8336,N_7976,N_7991);
or U8337 (N_8337,N_7572,N_7557);
or U8338 (N_8338,N_7813,N_7655);
xor U8339 (N_8339,N_7879,N_7944);
or U8340 (N_8340,N_7982,N_7674);
and U8341 (N_8341,N_7632,N_7559);
xor U8342 (N_8342,N_7725,N_7835);
and U8343 (N_8343,N_7848,N_7572);
xnor U8344 (N_8344,N_7509,N_7805);
xor U8345 (N_8345,N_7910,N_7916);
or U8346 (N_8346,N_7772,N_7967);
and U8347 (N_8347,N_7975,N_7761);
xnor U8348 (N_8348,N_7996,N_7767);
nor U8349 (N_8349,N_7516,N_7593);
and U8350 (N_8350,N_7779,N_7795);
nor U8351 (N_8351,N_7896,N_7759);
nor U8352 (N_8352,N_7779,N_7829);
xor U8353 (N_8353,N_7894,N_7687);
nand U8354 (N_8354,N_7541,N_7731);
and U8355 (N_8355,N_7902,N_7873);
or U8356 (N_8356,N_7908,N_7700);
nand U8357 (N_8357,N_7606,N_7963);
xnor U8358 (N_8358,N_7889,N_7554);
nand U8359 (N_8359,N_7805,N_7502);
and U8360 (N_8360,N_7903,N_7687);
nand U8361 (N_8361,N_7871,N_7506);
or U8362 (N_8362,N_7895,N_7567);
nor U8363 (N_8363,N_7519,N_7851);
nand U8364 (N_8364,N_7526,N_7947);
xor U8365 (N_8365,N_7719,N_7527);
nor U8366 (N_8366,N_7563,N_7721);
nor U8367 (N_8367,N_7708,N_7523);
nor U8368 (N_8368,N_7568,N_7947);
or U8369 (N_8369,N_7909,N_7679);
nand U8370 (N_8370,N_7653,N_7860);
nor U8371 (N_8371,N_7542,N_7794);
or U8372 (N_8372,N_7941,N_7932);
or U8373 (N_8373,N_7682,N_7766);
xnor U8374 (N_8374,N_7613,N_7813);
xor U8375 (N_8375,N_7883,N_7677);
and U8376 (N_8376,N_7753,N_7930);
or U8377 (N_8377,N_7580,N_7928);
or U8378 (N_8378,N_7982,N_7844);
nor U8379 (N_8379,N_7558,N_7914);
or U8380 (N_8380,N_7724,N_7741);
nand U8381 (N_8381,N_7567,N_7769);
xor U8382 (N_8382,N_7989,N_7959);
or U8383 (N_8383,N_7999,N_7898);
or U8384 (N_8384,N_7776,N_7779);
xor U8385 (N_8385,N_7707,N_7621);
nand U8386 (N_8386,N_7542,N_7789);
or U8387 (N_8387,N_7987,N_7511);
xnor U8388 (N_8388,N_7938,N_7939);
xor U8389 (N_8389,N_7838,N_7798);
nor U8390 (N_8390,N_7515,N_7572);
xor U8391 (N_8391,N_7931,N_7593);
nand U8392 (N_8392,N_7553,N_7505);
nor U8393 (N_8393,N_7758,N_7631);
xor U8394 (N_8394,N_7515,N_7646);
nand U8395 (N_8395,N_7594,N_7721);
nand U8396 (N_8396,N_7544,N_7531);
nor U8397 (N_8397,N_7571,N_7537);
xor U8398 (N_8398,N_7744,N_7537);
nor U8399 (N_8399,N_7650,N_7957);
xor U8400 (N_8400,N_7762,N_7835);
nor U8401 (N_8401,N_7558,N_7638);
and U8402 (N_8402,N_7649,N_7695);
and U8403 (N_8403,N_7910,N_7981);
nand U8404 (N_8404,N_7717,N_7575);
and U8405 (N_8405,N_7658,N_7795);
nand U8406 (N_8406,N_7728,N_7819);
nor U8407 (N_8407,N_7647,N_7669);
nor U8408 (N_8408,N_7734,N_7965);
or U8409 (N_8409,N_7872,N_7544);
and U8410 (N_8410,N_7687,N_7814);
nor U8411 (N_8411,N_7932,N_7717);
nand U8412 (N_8412,N_7549,N_7983);
nor U8413 (N_8413,N_7842,N_7758);
nand U8414 (N_8414,N_7940,N_7789);
and U8415 (N_8415,N_7944,N_7609);
and U8416 (N_8416,N_7562,N_7874);
nand U8417 (N_8417,N_7968,N_7571);
or U8418 (N_8418,N_7563,N_7749);
and U8419 (N_8419,N_7523,N_7861);
nand U8420 (N_8420,N_7696,N_7857);
or U8421 (N_8421,N_7798,N_7818);
nand U8422 (N_8422,N_7567,N_7699);
nand U8423 (N_8423,N_7822,N_7583);
nand U8424 (N_8424,N_7936,N_7606);
or U8425 (N_8425,N_7718,N_7617);
xnor U8426 (N_8426,N_7743,N_7810);
or U8427 (N_8427,N_7510,N_7824);
xnor U8428 (N_8428,N_7654,N_7910);
or U8429 (N_8429,N_7956,N_7560);
xnor U8430 (N_8430,N_7832,N_7938);
nand U8431 (N_8431,N_7843,N_7532);
or U8432 (N_8432,N_7530,N_7917);
or U8433 (N_8433,N_7717,N_7819);
nor U8434 (N_8434,N_7590,N_7722);
and U8435 (N_8435,N_7589,N_7733);
and U8436 (N_8436,N_7989,N_7646);
or U8437 (N_8437,N_7564,N_7664);
xor U8438 (N_8438,N_7986,N_7981);
nand U8439 (N_8439,N_7966,N_7533);
and U8440 (N_8440,N_7664,N_7807);
xor U8441 (N_8441,N_7705,N_7674);
or U8442 (N_8442,N_7595,N_7936);
xor U8443 (N_8443,N_7521,N_7722);
nor U8444 (N_8444,N_7971,N_7647);
nor U8445 (N_8445,N_7893,N_7542);
xor U8446 (N_8446,N_7651,N_7768);
and U8447 (N_8447,N_7946,N_7793);
xnor U8448 (N_8448,N_7947,N_7815);
xor U8449 (N_8449,N_7619,N_7663);
xor U8450 (N_8450,N_7939,N_7739);
nand U8451 (N_8451,N_7622,N_7973);
nor U8452 (N_8452,N_7921,N_7887);
and U8453 (N_8453,N_7644,N_7533);
nand U8454 (N_8454,N_7609,N_7639);
nand U8455 (N_8455,N_7913,N_7756);
nand U8456 (N_8456,N_7504,N_7862);
xnor U8457 (N_8457,N_7872,N_7702);
or U8458 (N_8458,N_7930,N_7766);
xor U8459 (N_8459,N_7828,N_7943);
nor U8460 (N_8460,N_7584,N_7877);
nand U8461 (N_8461,N_7784,N_7643);
and U8462 (N_8462,N_7927,N_7589);
nor U8463 (N_8463,N_7917,N_7836);
xor U8464 (N_8464,N_7944,N_7937);
nor U8465 (N_8465,N_7512,N_7713);
nand U8466 (N_8466,N_7618,N_7607);
nor U8467 (N_8467,N_7777,N_7851);
xor U8468 (N_8468,N_7906,N_7884);
nand U8469 (N_8469,N_7928,N_7669);
nor U8470 (N_8470,N_7792,N_7652);
nor U8471 (N_8471,N_7908,N_7666);
and U8472 (N_8472,N_7673,N_7975);
xor U8473 (N_8473,N_7617,N_7659);
and U8474 (N_8474,N_7843,N_7737);
nor U8475 (N_8475,N_7571,N_7564);
xnor U8476 (N_8476,N_7987,N_7765);
xor U8477 (N_8477,N_7813,N_7879);
nor U8478 (N_8478,N_7949,N_7649);
nand U8479 (N_8479,N_7644,N_7899);
or U8480 (N_8480,N_7909,N_7639);
or U8481 (N_8481,N_7512,N_7859);
or U8482 (N_8482,N_7668,N_7510);
xor U8483 (N_8483,N_7502,N_7850);
nand U8484 (N_8484,N_7522,N_7548);
xnor U8485 (N_8485,N_7653,N_7616);
and U8486 (N_8486,N_7597,N_7512);
or U8487 (N_8487,N_7967,N_7629);
and U8488 (N_8488,N_7650,N_7725);
nor U8489 (N_8489,N_7998,N_7970);
or U8490 (N_8490,N_7728,N_7860);
nor U8491 (N_8491,N_7997,N_7747);
nor U8492 (N_8492,N_7549,N_7543);
and U8493 (N_8493,N_7871,N_7587);
nand U8494 (N_8494,N_7544,N_7850);
nand U8495 (N_8495,N_7815,N_7994);
xor U8496 (N_8496,N_7744,N_7675);
xor U8497 (N_8497,N_7959,N_7901);
nand U8498 (N_8498,N_7919,N_7731);
xnor U8499 (N_8499,N_7612,N_7914);
and U8500 (N_8500,N_8177,N_8152);
nor U8501 (N_8501,N_8275,N_8041);
or U8502 (N_8502,N_8425,N_8002);
nor U8503 (N_8503,N_8304,N_8208);
nor U8504 (N_8504,N_8324,N_8056);
xor U8505 (N_8505,N_8154,N_8243);
nor U8506 (N_8506,N_8082,N_8386);
and U8507 (N_8507,N_8471,N_8367);
and U8508 (N_8508,N_8405,N_8232);
or U8509 (N_8509,N_8224,N_8058);
xor U8510 (N_8510,N_8246,N_8266);
xor U8511 (N_8511,N_8113,N_8206);
nand U8512 (N_8512,N_8273,N_8179);
and U8513 (N_8513,N_8492,N_8043);
and U8514 (N_8514,N_8466,N_8066);
or U8515 (N_8515,N_8469,N_8358);
nand U8516 (N_8516,N_8401,N_8191);
xor U8517 (N_8517,N_8253,N_8472);
xor U8518 (N_8518,N_8139,N_8402);
nor U8519 (N_8519,N_8292,N_8215);
or U8520 (N_8520,N_8359,N_8408);
or U8521 (N_8521,N_8474,N_8393);
nand U8522 (N_8522,N_8352,N_8419);
or U8523 (N_8523,N_8268,N_8487);
nand U8524 (N_8524,N_8259,N_8388);
and U8525 (N_8525,N_8060,N_8403);
or U8526 (N_8526,N_8396,N_8025);
or U8527 (N_8527,N_8449,N_8257);
nor U8528 (N_8528,N_8483,N_8424);
and U8529 (N_8529,N_8081,N_8184);
nand U8530 (N_8530,N_8315,N_8018);
or U8531 (N_8531,N_8050,N_8176);
and U8532 (N_8532,N_8497,N_8410);
and U8533 (N_8533,N_8490,N_8046);
or U8534 (N_8534,N_8207,N_8128);
nand U8535 (N_8535,N_8124,N_8015);
nor U8536 (N_8536,N_8332,N_8105);
nand U8537 (N_8537,N_8014,N_8013);
nor U8538 (N_8538,N_8297,N_8432);
or U8539 (N_8539,N_8159,N_8282);
nor U8540 (N_8540,N_8052,N_8075);
and U8541 (N_8541,N_8193,N_8278);
nand U8542 (N_8542,N_8155,N_8328);
nand U8543 (N_8543,N_8296,N_8476);
nor U8544 (N_8544,N_8054,N_8493);
and U8545 (N_8545,N_8484,N_8173);
xor U8546 (N_8546,N_8236,N_8106);
xnor U8547 (N_8547,N_8494,N_8016);
nor U8548 (N_8548,N_8241,N_8134);
xor U8549 (N_8549,N_8488,N_8391);
and U8550 (N_8550,N_8026,N_8376);
nor U8551 (N_8551,N_8011,N_8109);
nor U8552 (N_8552,N_8486,N_8069);
or U8553 (N_8553,N_8242,N_8086);
or U8554 (N_8554,N_8335,N_8024);
xor U8555 (N_8555,N_8100,N_8143);
nor U8556 (N_8556,N_8028,N_8174);
and U8557 (N_8557,N_8097,N_8355);
and U8558 (N_8558,N_8196,N_8204);
and U8559 (N_8559,N_8053,N_8478);
or U8560 (N_8560,N_8438,N_8460);
and U8561 (N_8561,N_8032,N_8063);
or U8562 (N_8562,N_8265,N_8140);
and U8563 (N_8563,N_8162,N_8192);
nor U8564 (N_8564,N_8302,N_8399);
nor U8565 (N_8565,N_8225,N_8163);
or U8566 (N_8566,N_8481,N_8338);
and U8567 (N_8567,N_8112,N_8446);
and U8568 (N_8568,N_8345,N_8299);
and U8569 (N_8569,N_8444,N_8330);
nor U8570 (N_8570,N_8489,N_8339);
xnor U8571 (N_8571,N_8360,N_8049);
or U8572 (N_8572,N_8323,N_8256);
nor U8573 (N_8573,N_8379,N_8167);
xnor U8574 (N_8574,N_8012,N_8228);
or U8575 (N_8575,N_8385,N_8321);
and U8576 (N_8576,N_8437,N_8305);
nor U8577 (N_8577,N_8217,N_8411);
and U8578 (N_8578,N_8423,N_8337);
and U8579 (N_8579,N_8095,N_8384);
xnor U8580 (N_8580,N_8482,N_8125);
nand U8581 (N_8581,N_8465,N_8222);
or U8582 (N_8582,N_8318,N_8198);
and U8583 (N_8583,N_8142,N_8205);
nor U8584 (N_8584,N_8145,N_8477);
and U8585 (N_8585,N_8195,N_8034);
nand U8586 (N_8586,N_8132,N_8348);
and U8587 (N_8587,N_8413,N_8197);
or U8588 (N_8588,N_8104,N_8291);
nor U8589 (N_8589,N_8447,N_8277);
nand U8590 (N_8590,N_8096,N_8290);
nor U8591 (N_8591,N_8064,N_8189);
xor U8592 (N_8592,N_8361,N_8045);
xor U8593 (N_8593,N_8209,N_8303);
nor U8594 (N_8594,N_8051,N_8480);
xor U8595 (N_8595,N_8312,N_8036);
xor U8596 (N_8596,N_8087,N_8168);
nand U8597 (N_8597,N_8107,N_8074);
and U8598 (N_8598,N_8377,N_8461);
nor U8599 (N_8599,N_8216,N_8427);
and U8600 (N_8600,N_8230,N_8412);
or U8601 (N_8601,N_8366,N_8457);
xor U8602 (N_8602,N_8071,N_8240);
or U8603 (N_8603,N_8153,N_8048);
nand U8604 (N_8604,N_8395,N_8373);
nor U8605 (N_8605,N_8283,N_8426);
xor U8606 (N_8606,N_8300,N_8033);
and U8607 (N_8607,N_8227,N_8148);
and U8608 (N_8608,N_8294,N_8418);
xor U8609 (N_8609,N_8059,N_8115);
and U8610 (N_8610,N_8284,N_8429);
xnor U8611 (N_8611,N_8185,N_8170);
and U8612 (N_8612,N_8433,N_8430);
xor U8613 (N_8613,N_8138,N_8368);
nor U8614 (N_8614,N_8378,N_8310);
and U8615 (N_8615,N_8311,N_8101);
nand U8616 (N_8616,N_8149,N_8194);
or U8617 (N_8617,N_8234,N_8037);
nand U8618 (N_8618,N_8350,N_8289);
xor U8619 (N_8619,N_8003,N_8091);
nor U8620 (N_8620,N_8004,N_8307);
and U8621 (N_8621,N_8027,N_8450);
or U8622 (N_8622,N_8021,N_8213);
or U8623 (N_8623,N_8333,N_8264);
or U8624 (N_8624,N_8130,N_8250);
nor U8625 (N_8625,N_8374,N_8137);
xnor U8626 (N_8626,N_8462,N_8431);
or U8627 (N_8627,N_8214,N_8279);
nor U8628 (N_8628,N_8070,N_8351);
xnor U8629 (N_8629,N_8404,N_8409);
or U8630 (N_8630,N_8165,N_8342);
xor U8631 (N_8631,N_8231,N_8147);
nand U8632 (N_8632,N_8455,N_8319);
xnor U8633 (N_8633,N_8201,N_8006);
xor U8634 (N_8634,N_8084,N_8451);
nor U8635 (N_8635,N_8326,N_8267);
and U8636 (N_8636,N_8336,N_8357);
xor U8637 (N_8637,N_8463,N_8262);
nor U8638 (N_8638,N_8072,N_8181);
nor U8639 (N_8639,N_8007,N_8245);
and U8640 (N_8640,N_8442,N_8023);
nand U8641 (N_8641,N_8369,N_8394);
xnor U8642 (N_8642,N_8479,N_8102);
nor U8643 (N_8643,N_8334,N_8382);
and U8644 (N_8644,N_8317,N_8035);
xnor U8645 (N_8645,N_8190,N_8151);
and U8646 (N_8646,N_8172,N_8473);
and U8647 (N_8647,N_8079,N_8235);
nor U8648 (N_8648,N_8040,N_8276);
xor U8649 (N_8649,N_8364,N_8448);
nor U8650 (N_8650,N_8067,N_8083);
xor U8651 (N_8651,N_8322,N_8252);
and U8652 (N_8652,N_8178,N_8415);
nand U8653 (N_8653,N_8491,N_8363);
or U8654 (N_8654,N_8287,N_8237);
or U8655 (N_8655,N_8212,N_8171);
nor U8656 (N_8656,N_8116,N_8261);
nand U8657 (N_8657,N_8325,N_8436);
and U8658 (N_8658,N_8248,N_8254);
nor U8659 (N_8659,N_8362,N_8293);
and U8660 (N_8660,N_8114,N_8440);
xor U8661 (N_8661,N_8380,N_8038);
xor U8662 (N_8662,N_8249,N_8286);
or U8663 (N_8663,N_8183,N_8009);
or U8664 (N_8664,N_8136,N_8270);
or U8665 (N_8665,N_8314,N_8498);
and U8666 (N_8666,N_8406,N_8202);
and U8667 (N_8667,N_8187,N_8200);
nand U8668 (N_8668,N_8381,N_8309);
xor U8669 (N_8669,N_8061,N_8397);
nor U8670 (N_8670,N_8306,N_8169);
nor U8671 (N_8671,N_8030,N_8094);
xor U8672 (N_8672,N_8260,N_8467);
xnor U8673 (N_8673,N_8416,N_8435);
xnor U8674 (N_8674,N_8042,N_8468);
and U8675 (N_8675,N_8392,N_8226);
nand U8676 (N_8676,N_8131,N_8055);
and U8677 (N_8677,N_8099,N_8400);
xnor U8678 (N_8678,N_8017,N_8414);
nor U8679 (N_8679,N_8085,N_8039);
and U8680 (N_8680,N_8499,N_8271);
xnor U8681 (N_8681,N_8164,N_8077);
or U8682 (N_8682,N_8120,N_8475);
nand U8683 (N_8683,N_8166,N_8210);
and U8684 (N_8684,N_8221,N_8090);
nand U8685 (N_8685,N_8135,N_8141);
nand U8686 (N_8686,N_8223,N_8255);
or U8687 (N_8687,N_8288,N_8441);
and U8688 (N_8688,N_8047,N_8272);
nand U8689 (N_8689,N_8160,N_8371);
xor U8690 (N_8690,N_8119,N_8301);
or U8691 (N_8691,N_8126,N_8496);
nor U8692 (N_8692,N_8244,N_8133);
nand U8693 (N_8693,N_8459,N_8199);
xnor U8694 (N_8694,N_8108,N_8111);
nand U8695 (N_8695,N_8331,N_8239);
xor U8696 (N_8696,N_8220,N_8110);
nor U8697 (N_8697,N_8356,N_8129);
or U8698 (N_8698,N_8158,N_8383);
nor U8699 (N_8699,N_8073,N_8103);
nor U8700 (N_8700,N_8057,N_8062);
nand U8701 (N_8701,N_8127,N_8161);
xor U8702 (N_8702,N_8452,N_8421);
or U8703 (N_8703,N_8233,N_8398);
or U8704 (N_8704,N_8008,N_8445);
nor U8705 (N_8705,N_8485,N_8258);
nor U8706 (N_8706,N_8005,N_8370);
or U8707 (N_8707,N_8443,N_8280);
xor U8708 (N_8708,N_8019,N_8247);
or U8709 (N_8709,N_8022,N_8308);
and U8710 (N_8710,N_8353,N_8347);
nor U8711 (N_8711,N_8121,N_8313);
xnor U8712 (N_8712,N_8001,N_8274);
nand U8713 (N_8713,N_8375,N_8117);
nand U8714 (N_8714,N_8320,N_8218);
nor U8715 (N_8715,N_8219,N_8118);
xnor U8716 (N_8716,N_8080,N_8093);
nor U8717 (N_8717,N_8044,N_8495);
xor U8718 (N_8718,N_8407,N_8156);
xor U8719 (N_8719,N_8175,N_8341);
nand U8720 (N_8720,N_8456,N_8417);
and U8721 (N_8721,N_8365,N_8150);
or U8722 (N_8722,N_8010,N_8470);
or U8723 (N_8723,N_8068,N_8434);
nor U8724 (N_8724,N_8186,N_8316);
nor U8725 (N_8725,N_8180,N_8029);
nand U8726 (N_8726,N_8387,N_8182);
xor U8727 (N_8727,N_8089,N_8065);
xnor U8728 (N_8728,N_8340,N_8123);
xnor U8729 (N_8729,N_8203,N_8251);
nand U8730 (N_8730,N_8454,N_8343);
and U8731 (N_8731,N_8098,N_8000);
nand U8732 (N_8732,N_8211,N_8031);
nand U8733 (N_8733,N_8020,N_8144);
nand U8734 (N_8734,N_8092,N_8389);
and U8735 (N_8735,N_8088,N_8188);
and U8736 (N_8736,N_8439,N_8146);
xnor U8737 (N_8737,N_8229,N_8428);
nor U8738 (N_8738,N_8458,N_8329);
and U8739 (N_8739,N_8238,N_8327);
xnor U8740 (N_8740,N_8464,N_8281);
nand U8741 (N_8741,N_8372,N_8422);
nor U8742 (N_8742,N_8346,N_8122);
nor U8743 (N_8743,N_8298,N_8157);
and U8744 (N_8744,N_8295,N_8354);
or U8745 (N_8745,N_8349,N_8285);
or U8746 (N_8746,N_8263,N_8076);
or U8747 (N_8747,N_8390,N_8453);
xor U8748 (N_8748,N_8078,N_8420);
or U8749 (N_8749,N_8344,N_8269);
and U8750 (N_8750,N_8069,N_8021);
and U8751 (N_8751,N_8363,N_8160);
nor U8752 (N_8752,N_8475,N_8366);
nand U8753 (N_8753,N_8016,N_8089);
nor U8754 (N_8754,N_8081,N_8458);
nor U8755 (N_8755,N_8164,N_8171);
nand U8756 (N_8756,N_8027,N_8406);
xnor U8757 (N_8757,N_8110,N_8071);
nor U8758 (N_8758,N_8183,N_8070);
nand U8759 (N_8759,N_8023,N_8464);
nor U8760 (N_8760,N_8272,N_8005);
or U8761 (N_8761,N_8157,N_8100);
or U8762 (N_8762,N_8184,N_8270);
nand U8763 (N_8763,N_8484,N_8416);
or U8764 (N_8764,N_8402,N_8460);
and U8765 (N_8765,N_8143,N_8164);
and U8766 (N_8766,N_8421,N_8478);
nor U8767 (N_8767,N_8454,N_8310);
or U8768 (N_8768,N_8262,N_8374);
nand U8769 (N_8769,N_8327,N_8159);
nand U8770 (N_8770,N_8448,N_8479);
xnor U8771 (N_8771,N_8444,N_8306);
nor U8772 (N_8772,N_8168,N_8029);
nor U8773 (N_8773,N_8139,N_8034);
and U8774 (N_8774,N_8101,N_8365);
nand U8775 (N_8775,N_8408,N_8400);
xor U8776 (N_8776,N_8301,N_8026);
xnor U8777 (N_8777,N_8183,N_8373);
and U8778 (N_8778,N_8378,N_8140);
nor U8779 (N_8779,N_8167,N_8361);
or U8780 (N_8780,N_8128,N_8413);
xor U8781 (N_8781,N_8168,N_8131);
nand U8782 (N_8782,N_8223,N_8363);
or U8783 (N_8783,N_8475,N_8221);
or U8784 (N_8784,N_8032,N_8319);
or U8785 (N_8785,N_8130,N_8236);
nor U8786 (N_8786,N_8294,N_8212);
nand U8787 (N_8787,N_8242,N_8022);
nor U8788 (N_8788,N_8452,N_8028);
or U8789 (N_8789,N_8201,N_8291);
nor U8790 (N_8790,N_8327,N_8354);
or U8791 (N_8791,N_8264,N_8108);
or U8792 (N_8792,N_8357,N_8044);
nand U8793 (N_8793,N_8211,N_8179);
nor U8794 (N_8794,N_8281,N_8048);
xor U8795 (N_8795,N_8447,N_8477);
or U8796 (N_8796,N_8276,N_8139);
nand U8797 (N_8797,N_8085,N_8213);
and U8798 (N_8798,N_8285,N_8484);
xnor U8799 (N_8799,N_8130,N_8379);
and U8800 (N_8800,N_8049,N_8083);
and U8801 (N_8801,N_8489,N_8103);
xor U8802 (N_8802,N_8180,N_8145);
and U8803 (N_8803,N_8083,N_8284);
and U8804 (N_8804,N_8356,N_8459);
or U8805 (N_8805,N_8383,N_8394);
and U8806 (N_8806,N_8249,N_8025);
xnor U8807 (N_8807,N_8103,N_8497);
xor U8808 (N_8808,N_8028,N_8495);
and U8809 (N_8809,N_8492,N_8351);
nand U8810 (N_8810,N_8178,N_8296);
nor U8811 (N_8811,N_8357,N_8237);
nand U8812 (N_8812,N_8240,N_8213);
and U8813 (N_8813,N_8299,N_8315);
or U8814 (N_8814,N_8163,N_8099);
and U8815 (N_8815,N_8048,N_8101);
and U8816 (N_8816,N_8236,N_8274);
and U8817 (N_8817,N_8485,N_8087);
xnor U8818 (N_8818,N_8291,N_8305);
or U8819 (N_8819,N_8070,N_8153);
nand U8820 (N_8820,N_8225,N_8145);
nand U8821 (N_8821,N_8310,N_8356);
or U8822 (N_8822,N_8015,N_8182);
nor U8823 (N_8823,N_8011,N_8226);
nor U8824 (N_8824,N_8321,N_8352);
nor U8825 (N_8825,N_8013,N_8117);
and U8826 (N_8826,N_8298,N_8141);
or U8827 (N_8827,N_8311,N_8002);
or U8828 (N_8828,N_8242,N_8255);
or U8829 (N_8829,N_8377,N_8436);
xor U8830 (N_8830,N_8022,N_8064);
or U8831 (N_8831,N_8087,N_8293);
or U8832 (N_8832,N_8278,N_8124);
nand U8833 (N_8833,N_8432,N_8034);
nor U8834 (N_8834,N_8289,N_8380);
xor U8835 (N_8835,N_8182,N_8478);
and U8836 (N_8836,N_8009,N_8177);
xor U8837 (N_8837,N_8073,N_8459);
xor U8838 (N_8838,N_8067,N_8137);
nand U8839 (N_8839,N_8482,N_8189);
nand U8840 (N_8840,N_8203,N_8468);
xor U8841 (N_8841,N_8369,N_8017);
and U8842 (N_8842,N_8339,N_8290);
nand U8843 (N_8843,N_8345,N_8026);
and U8844 (N_8844,N_8252,N_8019);
and U8845 (N_8845,N_8471,N_8094);
or U8846 (N_8846,N_8128,N_8047);
and U8847 (N_8847,N_8430,N_8382);
or U8848 (N_8848,N_8312,N_8488);
nand U8849 (N_8849,N_8067,N_8471);
or U8850 (N_8850,N_8119,N_8261);
nor U8851 (N_8851,N_8119,N_8453);
nor U8852 (N_8852,N_8052,N_8285);
nor U8853 (N_8853,N_8043,N_8405);
nor U8854 (N_8854,N_8177,N_8164);
or U8855 (N_8855,N_8369,N_8140);
nor U8856 (N_8856,N_8069,N_8308);
nor U8857 (N_8857,N_8145,N_8196);
xor U8858 (N_8858,N_8200,N_8089);
and U8859 (N_8859,N_8015,N_8418);
nand U8860 (N_8860,N_8354,N_8000);
xnor U8861 (N_8861,N_8466,N_8452);
or U8862 (N_8862,N_8237,N_8174);
and U8863 (N_8863,N_8106,N_8193);
or U8864 (N_8864,N_8246,N_8265);
or U8865 (N_8865,N_8213,N_8242);
or U8866 (N_8866,N_8051,N_8060);
nand U8867 (N_8867,N_8062,N_8209);
nand U8868 (N_8868,N_8211,N_8363);
or U8869 (N_8869,N_8356,N_8471);
nand U8870 (N_8870,N_8128,N_8466);
and U8871 (N_8871,N_8394,N_8291);
nand U8872 (N_8872,N_8447,N_8042);
xor U8873 (N_8873,N_8248,N_8152);
or U8874 (N_8874,N_8369,N_8356);
xor U8875 (N_8875,N_8413,N_8210);
nor U8876 (N_8876,N_8440,N_8310);
nand U8877 (N_8877,N_8374,N_8154);
xor U8878 (N_8878,N_8170,N_8404);
nor U8879 (N_8879,N_8154,N_8142);
or U8880 (N_8880,N_8420,N_8442);
nor U8881 (N_8881,N_8387,N_8395);
or U8882 (N_8882,N_8408,N_8397);
or U8883 (N_8883,N_8121,N_8079);
xnor U8884 (N_8884,N_8478,N_8134);
or U8885 (N_8885,N_8010,N_8267);
xor U8886 (N_8886,N_8088,N_8487);
nand U8887 (N_8887,N_8130,N_8406);
or U8888 (N_8888,N_8010,N_8158);
and U8889 (N_8889,N_8358,N_8082);
and U8890 (N_8890,N_8293,N_8185);
nor U8891 (N_8891,N_8095,N_8197);
or U8892 (N_8892,N_8005,N_8418);
nand U8893 (N_8893,N_8024,N_8215);
nor U8894 (N_8894,N_8119,N_8345);
nor U8895 (N_8895,N_8350,N_8474);
and U8896 (N_8896,N_8399,N_8059);
and U8897 (N_8897,N_8436,N_8246);
nor U8898 (N_8898,N_8057,N_8275);
xnor U8899 (N_8899,N_8181,N_8404);
or U8900 (N_8900,N_8361,N_8264);
nor U8901 (N_8901,N_8131,N_8144);
and U8902 (N_8902,N_8402,N_8201);
xnor U8903 (N_8903,N_8200,N_8004);
nor U8904 (N_8904,N_8330,N_8033);
and U8905 (N_8905,N_8135,N_8136);
and U8906 (N_8906,N_8091,N_8220);
nor U8907 (N_8907,N_8130,N_8145);
or U8908 (N_8908,N_8385,N_8340);
and U8909 (N_8909,N_8389,N_8442);
nor U8910 (N_8910,N_8092,N_8460);
and U8911 (N_8911,N_8285,N_8323);
or U8912 (N_8912,N_8076,N_8258);
xnor U8913 (N_8913,N_8333,N_8430);
or U8914 (N_8914,N_8031,N_8167);
nand U8915 (N_8915,N_8147,N_8036);
or U8916 (N_8916,N_8063,N_8112);
nand U8917 (N_8917,N_8277,N_8063);
or U8918 (N_8918,N_8145,N_8021);
nand U8919 (N_8919,N_8377,N_8240);
nor U8920 (N_8920,N_8068,N_8204);
and U8921 (N_8921,N_8047,N_8242);
nand U8922 (N_8922,N_8114,N_8312);
or U8923 (N_8923,N_8207,N_8472);
and U8924 (N_8924,N_8205,N_8328);
and U8925 (N_8925,N_8439,N_8086);
nand U8926 (N_8926,N_8330,N_8406);
nand U8927 (N_8927,N_8420,N_8111);
nor U8928 (N_8928,N_8269,N_8499);
and U8929 (N_8929,N_8222,N_8236);
nor U8930 (N_8930,N_8369,N_8111);
xor U8931 (N_8931,N_8236,N_8047);
nor U8932 (N_8932,N_8094,N_8392);
nand U8933 (N_8933,N_8112,N_8183);
or U8934 (N_8934,N_8325,N_8400);
xnor U8935 (N_8935,N_8382,N_8201);
nor U8936 (N_8936,N_8151,N_8092);
and U8937 (N_8937,N_8029,N_8491);
and U8938 (N_8938,N_8204,N_8417);
nor U8939 (N_8939,N_8362,N_8265);
and U8940 (N_8940,N_8238,N_8046);
xnor U8941 (N_8941,N_8003,N_8426);
nand U8942 (N_8942,N_8445,N_8329);
nor U8943 (N_8943,N_8375,N_8163);
nand U8944 (N_8944,N_8205,N_8414);
or U8945 (N_8945,N_8392,N_8447);
nand U8946 (N_8946,N_8316,N_8430);
nor U8947 (N_8947,N_8118,N_8426);
xnor U8948 (N_8948,N_8487,N_8499);
nand U8949 (N_8949,N_8275,N_8410);
nor U8950 (N_8950,N_8032,N_8422);
xor U8951 (N_8951,N_8043,N_8061);
nand U8952 (N_8952,N_8372,N_8055);
and U8953 (N_8953,N_8075,N_8110);
or U8954 (N_8954,N_8387,N_8009);
or U8955 (N_8955,N_8351,N_8265);
nand U8956 (N_8956,N_8092,N_8230);
nor U8957 (N_8957,N_8257,N_8245);
xor U8958 (N_8958,N_8333,N_8002);
xor U8959 (N_8959,N_8167,N_8001);
nor U8960 (N_8960,N_8036,N_8175);
nand U8961 (N_8961,N_8152,N_8093);
or U8962 (N_8962,N_8209,N_8147);
nor U8963 (N_8963,N_8310,N_8434);
and U8964 (N_8964,N_8411,N_8104);
nand U8965 (N_8965,N_8306,N_8043);
nor U8966 (N_8966,N_8269,N_8049);
or U8967 (N_8967,N_8364,N_8238);
xor U8968 (N_8968,N_8354,N_8254);
nor U8969 (N_8969,N_8236,N_8084);
nor U8970 (N_8970,N_8156,N_8050);
xor U8971 (N_8971,N_8496,N_8401);
and U8972 (N_8972,N_8267,N_8087);
nand U8973 (N_8973,N_8397,N_8077);
and U8974 (N_8974,N_8330,N_8341);
and U8975 (N_8975,N_8022,N_8101);
nand U8976 (N_8976,N_8425,N_8271);
nand U8977 (N_8977,N_8045,N_8228);
nor U8978 (N_8978,N_8329,N_8241);
and U8979 (N_8979,N_8177,N_8157);
nor U8980 (N_8980,N_8190,N_8335);
and U8981 (N_8981,N_8191,N_8153);
nand U8982 (N_8982,N_8194,N_8293);
nand U8983 (N_8983,N_8308,N_8447);
nor U8984 (N_8984,N_8144,N_8068);
xnor U8985 (N_8985,N_8250,N_8349);
nor U8986 (N_8986,N_8130,N_8154);
nand U8987 (N_8987,N_8438,N_8446);
xnor U8988 (N_8988,N_8217,N_8214);
and U8989 (N_8989,N_8365,N_8431);
or U8990 (N_8990,N_8482,N_8386);
xnor U8991 (N_8991,N_8010,N_8004);
nand U8992 (N_8992,N_8482,N_8342);
xnor U8993 (N_8993,N_8449,N_8347);
nor U8994 (N_8994,N_8285,N_8321);
nor U8995 (N_8995,N_8243,N_8098);
or U8996 (N_8996,N_8021,N_8066);
xnor U8997 (N_8997,N_8199,N_8294);
nand U8998 (N_8998,N_8164,N_8334);
or U8999 (N_8999,N_8443,N_8079);
nor U9000 (N_9000,N_8988,N_8511);
nor U9001 (N_9001,N_8981,N_8648);
and U9002 (N_9002,N_8880,N_8793);
nand U9003 (N_9003,N_8791,N_8612);
or U9004 (N_9004,N_8918,N_8805);
and U9005 (N_9005,N_8811,N_8937);
nor U9006 (N_9006,N_8570,N_8550);
nor U9007 (N_9007,N_8650,N_8777);
xnor U9008 (N_9008,N_8951,N_8718);
xnor U9009 (N_9009,N_8902,N_8929);
nor U9010 (N_9010,N_8606,N_8690);
or U9011 (N_9011,N_8595,N_8979);
xnor U9012 (N_9012,N_8700,N_8667);
and U9013 (N_9013,N_8707,N_8614);
or U9014 (N_9014,N_8655,N_8582);
or U9015 (N_9015,N_8523,N_8626);
nor U9016 (N_9016,N_8741,N_8512);
xor U9017 (N_9017,N_8543,N_8869);
and U9018 (N_9018,N_8607,N_8592);
xor U9019 (N_9019,N_8864,N_8965);
xnor U9020 (N_9020,N_8740,N_8598);
xor U9021 (N_9021,N_8708,N_8632);
or U9022 (N_9022,N_8733,N_8526);
and U9023 (N_9023,N_8802,N_8602);
or U9024 (N_9024,N_8853,N_8693);
and U9025 (N_9025,N_8521,N_8985);
nor U9026 (N_9026,N_8503,N_8754);
nor U9027 (N_9027,N_8509,N_8686);
xnor U9028 (N_9028,N_8987,N_8610);
xor U9029 (N_9029,N_8536,N_8659);
and U9030 (N_9030,N_8775,N_8574);
nand U9031 (N_9031,N_8761,N_8613);
xor U9032 (N_9032,N_8975,N_8564);
or U9033 (N_9033,N_8871,N_8563);
nor U9034 (N_9034,N_8720,N_8890);
and U9035 (N_9035,N_8762,N_8962);
xnor U9036 (N_9036,N_8580,N_8846);
nand U9037 (N_9037,N_8750,N_8668);
or U9038 (N_9038,N_8824,N_8528);
xor U9039 (N_9039,N_8591,N_8830);
or U9040 (N_9040,N_8784,N_8891);
and U9041 (N_9041,N_8866,N_8976);
or U9042 (N_9042,N_8944,N_8851);
or U9043 (N_9043,N_8705,N_8674);
and U9044 (N_9044,N_8692,N_8605);
nor U9045 (N_9045,N_8687,N_8747);
or U9046 (N_9046,N_8875,N_8813);
or U9047 (N_9047,N_8788,N_8816);
nor U9048 (N_9048,N_8546,N_8689);
nor U9049 (N_9049,N_8798,N_8653);
nor U9050 (N_9050,N_8746,N_8756);
and U9051 (N_9051,N_8801,N_8664);
nor U9052 (N_9052,N_8934,N_8993);
nand U9053 (N_9053,N_8537,N_8734);
xnor U9054 (N_9054,N_8634,N_8938);
nor U9055 (N_9055,N_8507,N_8919);
nand U9056 (N_9056,N_8646,N_8883);
xor U9057 (N_9057,N_8859,N_8948);
xor U9058 (N_9058,N_8994,N_8547);
or U9059 (N_9059,N_8554,N_8638);
xor U9060 (N_9060,N_8773,N_8709);
and U9061 (N_9061,N_8514,N_8921);
xor U9062 (N_9062,N_8819,N_8909);
or U9063 (N_9063,N_8889,N_8861);
xnor U9064 (N_9064,N_8518,N_8831);
xor U9065 (N_9065,N_8516,N_8914);
xnor U9066 (N_9066,N_8963,N_8641);
or U9067 (N_9067,N_8986,N_8669);
or U9068 (N_9068,N_8770,N_8779);
nor U9069 (N_9069,N_8695,N_8753);
nand U9070 (N_9070,N_8749,N_8623);
nor U9071 (N_9071,N_8942,N_8658);
nand U9072 (N_9072,N_8797,N_8678);
nand U9073 (N_9073,N_8862,N_8730);
nand U9074 (N_9074,N_8619,N_8844);
nand U9075 (N_9075,N_8616,N_8959);
nor U9076 (N_9076,N_8699,N_8631);
nor U9077 (N_9077,N_8838,N_8928);
nor U9078 (N_9078,N_8854,N_8728);
xnor U9079 (N_9079,N_8529,N_8751);
nand U9080 (N_9080,N_8897,N_8812);
and U9081 (N_9081,N_8737,N_8727);
nand U9082 (N_9082,N_8715,N_8886);
or U9083 (N_9083,N_8552,N_8571);
or U9084 (N_9084,N_8738,N_8917);
nor U9085 (N_9085,N_8639,N_8532);
nand U9086 (N_9086,N_8684,N_8561);
or U9087 (N_9087,N_8827,N_8873);
and U9088 (N_9088,N_8787,N_8723);
xor U9089 (N_9089,N_8618,N_8654);
and U9090 (N_9090,N_8596,N_8763);
nand U9091 (N_9091,N_8611,N_8531);
or U9092 (N_9092,N_8501,N_8939);
and U9093 (N_9093,N_8755,N_8556);
nor U9094 (N_9094,N_8573,N_8599);
and U9095 (N_9095,N_8587,N_8725);
xnor U9096 (N_9096,N_8583,N_8600);
xnor U9097 (N_9097,N_8577,N_8878);
or U9098 (N_9098,N_8527,N_8841);
xor U9099 (N_9099,N_8872,N_8832);
nand U9100 (N_9100,N_8767,N_8783);
nor U9101 (N_9101,N_8683,N_8676);
or U9102 (N_9102,N_8506,N_8964);
nor U9103 (N_9103,N_8636,N_8999);
or U9104 (N_9104,N_8984,N_8885);
nand U9105 (N_9105,N_8776,N_8996);
xnor U9106 (N_9106,N_8597,N_8967);
and U9107 (N_9107,N_8881,N_8804);
nand U9108 (N_9108,N_8814,N_8818);
nand U9109 (N_9109,N_8931,N_8796);
xnor U9110 (N_9110,N_8911,N_8661);
and U9111 (N_9111,N_8799,N_8961);
xnor U9112 (N_9112,N_8926,N_8500);
xor U9113 (N_9113,N_8863,N_8562);
and U9114 (N_9114,N_8820,N_8877);
or U9115 (N_9115,N_8666,N_8588);
nor U9116 (N_9116,N_8644,N_8790);
and U9117 (N_9117,N_8657,N_8515);
nor U9118 (N_9118,N_8968,N_8551);
and U9119 (N_9119,N_8713,N_8893);
xnor U9120 (N_9120,N_8558,N_8946);
nor U9121 (N_9121,N_8795,N_8789);
xor U9122 (N_9122,N_8604,N_8696);
nand U9123 (N_9123,N_8620,N_8945);
or U9124 (N_9124,N_8978,N_8935);
nor U9125 (N_9125,N_8868,N_8855);
and U9126 (N_9126,N_8936,N_8807);
xnor U9127 (N_9127,N_8972,N_8982);
and U9128 (N_9128,N_8545,N_8698);
or U9129 (N_9129,N_8840,N_8849);
nand U9130 (N_9130,N_8731,N_8785);
nand U9131 (N_9131,N_8736,N_8956);
or U9132 (N_9132,N_8989,N_8764);
xor U9133 (N_9133,N_8835,N_8508);
nor U9134 (N_9134,N_8702,N_8739);
and U9135 (N_9135,N_8930,N_8879);
nor U9136 (N_9136,N_8697,N_8924);
nand U9137 (N_9137,N_8679,N_8581);
xnor U9138 (N_9138,N_8887,N_8670);
and U9139 (N_9139,N_8912,N_8960);
xnor U9140 (N_9140,N_8572,N_8806);
nand U9141 (N_9141,N_8933,N_8958);
nand U9142 (N_9142,N_8565,N_8694);
and U9143 (N_9143,N_8732,N_8520);
xnor U9144 (N_9144,N_8557,N_8898);
and U9145 (N_9145,N_8836,N_8766);
or U9146 (N_9146,N_8566,N_8624);
and U9147 (N_9147,N_8932,N_8900);
nand U9148 (N_9148,N_8637,N_8651);
nand U9149 (N_9149,N_8895,N_8765);
and U9150 (N_9150,N_8829,N_8821);
xnor U9151 (N_9151,N_8815,N_8759);
nand U9152 (N_9152,N_8874,N_8622);
nand U9153 (N_9153,N_8839,N_8778);
or U9154 (N_9154,N_8822,N_8711);
or U9155 (N_9155,N_8649,N_8534);
xnor U9156 (N_9156,N_8792,N_8717);
or U9157 (N_9157,N_8685,N_8539);
xnor U9158 (N_9158,N_8782,N_8943);
nand U9159 (N_9159,N_8615,N_8860);
and U9160 (N_9160,N_8843,N_8823);
nor U9161 (N_9161,N_8995,N_8513);
and U9162 (N_9162,N_8553,N_8952);
nand U9163 (N_9163,N_8721,N_8809);
nand U9164 (N_9164,N_8991,N_8575);
nand U9165 (N_9165,N_8896,N_8768);
or U9166 (N_9166,N_8983,N_8970);
nor U9167 (N_9167,N_8927,N_8538);
xnor U9168 (N_9168,N_8635,N_8633);
nand U9169 (N_9169,N_8842,N_8542);
or U9170 (N_9170,N_8876,N_8540);
nand U9171 (N_9171,N_8541,N_8502);
and U9172 (N_9172,N_8524,N_8781);
and U9173 (N_9173,N_8601,N_8560);
or U9174 (N_9174,N_8567,N_8856);
and U9175 (N_9175,N_8701,N_8817);
nand U9176 (N_9176,N_8857,N_8892);
xor U9177 (N_9177,N_8533,N_8957);
nor U9178 (N_9178,N_8691,N_8833);
and U9179 (N_9179,N_8771,N_8998);
or U9180 (N_9180,N_8729,N_8714);
and U9181 (N_9181,N_8559,N_8735);
and U9182 (N_9182,N_8904,N_8954);
nand U9183 (N_9183,N_8915,N_8555);
and U9184 (N_9184,N_8758,N_8640);
and U9185 (N_9185,N_8584,N_8745);
xor U9186 (N_9186,N_8774,N_8752);
and U9187 (N_9187,N_8847,N_8834);
or U9188 (N_9188,N_8971,N_8769);
or U9189 (N_9189,N_8744,N_8660);
nand U9190 (N_9190,N_8585,N_8953);
nor U9191 (N_9191,N_8922,N_8688);
or U9192 (N_9192,N_8969,N_8672);
nand U9193 (N_9193,N_8913,N_8716);
and U9194 (N_9194,N_8704,N_8579);
or U9195 (N_9195,N_8621,N_8617);
nor U9196 (N_9196,N_8949,N_8522);
xor U9197 (N_9197,N_8907,N_8642);
xor U9198 (N_9198,N_8882,N_8825);
xnor U9199 (N_9199,N_8663,N_8858);
xor U9200 (N_9200,N_8643,N_8955);
nand U9201 (N_9201,N_8525,N_8810);
nand U9202 (N_9202,N_8808,N_8505);
xor U9203 (N_9203,N_8517,N_8760);
nor U9204 (N_9204,N_8677,N_8594);
and U9205 (N_9205,N_8530,N_8837);
and U9206 (N_9206,N_8652,N_8923);
nand U9207 (N_9207,N_8608,N_8681);
or U9208 (N_9208,N_8504,N_8908);
nor U9209 (N_9209,N_8903,N_8916);
or U9210 (N_9210,N_8724,N_8780);
nand U9211 (N_9211,N_8675,N_8910);
nand U9212 (N_9212,N_8710,N_8680);
nor U9213 (N_9213,N_8625,N_8662);
nor U9214 (N_9214,N_8647,N_8974);
xor U9215 (N_9215,N_8800,N_8656);
nor U9216 (N_9216,N_8941,N_8609);
or U9217 (N_9217,N_8757,N_8899);
xnor U9218 (N_9218,N_8645,N_8845);
or U9219 (N_9219,N_8627,N_8884);
nor U9220 (N_9220,N_8726,N_8870);
xnor U9221 (N_9221,N_8803,N_8888);
nor U9222 (N_9222,N_8629,N_8671);
xor U9223 (N_9223,N_8865,N_8980);
nor U9224 (N_9224,N_8920,N_8925);
nand U9225 (N_9225,N_8990,N_8535);
or U9226 (N_9226,N_8786,N_8850);
or U9227 (N_9227,N_8894,N_8682);
and U9228 (N_9228,N_8510,N_8901);
xor U9229 (N_9229,N_8576,N_8544);
or U9230 (N_9230,N_8548,N_8603);
nand U9231 (N_9231,N_8519,N_8719);
nand U9232 (N_9232,N_8947,N_8748);
and U9233 (N_9233,N_8673,N_8589);
nand U9234 (N_9234,N_8549,N_8706);
xor U9235 (N_9235,N_8992,N_8940);
nor U9236 (N_9236,N_8578,N_8997);
and U9237 (N_9237,N_8772,N_8867);
xor U9238 (N_9238,N_8712,N_8665);
nand U9239 (N_9239,N_8628,N_8569);
and U9240 (N_9240,N_8966,N_8973);
and U9241 (N_9241,N_8848,N_8906);
and U9242 (N_9242,N_8826,N_8905);
or U9243 (N_9243,N_8852,N_8586);
or U9244 (N_9244,N_8703,N_8722);
nor U9245 (N_9245,N_8742,N_8977);
or U9246 (N_9246,N_8590,N_8568);
or U9247 (N_9247,N_8828,N_8794);
nand U9248 (N_9248,N_8630,N_8743);
nor U9249 (N_9249,N_8593,N_8950);
or U9250 (N_9250,N_8948,N_8758);
xnor U9251 (N_9251,N_8904,N_8759);
xor U9252 (N_9252,N_8796,N_8717);
nand U9253 (N_9253,N_8786,N_8897);
nor U9254 (N_9254,N_8854,N_8700);
nor U9255 (N_9255,N_8522,N_8755);
or U9256 (N_9256,N_8730,N_8867);
nand U9257 (N_9257,N_8769,N_8551);
or U9258 (N_9258,N_8612,N_8599);
nor U9259 (N_9259,N_8713,N_8985);
and U9260 (N_9260,N_8719,N_8829);
or U9261 (N_9261,N_8665,N_8605);
xor U9262 (N_9262,N_8576,N_8951);
xnor U9263 (N_9263,N_8612,N_8774);
nand U9264 (N_9264,N_8947,N_8725);
nand U9265 (N_9265,N_8601,N_8730);
nand U9266 (N_9266,N_8898,N_8786);
and U9267 (N_9267,N_8946,N_8679);
and U9268 (N_9268,N_8627,N_8785);
nor U9269 (N_9269,N_8639,N_8663);
nand U9270 (N_9270,N_8950,N_8764);
or U9271 (N_9271,N_8737,N_8608);
xnor U9272 (N_9272,N_8798,N_8680);
nor U9273 (N_9273,N_8720,N_8735);
xnor U9274 (N_9274,N_8713,N_8576);
and U9275 (N_9275,N_8619,N_8829);
xnor U9276 (N_9276,N_8743,N_8656);
nor U9277 (N_9277,N_8742,N_8705);
and U9278 (N_9278,N_8588,N_8820);
nand U9279 (N_9279,N_8794,N_8813);
or U9280 (N_9280,N_8638,N_8750);
nor U9281 (N_9281,N_8527,N_8639);
or U9282 (N_9282,N_8592,N_8502);
xnor U9283 (N_9283,N_8505,N_8674);
nand U9284 (N_9284,N_8564,N_8941);
and U9285 (N_9285,N_8679,N_8701);
nand U9286 (N_9286,N_8719,N_8598);
nor U9287 (N_9287,N_8564,N_8701);
xnor U9288 (N_9288,N_8509,N_8608);
xor U9289 (N_9289,N_8808,N_8854);
nand U9290 (N_9290,N_8537,N_8681);
or U9291 (N_9291,N_8700,N_8961);
nor U9292 (N_9292,N_8730,N_8690);
xor U9293 (N_9293,N_8546,N_8656);
and U9294 (N_9294,N_8930,N_8884);
and U9295 (N_9295,N_8619,N_8639);
or U9296 (N_9296,N_8840,N_8731);
and U9297 (N_9297,N_8814,N_8936);
and U9298 (N_9298,N_8539,N_8658);
xnor U9299 (N_9299,N_8883,N_8988);
nor U9300 (N_9300,N_8689,N_8743);
nand U9301 (N_9301,N_8900,N_8614);
or U9302 (N_9302,N_8536,N_8779);
or U9303 (N_9303,N_8944,N_8544);
xnor U9304 (N_9304,N_8828,N_8841);
xor U9305 (N_9305,N_8604,N_8965);
nand U9306 (N_9306,N_8660,N_8918);
and U9307 (N_9307,N_8994,N_8945);
nand U9308 (N_9308,N_8538,N_8544);
and U9309 (N_9309,N_8583,N_8851);
and U9310 (N_9310,N_8886,N_8942);
or U9311 (N_9311,N_8670,N_8651);
and U9312 (N_9312,N_8642,N_8661);
xnor U9313 (N_9313,N_8785,N_8994);
and U9314 (N_9314,N_8888,N_8604);
xnor U9315 (N_9315,N_8949,N_8927);
nand U9316 (N_9316,N_8799,N_8866);
nand U9317 (N_9317,N_8759,N_8649);
or U9318 (N_9318,N_8635,N_8772);
and U9319 (N_9319,N_8823,N_8606);
xnor U9320 (N_9320,N_8921,N_8911);
xor U9321 (N_9321,N_8890,N_8702);
or U9322 (N_9322,N_8873,N_8848);
nor U9323 (N_9323,N_8788,N_8605);
nand U9324 (N_9324,N_8891,N_8969);
and U9325 (N_9325,N_8546,N_8734);
nand U9326 (N_9326,N_8891,N_8874);
nand U9327 (N_9327,N_8556,N_8865);
nand U9328 (N_9328,N_8995,N_8778);
nand U9329 (N_9329,N_8699,N_8653);
nand U9330 (N_9330,N_8557,N_8952);
or U9331 (N_9331,N_8956,N_8702);
nor U9332 (N_9332,N_8917,N_8574);
nand U9333 (N_9333,N_8786,N_8509);
xnor U9334 (N_9334,N_8520,N_8836);
or U9335 (N_9335,N_8818,N_8657);
and U9336 (N_9336,N_8501,N_8641);
nor U9337 (N_9337,N_8713,N_8556);
xor U9338 (N_9338,N_8707,N_8916);
nand U9339 (N_9339,N_8539,N_8687);
or U9340 (N_9340,N_8845,N_8573);
nand U9341 (N_9341,N_8908,N_8812);
and U9342 (N_9342,N_8856,N_8811);
xor U9343 (N_9343,N_8590,N_8594);
or U9344 (N_9344,N_8663,N_8539);
and U9345 (N_9345,N_8752,N_8720);
xnor U9346 (N_9346,N_8992,N_8728);
or U9347 (N_9347,N_8765,N_8634);
nand U9348 (N_9348,N_8964,N_8670);
and U9349 (N_9349,N_8751,N_8637);
xnor U9350 (N_9350,N_8758,N_8731);
nor U9351 (N_9351,N_8586,N_8767);
or U9352 (N_9352,N_8632,N_8671);
or U9353 (N_9353,N_8998,N_8745);
nor U9354 (N_9354,N_8850,N_8875);
nor U9355 (N_9355,N_8772,N_8528);
xor U9356 (N_9356,N_8977,N_8806);
nor U9357 (N_9357,N_8754,N_8931);
or U9358 (N_9358,N_8596,N_8779);
or U9359 (N_9359,N_8645,N_8762);
and U9360 (N_9360,N_8586,N_8803);
xor U9361 (N_9361,N_8627,N_8943);
and U9362 (N_9362,N_8858,N_8547);
nor U9363 (N_9363,N_8876,N_8820);
nor U9364 (N_9364,N_8718,N_8822);
and U9365 (N_9365,N_8619,N_8520);
xnor U9366 (N_9366,N_8928,N_8987);
nor U9367 (N_9367,N_8900,N_8690);
or U9368 (N_9368,N_8950,N_8827);
xnor U9369 (N_9369,N_8511,N_8700);
and U9370 (N_9370,N_8838,N_8945);
nand U9371 (N_9371,N_8815,N_8605);
nor U9372 (N_9372,N_8672,N_8838);
nand U9373 (N_9373,N_8802,N_8827);
or U9374 (N_9374,N_8932,N_8911);
and U9375 (N_9375,N_8997,N_8651);
nor U9376 (N_9376,N_8913,N_8554);
and U9377 (N_9377,N_8831,N_8717);
xnor U9378 (N_9378,N_8972,N_8735);
xor U9379 (N_9379,N_8639,N_8807);
or U9380 (N_9380,N_8591,N_8923);
xnor U9381 (N_9381,N_8942,N_8835);
and U9382 (N_9382,N_8645,N_8932);
xnor U9383 (N_9383,N_8649,N_8655);
and U9384 (N_9384,N_8693,N_8570);
nand U9385 (N_9385,N_8925,N_8546);
nor U9386 (N_9386,N_8726,N_8909);
xor U9387 (N_9387,N_8990,N_8656);
or U9388 (N_9388,N_8504,N_8526);
or U9389 (N_9389,N_8522,N_8575);
nand U9390 (N_9390,N_8690,N_8863);
nand U9391 (N_9391,N_8646,N_8880);
or U9392 (N_9392,N_8996,N_8666);
xor U9393 (N_9393,N_8869,N_8934);
xnor U9394 (N_9394,N_8819,N_8970);
nor U9395 (N_9395,N_8896,N_8557);
xnor U9396 (N_9396,N_8660,N_8809);
xor U9397 (N_9397,N_8712,N_8895);
nand U9398 (N_9398,N_8971,N_8974);
nor U9399 (N_9399,N_8992,N_8526);
xor U9400 (N_9400,N_8674,N_8947);
nand U9401 (N_9401,N_8708,N_8962);
and U9402 (N_9402,N_8784,N_8838);
nor U9403 (N_9403,N_8853,N_8575);
nand U9404 (N_9404,N_8678,N_8682);
nor U9405 (N_9405,N_8925,N_8534);
nand U9406 (N_9406,N_8721,N_8734);
and U9407 (N_9407,N_8730,N_8815);
nand U9408 (N_9408,N_8885,N_8558);
xnor U9409 (N_9409,N_8511,N_8701);
nand U9410 (N_9410,N_8958,N_8658);
or U9411 (N_9411,N_8936,N_8674);
nor U9412 (N_9412,N_8559,N_8728);
nor U9413 (N_9413,N_8822,N_8906);
nor U9414 (N_9414,N_8780,N_8776);
xor U9415 (N_9415,N_8996,N_8661);
xor U9416 (N_9416,N_8769,N_8709);
nor U9417 (N_9417,N_8757,N_8959);
nor U9418 (N_9418,N_8686,N_8895);
or U9419 (N_9419,N_8583,N_8598);
or U9420 (N_9420,N_8631,N_8883);
and U9421 (N_9421,N_8733,N_8609);
or U9422 (N_9422,N_8611,N_8914);
and U9423 (N_9423,N_8646,N_8809);
or U9424 (N_9424,N_8610,N_8756);
and U9425 (N_9425,N_8628,N_8518);
nor U9426 (N_9426,N_8939,N_8753);
xor U9427 (N_9427,N_8768,N_8682);
or U9428 (N_9428,N_8861,N_8714);
nor U9429 (N_9429,N_8727,N_8547);
or U9430 (N_9430,N_8565,N_8648);
nor U9431 (N_9431,N_8567,N_8606);
xnor U9432 (N_9432,N_8983,N_8619);
nor U9433 (N_9433,N_8757,N_8812);
or U9434 (N_9434,N_8641,N_8819);
and U9435 (N_9435,N_8736,N_8582);
and U9436 (N_9436,N_8981,N_8730);
nor U9437 (N_9437,N_8918,N_8547);
xnor U9438 (N_9438,N_8613,N_8731);
or U9439 (N_9439,N_8581,N_8550);
and U9440 (N_9440,N_8919,N_8728);
and U9441 (N_9441,N_8568,N_8760);
and U9442 (N_9442,N_8523,N_8957);
and U9443 (N_9443,N_8814,N_8852);
xnor U9444 (N_9444,N_8992,N_8552);
and U9445 (N_9445,N_8767,N_8755);
xor U9446 (N_9446,N_8720,N_8946);
xnor U9447 (N_9447,N_8903,N_8530);
or U9448 (N_9448,N_8564,N_8860);
nand U9449 (N_9449,N_8592,N_8603);
and U9450 (N_9450,N_8644,N_8859);
xnor U9451 (N_9451,N_8532,N_8929);
xor U9452 (N_9452,N_8500,N_8643);
nand U9453 (N_9453,N_8847,N_8761);
nand U9454 (N_9454,N_8996,N_8893);
nor U9455 (N_9455,N_8530,N_8842);
nor U9456 (N_9456,N_8931,N_8762);
nor U9457 (N_9457,N_8993,N_8624);
xor U9458 (N_9458,N_8633,N_8759);
xnor U9459 (N_9459,N_8564,N_8824);
and U9460 (N_9460,N_8667,N_8773);
and U9461 (N_9461,N_8700,N_8680);
or U9462 (N_9462,N_8620,N_8662);
xor U9463 (N_9463,N_8591,N_8936);
or U9464 (N_9464,N_8527,N_8979);
xor U9465 (N_9465,N_8750,N_8945);
nand U9466 (N_9466,N_8969,N_8547);
nor U9467 (N_9467,N_8780,N_8700);
nor U9468 (N_9468,N_8903,N_8841);
and U9469 (N_9469,N_8813,N_8996);
and U9470 (N_9470,N_8887,N_8504);
xor U9471 (N_9471,N_8886,N_8884);
nand U9472 (N_9472,N_8776,N_8608);
nor U9473 (N_9473,N_8688,N_8701);
nand U9474 (N_9474,N_8906,N_8570);
nand U9475 (N_9475,N_8506,N_8610);
xor U9476 (N_9476,N_8609,N_8927);
or U9477 (N_9477,N_8979,N_8965);
or U9478 (N_9478,N_8791,N_8579);
and U9479 (N_9479,N_8594,N_8583);
or U9480 (N_9480,N_8945,N_8950);
nor U9481 (N_9481,N_8795,N_8769);
or U9482 (N_9482,N_8636,N_8909);
nand U9483 (N_9483,N_8702,N_8737);
xnor U9484 (N_9484,N_8598,N_8859);
or U9485 (N_9485,N_8985,N_8838);
and U9486 (N_9486,N_8807,N_8737);
nor U9487 (N_9487,N_8875,N_8712);
nand U9488 (N_9488,N_8563,N_8968);
nor U9489 (N_9489,N_8657,N_8622);
xor U9490 (N_9490,N_8963,N_8896);
nand U9491 (N_9491,N_8953,N_8932);
nor U9492 (N_9492,N_8694,N_8753);
or U9493 (N_9493,N_8810,N_8539);
nor U9494 (N_9494,N_8544,N_8503);
nor U9495 (N_9495,N_8751,N_8562);
and U9496 (N_9496,N_8905,N_8838);
nand U9497 (N_9497,N_8700,N_8804);
or U9498 (N_9498,N_8875,N_8537);
nor U9499 (N_9499,N_8807,N_8992);
and U9500 (N_9500,N_9328,N_9458);
and U9501 (N_9501,N_9412,N_9290);
or U9502 (N_9502,N_9184,N_9371);
nor U9503 (N_9503,N_9124,N_9359);
nor U9504 (N_9504,N_9122,N_9394);
nand U9505 (N_9505,N_9248,N_9486);
xor U9506 (N_9506,N_9396,N_9078);
xnor U9507 (N_9507,N_9188,N_9229);
nand U9508 (N_9508,N_9464,N_9120);
and U9509 (N_9509,N_9215,N_9024);
xnor U9510 (N_9510,N_9360,N_9468);
nand U9511 (N_9511,N_9212,N_9279);
and U9512 (N_9512,N_9146,N_9138);
xnor U9513 (N_9513,N_9071,N_9154);
nand U9514 (N_9514,N_9075,N_9079);
nor U9515 (N_9515,N_9128,N_9048);
nor U9516 (N_9516,N_9339,N_9186);
xnor U9517 (N_9517,N_9220,N_9352);
xor U9518 (N_9518,N_9305,N_9253);
nor U9519 (N_9519,N_9424,N_9281);
nand U9520 (N_9520,N_9152,N_9293);
xnor U9521 (N_9521,N_9441,N_9264);
xnor U9522 (N_9522,N_9145,N_9170);
nor U9523 (N_9523,N_9387,N_9002);
nand U9524 (N_9524,N_9289,N_9231);
nor U9525 (N_9525,N_9208,N_9066);
nand U9526 (N_9526,N_9378,N_9385);
or U9527 (N_9527,N_9337,N_9237);
xnor U9528 (N_9528,N_9295,N_9272);
xnor U9529 (N_9529,N_9038,N_9020);
or U9530 (N_9530,N_9044,N_9327);
nand U9531 (N_9531,N_9018,N_9347);
nand U9532 (N_9532,N_9420,N_9318);
and U9533 (N_9533,N_9452,N_9217);
or U9534 (N_9534,N_9454,N_9057);
and U9535 (N_9535,N_9368,N_9285);
or U9536 (N_9536,N_9251,N_9287);
xnor U9537 (N_9537,N_9111,N_9160);
xnor U9538 (N_9538,N_9045,N_9003);
and U9539 (N_9539,N_9123,N_9241);
xnor U9540 (N_9540,N_9398,N_9422);
xnor U9541 (N_9541,N_9351,N_9275);
nor U9542 (N_9542,N_9306,N_9076);
nand U9543 (N_9543,N_9322,N_9291);
xor U9544 (N_9544,N_9479,N_9175);
or U9545 (N_9545,N_9397,N_9187);
and U9546 (N_9546,N_9246,N_9384);
nand U9547 (N_9547,N_9349,N_9069);
nand U9548 (N_9548,N_9206,N_9029);
nand U9549 (N_9549,N_9365,N_9047);
and U9550 (N_9550,N_9164,N_9004);
or U9551 (N_9551,N_9098,N_9153);
nand U9552 (N_9552,N_9355,N_9483);
nand U9553 (N_9553,N_9090,N_9114);
nand U9554 (N_9554,N_9340,N_9086);
and U9555 (N_9555,N_9294,N_9453);
nor U9556 (N_9556,N_9249,N_9406);
and U9557 (N_9557,N_9165,N_9174);
or U9558 (N_9558,N_9162,N_9299);
xor U9559 (N_9559,N_9068,N_9133);
and U9560 (N_9560,N_9429,N_9207);
or U9561 (N_9561,N_9242,N_9457);
nand U9562 (N_9562,N_9224,N_9159);
nand U9563 (N_9563,N_9271,N_9459);
nand U9564 (N_9564,N_9041,N_9277);
nor U9565 (N_9565,N_9150,N_9151);
xor U9566 (N_9566,N_9116,N_9223);
nor U9567 (N_9567,N_9017,N_9383);
nand U9568 (N_9568,N_9324,N_9490);
nand U9569 (N_9569,N_9094,N_9315);
or U9570 (N_9570,N_9370,N_9303);
nor U9571 (N_9571,N_9178,N_9497);
xor U9572 (N_9572,N_9445,N_9115);
xor U9573 (N_9573,N_9230,N_9260);
xnor U9574 (N_9574,N_9301,N_9407);
nand U9575 (N_9575,N_9052,N_9390);
and U9576 (N_9576,N_9252,N_9037);
xnor U9577 (N_9577,N_9030,N_9088);
and U9578 (N_9578,N_9369,N_9395);
nor U9579 (N_9579,N_9101,N_9286);
nor U9580 (N_9580,N_9434,N_9307);
nand U9581 (N_9581,N_9200,N_9028);
or U9582 (N_9582,N_9411,N_9491);
or U9583 (N_9583,N_9012,N_9319);
or U9584 (N_9584,N_9334,N_9344);
xor U9585 (N_9585,N_9225,N_9102);
xnor U9586 (N_9586,N_9209,N_9167);
and U9587 (N_9587,N_9494,N_9130);
or U9588 (N_9588,N_9325,N_9110);
xor U9589 (N_9589,N_9269,N_9134);
xnor U9590 (N_9590,N_9067,N_9320);
and U9591 (N_9591,N_9182,N_9080);
and U9592 (N_9592,N_9191,N_9027);
or U9593 (N_9593,N_9058,N_9033);
nor U9594 (N_9594,N_9485,N_9064);
xnor U9595 (N_9595,N_9021,N_9274);
and U9596 (N_9596,N_9373,N_9423);
xor U9597 (N_9597,N_9268,N_9444);
xor U9598 (N_9598,N_9427,N_9391);
nand U9599 (N_9599,N_9205,N_9019);
nor U9600 (N_9600,N_9006,N_9478);
or U9601 (N_9601,N_9119,N_9400);
and U9602 (N_9602,N_9065,N_9085);
and U9603 (N_9603,N_9488,N_9345);
nor U9604 (N_9604,N_9392,N_9292);
and U9605 (N_9605,N_9034,N_9399);
and U9606 (N_9606,N_9129,N_9117);
or U9607 (N_9607,N_9432,N_9022);
or U9608 (N_9608,N_9449,N_9354);
and U9609 (N_9609,N_9317,N_9192);
nand U9610 (N_9610,N_9202,N_9240);
or U9611 (N_9611,N_9031,N_9196);
and U9612 (N_9612,N_9297,N_9131);
nor U9613 (N_9613,N_9127,N_9042);
nand U9614 (N_9614,N_9216,N_9061);
or U9615 (N_9615,N_9036,N_9198);
xnor U9616 (N_9616,N_9487,N_9415);
xnor U9617 (N_9617,N_9163,N_9176);
nor U9618 (N_9618,N_9109,N_9336);
or U9619 (N_9619,N_9435,N_9469);
and U9620 (N_9620,N_9335,N_9084);
and U9621 (N_9621,N_9189,N_9376);
xor U9622 (N_9622,N_9169,N_9092);
and U9623 (N_9623,N_9257,N_9363);
nand U9624 (N_9624,N_9179,N_9032);
or U9625 (N_9625,N_9149,N_9227);
and U9626 (N_9626,N_9462,N_9155);
nand U9627 (N_9627,N_9380,N_9346);
nand U9628 (N_9628,N_9136,N_9498);
xnor U9629 (N_9629,N_9342,N_9470);
xor U9630 (N_9630,N_9461,N_9473);
and U9631 (N_9631,N_9472,N_9460);
or U9632 (N_9632,N_9244,N_9245);
and U9633 (N_9633,N_9439,N_9323);
nand U9634 (N_9634,N_9266,N_9330);
nand U9635 (N_9635,N_9144,N_9262);
nand U9636 (N_9636,N_9063,N_9433);
nand U9637 (N_9637,N_9353,N_9492);
or U9638 (N_9638,N_9118,N_9425);
or U9639 (N_9639,N_9157,N_9414);
nand U9640 (N_9640,N_9446,N_9161);
nand U9641 (N_9641,N_9300,N_9333);
nand U9642 (N_9642,N_9168,N_9280);
or U9643 (N_9643,N_9309,N_9005);
xnor U9644 (N_9644,N_9405,N_9180);
nor U9645 (N_9645,N_9082,N_9476);
nor U9646 (N_9646,N_9059,N_9493);
nor U9647 (N_9647,N_9147,N_9402);
nand U9648 (N_9648,N_9475,N_9357);
nand U9649 (N_9649,N_9233,N_9421);
xor U9650 (N_9650,N_9093,N_9386);
xnor U9651 (N_9651,N_9308,N_9338);
or U9652 (N_9652,N_9097,N_9204);
or U9653 (N_9653,N_9190,N_9350);
nand U9654 (N_9654,N_9374,N_9073);
or U9655 (N_9655,N_9104,N_9053);
and U9656 (N_9656,N_9331,N_9055);
xnor U9657 (N_9657,N_9213,N_9426);
nor U9658 (N_9658,N_9141,N_9143);
or U9659 (N_9659,N_9077,N_9410);
and U9660 (N_9660,N_9070,N_9362);
and U9661 (N_9661,N_9142,N_9329);
nor U9662 (N_9662,N_9437,N_9232);
xnor U9663 (N_9663,N_9183,N_9100);
nor U9664 (N_9664,N_9443,N_9238);
xnor U9665 (N_9665,N_9348,N_9393);
and U9666 (N_9666,N_9276,N_9218);
nand U9667 (N_9667,N_9107,N_9364);
or U9668 (N_9668,N_9015,N_9312);
nand U9669 (N_9669,N_9288,N_9332);
and U9670 (N_9670,N_9171,N_9259);
and U9671 (N_9671,N_9025,N_9417);
xor U9672 (N_9672,N_9001,N_9148);
and U9673 (N_9673,N_9263,N_9239);
nand U9674 (N_9674,N_9377,N_9408);
xor U9675 (N_9675,N_9236,N_9014);
or U9676 (N_9676,N_9382,N_9404);
or U9677 (N_9677,N_9105,N_9416);
nand U9678 (N_9678,N_9440,N_9228);
nand U9679 (N_9679,N_9140,N_9375);
nand U9680 (N_9680,N_9010,N_9035);
xor U9681 (N_9681,N_9480,N_9273);
nand U9682 (N_9682,N_9298,N_9210);
and U9683 (N_9683,N_9283,N_9413);
and U9684 (N_9684,N_9139,N_9051);
xnor U9685 (N_9685,N_9087,N_9096);
and U9686 (N_9686,N_9282,N_9467);
and U9687 (N_9687,N_9026,N_9050);
nand U9688 (N_9688,N_9040,N_9296);
and U9689 (N_9689,N_9270,N_9489);
or U9690 (N_9690,N_9091,N_9284);
and U9691 (N_9691,N_9341,N_9495);
nand U9692 (N_9692,N_9356,N_9234);
nand U9693 (N_9693,N_9103,N_9194);
xnor U9694 (N_9694,N_9361,N_9023);
nand U9695 (N_9695,N_9372,N_9316);
nor U9696 (N_9696,N_9166,N_9197);
nor U9697 (N_9697,N_9013,N_9177);
xnor U9698 (N_9698,N_9267,N_9173);
nor U9699 (N_9699,N_9056,N_9049);
and U9700 (N_9700,N_9172,N_9313);
nor U9701 (N_9701,N_9403,N_9448);
nand U9702 (N_9702,N_9302,N_9314);
or U9703 (N_9703,N_9442,N_9009);
nor U9704 (N_9704,N_9256,N_9447);
and U9705 (N_9705,N_9326,N_9254);
nor U9706 (N_9706,N_9438,N_9258);
or U9707 (N_9707,N_9121,N_9226);
xnor U9708 (N_9708,N_9247,N_9428);
nand U9709 (N_9709,N_9074,N_9113);
or U9710 (N_9710,N_9203,N_9465);
or U9711 (N_9711,N_9039,N_9137);
nand U9712 (N_9712,N_9158,N_9060);
nor U9713 (N_9713,N_9126,N_9471);
nor U9714 (N_9714,N_9000,N_9481);
or U9715 (N_9715,N_9455,N_9211);
nand U9716 (N_9716,N_9484,N_9156);
xor U9717 (N_9717,N_9451,N_9409);
nand U9718 (N_9718,N_9343,N_9219);
nor U9719 (N_9719,N_9311,N_9089);
xor U9720 (N_9720,N_9108,N_9199);
and U9721 (N_9721,N_9358,N_9201);
nand U9722 (N_9722,N_9072,N_9255);
xor U9723 (N_9723,N_9321,N_9054);
xor U9724 (N_9724,N_9366,N_9008);
nor U9725 (N_9725,N_9099,N_9450);
nor U9726 (N_9726,N_9401,N_9222);
nand U9727 (N_9727,N_9431,N_9310);
or U9728 (N_9728,N_9367,N_9388);
xor U9729 (N_9729,N_9046,N_9132);
xnor U9730 (N_9730,N_9062,N_9193);
and U9731 (N_9731,N_9477,N_9016);
xnor U9732 (N_9732,N_9499,N_9265);
nor U9733 (N_9733,N_9083,N_9243);
nand U9734 (N_9734,N_9379,N_9474);
or U9735 (N_9735,N_9181,N_9466);
xnor U9736 (N_9736,N_9389,N_9496);
xnor U9737 (N_9737,N_9007,N_9381);
or U9738 (N_9738,N_9278,N_9463);
or U9739 (N_9739,N_9221,N_9250);
xor U9740 (N_9740,N_9043,N_9135);
nor U9741 (N_9741,N_9112,N_9195);
nand U9742 (N_9742,N_9125,N_9436);
nor U9743 (N_9743,N_9418,N_9106);
xnor U9744 (N_9744,N_9235,N_9081);
or U9745 (N_9745,N_9011,N_9419);
and U9746 (N_9746,N_9482,N_9185);
and U9747 (N_9747,N_9456,N_9214);
or U9748 (N_9748,N_9304,N_9430);
nor U9749 (N_9749,N_9261,N_9095);
and U9750 (N_9750,N_9396,N_9066);
and U9751 (N_9751,N_9069,N_9466);
and U9752 (N_9752,N_9298,N_9382);
or U9753 (N_9753,N_9157,N_9223);
nand U9754 (N_9754,N_9119,N_9289);
and U9755 (N_9755,N_9028,N_9023);
nor U9756 (N_9756,N_9350,N_9229);
or U9757 (N_9757,N_9251,N_9254);
and U9758 (N_9758,N_9384,N_9271);
and U9759 (N_9759,N_9411,N_9077);
or U9760 (N_9760,N_9273,N_9108);
and U9761 (N_9761,N_9169,N_9463);
xor U9762 (N_9762,N_9026,N_9294);
nand U9763 (N_9763,N_9355,N_9135);
or U9764 (N_9764,N_9197,N_9222);
or U9765 (N_9765,N_9416,N_9380);
nand U9766 (N_9766,N_9437,N_9184);
nor U9767 (N_9767,N_9096,N_9315);
nand U9768 (N_9768,N_9411,N_9166);
or U9769 (N_9769,N_9057,N_9177);
nor U9770 (N_9770,N_9441,N_9043);
or U9771 (N_9771,N_9168,N_9016);
and U9772 (N_9772,N_9415,N_9385);
nor U9773 (N_9773,N_9340,N_9294);
and U9774 (N_9774,N_9217,N_9376);
xor U9775 (N_9775,N_9148,N_9306);
and U9776 (N_9776,N_9061,N_9257);
xnor U9777 (N_9777,N_9436,N_9191);
nand U9778 (N_9778,N_9357,N_9486);
and U9779 (N_9779,N_9457,N_9368);
or U9780 (N_9780,N_9349,N_9198);
xnor U9781 (N_9781,N_9122,N_9439);
nor U9782 (N_9782,N_9220,N_9290);
and U9783 (N_9783,N_9229,N_9230);
nand U9784 (N_9784,N_9284,N_9212);
or U9785 (N_9785,N_9383,N_9029);
nor U9786 (N_9786,N_9318,N_9306);
nor U9787 (N_9787,N_9314,N_9020);
and U9788 (N_9788,N_9338,N_9331);
or U9789 (N_9789,N_9125,N_9400);
nand U9790 (N_9790,N_9033,N_9422);
or U9791 (N_9791,N_9042,N_9045);
nand U9792 (N_9792,N_9287,N_9183);
and U9793 (N_9793,N_9093,N_9257);
nor U9794 (N_9794,N_9073,N_9030);
or U9795 (N_9795,N_9202,N_9314);
xor U9796 (N_9796,N_9304,N_9099);
or U9797 (N_9797,N_9108,N_9319);
or U9798 (N_9798,N_9108,N_9162);
or U9799 (N_9799,N_9366,N_9297);
and U9800 (N_9800,N_9247,N_9006);
xnor U9801 (N_9801,N_9087,N_9013);
nor U9802 (N_9802,N_9454,N_9013);
or U9803 (N_9803,N_9423,N_9269);
nand U9804 (N_9804,N_9011,N_9328);
nor U9805 (N_9805,N_9126,N_9138);
and U9806 (N_9806,N_9489,N_9036);
xnor U9807 (N_9807,N_9156,N_9006);
nor U9808 (N_9808,N_9206,N_9441);
nor U9809 (N_9809,N_9026,N_9325);
xnor U9810 (N_9810,N_9287,N_9283);
xnor U9811 (N_9811,N_9275,N_9121);
nand U9812 (N_9812,N_9040,N_9432);
and U9813 (N_9813,N_9136,N_9414);
xnor U9814 (N_9814,N_9413,N_9470);
or U9815 (N_9815,N_9190,N_9149);
nand U9816 (N_9816,N_9172,N_9216);
and U9817 (N_9817,N_9146,N_9254);
xor U9818 (N_9818,N_9263,N_9074);
nor U9819 (N_9819,N_9004,N_9406);
and U9820 (N_9820,N_9134,N_9198);
xnor U9821 (N_9821,N_9388,N_9356);
and U9822 (N_9822,N_9396,N_9068);
xor U9823 (N_9823,N_9265,N_9303);
nor U9824 (N_9824,N_9298,N_9172);
nand U9825 (N_9825,N_9477,N_9257);
nand U9826 (N_9826,N_9366,N_9244);
nand U9827 (N_9827,N_9109,N_9415);
xnor U9828 (N_9828,N_9309,N_9181);
or U9829 (N_9829,N_9104,N_9390);
and U9830 (N_9830,N_9270,N_9116);
or U9831 (N_9831,N_9176,N_9369);
nand U9832 (N_9832,N_9111,N_9315);
or U9833 (N_9833,N_9316,N_9208);
xnor U9834 (N_9834,N_9216,N_9067);
nand U9835 (N_9835,N_9128,N_9115);
xnor U9836 (N_9836,N_9118,N_9423);
and U9837 (N_9837,N_9441,N_9151);
nor U9838 (N_9838,N_9299,N_9086);
and U9839 (N_9839,N_9106,N_9142);
xnor U9840 (N_9840,N_9391,N_9312);
or U9841 (N_9841,N_9165,N_9479);
nand U9842 (N_9842,N_9084,N_9257);
or U9843 (N_9843,N_9382,N_9280);
and U9844 (N_9844,N_9087,N_9111);
nor U9845 (N_9845,N_9498,N_9427);
xor U9846 (N_9846,N_9411,N_9389);
or U9847 (N_9847,N_9018,N_9045);
and U9848 (N_9848,N_9138,N_9482);
nor U9849 (N_9849,N_9235,N_9027);
nor U9850 (N_9850,N_9321,N_9000);
nand U9851 (N_9851,N_9088,N_9194);
or U9852 (N_9852,N_9299,N_9276);
nor U9853 (N_9853,N_9343,N_9464);
nand U9854 (N_9854,N_9332,N_9453);
or U9855 (N_9855,N_9176,N_9368);
xor U9856 (N_9856,N_9381,N_9318);
nor U9857 (N_9857,N_9296,N_9260);
nor U9858 (N_9858,N_9256,N_9414);
and U9859 (N_9859,N_9298,N_9233);
and U9860 (N_9860,N_9009,N_9414);
and U9861 (N_9861,N_9164,N_9425);
or U9862 (N_9862,N_9460,N_9348);
nand U9863 (N_9863,N_9007,N_9373);
nand U9864 (N_9864,N_9119,N_9387);
xor U9865 (N_9865,N_9011,N_9264);
xnor U9866 (N_9866,N_9207,N_9388);
or U9867 (N_9867,N_9089,N_9400);
nor U9868 (N_9868,N_9343,N_9489);
or U9869 (N_9869,N_9494,N_9354);
or U9870 (N_9870,N_9371,N_9238);
nor U9871 (N_9871,N_9130,N_9033);
and U9872 (N_9872,N_9067,N_9460);
or U9873 (N_9873,N_9059,N_9300);
or U9874 (N_9874,N_9013,N_9193);
and U9875 (N_9875,N_9452,N_9230);
and U9876 (N_9876,N_9083,N_9392);
or U9877 (N_9877,N_9393,N_9479);
nand U9878 (N_9878,N_9445,N_9116);
xor U9879 (N_9879,N_9050,N_9055);
and U9880 (N_9880,N_9349,N_9476);
nand U9881 (N_9881,N_9306,N_9372);
nor U9882 (N_9882,N_9288,N_9103);
or U9883 (N_9883,N_9202,N_9367);
or U9884 (N_9884,N_9416,N_9098);
and U9885 (N_9885,N_9206,N_9484);
and U9886 (N_9886,N_9470,N_9062);
nor U9887 (N_9887,N_9030,N_9347);
or U9888 (N_9888,N_9023,N_9490);
nor U9889 (N_9889,N_9468,N_9264);
and U9890 (N_9890,N_9354,N_9467);
nor U9891 (N_9891,N_9008,N_9291);
or U9892 (N_9892,N_9462,N_9387);
xor U9893 (N_9893,N_9227,N_9170);
nor U9894 (N_9894,N_9429,N_9002);
nand U9895 (N_9895,N_9113,N_9378);
xor U9896 (N_9896,N_9195,N_9040);
nor U9897 (N_9897,N_9419,N_9018);
or U9898 (N_9898,N_9178,N_9053);
nor U9899 (N_9899,N_9077,N_9214);
and U9900 (N_9900,N_9200,N_9319);
xnor U9901 (N_9901,N_9291,N_9162);
nand U9902 (N_9902,N_9110,N_9061);
or U9903 (N_9903,N_9155,N_9253);
nand U9904 (N_9904,N_9333,N_9224);
or U9905 (N_9905,N_9097,N_9413);
nor U9906 (N_9906,N_9026,N_9006);
nand U9907 (N_9907,N_9446,N_9151);
xnor U9908 (N_9908,N_9281,N_9470);
xor U9909 (N_9909,N_9435,N_9492);
and U9910 (N_9910,N_9205,N_9199);
xnor U9911 (N_9911,N_9489,N_9156);
or U9912 (N_9912,N_9187,N_9216);
and U9913 (N_9913,N_9025,N_9413);
xor U9914 (N_9914,N_9183,N_9488);
and U9915 (N_9915,N_9402,N_9400);
and U9916 (N_9916,N_9277,N_9383);
or U9917 (N_9917,N_9484,N_9395);
xor U9918 (N_9918,N_9365,N_9261);
xor U9919 (N_9919,N_9407,N_9156);
nor U9920 (N_9920,N_9086,N_9175);
nor U9921 (N_9921,N_9350,N_9162);
and U9922 (N_9922,N_9362,N_9158);
and U9923 (N_9923,N_9208,N_9198);
or U9924 (N_9924,N_9288,N_9160);
nor U9925 (N_9925,N_9208,N_9175);
nand U9926 (N_9926,N_9322,N_9124);
or U9927 (N_9927,N_9385,N_9222);
xnor U9928 (N_9928,N_9457,N_9138);
or U9929 (N_9929,N_9000,N_9210);
or U9930 (N_9930,N_9233,N_9104);
nor U9931 (N_9931,N_9246,N_9263);
nor U9932 (N_9932,N_9011,N_9458);
nand U9933 (N_9933,N_9172,N_9343);
and U9934 (N_9934,N_9209,N_9393);
or U9935 (N_9935,N_9326,N_9192);
xnor U9936 (N_9936,N_9225,N_9471);
or U9937 (N_9937,N_9337,N_9021);
nand U9938 (N_9938,N_9103,N_9240);
nor U9939 (N_9939,N_9127,N_9084);
and U9940 (N_9940,N_9188,N_9161);
or U9941 (N_9941,N_9010,N_9033);
or U9942 (N_9942,N_9405,N_9419);
and U9943 (N_9943,N_9276,N_9005);
xnor U9944 (N_9944,N_9089,N_9194);
nand U9945 (N_9945,N_9444,N_9384);
xnor U9946 (N_9946,N_9110,N_9177);
nor U9947 (N_9947,N_9121,N_9187);
or U9948 (N_9948,N_9017,N_9488);
and U9949 (N_9949,N_9053,N_9441);
and U9950 (N_9950,N_9224,N_9153);
or U9951 (N_9951,N_9425,N_9312);
nand U9952 (N_9952,N_9153,N_9263);
or U9953 (N_9953,N_9298,N_9160);
or U9954 (N_9954,N_9477,N_9275);
nand U9955 (N_9955,N_9071,N_9290);
nor U9956 (N_9956,N_9051,N_9270);
xnor U9957 (N_9957,N_9015,N_9001);
and U9958 (N_9958,N_9418,N_9241);
nor U9959 (N_9959,N_9172,N_9448);
nand U9960 (N_9960,N_9131,N_9487);
or U9961 (N_9961,N_9173,N_9133);
and U9962 (N_9962,N_9315,N_9261);
and U9963 (N_9963,N_9398,N_9034);
nor U9964 (N_9964,N_9240,N_9138);
xor U9965 (N_9965,N_9446,N_9473);
xor U9966 (N_9966,N_9159,N_9408);
or U9967 (N_9967,N_9172,N_9450);
xnor U9968 (N_9968,N_9423,N_9382);
nand U9969 (N_9969,N_9061,N_9400);
nor U9970 (N_9970,N_9158,N_9209);
and U9971 (N_9971,N_9354,N_9497);
and U9972 (N_9972,N_9257,N_9300);
or U9973 (N_9973,N_9348,N_9054);
or U9974 (N_9974,N_9340,N_9346);
nor U9975 (N_9975,N_9075,N_9071);
or U9976 (N_9976,N_9252,N_9080);
and U9977 (N_9977,N_9188,N_9051);
or U9978 (N_9978,N_9241,N_9245);
and U9979 (N_9979,N_9407,N_9061);
nand U9980 (N_9980,N_9055,N_9382);
xnor U9981 (N_9981,N_9476,N_9035);
or U9982 (N_9982,N_9273,N_9276);
nor U9983 (N_9983,N_9104,N_9317);
and U9984 (N_9984,N_9399,N_9326);
xor U9985 (N_9985,N_9185,N_9068);
xnor U9986 (N_9986,N_9169,N_9288);
or U9987 (N_9987,N_9068,N_9072);
xor U9988 (N_9988,N_9478,N_9325);
nor U9989 (N_9989,N_9333,N_9153);
xnor U9990 (N_9990,N_9319,N_9119);
and U9991 (N_9991,N_9031,N_9137);
and U9992 (N_9992,N_9368,N_9267);
nand U9993 (N_9993,N_9213,N_9218);
or U9994 (N_9994,N_9081,N_9395);
or U9995 (N_9995,N_9439,N_9258);
or U9996 (N_9996,N_9224,N_9401);
nor U9997 (N_9997,N_9320,N_9240);
xor U9998 (N_9998,N_9352,N_9225);
xnor U9999 (N_9999,N_9427,N_9402);
nand U10000 (N_10000,N_9764,N_9968);
or U10001 (N_10001,N_9563,N_9709);
nand U10002 (N_10002,N_9502,N_9575);
xor U10003 (N_10003,N_9790,N_9545);
xnor U10004 (N_10004,N_9802,N_9566);
nor U10005 (N_10005,N_9684,N_9945);
nand U10006 (N_10006,N_9973,N_9985);
nand U10007 (N_10007,N_9662,N_9801);
nand U10008 (N_10008,N_9653,N_9839);
or U10009 (N_10009,N_9553,N_9676);
or U10010 (N_10010,N_9842,N_9792);
and U10011 (N_10011,N_9648,N_9503);
xnor U10012 (N_10012,N_9959,N_9532);
xor U10013 (N_10013,N_9810,N_9706);
xor U10014 (N_10014,N_9865,N_9844);
nor U10015 (N_10015,N_9965,N_9716);
and U10016 (N_10016,N_9962,N_9907);
or U10017 (N_10017,N_9585,N_9953);
xnor U10018 (N_10018,N_9657,N_9586);
nand U10019 (N_10019,N_9666,N_9917);
and U10020 (N_10020,N_9971,N_9649);
and U10021 (N_10021,N_9938,N_9853);
xnor U10022 (N_10022,N_9602,N_9698);
nand U10023 (N_10023,N_9685,N_9550);
or U10024 (N_10024,N_9882,N_9674);
and U10025 (N_10025,N_9847,N_9978);
xnor U10026 (N_10026,N_9683,N_9607);
or U10027 (N_10027,N_9687,N_9606);
xnor U10028 (N_10028,N_9824,N_9769);
xnor U10029 (N_10029,N_9901,N_9956);
and U10030 (N_10030,N_9808,N_9871);
nand U10031 (N_10031,N_9535,N_9568);
xor U10032 (N_10032,N_9711,N_9936);
and U10033 (N_10033,N_9788,N_9919);
or U10034 (N_10034,N_9988,N_9745);
and U10035 (N_10035,N_9722,N_9806);
and U10036 (N_10036,N_9610,N_9644);
nor U10037 (N_10037,N_9759,N_9900);
or U10038 (N_10038,N_9558,N_9887);
xor U10039 (N_10039,N_9534,N_9598);
xnor U10040 (N_10040,N_9693,N_9567);
or U10041 (N_10041,N_9647,N_9856);
xor U10042 (N_10042,N_9692,N_9737);
or U10043 (N_10043,N_9739,N_9754);
xor U10044 (N_10044,N_9541,N_9705);
and U10045 (N_10045,N_9512,N_9990);
nor U10046 (N_10046,N_9951,N_9794);
xor U10047 (N_10047,N_9542,N_9531);
or U10048 (N_10048,N_9569,N_9899);
and U10049 (N_10049,N_9741,N_9616);
and U10050 (N_10050,N_9556,N_9646);
xnor U10051 (N_10051,N_9609,N_9690);
and U10052 (N_10052,N_9633,N_9715);
nand U10053 (N_10053,N_9580,N_9755);
nand U10054 (N_10054,N_9735,N_9537);
or U10055 (N_10055,N_9520,N_9934);
and U10056 (N_10056,N_9869,N_9504);
xnor U10057 (N_10057,N_9601,N_9798);
nor U10058 (N_10058,N_9584,N_9819);
nand U10059 (N_10059,N_9855,N_9564);
xnor U10060 (N_10060,N_9944,N_9719);
nor U10061 (N_10061,N_9667,N_9822);
and U10062 (N_10062,N_9757,N_9786);
nor U10063 (N_10063,N_9866,N_9695);
xor U10064 (N_10064,N_9659,N_9526);
nand U10065 (N_10065,N_9500,N_9993);
nand U10066 (N_10066,N_9797,N_9777);
nand U10067 (N_10067,N_9625,N_9572);
or U10068 (N_10068,N_9758,N_9913);
xor U10069 (N_10069,N_9997,N_9549);
and U10070 (N_10070,N_9591,N_9821);
nand U10071 (N_10071,N_9989,N_9961);
and U10072 (N_10072,N_9544,N_9574);
nand U10073 (N_10073,N_9561,N_9589);
and U10074 (N_10074,N_9884,N_9579);
and U10075 (N_10075,N_9783,N_9700);
and U10076 (N_10076,N_9603,N_9614);
nor U10077 (N_10077,N_9704,N_9582);
nor U10078 (N_10078,N_9778,N_9630);
or U10079 (N_10079,N_9905,N_9519);
nor U10080 (N_10080,N_9546,N_9779);
and U10081 (N_10081,N_9833,N_9599);
nor U10082 (N_10082,N_9627,N_9636);
or U10083 (N_10083,N_9966,N_9686);
xnor U10084 (N_10084,N_9986,N_9923);
or U10085 (N_10085,N_9734,N_9748);
nand U10086 (N_10086,N_9509,N_9817);
and U10087 (N_10087,N_9896,N_9639);
and U10088 (N_10088,N_9780,N_9694);
nor U10089 (N_10089,N_9789,N_9624);
xor U10090 (N_10090,N_9729,N_9845);
nand U10091 (N_10091,N_9916,N_9728);
or U10092 (N_10092,N_9540,N_9726);
or U10093 (N_10093,N_9577,N_9708);
nand U10094 (N_10094,N_9909,N_9820);
xor U10095 (N_10095,N_9524,N_9725);
and U10096 (N_10096,N_9751,N_9656);
nor U10097 (N_10097,N_9892,N_9514);
nor U10098 (N_10098,N_9890,N_9620);
or U10099 (N_10099,N_9756,N_9581);
nor U10100 (N_10100,N_9940,N_9795);
xor U10101 (N_10101,N_9781,N_9912);
nand U10102 (N_10102,N_9860,N_9511);
and U10103 (N_10103,N_9927,N_9628);
or U10104 (N_10104,N_9947,N_9730);
or U10105 (N_10105,N_9749,N_9731);
and U10106 (N_10106,N_9861,N_9999);
nand U10107 (N_10107,N_9623,N_9902);
or U10108 (N_10108,N_9634,N_9618);
nor U10109 (N_10109,N_9987,N_9642);
or U10110 (N_10110,N_9652,N_9727);
and U10111 (N_10111,N_9931,N_9689);
or U10112 (N_10112,N_9736,N_9782);
or U10113 (N_10113,N_9600,N_9576);
or U10114 (N_10114,N_9939,N_9660);
or U10115 (N_10115,N_9641,N_9984);
xnor U10116 (N_10116,N_9981,N_9932);
xor U10117 (N_10117,N_9772,N_9594);
nor U10118 (N_10118,N_9992,N_9738);
and U10119 (N_10119,N_9710,N_9681);
nor U10120 (N_10120,N_9527,N_9721);
and U10121 (N_10121,N_9617,N_9565);
and U10122 (N_10122,N_9638,N_9508);
or U10123 (N_10123,N_9889,N_9925);
nor U10124 (N_10124,N_9793,N_9843);
nor U10125 (N_10125,N_9977,N_9744);
and U10126 (N_10126,N_9562,N_9891);
xnor U10127 (N_10127,N_9870,N_9631);
nand U10128 (N_10128,N_9807,N_9650);
or U10129 (N_10129,N_9543,N_9615);
nand U10130 (N_10130,N_9611,N_9643);
nand U10131 (N_10131,N_9516,N_9935);
xnor U10132 (N_10132,N_9864,N_9950);
nor U10133 (N_10133,N_9863,N_9828);
and U10134 (N_10134,N_9626,N_9943);
or U10135 (N_10135,N_9813,N_9661);
and U10136 (N_10136,N_9895,N_9505);
nand U10137 (N_10137,N_9829,N_9547);
and U10138 (N_10138,N_9560,N_9678);
xnor U10139 (N_10139,N_9873,N_9818);
nor U10140 (N_10140,N_9964,N_9852);
nand U10141 (N_10141,N_9960,N_9885);
nor U10142 (N_10142,N_9823,N_9770);
and U10143 (N_10143,N_9904,N_9752);
and U10144 (N_10144,N_9530,N_9906);
or U10145 (N_10145,N_9812,N_9976);
or U10146 (N_10146,N_9980,N_9982);
xor U10147 (N_10147,N_9991,N_9557);
nand U10148 (N_10148,N_9548,N_9903);
nand U10149 (N_10149,N_9697,N_9867);
and U10150 (N_10150,N_9688,N_9761);
xnor U10151 (N_10151,N_9814,N_9604);
and U10152 (N_10152,N_9879,N_9791);
and U10153 (N_10153,N_9803,N_9868);
xor U10154 (N_10154,N_9523,N_9773);
and U10155 (N_10155,N_9994,N_9529);
nor U10156 (N_10156,N_9654,N_9522);
or U10157 (N_10157,N_9664,N_9894);
nor U10158 (N_10158,N_9714,N_9655);
xnor U10159 (N_10159,N_9637,N_9827);
xor U10160 (N_10160,N_9877,N_9703);
and U10161 (N_10161,N_9910,N_9525);
and U10162 (N_10162,N_9858,N_9753);
or U10163 (N_10163,N_9929,N_9501);
or U10164 (N_10164,N_9914,N_9670);
and U10165 (N_10165,N_9679,N_9713);
xnor U10166 (N_10166,N_9672,N_9521);
nor U10167 (N_10167,N_9775,N_9857);
or U10168 (N_10168,N_9608,N_9588);
nand U10169 (N_10169,N_9846,N_9538);
nor U10170 (N_10170,N_9876,N_9799);
nand U10171 (N_10171,N_9732,N_9671);
nand U10172 (N_10172,N_9510,N_9831);
nor U10173 (N_10173,N_9613,N_9570);
nand U10174 (N_10174,N_9733,N_9513);
nor U10175 (N_10175,N_9677,N_9645);
and U10176 (N_10176,N_9804,N_9922);
nand U10177 (N_10177,N_9629,N_9724);
nand U10178 (N_10178,N_9924,N_9893);
and U10179 (N_10179,N_9663,N_9963);
or U10180 (N_10180,N_9969,N_9528);
and U10181 (N_10181,N_9699,N_9878);
xor U10182 (N_10182,N_9949,N_9768);
nand U10183 (N_10183,N_9880,N_9702);
nand U10184 (N_10184,N_9918,N_9958);
xor U10185 (N_10185,N_9838,N_9762);
and U10186 (N_10186,N_9701,N_9974);
nand U10187 (N_10187,N_9948,N_9849);
nand U10188 (N_10188,N_9536,N_9928);
nand U10189 (N_10189,N_9712,N_9825);
xnor U10190 (N_10190,N_9665,N_9595);
or U10191 (N_10191,N_9800,N_9826);
and U10192 (N_10192,N_9952,N_9590);
and U10193 (N_10193,N_9747,N_9740);
nor U10194 (N_10194,N_9957,N_9785);
nor U10195 (N_10195,N_9811,N_9658);
and U10196 (N_10196,N_9539,N_9983);
or U10197 (N_10197,N_9837,N_9888);
nand U10198 (N_10198,N_9743,N_9597);
nor U10199 (N_10199,N_9612,N_9533);
xor U10200 (N_10200,N_9854,N_9809);
and U10201 (N_10201,N_9651,N_9517);
or U10202 (N_10202,N_9834,N_9796);
or U10203 (N_10203,N_9787,N_9859);
nor U10204 (N_10204,N_9998,N_9967);
nand U10205 (N_10205,N_9621,N_9552);
xnor U10206 (N_10206,N_9571,N_9954);
nor U10207 (N_10207,N_9805,N_9862);
or U10208 (N_10208,N_9765,N_9933);
nor U10209 (N_10209,N_9691,N_9955);
and U10210 (N_10210,N_9816,N_9559);
xnor U10211 (N_10211,N_9763,N_9682);
nand U10212 (N_10212,N_9515,N_9605);
nor U10213 (N_10213,N_9851,N_9832);
xor U10214 (N_10214,N_9596,N_9723);
or U10215 (N_10215,N_9883,N_9675);
and U10216 (N_10216,N_9937,N_9680);
or U10217 (N_10217,N_9995,N_9746);
or U10218 (N_10218,N_9920,N_9996);
nand U10219 (N_10219,N_9921,N_9946);
xnor U10220 (N_10220,N_9942,N_9897);
or U10221 (N_10221,N_9908,N_9970);
and U10222 (N_10222,N_9668,N_9926);
nor U10223 (N_10223,N_9593,N_9881);
nand U10224 (N_10224,N_9841,N_9506);
and U10225 (N_10225,N_9972,N_9930);
nor U10226 (N_10226,N_9840,N_9815);
nand U10227 (N_10227,N_9592,N_9941);
or U10228 (N_10228,N_9836,N_9573);
xor U10229 (N_10229,N_9886,N_9507);
nor U10230 (N_10230,N_9717,N_9622);
and U10231 (N_10231,N_9742,N_9979);
and U10232 (N_10232,N_9555,N_9850);
nand U10233 (N_10233,N_9872,N_9975);
xnor U10234 (N_10234,N_9554,N_9583);
and U10235 (N_10235,N_9774,N_9771);
nand U10236 (N_10236,N_9578,N_9640);
nor U10237 (N_10237,N_9696,N_9915);
and U10238 (N_10238,N_9875,N_9720);
or U10239 (N_10239,N_9551,N_9767);
nand U10240 (N_10240,N_9784,N_9619);
nor U10241 (N_10241,N_9830,N_9673);
and U10242 (N_10242,N_9707,N_9518);
xor U10243 (N_10243,N_9635,N_9632);
nor U10244 (N_10244,N_9911,N_9760);
or U10245 (N_10245,N_9776,N_9718);
and U10246 (N_10246,N_9587,N_9848);
or U10247 (N_10247,N_9874,N_9766);
or U10248 (N_10248,N_9898,N_9835);
nor U10249 (N_10249,N_9669,N_9750);
and U10250 (N_10250,N_9685,N_9651);
xnor U10251 (N_10251,N_9572,N_9850);
and U10252 (N_10252,N_9566,N_9699);
or U10253 (N_10253,N_9873,N_9642);
and U10254 (N_10254,N_9635,N_9534);
nand U10255 (N_10255,N_9890,N_9714);
and U10256 (N_10256,N_9731,N_9501);
and U10257 (N_10257,N_9870,N_9845);
and U10258 (N_10258,N_9738,N_9804);
nand U10259 (N_10259,N_9657,N_9998);
nand U10260 (N_10260,N_9756,N_9799);
nor U10261 (N_10261,N_9910,N_9852);
xor U10262 (N_10262,N_9761,N_9795);
or U10263 (N_10263,N_9527,N_9919);
and U10264 (N_10264,N_9649,N_9949);
nor U10265 (N_10265,N_9866,N_9616);
and U10266 (N_10266,N_9941,N_9583);
xnor U10267 (N_10267,N_9608,N_9770);
and U10268 (N_10268,N_9746,N_9649);
nand U10269 (N_10269,N_9944,N_9856);
and U10270 (N_10270,N_9630,N_9793);
nand U10271 (N_10271,N_9912,N_9558);
or U10272 (N_10272,N_9942,N_9908);
or U10273 (N_10273,N_9752,N_9598);
or U10274 (N_10274,N_9794,N_9978);
and U10275 (N_10275,N_9561,N_9897);
nor U10276 (N_10276,N_9960,N_9874);
nor U10277 (N_10277,N_9674,N_9509);
nand U10278 (N_10278,N_9925,N_9733);
nor U10279 (N_10279,N_9603,N_9786);
nand U10280 (N_10280,N_9780,N_9608);
and U10281 (N_10281,N_9969,N_9798);
or U10282 (N_10282,N_9921,N_9523);
xnor U10283 (N_10283,N_9738,N_9813);
nand U10284 (N_10284,N_9737,N_9677);
xnor U10285 (N_10285,N_9841,N_9542);
or U10286 (N_10286,N_9585,N_9529);
or U10287 (N_10287,N_9513,N_9673);
nor U10288 (N_10288,N_9765,N_9595);
or U10289 (N_10289,N_9725,N_9621);
and U10290 (N_10290,N_9974,N_9541);
nand U10291 (N_10291,N_9627,N_9582);
nor U10292 (N_10292,N_9729,N_9897);
and U10293 (N_10293,N_9690,N_9530);
and U10294 (N_10294,N_9780,N_9965);
nand U10295 (N_10295,N_9969,N_9728);
nand U10296 (N_10296,N_9905,N_9907);
or U10297 (N_10297,N_9839,N_9865);
and U10298 (N_10298,N_9882,N_9748);
nand U10299 (N_10299,N_9736,N_9713);
or U10300 (N_10300,N_9701,N_9784);
xnor U10301 (N_10301,N_9928,N_9678);
nor U10302 (N_10302,N_9782,N_9587);
or U10303 (N_10303,N_9734,N_9784);
xor U10304 (N_10304,N_9542,N_9519);
nand U10305 (N_10305,N_9834,N_9506);
or U10306 (N_10306,N_9607,N_9630);
nand U10307 (N_10307,N_9991,N_9631);
and U10308 (N_10308,N_9671,N_9765);
nor U10309 (N_10309,N_9571,N_9653);
xnor U10310 (N_10310,N_9515,N_9708);
and U10311 (N_10311,N_9613,N_9834);
or U10312 (N_10312,N_9640,N_9854);
nand U10313 (N_10313,N_9983,N_9792);
nor U10314 (N_10314,N_9721,N_9570);
nor U10315 (N_10315,N_9579,N_9922);
nor U10316 (N_10316,N_9874,N_9942);
xor U10317 (N_10317,N_9859,N_9931);
nand U10318 (N_10318,N_9607,N_9840);
and U10319 (N_10319,N_9509,N_9601);
or U10320 (N_10320,N_9878,N_9860);
nor U10321 (N_10321,N_9939,N_9757);
or U10322 (N_10322,N_9667,N_9599);
nand U10323 (N_10323,N_9603,N_9583);
xor U10324 (N_10324,N_9962,N_9564);
and U10325 (N_10325,N_9982,N_9596);
nand U10326 (N_10326,N_9922,N_9996);
nand U10327 (N_10327,N_9940,N_9966);
nand U10328 (N_10328,N_9687,N_9870);
nor U10329 (N_10329,N_9577,N_9728);
and U10330 (N_10330,N_9607,N_9515);
nand U10331 (N_10331,N_9819,N_9637);
and U10332 (N_10332,N_9784,N_9739);
or U10333 (N_10333,N_9729,N_9771);
nor U10334 (N_10334,N_9640,N_9661);
and U10335 (N_10335,N_9685,N_9737);
nand U10336 (N_10336,N_9591,N_9627);
and U10337 (N_10337,N_9970,N_9649);
nand U10338 (N_10338,N_9563,N_9541);
and U10339 (N_10339,N_9501,N_9679);
xor U10340 (N_10340,N_9742,N_9906);
and U10341 (N_10341,N_9833,N_9829);
nor U10342 (N_10342,N_9937,N_9798);
nor U10343 (N_10343,N_9815,N_9687);
nand U10344 (N_10344,N_9746,N_9611);
and U10345 (N_10345,N_9852,N_9797);
nor U10346 (N_10346,N_9797,N_9745);
or U10347 (N_10347,N_9959,N_9739);
nor U10348 (N_10348,N_9829,N_9776);
or U10349 (N_10349,N_9787,N_9752);
xnor U10350 (N_10350,N_9520,N_9787);
and U10351 (N_10351,N_9546,N_9567);
nand U10352 (N_10352,N_9754,N_9667);
and U10353 (N_10353,N_9864,N_9712);
and U10354 (N_10354,N_9707,N_9968);
nand U10355 (N_10355,N_9683,N_9742);
or U10356 (N_10356,N_9566,N_9826);
or U10357 (N_10357,N_9834,N_9649);
xor U10358 (N_10358,N_9874,N_9830);
or U10359 (N_10359,N_9511,N_9890);
xor U10360 (N_10360,N_9958,N_9767);
nand U10361 (N_10361,N_9531,N_9559);
nor U10362 (N_10362,N_9792,N_9766);
nand U10363 (N_10363,N_9643,N_9821);
nor U10364 (N_10364,N_9881,N_9521);
and U10365 (N_10365,N_9917,N_9866);
nor U10366 (N_10366,N_9914,N_9719);
or U10367 (N_10367,N_9706,N_9656);
and U10368 (N_10368,N_9686,N_9520);
nand U10369 (N_10369,N_9809,N_9682);
or U10370 (N_10370,N_9973,N_9941);
or U10371 (N_10371,N_9902,N_9711);
nand U10372 (N_10372,N_9897,N_9858);
nor U10373 (N_10373,N_9844,N_9764);
nor U10374 (N_10374,N_9881,N_9675);
nor U10375 (N_10375,N_9594,N_9584);
nor U10376 (N_10376,N_9729,N_9955);
nand U10377 (N_10377,N_9936,N_9714);
nor U10378 (N_10378,N_9819,N_9982);
or U10379 (N_10379,N_9787,N_9709);
nand U10380 (N_10380,N_9583,N_9903);
and U10381 (N_10381,N_9879,N_9591);
nand U10382 (N_10382,N_9631,N_9886);
nand U10383 (N_10383,N_9902,N_9878);
or U10384 (N_10384,N_9640,N_9803);
nand U10385 (N_10385,N_9571,N_9792);
nor U10386 (N_10386,N_9695,N_9629);
nor U10387 (N_10387,N_9577,N_9700);
and U10388 (N_10388,N_9790,N_9638);
xnor U10389 (N_10389,N_9803,N_9765);
and U10390 (N_10390,N_9622,N_9785);
xnor U10391 (N_10391,N_9616,N_9733);
xnor U10392 (N_10392,N_9722,N_9866);
nand U10393 (N_10393,N_9520,N_9524);
xnor U10394 (N_10394,N_9922,N_9805);
xnor U10395 (N_10395,N_9937,N_9670);
or U10396 (N_10396,N_9737,N_9628);
xor U10397 (N_10397,N_9720,N_9700);
or U10398 (N_10398,N_9575,N_9703);
nand U10399 (N_10399,N_9850,N_9608);
and U10400 (N_10400,N_9728,N_9822);
and U10401 (N_10401,N_9675,N_9741);
and U10402 (N_10402,N_9872,N_9842);
xor U10403 (N_10403,N_9806,N_9691);
xor U10404 (N_10404,N_9811,N_9890);
and U10405 (N_10405,N_9981,N_9660);
nor U10406 (N_10406,N_9854,N_9876);
and U10407 (N_10407,N_9914,N_9502);
nor U10408 (N_10408,N_9826,N_9513);
nand U10409 (N_10409,N_9995,N_9627);
nor U10410 (N_10410,N_9880,N_9500);
and U10411 (N_10411,N_9643,N_9989);
nand U10412 (N_10412,N_9760,N_9774);
or U10413 (N_10413,N_9790,N_9507);
nand U10414 (N_10414,N_9920,N_9959);
and U10415 (N_10415,N_9755,N_9968);
or U10416 (N_10416,N_9900,N_9587);
nor U10417 (N_10417,N_9992,N_9501);
nand U10418 (N_10418,N_9780,N_9506);
nand U10419 (N_10419,N_9604,N_9667);
xor U10420 (N_10420,N_9658,N_9607);
or U10421 (N_10421,N_9987,N_9591);
xnor U10422 (N_10422,N_9851,N_9828);
xor U10423 (N_10423,N_9948,N_9585);
or U10424 (N_10424,N_9879,N_9878);
xnor U10425 (N_10425,N_9756,N_9917);
or U10426 (N_10426,N_9901,N_9962);
nand U10427 (N_10427,N_9603,N_9868);
xnor U10428 (N_10428,N_9610,N_9510);
and U10429 (N_10429,N_9597,N_9846);
xor U10430 (N_10430,N_9910,N_9533);
or U10431 (N_10431,N_9803,N_9731);
or U10432 (N_10432,N_9758,N_9870);
nand U10433 (N_10433,N_9864,N_9656);
xnor U10434 (N_10434,N_9512,N_9877);
or U10435 (N_10435,N_9754,N_9702);
xor U10436 (N_10436,N_9913,N_9922);
nand U10437 (N_10437,N_9587,N_9556);
nand U10438 (N_10438,N_9943,N_9756);
nand U10439 (N_10439,N_9708,N_9758);
or U10440 (N_10440,N_9771,N_9857);
and U10441 (N_10441,N_9836,N_9876);
nand U10442 (N_10442,N_9686,N_9621);
xnor U10443 (N_10443,N_9978,N_9536);
and U10444 (N_10444,N_9877,N_9807);
nand U10445 (N_10445,N_9841,N_9787);
and U10446 (N_10446,N_9529,N_9872);
xnor U10447 (N_10447,N_9907,N_9692);
or U10448 (N_10448,N_9829,N_9728);
or U10449 (N_10449,N_9895,N_9922);
nor U10450 (N_10450,N_9688,N_9863);
nor U10451 (N_10451,N_9507,N_9773);
xor U10452 (N_10452,N_9763,N_9721);
or U10453 (N_10453,N_9994,N_9749);
nor U10454 (N_10454,N_9917,N_9575);
and U10455 (N_10455,N_9877,N_9907);
nor U10456 (N_10456,N_9645,N_9957);
nand U10457 (N_10457,N_9892,N_9680);
or U10458 (N_10458,N_9946,N_9830);
nand U10459 (N_10459,N_9608,N_9703);
nor U10460 (N_10460,N_9554,N_9859);
nor U10461 (N_10461,N_9739,N_9808);
or U10462 (N_10462,N_9625,N_9704);
xnor U10463 (N_10463,N_9815,N_9614);
or U10464 (N_10464,N_9901,N_9846);
or U10465 (N_10465,N_9974,N_9545);
nand U10466 (N_10466,N_9698,N_9944);
nor U10467 (N_10467,N_9886,N_9775);
nand U10468 (N_10468,N_9612,N_9670);
nand U10469 (N_10469,N_9587,N_9840);
xnor U10470 (N_10470,N_9874,N_9834);
nor U10471 (N_10471,N_9830,N_9976);
nor U10472 (N_10472,N_9688,N_9556);
nand U10473 (N_10473,N_9632,N_9521);
nor U10474 (N_10474,N_9640,N_9648);
nor U10475 (N_10475,N_9739,N_9731);
or U10476 (N_10476,N_9843,N_9748);
nand U10477 (N_10477,N_9901,N_9511);
nor U10478 (N_10478,N_9607,N_9990);
xnor U10479 (N_10479,N_9589,N_9603);
xnor U10480 (N_10480,N_9769,N_9609);
nand U10481 (N_10481,N_9589,N_9597);
nand U10482 (N_10482,N_9727,N_9632);
and U10483 (N_10483,N_9761,N_9971);
or U10484 (N_10484,N_9920,N_9800);
nand U10485 (N_10485,N_9655,N_9948);
nor U10486 (N_10486,N_9556,N_9667);
nand U10487 (N_10487,N_9778,N_9529);
nor U10488 (N_10488,N_9898,N_9636);
or U10489 (N_10489,N_9757,N_9506);
and U10490 (N_10490,N_9523,N_9795);
nor U10491 (N_10491,N_9581,N_9815);
xnor U10492 (N_10492,N_9732,N_9871);
nand U10493 (N_10493,N_9859,N_9510);
and U10494 (N_10494,N_9944,N_9697);
nor U10495 (N_10495,N_9889,N_9919);
or U10496 (N_10496,N_9514,N_9615);
or U10497 (N_10497,N_9815,N_9960);
or U10498 (N_10498,N_9708,N_9679);
nand U10499 (N_10499,N_9681,N_9651);
nand U10500 (N_10500,N_10223,N_10451);
nand U10501 (N_10501,N_10140,N_10022);
nor U10502 (N_10502,N_10007,N_10214);
xor U10503 (N_10503,N_10490,N_10183);
xnor U10504 (N_10504,N_10295,N_10073);
nor U10505 (N_10505,N_10054,N_10409);
or U10506 (N_10506,N_10215,N_10219);
nand U10507 (N_10507,N_10333,N_10043);
nor U10508 (N_10508,N_10370,N_10011);
or U10509 (N_10509,N_10013,N_10345);
and U10510 (N_10510,N_10119,N_10312);
nor U10511 (N_10511,N_10423,N_10390);
or U10512 (N_10512,N_10006,N_10252);
and U10513 (N_10513,N_10026,N_10275);
nor U10514 (N_10514,N_10354,N_10014);
nor U10515 (N_10515,N_10415,N_10466);
nor U10516 (N_10516,N_10401,N_10450);
or U10517 (N_10517,N_10260,N_10138);
nor U10518 (N_10518,N_10303,N_10489);
nor U10519 (N_10519,N_10123,N_10281);
nand U10520 (N_10520,N_10015,N_10055);
or U10521 (N_10521,N_10030,N_10291);
or U10522 (N_10522,N_10129,N_10106);
and U10523 (N_10523,N_10367,N_10320);
nor U10524 (N_10524,N_10066,N_10203);
nand U10525 (N_10525,N_10440,N_10216);
nor U10526 (N_10526,N_10372,N_10062);
nor U10527 (N_10527,N_10114,N_10069);
nand U10528 (N_10528,N_10381,N_10078);
nor U10529 (N_10529,N_10137,N_10156);
xor U10530 (N_10530,N_10096,N_10496);
and U10531 (N_10531,N_10128,N_10249);
xor U10532 (N_10532,N_10202,N_10186);
or U10533 (N_10533,N_10135,N_10087);
nand U10534 (N_10534,N_10158,N_10472);
and U10535 (N_10535,N_10448,N_10000);
and U10536 (N_10536,N_10175,N_10155);
and U10537 (N_10537,N_10072,N_10082);
xnor U10538 (N_10538,N_10459,N_10134);
xnor U10539 (N_10539,N_10263,N_10467);
xnor U10540 (N_10540,N_10031,N_10171);
xnor U10541 (N_10541,N_10361,N_10301);
and U10542 (N_10542,N_10360,N_10093);
and U10543 (N_10543,N_10331,N_10003);
and U10544 (N_10544,N_10427,N_10235);
nor U10545 (N_10545,N_10244,N_10461);
or U10546 (N_10546,N_10439,N_10229);
and U10547 (N_10547,N_10420,N_10413);
nor U10548 (N_10548,N_10110,N_10391);
xnor U10549 (N_10549,N_10435,N_10288);
and U10550 (N_10550,N_10456,N_10454);
xor U10551 (N_10551,N_10330,N_10233);
nor U10552 (N_10552,N_10463,N_10120);
and U10553 (N_10553,N_10132,N_10254);
nand U10554 (N_10554,N_10259,N_10197);
nand U10555 (N_10555,N_10144,N_10028);
and U10556 (N_10556,N_10111,N_10002);
nand U10557 (N_10557,N_10341,N_10227);
nand U10558 (N_10558,N_10284,N_10344);
and U10559 (N_10559,N_10104,N_10040);
xnor U10560 (N_10560,N_10404,N_10443);
nor U10561 (N_10561,N_10188,N_10178);
or U10562 (N_10562,N_10160,N_10060);
or U10563 (N_10563,N_10152,N_10092);
and U10564 (N_10564,N_10469,N_10280);
nand U10565 (N_10565,N_10416,N_10098);
or U10566 (N_10566,N_10187,N_10293);
or U10567 (N_10567,N_10462,N_10099);
xor U10568 (N_10568,N_10204,N_10185);
and U10569 (N_10569,N_10425,N_10497);
nor U10570 (N_10570,N_10090,N_10273);
xnor U10571 (N_10571,N_10211,N_10327);
or U10572 (N_10572,N_10256,N_10148);
xnor U10573 (N_10573,N_10348,N_10217);
or U10574 (N_10574,N_10210,N_10083);
nand U10575 (N_10575,N_10480,N_10172);
and U10576 (N_10576,N_10085,N_10397);
xnor U10577 (N_10577,N_10473,N_10323);
nor U10578 (N_10578,N_10436,N_10195);
or U10579 (N_10579,N_10097,N_10412);
or U10580 (N_10580,N_10136,N_10116);
nand U10581 (N_10581,N_10200,N_10258);
nor U10582 (N_10582,N_10447,N_10336);
and U10583 (N_10583,N_10351,N_10118);
or U10584 (N_10584,N_10269,N_10322);
and U10585 (N_10585,N_10405,N_10105);
and U10586 (N_10586,N_10262,N_10222);
or U10587 (N_10587,N_10408,N_10292);
nor U10588 (N_10588,N_10008,N_10488);
xnor U10589 (N_10589,N_10154,N_10418);
xor U10590 (N_10590,N_10166,N_10304);
and U10591 (N_10591,N_10316,N_10426);
xnor U10592 (N_10592,N_10274,N_10133);
nor U10593 (N_10593,N_10342,N_10431);
or U10594 (N_10594,N_10143,N_10414);
or U10595 (N_10595,N_10302,N_10057);
and U10596 (N_10596,N_10283,N_10108);
xor U10597 (N_10597,N_10241,N_10368);
and U10598 (N_10598,N_10474,N_10359);
nand U10599 (N_10599,N_10117,N_10220);
nor U10600 (N_10600,N_10061,N_10386);
nor U10601 (N_10601,N_10387,N_10168);
or U10602 (N_10602,N_10430,N_10261);
and U10603 (N_10603,N_10130,N_10157);
and U10604 (N_10604,N_10159,N_10242);
xnor U10605 (N_10605,N_10356,N_10240);
nor U10606 (N_10606,N_10406,N_10319);
or U10607 (N_10607,N_10221,N_10079);
and U10608 (N_10608,N_10433,N_10286);
nand U10609 (N_10609,N_10045,N_10245);
and U10610 (N_10610,N_10324,N_10476);
nand U10611 (N_10611,N_10493,N_10034);
xor U10612 (N_10612,N_10201,N_10174);
nand U10613 (N_10613,N_10306,N_10428);
or U10614 (N_10614,N_10024,N_10343);
or U10615 (N_10615,N_10165,N_10475);
xor U10616 (N_10616,N_10296,N_10206);
nand U10617 (N_10617,N_10021,N_10371);
xor U10618 (N_10618,N_10184,N_10355);
nand U10619 (N_10619,N_10257,N_10094);
or U10620 (N_10620,N_10495,N_10334);
xor U10621 (N_10621,N_10004,N_10102);
nand U10622 (N_10622,N_10470,N_10207);
and U10623 (N_10623,N_10308,N_10363);
and U10624 (N_10624,N_10396,N_10010);
and U10625 (N_10625,N_10032,N_10075);
or U10626 (N_10626,N_10067,N_10246);
or U10627 (N_10627,N_10478,N_10023);
xor U10628 (N_10628,N_10453,N_10411);
nor U10629 (N_10629,N_10176,N_10335);
nor U10630 (N_10630,N_10383,N_10272);
and U10631 (N_10631,N_10276,N_10389);
xor U10632 (N_10632,N_10310,N_10394);
nor U10633 (N_10633,N_10253,N_10100);
and U10634 (N_10634,N_10358,N_10270);
or U10635 (N_10635,N_10374,N_10047);
and U10636 (N_10636,N_10267,N_10329);
xor U10637 (N_10637,N_10499,N_10049);
nor U10638 (N_10638,N_10224,N_10001);
nor U10639 (N_10639,N_10264,N_10337);
nand U10640 (N_10640,N_10313,N_10350);
xnor U10641 (N_10641,N_10321,N_10289);
xor U10642 (N_10642,N_10036,N_10305);
nor U10643 (N_10643,N_10056,N_10027);
nor U10644 (N_10644,N_10146,N_10437);
nor U10645 (N_10645,N_10125,N_10121);
xnor U10646 (N_10646,N_10382,N_10452);
nand U10647 (N_10647,N_10471,N_10053);
and U10648 (N_10648,N_10378,N_10189);
nor U10649 (N_10649,N_10018,N_10194);
and U10650 (N_10650,N_10208,N_10477);
or U10651 (N_10651,N_10226,N_10081);
xor U10652 (N_10652,N_10145,N_10161);
xnor U10653 (N_10653,N_10464,N_10112);
xnor U10654 (N_10654,N_10353,N_10379);
nand U10655 (N_10655,N_10434,N_10277);
nor U10656 (N_10656,N_10339,N_10153);
nor U10657 (N_10657,N_10239,N_10347);
or U10658 (N_10658,N_10063,N_10362);
xnor U10659 (N_10659,N_10167,N_10332);
nor U10660 (N_10660,N_10457,N_10065);
or U10661 (N_10661,N_10050,N_10309);
xor U10662 (N_10662,N_10012,N_10432);
xor U10663 (N_10663,N_10492,N_10016);
nand U10664 (N_10664,N_10460,N_10163);
and U10665 (N_10665,N_10298,N_10248);
and U10666 (N_10666,N_10278,N_10033);
and U10667 (N_10667,N_10421,N_10369);
or U10668 (N_10668,N_10266,N_10046);
xnor U10669 (N_10669,N_10458,N_10131);
and U10670 (N_10670,N_10441,N_10009);
nor U10671 (N_10671,N_10349,N_10212);
xnor U10672 (N_10672,N_10398,N_10044);
nor U10673 (N_10673,N_10429,N_10290);
nand U10674 (N_10674,N_10041,N_10243);
xnor U10675 (N_10675,N_10483,N_10395);
nor U10676 (N_10676,N_10445,N_10139);
nor U10677 (N_10677,N_10232,N_10019);
xor U10678 (N_10678,N_10251,N_10020);
nor U10679 (N_10679,N_10084,N_10279);
nand U10680 (N_10680,N_10255,N_10029);
or U10681 (N_10681,N_10377,N_10237);
or U10682 (N_10682,N_10052,N_10315);
or U10683 (N_10683,N_10205,N_10095);
nand U10684 (N_10684,N_10352,N_10113);
and U10685 (N_10685,N_10268,N_10170);
or U10686 (N_10686,N_10230,N_10192);
and U10687 (N_10687,N_10231,N_10042);
nor U10688 (N_10688,N_10025,N_10228);
xnor U10689 (N_10689,N_10035,N_10070);
and U10690 (N_10690,N_10384,N_10109);
nand U10691 (N_10691,N_10482,N_10039);
nor U10692 (N_10692,N_10299,N_10326);
nand U10693 (N_10693,N_10150,N_10364);
nor U10694 (N_10694,N_10287,N_10058);
xor U10695 (N_10695,N_10089,N_10338);
or U10696 (N_10696,N_10402,N_10051);
nand U10697 (N_10697,N_10271,N_10124);
nand U10698 (N_10698,N_10307,N_10068);
xor U10699 (N_10699,N_10422,N_10455);
and U10700 (N_10700,N_10407,N_10141);
or U10701 (N_10701,N_10285,N_10481);
xor U10702 (N_10702,N_10376,N_10357);
nand U10703 (N_10703,N_10468,N_10325);
xor U10704 (N_10704,N_10162,N_10314);
nand U10705 (N_10705,N_10375,N_10218);
nor U10706 (N_10706,N_10236,N_10196);
and U10707 (N_10707,N_10151,N_10300);
xor U10708 (N_10708,N_10179,N_10126);
and U10709 (N_10709,N_10494,N_10127);
nand U10710 (N_10710,N_10209,N_10080);
xor U10711 (N_10711,N_10449,N_10328);
nor U10712 (N_10712,N_10182,N_10318);
nor U10713 (N_10713,N_10250,N_10380);
and U10714 (N_10714,N_10400,N_10388);
and U10715 (N_10715,N_10142,N_10417);
nor U10716 (N_10716,N_10410,N_10169);
or U10717 (N_10717,N_10491,N_10297);
nor U10718 (N_10718,N_10064,N_10419);
or U10719 (N_10719,N_10190,N_10234);
or U10720 (N_10720,N_10091,N_10446);
or U10721 (N_10721,N_10198,N_10238);
nor U10722 (N_10722,N_10038,N_10294);
and U10723 (N_10723,N_10103,N_10444);
nor U10724 (N_10724,N_10177,N_10115);
nor U10725 (N_10725,N_10181,N_10247);
nor U10726 (N_10726,N_10048,N_10487);
xnor U10727 (N_10727,N_10282,N_10173);
xor U10728 (N_10728,N_10071,N_10191);
nand U10729 (N_10729,N_10346,N_10037);
nor U10730 (N_10730,N_10164,N_10424);
nand U10731 (N_10731,N_10199,N_10147);
nor U10732 (N_10732,N_10442,N_10403);
xnor U10733 (N_10733,N_10393,N_10265);
xor U10734 (N_10734,N_10438,N_10484);
or U10735 (N_10735,N_10465,N_10193);
and U10736 (N_10736,N_10366,N_10373);
xnor U10737 (N_10737,N_10392,N_10017);
nor U10738 (N_10738,N_10479,N_10076);
xor U10739 (N_10739,N_10059,N_10498);
or U10740 (N_10740,N_10213,N_10086);
nor U10741 (N_10741,N_10107,N_10385);
or U10742 (N_10742,N_10122,N_10311);
and U10743 (N_10743,N_10149,N_10340);
and U10744 (N_10744,N_10005,N_10485);
nand U10745 (N_10745,N_10486,N_10399);
nor U10746 (N_10746,N_10074,N_10365);
xor U10747 (N_10747,N_10180,N_10317);
nor U10748 (N_10748,N_10225,N_10088);
xnor U10749 (N_10749,N_10077,N_10101);
and U10750 (N_10750,N_10292,N_10156);
or U10751 (N_10751,N_10132,N_10094);
nand U10752 (N_10752,N_10287,N_10156);
xnor U10753 (N_10753,N_10113,N_10292);
nand U10754 (N_10754,N_10306,N_10285);
xnor U10755 (N_10755,N_10308,N_10052);
nand U10756 (N_10756,N_10089,N_10398);
or U10757 (N_10757,N_10171,N_10211);
xnor U10758 (N_10758,N_10285,N_10240);
nor U10759 (N_10759,N_10287,N_10071);
or U10760 (N_10760,N_10086,N_10130);
or U10761 (N_10761,N_10464,N_10237);
xor U10762 (N_10762,N_10084,N_10217);
and U10763 (N_10763,N_10120,N_10220);
nor U10764 (N_10764,N_10069,N_10415);
or U10765 (N_10765,N_10202,N_10227);
xor U10766 (N_10766,N_10353,N_10014);
and U10767 (N_10767,N_10352,N_10449);
xnor U10768 (N_10768,N_10046,N_10027);
or U10769 (N_10769,N_10317,N_10321);
nor U10770 (N_10770,N_10241,N_10151);
xor U10771 (N_10771,N_10053,N_10042);
xor U10772 (N_10772,N_10013,N_10298);
nand U10773 (N_10773,N_10401,N_10438);
or U10774 (N_10774,N_10173,N_10279);
or U10775 (N_10775,N_10466,N_10024);
nor U10776 (N_10776,N_10029,N_10488);
nand U10777 (N_10777,N_10007,N_10047);
nor U10778 (N_10778,N_10492,N_10290);
nand U10779 (N_10779,N_10443,N_10406);
nand U10780 (N_10780,N_10408,N_10435);
or U10781 (N_10781,N_10030,N_10407);
xor U10782 (N_10782,N_10177,N_10404);
nand U10783 (N_10783,N_10005,N_10310);
or U10784 (N_10784,N_10332,N_10429);
nor U10785 (N_10785,N_10107,N_10095);
xnor U10786 (N_10786,N_10118,N_10110);
and U10787 (N_10787,N_10134,N_10058);
and U10788 (N_10788,N_10434,N_10417);
nand U10789 (N_10789,N_10173,N_10248);
and U10790 (N_10790,N_10327,N_10102);
nor U10791 (N_10791,N_10343,N_10161);
xnor U10792 (N_10792,N_10365,N_10321);
or U10793 (N_10793,N_10292,N_10008);
nor U10794 (N_10794,N_10156,N_10047);
or U10795 (N_10795,N_10219,N_10099);
xnor U10796 (N_10796,N_10019,N_10423);
and U10797 (N_10797,N_10499,N_10391);
nor U10798 (N_10798,N_10391,N_10400);
or U10799 (N_10799,N_10055,N_10160);
nor U10800 (N_10800,N_10422,N_10290);
or U10801 (N_10801,N_10031,N_10002);
or U10802 (N_10802,N_10058,N_10140);
nor U10803 (N_10803,N_10362,N_10008);
nor U10804 (N_10804,N_10310,N_10499);
nand U10805 (N_10805,N_10056,N_10013);
nor U10806 (N_10806,N_10233,N_10488);
nor U10807 (N_10807,N_10147,N_10005);
xor U10808 (N_10808,N_10143,N_10215);
or U10809 (N_10809,N_10455,N_10213);
and U10810 (N_10810,N_10407,N_10064);
or U10811 (N_10811,N_10240,N_10208);
nand U10812 (N_10812,N_10145,N_10284);
and U10813 (N_10813,N_10060,N_10213);
and U10814 (N_10814,N_10455,N_10251);
or U10815 (N_10815,N_10371,N_10264);
nand U10816 (N_10816,N_10215,N_10239);
or U10817 (N_10817,N_10006,N_10371);
nor U10818 (N_10818,N_10299,N_10423);
nand U10819 (N_10819,N_10472,N_10171);
nor U10820 (N_10820,N_10049,N_10165);
or U10821 (N_10821,N_10250,N_10435);
and U10822 (N_10822,N_10144,N_10150);
nor U10823 (N_10823,N_10234,N_10059);
or U10824 (N_10824,N_10276,N_10322);
or U10825 (N_10825,N_10077,N_10451);
nor U10826 (N_10826,N_10193,N_10071);
xnor U10827 (N_10827,N_10042,N_10339);
or U10828 (N_10828,N_10058,N_10342);
nand U10829 (N_10829,N_10198,N_10393);
xor U10830 (N_10830,N_10098,N_10102);
nand U10831 (N_10831,N_10163,N_10195);
or U10832 (N_10832,N_10108,N_10030);
xor U10833 (N_10833,N_10030,N_10406);
nor U10834 (N_10834,N_10014,N_10381);
and U10835 (N_10835,N_10258,N_10087);
nand U10836 (N_10836,N_10464,N_10275);
and U10837 (N_10837,N_10073,N_10442);
and U10838 (N_10838,N_10427,N_10161);
xnor U10839 (N_10839,N_10089,N_10008);
nand U10840 (N_10840,N_10460,N_10226);
or U10841 (N_10841,N_10053,N_10073);
nor U10842 (N_10842,N_10374,N_10193);
nand U10843 (N_10843,N_10165,N_10323);
and U10844 (N_10844,N_10376,N_10420);
xor U10845 (N_10845,N_10381,N_10283);
nand U10846 (N_10846,N_10044,N_10075);
xnor U10847 (N_10847,N_10158,N_10389);
and U10848 (N_10848,N_10318,N_10123);
and U10849 (N_10849,N_10364,N_10279);
or U10850 (N_10850,N_10487,N_10342);
nand U10851 (N_10851,N_10444,N_10062);
xnor U10852 (N_10852,N_10317,N_10490);
nand U10853 (N_10853,N_10280,N_10255);
nand U10854 (N_10854,N_10454,N_10143);
and U10855 (N_10855,N_10386,N_10137);
and U10856 (N_10856,N_10046,N_10146);
nand U10857 (N_10857,N_10126,N_10210);
or U10858 (N_10858,N_10492,N_10165);
and U10859 (N_10859,N_10303,N_10398);
or U10860 (N_10860,N_10202,N_10077);
or U10861 (N_10861,N_10017,N_10470);
nor U10862 (N_10862,N_10033,N_10486);
or U10863 (N_10863,N_10151,N_10265);
or U10864 (N_10864,N_10311,N_10043);
xor U10865 (N_10865,N_10303,N_10323);
and U10866 (N_10866,N_10315,N_10107);
and U10867 (N_10867,N_10448,N_10176);
and U10868 (N_10868,N_10414,N_10299);
and U10869 (N_10869,N_10281,N_10211);
nor U10870 (N_10870,N_10392,N_10220);
nand U10871 (N_10871,N_10357,N_10284);
or U10872 (N_10872,N_10457,N_10171);
and U10873 (N_10873,N_10261,N_10121);
nand U10874 (N_10874,N_10399,N_10060);
nor U10875 (N_10875,N_10346,N_10306);
and U10876 (N_10876,N_10058,N_10375);
nand U10877 (N_10877,N_10393,N_10132);
or U10878 (N_10878,N_10155,N_10325);
and U10879 (N_10879,N_10435,N_10240);
nor U10880 (N_10880,N_10109,N_10458);
xnor U10881 (N_10881,N_10408,N_10011);
or U10882 (N_10882,N_10217,N_10137);
nor U10883 (N_10883,N_10465,N_10203);
xnor U10884 (N_10884,N_10113,N_10296);
nand U10885 (N_10885,N_10292,N_10047);
xor U10886 (N_10886,N_10370,N_10055);
xnor U10887 (N_10887,N_10328,N_10306);
nand U10888 (N_10888,N_10363,N_10101);
and U10889 (N_10889,N_10168,N_10421);
nand U10890 (N_10890,N_10498,N_10455);
or U10891 (N_10891,N_10322,N_10377);
and U10892 (N_10892,N_10352,N_10437);
nor U10893 (N_10893,N_10022,N_10071);
and U10894 (N_10894,N_10343,N_10205);
nand U10895 (N_10895,N_10382,N_10332);
nand U10896 (N_10896,N_10162,N_10434);
xor U10897 (N_10897,N_10470,N_10310);
nand U10898 (N_10898,N_10402,N_10221);
or U10899 (N_10899,N_10250,N_10106);
nand U10900 (N_10900,N_10137,N_10032);
nor U10901 (N_10901,N_10473,N_10284);
and U10902 (N_10902,N_10421,N_10125);
nand U10903 (N_10903,N_10096,N_10358);
xnor U10904 (N_10904,N_10377,N_10253);
and U10905 (N_10905,N_10275,N_10073);
and U10906 (N_10906,N_10150,N_10138);
and U10907 (N_10907,N_10020,N_10039);
and U10908 (N_10908,N_10428,N_10497);
nor U10909 (N_10909,N_10362,N_10125);
or U10910 (N_10910,N_10340,N_10043);
xnor U10911 (N_10911,N_10364,N_10382);
nand U10912 (N_10912,N_10357,N_10417);
xor U10913 (N_10913,N_10030,N_10362);
nand U10914 (N_10914,N_10019,N_10122);
and U10915 (N_10915,N_10361,N_10338);
nor U10916 (N_10916,N_10499,N_10444);
and U10917 (N_10917,N_10053,N_10485);
and U10918 (N_10918,N_10332,N_10197);
and U10919 (N_10919,N_10363,N_10236);
and U10920 (N_10920,N_10007,N_10305);
xor U10921 (N_10921,N_10393,N_10018);
or U10922 (N_10922,N_10042,N_10257);
xor U10923 (N_10923,N_10134,N_10398);
nor U10924 (N_10924,N_10051,N_10417);
nor U10925 (N_10925,N_10117,N_10392);
and U10926 (N_10926,N_10347,N_10147);
xor U10927 (N_10927,N_10346,N_10220);
and U10928 (N_10928,N_10036,N_10083);
nor U10929 (N_10929,N_10004,N_10058);
xnor U10930 (N_10930,N_10147,N_10382);
xor U10931 (N_10931,N_10005,N_10054);
or U10932 (N_10932,N_10315,N_10392);
nand U10933 (N_10933,N_10063,N_10489);
nand U10934 (N_10934,N_10098,N_10020);
xor U10935 (N_10935,N_10451,N_10003);
nor U10936 (N_10936,N_10248,N_10425);
xnor U10937 (N_10937,N_10498,N_10335);
nand U10938 (N_10938,N_10043,N_10138);
and U10939 (N_10939,N_10324,N_10400);
or U10940 (N_10940,N_10133,N_10293);
and U10941 (N_10941,N_10261,N_10314);
nor U10942 (N_10942,N_10111,N_10389);
and U10943 (N_10943,N_10294,N_10234);
and U10944 (N_10944,N_10455,N_10032);
or U10945 (N_10945,N_10108,N_10214);
nand U10946 (N_10946,N_10277,N_10293);
and U10947 (N_10947,N_10471,N_10475);
nor U10948 (N_10948,N_10202,N_10098);
xnor U10949 (N_10949,N_10465,N_10178);
nor U10950 (N_10950,N_10216,N_10123);
and U10951 (N_10951,N_10424,N_10440);
xnor U10952 (N_10952,N_10382,N_10198);
xor U10953 (N_10953,N_10432,N_10410);
or U10954 (N_10954,N_10231,N_10326);
or U10955 (N_10955,N_10265,N_10298);
and U10956 (N_10956,N_10000,N_10304);
nand U10957 (N_10957,N_10275,N_10413);
and U10958 (N_10958,N_10422,N_10176);
and U10959 (N_10959,N_10354,N_10383);
nand U10960 (N_10960,N_10490,N_10428);
xor U10961 (N_10961,N_10254,N_10283);
and U10962 (N_10962,N_10119,N_10092);
nand U10963 (N_10963,N_10465,N_10397);
nor U10964 (N_10964,N_10449,N_10388);
nor U10965 (N_10965,N_10212,N_10074);
or U10966 (N_10966,N_10010,N_10335);
and U10967 (N_10967,N_10102,N_10220);
or U10968 (N_10968,N_10158,N_10185);
nand U10969 (N_10969,N_10270,N_10276);
and U10970 (N_10970,N_10464,N_10480);
nand U10971 (N_10971,N_10092,N_10389);
and U10972 (N_10972,N_10263,N_10214);
and U10973 (N_10973,N_10207,N_10178);
and U10974 (N_10974,N_10376,N_10390);
and U10975 (N_10975,N_10394,N_10079);
nand U10976 (N_10976,N_10236,N_10388);
and U10977 (N_10977,N_10253,N_10416);
nand U10978 (N_10978,N_10022,N_10498);
nand U10979 (N_10979,N_10069,N_10381);
or U10980 (N_10980,N_10475,N_10110);
nand U10981 (N_10981,N_10429,N_10105);
nor U10982 (N_10982,N_10154,N_10489);
nor U10983 (N_10983,N_10092,N_10062);
nand U10984 (N_10984,N_10066,N_10241);
nand U10985 (N_10985,N_10483,N_10002);
nand U10986 (N_10986,N_10415,N_10208);
nor U10987 (N_10987,N_10085,N_10103);
nand U10988 (N_10988,N_10267,N_10268);
xor U10989 (N_10989,N_10301,N_10407);
nor U10990 (N_10990,N_10267,N_10424);
nand U10991 (N_10991,N_10405,N_10110);
nor U10992 (N_10992,N_10010,N_10077);
xnor U10993 (N_10993,N_10094,N_10118);
nor U10994 (N_10994,N_10414,N_10106);
nor U10995 (N_10995,N_10214,N_10382);
nand U10996 (N_10996,N_10012,N_10283);
or U10997 (N_10997,N_10111,N_10284);
nor U10998 (N_10998,N_10128,N_10445);
and U10999 (N_10999,N_10463,N_10438);
nand U11000 (N_11000,N_10660,N_10911);
or U11001 (N_11001,N_10916,N_10574);
xnor U11002 (N_11002,N_10745,N_10625);
and U11003 (N_11003,N_10606,N_10759);
nand U11004 (N_11004,N_10630,N_10912);
nand U11005 (N_11005,N_10835,N_10667);
nand U11006 (N_11006,N_10866,N_10734);
nor U11007 (N_11007,N_10590,N_10615);
and U11008 (N_11008,N_10897,N_10949);
nor U11009 (N_11009,N_10594,N_10683);
nand U11010 (N_11010,N_10885,N_10591);
xor U11011 (N_11011,N_10570,N_10658);
or U11012 (N_11012,N_10882,N_10635);
and U11013 (N_11013,N_10676,N_10934);
nand U11014 (N_11014,N_10673,N_10741);
nand U11015 (N_11015,N_10604,N_10889);
xnor U11016 (N_11016,N_10770,N_10657);
or U11017 (N_11017,N_10565,N_10593);
nor U11018 (N_11018,N_10808,N_10905);
or U11019 (N_11019,N_10785,N_10776);
nand U11020 (N_11020,N_10787,N_10925);
nand U11021 (N_11021,N_10620,N_10576);
nor U11022 (N_11022,N_10645,N_10842);
xor U11023 (N_11023,N_10730,N_10780);
xnor U11024 (N_11024,N_10709,N_10539);
xor U11025 (N_11025,N_10598,N_10840);
and U11026 (N_11026,N_10806,N_10633);
and U11027 (N_11027,N_10874,N_10860);
nor U11028 (N_11028,N_10611,N_10650);
or U11029 (N_11029,N_10551,N_10777);
nor U11030 (N_11030,N_10967,N_10568);
nand U11031 (N_11031,N_10783,N_10721);
nand U11032 (N_11032,N_10970,N_10861);
and U11033 (N_11033,N_10933,N_10750);
and U11034 (N_11034,N_10548,N_10671);
nand U11035 (N_11035,N_10538,N_10752);
or U11036 (N_11036,N_10743,N_10838);
or U11037 (N_11037,N_10832,N_10844);
xnor U11038 (N_11038,N_10554,N_10731);
and U11039 (N_11039,N_10940,N_10772);
and U11040 (N_11040,N_10955,N_10631);
xnor U11041 (N_11041,N_10675,N_10899);
nand U11042 (N_11042,N_10792,N_10690);
xnor U11043 (N_11043,N_10504,N_10677);
or U11044 (N_11044,N_10978,N_10878);
nor U11045 (N_11045,N_10917,N_10961);
or U11046 (N_11046,N_10986,N_10900);
nor U11047 (N_11047,N_10999,N_10754);
xnor U11048 (N_11048,N_10960,N_10664);
nor U11049 (N_11049,N_10649,N_10848);
nor U11050 (N_11050,N_10890,N_10722);
and U11051 (N_11051,N_10951,N_10699);
and U11052 (N_11052,N_10821,N_10617);
and U11053 (N_11053,N_10862,N_10627);
nand U11054 (N_11054,N_10869,N_10796);
xor U11055 (N_11055,N_10875,N_10534);
and U11056 (N_11056,N_10541,N_10725);
nor U11057 (N_11057,N_10510,N_10863);
nor U11058 (N_11058,N_10995,N_10597);
or U11059 (N_11059,N_10872,N_10605);
and U11060 (N_11060,N_10518,N_10910);
nor U11061 (N_11061,N_10589,N_10527);
nor U11062 (N_11062,N_10824,N_10540);
or U11063 (N_11063,N_10585,N_10569);
and U11064 (N_11064,N_10566,N_10798);
nor U11065 (N_11065,N_10942,N_10966);
nor U11066 (N_11066,N_10694,N_10713);
nand U11067 (N_11067,N_10572,N_10755);
nand U11068 (N_11068,N_10523,N_10877);
nor U11069 (N_11069,N_10564,N_10829);
or U11070 (N_11070,N_10624,N_10950);
xor U11071 (N_11071,N_10791,N_10653);
or U11072 (N_11072,N_10674,N_10853);
nor U11073 (N_11073,N_10610,N_10517);
xnor U11074 (N_11074,N_10632,N_10825);
nor U11075 (N_11075,N_10726,N_10507);
nand U11076 (N_11076,N_10827,N_10904);
nor U11077 (N_11077,N_10662,N_10758);
nor U11078 (N_11078,N_10747,N_10854);
nor U11079 (N_11079,N_10587,N_10839);
or U11080 (N_11080,N_10810,N_10544);
or U11081 (N_11081,N_10719,N_10663);
nor U11082 (N_11082,N_10710,N_10870);
or U11083 (N_11083,N_10816,N_10828);
or U11084 (N_11084,N_10814,N_10740);
or U11085 (N_11085,N_10919,N_10707);
xnor U11086 (N_11086,N_10943,N_10580);
nor U11087 (N_11087,N_10879,N_10998);
xnor U11088 (N_11088,N_10833,N_10962);
or U11089 (N_11089,N_10815,N_10669);
nand U11090 (N_11090,N_10773,N_10644);
and U11091 (N_11091,N_10898,N_10531);
nor U11092 (N_11092,N_10646,N_10768);
and U11093 (N_11093,N_10502,N_10621);
nand U11094 (N_11094,N_10774,N_10603);
nand U11095 (N_11095,N_10855,N_10928);
or U11096 (N_11096,N_10563,N_10948);
and U11097 (N_11097,N_10931,N_10884);
and U11098 (N_11098,N_10636,N_10975);
nor U11099 (N_11099,N_10913,N_10915);
xor U11100 (N_11100,N_10512,N_10926);
nand U11101 (N_11101,N_10573,N_10953);
and U11102 (N_11102,N_10515,N_10584);
or U11103 (N_11103,N_10642,N_10562);
and U11104 (N_11104,N_10845,N_10641);
nor U11105 (N_11105,N_10972,N_10764);
nand U11106 (N_11106,N_10763,N_10516);
xnor U11107 (N_11107,N_10982,N_10742);
nor U11108 (N_11108,N_10880,N_10537);
nand U11109 (N_11109,N_10823,N_10588);
and U11110 (N_11110,N_10685,N_10684);
nand U11111 (N_11111,N_10647,N_10968);
or U11112 (N_11112,N_10867,N_10729);
and U11113 (N_11113,N_10756,N_10766);
and U11114 (N_11114,N_10637,N_10914);
or U11115 (N_11115,N_10638,N_10891);
nand U11116 (N_11116,N_10571,N_10530);
or U11117 (N_11117,N_10941,N_10733);
nand U11118 (N_11118,N_10993,N_10822);
and U11119 (N_11119,N_10689,N_10586);
nor U11120 (N_11120,N_10503,N_10757);
nand U11121 (N_11121,N_10522,N_10618);
nand U11122 (N_11122,N_10944,N_10918);
xnor U11123 (N_11123,N_10923,N_10679);
or U11124 (N_11124,N_10697,N_10672);
or U11125 (N_11125,N_10850,N_10909);
nand U11126 (N_11126,N_10881,N_10558);
nor U11127 (N_11127,N_10991,N_10852);
and U11128 (N_11128,N_10996,N_10871);
and U11129 (N_11129,N_10578,N_10985);
nor U11130 (N_11130,N_10612,N_10864);
nor U11131 (N_11131,N_10989,N_10629);
or U11132 (N_11132,N_10924,N_10525);
nor U11133 (N_11133,N_10920,N_10681);
nor U11134 (N_11134,N_10735,N_10765);
nand U11135 (N_11135,N_10847,N_10997);
nand U11136 (N_11136,N_10784,N_10983);
nand U11137 (N_11137,N_10720,N_10686);
xnor U11138 (N_11138,N_10805,N_10936);
and U11139 (N_11139,N_10728,N_10732);
and U11140 (N_11140,N_10818,N_10809);
and U11141 (N_11141,N_10526,N_10797);
and U11142 (N_11142,N_10979,N_10613);
xor U11143 (N_11143,N_10813,N_10581);
or U11144 (N_11144,N_10939,N_10654);
nor U11145 (N_11145,N_10511,N_10799);
nor U11146 (N_11146,N_10557,N_10521);
nand U11147 (N_11147,N_10789,N_10536);
xnor U11148 (N_11148,N_10836,N_10958);
and U11149 (N_11149,N_10746,N_10807);
or U11150 (N_11150,N_10820,N_10841);
xor U11151 (N_11151,N_10906,N_10856);
xor U11152 (N_11152,N_10506,N_10665);
or U11153 (N_11153,N_10990,N_10802);
nand U11154 (N_11154,N_10577,N_10894);
and U11155 (N_11155,N_10553,N_10737);
nor U11156 (N_11156,N_10529,N_10701);
nor U11157 (N_11157,N_10753,N_10937);
and U11158 (N_11158,N_10984,N_10930);
or U11159 (N_11159,N_10819,N_10851);
nand U11160 (N_11160,N_10767,N_10843);
nand U11161 (N_11161,N_10678,N_10692);
xnor U11162 (N_11162,N_10771,N_10501);
or U11163 (N_11163,N_10602,N_10609);
or U11164 (N_11164,N_10957,N_10668);
and U11165 (N_11165,N_10691,N_10727);
or U11166 (N_11166,N_10788,N_10542);
or U11167 (N_11167,N_10888,N_10932);
xor U11168 (N_11168,N_10579,N_10549);
xor U11169 (N_11169,N_10831,N_10801);
nand U11170 (N_11170,N_10670,N_10688);
xor U11171 (N_11171,N_10698,N_10849);
or U11172 (N_11172,N_10595,N_10626);
nand U11173 (N_11173,N_10896,N_10723);
nand U11174 (N_11174,N_10552,N_10736);
or U11175 (N_11175,N_10859,N_10614);
nand U11176 (N_11176,N_10706,N_10708);
xor U11177 (N_11177,N_10519,N_10976);
or U11178 (N_11178,N_10945,N_10546);
nand U11179 (N_11179,N_10769,N_10837);
and U11180 (N_11180,N_10744,N_10717);
and U11181 (N_11181,N_10971,N_10956);
nand U11182 (N_11182,N_10718,N_10892);
nor U11183 (N_11183,N_10600,N_10749);
nor U11184 (N_11184,N_10596,N_10508);
nor U11185 (N_11185,N_10947,N_10651);
nand U11186 (N_11186,N_10927,N_10567);
nand U11187 (N_11187,N_10704,N_10500);
and U11188 (N_11188,N_10703,N_10908);
and U11189 (N_11189,N_10994,N_10607);
nand U11190 (N_11190,N_10505,N_10830);
nand U11191 (N_11191,N_10693,N_10560);
and U11192 (N_11192,N_10901,N_10963);
xnor U11193 (N_11193,N_10616,N_10778);
nor U11194 (N_11194,N_10826,N_10751);
nand U11195 (N_11195,N_10846,N_10887);
nand U11196 (N_11196,N_10700,N_10652);
nor U11197 (N_11197,N_10903,N_10550);
and U11198 (N_11198,N_10643,N_10938);
xnor U11199 (N_11199,N_10781,N_10795);
nor U11200 (N_11200,N_10954,N_10794);
nand U11201 (N_11201,N_10812,N_10648);
nor U11202 (N_11202,N_10582,N_10779);
nor U11203 (N_11203,N_10682,N_10858);
nor U11204 (N_11204,N_10992,N_10680);
and U11205 (N_11205,N_10656,N_10528);
or U11206 (N_11206,N_10974,N_10738);
nor U11207 (N_11207,N_10661,N_10556);
or U11208 (N_11208,N_10599,N_10760);
nor U11209 (N_11209,N_10705,N_10762);
or U11210 (N_11210,N_10714,N_10639);
nor U11211 (N_11211,N_10561,N_10761);
xnor U11212 (N_11212,N_10575,N_10748);
xor U11213 (N_11213,N_10817,N_10811);
nand U11214 (N_11214,N_10775,N_10868);
nand U11215 (N_11215,N_10702,N_10634);
xnor U11216 (N_11216,N_10907,N_10782);
xnor U11217 (N_11217,N_10977,N_10959);
nand U11218 (N_11218,N_10623,N_10902);
nand U11219 (N_11219,N_10659,N_10524);
or U11220 (N_11220,N_10793,N_10886);
nand U11221 (N_11221,N_10592,N_10724);
xnor U11222 (N_11222,N_10981,N_10922);
nor U11223 (N_11223,N_10895,N_10969);
and U11224 (N_11224,N_10695,N_10987);
nor U11225 (N_11225,N_10543,N_10857);
or U11226 (N_11226,N_10804,N_10622);
and U11227 (N_11227,N_10555,N_10559);
nor U11228 (N_11228,N_10883,N_10952);
and U11229 (N_11229,N_10964,N_10973);
nand U11230 (N_11230,N_10535,N_10965);
xnor U11231 (N_11231,N_10929,N_10696);
nor U11232 (N_11232,N_10786,N_10865);
nand U11233 (N_11233,N_10800,N_10790);
xnor U11234 (N_11234,N_10980,N_10509);
nor U11235 (N_11235,N_10715,N_10514);
and U11236 (N_11236,N_10988,N_10608);
nor U11237 (N_11237,N_10946,N_10834);
xnor U11238 (N_11238,N_10712,N_10921);
xnor U11239 (N_11239,N_10666,N_10628);
nand U11240 (N_11240,N_10532,N_10545);
or U11241 (N_11241,N_10533,N_10655);
nand U11242 (N_11242,N_10803,N_10520);
or U11243 (N_11243,N_10547,N_10876);
and U11244 (N_11244,N_10711,N_10687);
nor U11245 (N_11245,N_10873,N_10640);
or U11246 (N_11246,N_10935,N_10601);
and U11247 (N_11247,N_10716,N_10619);
xor U11248 (N_11248,N_10513,N_10583);
or U11249 (N_11249,N_10739,N_10893);
or U11250 (N_11250,N_10635,N_10582);
nand U11251 (N_11251,N_10636,N_10752);
and U11252 (N_11252,N_10825,N_10789);
or U11253 (N_11253,N_10671,N_10880);
and U11254 (N_11254,N_10963,N_10713);
nand U11255 (N_11255,N_10538,N_10942);
or U11256 (N_11256,N_10624,N_10513);
nand U11257 (N_11257,N_10670,N_10570);
nand U11258 (N_11258,N_10579,N_10671);
nor U11259 (N_11259,N_10573,N_10777);
and U11260 (N_11260,N_10620,N_10662);
nor U11261 (N_11261,N_10775,N_10897);
or U11262 (N_11262,N_10537,N_10581);
xor U11263 (N_11263,N_10520,N_10693);
xnor U11264 (N_11264,N_10949,N_10839);
xnor U11265 (N_11265,N_10751,N_10894);
and U11266 (N_11266,N_10620,N_10505);
and U11267 (N_11267,N_10918,N_10853);
or U11268 (N_11268,N_10694,N_10886);
or U11269 (N_11269,N_10537,N_10913);
and U11270 (N_11270,N_10879,N_10985);
nand U11271 (N_11271,N_10639,N_10687);
nand U11272 (N_11272,N_10919,N_10802);
and U11273 (N_11273,N_10712,N_10573);
nor U11274 (N_11274,N_10573,N_10921);
nor U11275 (N_11275,N_10694,N_10541);
or U11276 (N_11276,N_10790,N_10987);
nand U11277 (N_11277,N_10740,N_10910);
nor U11278 (N_11278,N_10975,N_10695);
nor U11279 (N_11279,N_10923,N_10654);
xnor U11280 (N_11280,N_10944,N_10517);
nor U11281 (N_11281,N_10740,N_10792);
and U11282 (N_11282,N_10822,N_10911);
nor U11283 (N_11283,N_10649,N_10911);
nor U11284 (N_11284,N_10527,N_10795);
nor U11285 (N_11285,N_10825,N_10853);
nand U11286 (N_11286,N_10844,N_10648);
nand U11287 (N_11287,N_10609,N_10643);
or U11288 (N_11288,N_10675,N_10755);
nand U11289 (N_11289,N_10993,N_10584);
and U11290 (N_11290,N_10939,N_10824);
nand U11291 (N_11291,N_10537,N_10577);
and U11292 (N_11292,N_10719,N_10965);
nor U11293 (N_11293,N_10796,N_10541);
nand U11294 (N_11294,N_10560,N_10847);
xor U11295 (N_11295,N_10650,N_10606);
and U11296 (N_11296,N_10540,N_10502);
or U11297 (N_11297,N_10816,N_10982);
xor U11298 (N_11298,N_10856,N_10615);
and U11299 (N_11299,N_10913,N_10811);
nand U11300 (N_11300,N_10549,N_10956);
or U11301 (N_11301,N_10719,N_10850);
xnor U11302 (N_11302,N_10745,N_10608);
nor U11303 (N_11303,N_10942,N_10607);
nand U11304 (N_11304,N_10961,N_10880);
nand U11305 (N_11305,N_10921,N_10525);
nor U11306 (N_11306,N_10766,N_10734);
and U11307 (N_11307,N_10690,N_10912);
and U11308 (N_11308,N_10653,N_10575);
nand U11309 (N_11309,N_10632,N_10730);
xnor U11310 (N_11310,N_10533,N_10836);
nor U11311 (N_11311,N_10740,N_10698);
nor U11312 (N_11312,N_10717,N_10500);
or U11313 (N_11313,N_10841,N_10516);
xor U11314 (N_11314,N_10813,N_10903);
nand U11315 (N_11315,N_10996,N_10525);
xnor U11316 (N_11316,N_10537,N_10601);
xor U11317 (N_11317,N_10939,N_10883);
nor U11318 (N_11318,N_10668,N_10992);
and U11319 (N_11319,N_10878,N_10706);
xnor U11320 (N_11320,N_10685,N_10746);
and U11321 (N_11321,N_10880,N_10802);
and U11322 (N_11322,N_10795,N_10565);
or U11323 (N_11323,N_10569,N_10784);
and U11324 (N_11324,N_10537,N_10630);
nand U11325 (N_11325,N_10917,N_10697);
or U11326 (N_11326,N_10976,N_10623);
nor U11327 (N_11327,N_10616,N_10793);
nand U11328 (N_11328,N_10714,N_10758);
and U11329 (N_11329,N_10673,N_10755);
nand U11330 (N_11330,N_10607,N_10740);
nor U11331 (N_11331,N_10769,N_10605);
nor U11332 (N_11332,N_10827,N_10552);
and U11333 (N_11333,N_10878,N_10686);
xnor U11334 (N_11334,N_10502,N_10748);
xor U11335 (N_11335,N_10948,N_10884);
xnor U11336 (N_11336,N_10909,N_10647);
and U11337 (N_11337,N_10876,N_10772);
or U11338 (N_11338,N_10711,N_10591);
and U11339 (N_11339,N_10784,N_10714);
and U11340 (N_11340,N_10784,N_10655);
and U11341 (N_11341,N_10901,N_10528);
nand U11342 (N_11342,N_10595,N_10814);
nor U11343 (N_11343,N_10760,N_10948);
xnor U11344 (N_11344,N_10950,N_10519);
nor U11345 (N_11345,N_10672,N_10614);
or U11346 (N_11346,N_10857,N_10509);
nand U11347 (N_11347,N_10886,N_10950);
xnor U11348 (N_11348,N_10980,N_10783);
nand U11349 (N_11349,N_10935,N_10837);
or U11350 (N_11350,N_10935,N_10575);
and U11351 (N_11351,N_10665,N_10974);
xor U11352 (N_11352,N_10600,N_10912);
nand U11353 (N_11353,N_10951,N_10604);
nand U11354 (N_11354,N_10727,N_10794);
or U11355 (N_11355,N_10583,N_10813);
nor U11356 (N_11356,N_10664,N_10760);
or U11357 (N_11357,N_10858,N_10805);
nor U11358 (N_11358,N_10752,N_10829);
or U11359 (N_11359,N_10955,N_10777);
nor U11360 (N_11360,N_10760,N_10657);
or U11361 (N_11361,N_10907,N_10816);
xor U11362 (N_11362,N_10671,N_10876);
nor U11363 (N_11363,N_10770,N_10939);
nand U11364 (N_11364,N_10993,N_10918);
nand U11365 (N_11365,N_10889,N_10539);
and U11366 (N_11366,N_10510,N_10859);
xor U11367 (N_11367,N_10715,N_10862);
and U11368 (N_11368,N_10851,N_10839);
nor U11369 (N_11369,N_10803,N_10784);
and U11370 (N_11370,N_10832,N_10554);
nand U11371 (N_11371,N_10834,N_10615);
and U11372 (N_11372,N_10671,N_10739);
or U11373 (N_11373,N_10672,N_10781);
and U11374 (N_11374,N_10980,N_10590);
xnor U11375 (N_11375,N_10967,N_10575);
xnor U11376 (N_11376,N_10861,N_10876);
xnor U11377 (N_11377,N_10608,N_10808);
nand U11378 (N_11378,N_10847,N_10635);
xor U11379 (N_11379,N_10819,N_10729);
nand U11380 (N_11380,N_10755,N_10720);
nor U11381 (N_11381,N_10853,N_10901);
nand U11382 (N_11382,N_10547,N_10987);
xor U11383 (N_11383,N_10685,N_10760);
and U11384 (N_11384,N_10710,N_10704);
nand U11385 (N_11385,N_10711,N_10558);
xnor U11386 (N_11386,N_10563,N_10607);
xor U11387 (N_11387,N_10647,N_10605);
or U11388 (N_11388,N_10594,N_10612);
nand U11389 (N_11389,N_10849,N_10510);
xor U11390 (N_11390,N_10665,N_10840);
and U11391 (N_11391,N_10703,N_10869);
nor U11392 (N_11392,N_10713,N_10601);
nor U11393 (N_11393,N_10780,N_10556);
and U11394 (N_11394,N_10929,N_10897);
nor U11395 (N_11395,N_10992,N_10595);
or U11396 (N_11396,N_10514,N_10993);
nor U11397 (N_11397,N_10997,N_10564);
and U11398 (N_11398,N_10637,N_10857);
or U11399 (N_11399,N_10537,N_10639);
nor U11400 (N_11400,N_10576,N_10756);
xor U11401 (N_11401,N_10760,N_10892);
nor U11402 (N_11402,N_10653,N_10546);
nand U11403 (N_11403,N_10938,N_10729);
xnor U11404 (N_11404,N_10860,N_10986);
xnor U11405 (N_11405,N_10955,N_10618);
and U11406 (N_11406,N_10939,N_10992);
or U11407 (N_11407,N_10555,N_10921);
nor U11408 (N_11408,N_10771,N_10990);
xnor U11409 (N_11409,N_10758,N_10844);
or U11410 (N_11410,N_10749,N_10755);
and U11411 (N_11411,N_10652,N_10715);
xnor U11412 (N_11412,N_10710,N_10902);
xor U11413 (N_11413,N_10608,N_10559);
nor U11414 (N_11414,N_10960,N_10733);
xor U11415 (N_11415,N_10873,N_10569);
and U11416 (N_11416,N_10775,N_10661);
and U11417 (N_11417,N_10954,N_10618);
nand U11418 (N_11418,N_10632,N_10560);
xnor U11419 (N_11419,N_10541,N_10517);
xnor U11420 (N_11420,N_10888,N_10599);
and U11421 (N_11421,N_10580,N_10863);
or U11422 (N_11422,N_10874,N_10627);
nand U11423 (N_11423,N_10659,N_10699);
xor U11424 (N_11424,N_10677,N_10685);
or U11425 (N_11425,N_10811,N_10814);
or U11426 (N_11426,N_10518,N_10628);
nand U11427 (N_11427,N_10509,N_10591);
xnor U11428 (N_11428,N_10606,N_10909);
nand U11429 (N_11429,N_10965,N_10775);
or U11430 (N_11430,N_10961,N_10661);
and U11431 (N_11431,N_10608,N_10863);
nor U11432 (N_11432,N_10859,N_10787);
and U11433 (N_11433,N_10635,N_10934);
nor U11434 (N_11434,N_10729,N_10801);
or U11435 (N_11435,N_10603,N_10820);
or U11436 (N_11436,N_10826,N_10691);
and U11437 (N_11437,N_10666,N_10703);
and U11438 (N_11438,N_10544,N_10662);
and U11439 (N_11439,N_10537,N_10621);
xor U11440 (N_11440,N_10629,N_10797);
or U11441 (N_11441,N_10751,N_10524);
nand U11442 (N_11442,N_10830,N_10724);
or U11443 (N_11443,N_10621,N_10963);
xor U11444 (N_11444,N_10627,N_10938);
or U11445 (N_11445,N_10844,N_10789);
nand U11446 (N_11446,N_10996,N_10595);
nor U11447 (N_11447,N_10933,N_10514);
xnor U11448 (N_11448,N_10658,N_10602);
or U11449 (N_11449,N_10871,N_10808);
xnor U11450 (N_11450,N_10535,N_10576);
or U11451 (N_11451,N_10864,N_10821);
xor U11452 (N_11452,N_10599,N_10913);
nand U11453 (N_11453,N_10766,N_10730);
and U11454 (N_11454,N_10953,N_10593);
and U11455 (N_11455,N_10689,N_10842);
and U11456 (N_11456,N_10505,N_10791);
xor U11457 (N_11457,N_10546,N_10778);
xnor U11458 (N_11458,N_10872,N_10916);
nor U11459 (N_11459,N_10542,N_10633);
nor U11460 (N_11460,N_10598,N_10543);
or U11461 (N_11461,N_10601,N_10715);
nor U11462 (N_11462,N_10811,N_10746);
nor U11463 (N_11463,N_10977,N_10596);
nor U11464 (N_11464,N_10909,N_10875);
nor U11465 (N_11465,N_10665,N_10543);
or U11466 (N_11466,N_10730,N_10744);
or U11467 (N_11467,N_10529,N_10541);
xnor U11468 (N_11468,N_10655,N_10689);
or U11469 (N_11469,N_10619,N_10863);
or U11470 (N_11470,N_10724,N_10617);
nor U11471 (N_11471,N_10770,N_10832);
xor U11472 (N_11472,N_10970,N_10723);
or U11473 (N_11473,N_10815,N_10510);
nor U11474 (N_11474,N_10704,N_10675);
and U11475 (N_11475,N_10525,N_10768);
and U11476 (N_11476,N_10942,N_10653);
or U11477 (N_11477,N_10905,N_10916);
xor U11478 (N_11478,N_10808,N_10615);
xnor U11479 (N_11479,N_10606,N_10754);
or U11480 (N_11480,N_10959,N_10915);
nor U11481 (N_11481,N_10940,N_10660);
and U11482 (N_11482,N_10700,N_10661);
or U11483 (N_11483,N_10583,N_10922);
and U11484 (N_11484,N_10939,N_10680);
and U11485 (N_11485,N_10662,N_10731);
nand U11486 (N_11486,N_10582,N_10749);
or U11487 (N_11487,N_10824,N_10619);
nand U11488 (N_11488,N_10705,N_10685);
xor U11489 (N_11489,N_10889,N_10514);
and U11490 (N_11490,N_10600,N_10826);
or U11491 (N_11491,N_10840,N_10553);
nand U11492 (N_11492,N_10929,N_10883);
or U11493 (N_11493,N_10502,N_10830);
and U11494 (N_11494,N_10844,N_10681);
nand U11495 (N_11495,N_10939,N_10629);
and U11496 (N_11496,N_10978,N_10633);
or U11497 (N_11497,N_10884,N_10772);
nand U11498 (N_11498,N_10618,N_10857);
nand U11499 (N_11499,N_10802,N_10797);
or U11500 (N_11500,N_11140,N_11065);
or U11501 (N_11501,N_11024,N_11409);
xnor U11502 (N_11502,N_11273,N_11298);
and U11503 (N_11503,N_11057,N_11306);
or U11504 (N_11504,N_11494,N_11170);
xnor U11505 (N_11505,N_11437,N_11233);
nor U11506 (N_11506,N_11261,N_11412);
and U11507 (N_11507,N_11434,N_11142);
nor U11508 (N_11508,N_11270,N_11439);
nor U11509 (N_11509,N_11429,N_11042);
or U11510 (N_11510,N_11080,N_11128);
nor U11511 (N_11511,N_11077,N_11256);
xor U11512 (N_11512,N_11375,N_11364);
xnor U11513 (N_11513,N_11352,N_11118);
xnor U11514 (N_11514,N_11351,N_11154);
or U11515 (N_11515,N_11000,N_11411);
xnor U11516 (N_11516,N_11368,N_11038);
xnor U11517 (N_11517,N_11201,N_11378);
nand U11518 (N_11518,N_11067,N_11497);
and U11519 (N_11519,N_11468,N_11059);
nand U11520 (N_11520,N_11149,N_11204);
nor U11521 (N_11521,N_11056,N_11480);
or U11522 (N_11522,N_11123,N_11459);
and U11523 (N_11523,N_11147,N_11444);
and U11524 (N_11524,N_11373,N_11258);
or U11525 (N_11525,N_11071,N_11338);
and U11526 (N_11526,N_11407,N_11075);
or U11527 (N_11527,N_11010,N_11166);
nand U11528 (N_11528,N_11453,N_11356);
or U11529 (N_11529,N_11357,N_11168);
nor U11530 (N_11530,N_11105,N_11241);
xor U11531 (N_11531,N_11287,N_11249);
and U11532 (N_11532,N_11322,N_11470);
nor U11533 (N_11533,N_11353,N_11167);
nor U11534 (N_11534,N_11052,N_11033);
nand U11535 (N_11535,N_11019,N_11485);
nor U11536 (N_11536,N_11321,N_11387);
nor U11537 (N_11537,N_11224,N_11349);
nor U11538 (N_11538,N_11163,N_11223);
and U11539 (N_11539,N_11164,N_11126);
nor U11540 (N_11540,N_11145,N_11236);
nor U11541 (N_11541,N_11127,N_11451);
xor U11542 (N_11542,N_11324,N_11394);
nand U11543 (N_11543,N_11002,N_11441);
nand U11544 (N_11544,N_11331,N_11187);
nor U11545 (N_11545,N_11202,N_11252);
or U11546 (N_11546,N_11427,N_11291);
nor U11547 (N_11547,N_11469,N_11104);
xor U11548 (N_11548,N_11173,N_11443);
xor U11549 (N_11549,N_11035,N_11440);
nor U11550 (N_11550,N_11212,N_11216);
nand U11551 (N_11551,N_11304,N_11445);
nor U11552 (N_11552,N_11228,N_11395);
and U11553 (N_11553,N_11015,N_11141);
and U11554 (N_11554,N_11060,N_11276);
and U11555 (N_11555,N_11405,N_11272);
nand U11556 (N_11556,N_11121,N_11205);
nor U11557 (N_11557,N_11450,N_11243);
or U11558 (N_11558,N_11169,N_11380);
and U11559 (N_11559,N_11054,N_11420);
and U11560 (N_11560,N_11152,N_11458);
nor U11561 (N_11561,N_11006,N_11442);
and U11562 (N_11562,N_11242,N_11234);
nand U11563 (N_11563,N_11131,N_11089);
nor U11564 (N_11564,N_11221,N_11136);
or U11565 (N_11565,N_11174,N_11436);
nor U11566 (N_11566,N_11397,N_11225);
and U11567 (N_11567,N_11007,N_11044);
nand U11568 (N_11568,N_11172,N_11425);
nor U11569 (N_11569,N_11008,N_11078);
nor U11570 (N_11570,N_11328,N_11031);
nand U11571 (N_11571,N_11301,N_11426);
or U11572 (N_11572,N_11327,N_11367);
and U11573 (N_11573,N_11274,N_11063);
nor U11574 (N_11574,N_11218,N_11004);
or U11575 (N_11575,N_11277,N_11160);
nor U11576 (N_11576,N_11460,N_11198);
nor U11577 (N_11577,N_11239,N_11210);
xor U11578 (N_11578,N_11058,N_11398);
nand U11579 (N_11579,N_11133,N_11354);
or U11580 (N_11580,N_11259,N_11325);
and U11581 (N_11581,N_11208,N_11487);
xnor U11582 (N_11582,N_11064,N_11361);
nand U11583 (N_11583,N_11101,N_11120);
xor U11584 (N_11584,N_11157,N_11314);
or U11585 (N_11585,N_11475,N_11176);
and U11586 (N_11586,N_11413,N_11286);
nand U11587 (N_11587,N_11390,N_11399);
or U11588 (N_11588,N_11417,N_11307);
nand U11589 (N_11589,N_11416,N_11247);
nor U11590 (N_11590,N_11384,N_11358);
or U11591 (N_11591,N_11408,N_11194);
and U11592 (N_11592,N_11043,N_11098);
nand U11593 (N_11593,N_11014,N_11271);
and U11594 (N_11594,N_11448,N_11222);
nand U11595 (N_11595,N_11496,N_11396);
or U11596 (N_11596,N_11207,N_11269);
and U11597 (N_11597,N_11192,N_11340);
nand U11598 (N_11598,N_11464,N_11171);
nand U11599 (N_11599,N_11251,N_11144);
and U11600 (N_11600,N_11250,N_11438);
xnor U11601 (N_11601,N_11435,N_11099);
xor U11602 (N_11602,N_11386,N_11323);
and U11603 (N_11603,N_11045,N_11418);
and U11604 (N_11604,N_11492,N_11090);
or U11605 (N_11605,N_11103,N_11148);
xnor U11606 (N_11606,N_11203,N_11454);
and U11607 (N_11607,N_11153,N_11481);
and U11608 (N_11608,N_11095,N_11263);
nor U11609 (N_11609,N_11074,N_11283);
or U11610 (N_11610,N_11217,N_11486);
and U11611 (N_11611,N_11404,N_11027);
nand U11612 (N_11612,N_11053,N_11490);
nand U11613 (N_11613,N_11318,N_11433);
or U11614 (N_11614,N_11191,N_11230);
nor U11615 (N_11615,N_11483,N_11041);
and U11616 (N_11616,N_11360,N_11343);
and U11617 (N_11617,N_11359,N_11262);
or U11618 (N_11618,N_11461,N_11350);
nand U11619 (N_11619,N_11206,N_11051);
or U11620 (N_11620,N_11190,N_11288);
or U11621 (N_11621,N_11320,N_11345);
xnor U11622 (N_11622,N_11267,N_11185);
nor U11623 (N_11623,N_11299,N_11482);
and U11624 (N_11624,N_11165,N_11312);
nand U11625 (N_11625,N_11430,N_11319);
xnor U11626 (N_11626,N_11290,N_11189);
or U11627 (N_11627,N_11130,N_11294);
and U11628 (N_11628,N_11134,N_11334);
and U11629 (N_11629,N_11363,N_11085);
nor U11630 (N_11630,N_11421,N_11342);
and U11631 (N_11631,N_11178,N_11048);
or U11632 (N_11632,N_11339,N_11248);
xor U11633 (N_11633,N_11215,N_11235);
or U11634 (N_11634,N_11061,N_11009);
nand U11635 (N_11635,N_11220,N_11452);
or U11636 (N_11636,N_11385,N_11158);
and U11637 (N_11637,N_11428,N_11050);
nor U11638 (N_11638,N_11335,N_11110);
nor U11639 (N_11639,N_11083,N_11293);
xnor U11640 (N_11640,N_11406,N_11034);
xor U11641 (N_11641,N_11072,N_11232);
nand U11642 (N_11642,N_11474,N_11280);
xnor U11643 (N_11643,N_11382,N_11477);
or U11644 (N_11644,N_11200,N_11374);
and U11645 (N_11645,N_11295,N_11484);
and U11646 (N_11646,N_11111,N_11400);
nor U11647 (N_11647,N_11316,N_11037);
nand U11648 (N_11648,N_11457,N_11296);
or U11649 (N_11649,N_11186,N_11467);
nor U11650 (N_11650,N_11070,N_11137);
or U11651 (N_11651,N_11237,N_11161);
nor U11652 (N_11652,N_11300,N_11117);
and U11653 (N_11653,N_11278,N_11389);
nor U11654 (N_11654,N_11046,N_11254);
or U11655 (N_11655,N_11371,N_11183);
nor U11656 (N_11656,N_11022,N_11303);
and U11657 (N_11657,N_11087,N_11313);
nand U11658 (N_11658,N_11138,N_11143);
xnor U11659 (N_11659,N_11003,N_11377);
and U11660 (N_11660,N_11119,N_11036);
xnor U11661 (N_11661,N_11253,N_11370);
and U11662 (N_11662,N_11102,N_11011);
nand U11663 (N_11663,N_11344,N_11476);
nor U11664 (N_11664,N_11336,N_11238);
xnor U11665 (N_11665,N_11092,N_11446);
or U11666 (N_11666,N_11348,N_11069);
nor U11667 (N_11667,N_11379,N_11181);
and U11668 (N_11668,N_11260,N_11195);
and U11669 (N_11669,N_11155,N_11424);
and U11670 (N_11670,N_11240,N_11284);
xor U11671 (N_11671,N_11499,N_11179);
and U11672 (N_11672,N_11310,N_11062);
and U11673 (N_11673,N_11175,N_11432);
nor U11674 (N_11674,N_11100,N_11403);
nor U11675 (N_11675,N_11018,N_11135);
nand U11676 (N_11676,N_11422,N_11226);
nand U11677 (N_11677,N_11268,N_11026);
and U11678 (N_11678,N_11199,N_11473);
xor U11679 (N_11679,N_11392,N_11094);
nand U11680 (N_11680,N_11495,N_11193);
nand U11681 (N_11681,N_11297,N_11292);
and U11682 (N_11682,N_11023,N_11016);
nand U11683 (N_11683,N_11463,N_11017);
or U11684 (N_11684,N_11419,N_11214);
and U11685 (N_11685,N_11455,N_11456);
nand U11686 (N_11686,N_11381,N_11329);
nand U11687 (N_11687,N_11055,N_11229);
xor U11688 (N_11688,N_11182,N_11088);
nand U11689 (N_11689,N_11097,N_11423);
nor U11690 (N_11690,N_11479,N_11219);
xnor U11691 (N_11691,N_11466,N_11330);
and U11692 (N_11692,N_11106,N_11115);
nor U11693 (N_11693,N_11346,N_11401);
or U11694 (N_11694,N_11391,N_11040);
nand U11695 (N_11695,N_11279,N_11383);
nor U11696 (N_11696,N_11122,N_11255);
xor U11697 (N_11697,N_11305,N_11073);
nor U11698 (N_11698,N_11049,N_11326);
xor U11699 (N_11699,N_11197,N_11369);
nor U11700 (N_11700,N_11347,N_11030);
and U11701 (N_11701,N_11245,N_11415);
nor U11702 (N_11702,N_11431,N_11315);
nor U11703 (N_11703,N_11159,N_11465);
nand U11704 (N_11704,N_11489,N_11414);
xor U11705 (N_11705,N_11112,N_11076);
xor U11706 (N_11706,N_11333,N_11093);
xor U11707 (N_11707,N_11244,N_11084);
and U11708 (N_11708,N_11341,N_11209);
xor U11709 (N_11709,N_11498,N_11177);
nor U11710 (N_11710,N_11410,N_11107);
nor U11711 (N_11711,N_11151,N_11355);
xnor U11712 (N_11712,N_11025,N_11488);
xnor U11713 (N_11713,N_11086,N_11317);
nand U11714 (N_11714,N_11012,N_11028);
and U11715 (N_11715,N_11082,N_11289);
or U11716 (N_11716,N_11309,N_11047);
nand U11717 (N_11717,N_11362,N_11013);
and U11718 (N_11718,N_11462,N_11332);
xor U11719 (N_11719,N_11139,N_11264);
nor U11720 (N_11720,N_11196,N_11302);
xnor U11721 (N_11721,N_11162,N_11447);
xnor U11722 (N_11722,N_11032,N_11366);
xnor U11723 (N_11723,N_11132,N_11472);
or U11724 (N_11724,N_11372,N_11184);
nor U11725 (N_11725,N_11146,N_11337);
nand U11726 (N_11726,N_11231,N_11113);
nor U11727 (N_11727,N_11150,N_11109);
or U11728 (N_11728,N_11211,N_11265);
nor U11729 (N_11729,N_11478,N_11091);
or U11730 (N_11730,N_11491,N_11068);
and U11731 (N_11731,N_11129,N_11020);
and U11732 (N_11732,N_11081,N_11188);
nand U11733 (N_11733,N_11213,N_11376);
nor U11734 (N_11734,N_11281,N_11266);
nand U11735 (N_11735,N_11257,N_11039);
nor U11736 (N_11736,N_11066,N_11114);
and U11737 (N_11737,N_11449,N_11311);
nand U11738 (N_11738,N_11156,N_11180);
nand U11739 (N_11739,N_11365,N_11388);
or U11740 (N_11740,N_11125,N_11029);
xnor U11741 (N_11741,N_11227,N_11493);
nand U11742 (N_11742,N_11079,N_11308);
xor U11743 (N_11743,N_11285,N_11402);
nand U11744 (N_11744,N_11282,N_11116);
nor U11745 (N_11745,N_11124,N_11108);
nand U11746 (N_11746,N_11275,N_11096);
or U11747 (N_11747,N_11001,N_11246);
nor U11748 (N_11748,N_11021,N_11005);
xnor U11749 (N_11749,N_11471,N_11393);
nand U11750 (N_11750,N_11130,N_11176);
or U11751 (N_11751,N_11498,N_11128);
nor U11752 (N_11752,N_11405,N_11104);
or U11753 (N_11753,N_11400,N_11486);
xor U11754 (N_11754,N_11419,N_11291);
and U11755 (N_11755,N_11481,N_11340);
or U11756 (N_11756,N_11291,N_11261);
or U11757 (N_11757,N_11408,N_11222);
or U11758 (N_11758,N_11468,N_11390);
nand U11759 (N_11759,N_11454,N_11032);
nor U11760 (N_11760,N_11058,N_11242);
and U11761 (N_11761,N_11129,N_11077);
nor U11762 (N_11762,N_11105,N_11301);
xnor U11763 (N_11763,N_11457,N_11033);
or U11764 (N_11764,N_11478,N_11020);
nor U11765 (N_11765,N_11141,N_11494);
or U11766 (N_11766,N_11197,N_11463);
nand U11767 (N_11767,N_11225,N_11075);
nand U11768 (N_11768,N_11019,N_11436);
xnor U11769 (N_11769,N_11297,N_11396);
xnor U11770 (N_11770,N_11340,N_11071);
or U11771 (N_11771,N_11483,N_11110);
nor U11772 (N_11772,N_11141,N_11295);
nor U11773 (N_11773,N_11154,N_11078);
or U11774 (N_11774,N_11468,N_11241);
and U11775 (N_11775,N_11259,N_11092);
xnor U11776 (N_11776,N_11461,N_11378);
xnor U11777 (N_11777,N_11174,N_11210);
xnor U11778 (N_11778,N_11422,N_11362);
nand U11779 (N_11779,N_11162,N_11218);
and U11780 (N_11780,N_11149,N_11099);
or U11781 (N_11781,N_11474,N_11471);
xor U11782 (N_11782,N_11190,N_11053);
xnor U11783 (N_11783,N_11205,N_11298);
nand U11784 (N_11784,N_11061,N_11470);
xnor U11785 (N_11785,N_11378,N_11476);
nor U11786 (N_11786,N_11088,N_11370);
and U11787 (N_11787,N_11377,N_11233);
nand U11788 (N_11788,N_11323,N_11312);
xor U11789 (N_11789,N_11194,N_11243);
nand U11790 (N_11790,N_11499,N_11212);
nor U11791 (N_11791,N_11160,N_11450);
nand U11792 (N_11792,N_11232,N_11209);
nand U11793 (N_11793,N_11030,N_11437);
xor U11794 (N_11794,N_11337,N_11205);
xnor U11795 (N_11795,N_11239,N_11313);
xnor U11796 (N_11796,N_11494,N_11183);
nand U11797 (N_11797,N_11413,N_11376);
nor U11798 (N_11798,N_11069,N_11090);
nand U11799 (N_11799,N_11352,N_11190);
nand U11800 (N_11800,N_11142,N_11300);
nand U11801 (N_11801,N_11193,N_11061);
nand U11802 (N_11802,N_11084,N_11398);
xor U11803 (N_11803,N_11042,N_11139);
nor U11804 (N_11804,N_11156,N_11137);
nand U11805 (N_11805,N_11383,N_11369);
xnor U11806 (N_11806,N_11436,N_11297);
or U11807 (N_11807,N_11102,N_11311);
xnor U11808 (N_11808,N_11130,N_11137);
or U11809 (N_11809,N_11458,N_11466);
nand U11810 (N_11810,N_11417,N_11042);
or U11811 (N_11811,N_11332,N_11148);
nand U11812 (N_11812,N_11127,N_11295);
nand U11813 (N_11813,N_11357,N_11493);
nand U11814 (N_11814,N_11134,N_11243);
or U11815 (N_11815,N_11005,N_11013);
or U11816 (N_11816,N_11248,N_11046);
or U11817 (N_11817,N_11338,N_11394);
nor U11818 (N_11818,N_11381,N_11048);
nand U11819 (N_11819,N_11069,N_11242);
nor U11820 (N_11820,N_11123,N_11103);
and U11821 (N_11821,N_11068,N_11038);
nor U11822 (N_11822,N_11352,N_11380);
xnor U11823 (N_11823,N_11076,N_11003);
or U11824 (N_11824,N_11167,N_11497);
nand U11825 (N_11825,N_11032,N_11463);
and U11826 (N_11826,N_11300,N_11057);
or U11827 (N_11827,N_11246,N_11166);
nor U11828 (N_11828,N_11219,N_11437);
and U11829 (N_11829,N_11153,N_11120);
and U11830 (N_11830,N_11422,N_11258);
nand U11831 (N_11831,N_11067,N_11313);
and U11832 (N_11832,N_11383,N_11333);
xor U11833 (N_11833,N_11408,N_11377);
xor U11834 (N_11834,N_11442,N_11221);
nand U11835 (N_11835,N_11359,N_11153);
and U11836 (N_11836,N_11214,N_11171);
nand U11837 (N_11837,N_11109,N_11199);
nor U11838 (N_11838,N_11298,N_11437);
nand U11839 (N_11839,N_11383,N_11001);
nand U11840 (N_11840,N_11065,N_11300);
or U11841 (N_11841,N_11001,N_11004);
nor U11842 (N_11842,N_11019,N_11468);
nand U11843 (N_11843,N_11289,N_11226);
nor U11844 (N_11844,N_11343,N_11051);
nor U11845 (N_11845,N_11281,N_11484);
nand U11846 (N_11846,N_11368,N_11331);
xor U11847 (N_11847,N_11183,N_11412);
xnor U11848 (N_11848,N_11196,N_11296);
nand U11849 (N_11849,N_11339,N_11167);
or U11850 (N_11850,N_11287,N_11179);
xnor U11851 (N_11851,N_11131,N_11150);
nand U11852 (N_11852,N_11225,N_11044);
nor U11853 (N_11853,N_11485,N_11401);
nor U11854 (N_11854,N_11050,N_11356);
nand U11855 (N_11855,N_11406,N_11015);
xor U11856 (N_11856,N_11003,N_11439);
xnor U11857 (N_11857,N_11254,N_11252);
nor U11858 (N_11858,N_11082,N_11094);
xnor U11859 (N_11859,N_11459,N_11471);
and U11860 (N_11860,N_11126,N_11385);
xor U11861 (N_11861,N_11250,N_11189);
nor U11862 (N_11862,N_11209,N_11044);
or U11863 (N_11863,N_11150,N_11172);
nor U11864 (N_11864,N_11021,N_11271);
nand U11865 (N_11865,N_11143,N_11090);
or U11866 (N_11866,N_11476,N_11238);
nor U11867 (N_11867,N_11355,N_11197);
nor U11868 (N_11868,N_11308,N_11061);
and U11869 (N_11869,N_11296,N_11382);
xor U11870 (N_11870,N_11100,N_11039);
nor U11871 (N_11871,N_11178,N_11298);
nand U11872 (N_11872,N_11419,N_11347);
or U11873 (N_11873,N_11223,N_11482);
and U11874 (N_11874,N_11462,N_11001);
or U11875 (N_11875,N_11471,N_11173);
nor U11876 (N_11876,N_11312,N_11129);
or U11877 (N_11877,N_11478,N_11075);
nand U11878 (N_11878,N_11499,N_11477);
nand U11879 (N_11879,N_11387,N_11028);
xor U11880 (N_11880,N_11306,N_11322);
xor U11881 (N_11881,N_11392,N_11104);
xnor U11882 (N_11882,N_11044,N_11058);
or U11883 (N_11883,N_11499,N_11199);
and U11884 (N_11884,N_11288,N_11312);
nand U11885 (N_11885,N_11351,N_11374);
nand U11886 (N_11886,N_11437,N_11289);
or U11887 (N_11887,N_11317,N_11366);
and U11888 (N_11888,N_11259,N_11357);
and U11889 (N_11889,N_11134,N_11415);
xor U11890 (N_11890,N_11335,N_11413);
or U11891 (N_11891,N_11256,N_11132);
nand U11892 (N_11892,N_11170,N_11276);
xnor U11893 (N_11893,N_11261,N_11435);
nor U11894 (N_11894,N_11208,N_11243);
nand U11895 (N_11895,N_11210,N_11267);
or U11896 (N_11896,N_11333,N_11415);
or U11897 (N_11897,N_11139,N_11324);
nor U11898 (N_11898,N_11234,N_11495);
nor U11899 (N_11899,N_11111,N_11232);
or U11900 (N_11900,N_11474,N_11224);
nand U11901 (N_11901,N_11175,N_11168);
xor U11902 (N_11902,N_11100,N_11064);
xnor U11903 (N_11903,N_11165,N_11055);
or U11904 (N_11904,N_11386,N_11061);
or U11905 (N_11905,N_11297,N_11184);
nor U11906 (N_11906,N_11302,N_11448);
or U11907 (N_11907,N_11283,N_11362);
nand U11908 (N_11908,N_11498,N_11071);
or U11909 (N_11909,N_11321,N_11246);
xor U11910 (N_11910,N_11224,N_11172);
xnor U11911 (N_11911,N_11040,N_11133);
and U11912 (N_11912,N_11341,N_11354);
xnor U11913 (N_11913,N_11166,N_11474);
and U11914 (N_11914,N_11261,N_11133);
and U11915 (N_11915,N_11301,N_11249);
and U11916 (N_11916,N_11461,N_11053);
or U11917 (N_11917,N_11317,N_11396);
nor U11918 (N_11918,N_11151,N_11270);
xor U11919 (N_11919,N_11495,N_11435);
nor U11920 (N_11920,N_11433,N_11490);
xor U11921 (N_11921,N_11490,N_11155);
nor U11922 (N_11922,N_11230,N_11008);
xor U11923 (N_11923,N_11032,N_11355);
or U11924 (N_11924,N_11026,N_11078);
nor U11925 (N_11925,N_11260,N_11230);
and U11926 (N_11926,N_11035,N_11453);
xnor U11927 (N_11927,N_11021,N_11350);
nor U11928 (N_11928,N_11020,N_11150);
nand U11929 (N_11929,N_11171,N_11048);
or U11930 (N_11930,N_11477,N_11474);
xnor U11931 (N_11931,N_11498,N_11083);
nand U11932 (N_11932,N_11160,N_11155);
nand U11933 (N_11933,N_11035,N_11322);
xnor U11934 (N_11934,N_11461,N_11259);
xnor U11935 (N_11935,N_11157,N_11280);
nand U11936 (N_11936,N_11030,N_11455);
nand U11937 (N_11937,N_11307,N_11126);
or U11938 (N_11938,N_11205,N_11250);
nor U11939 (N_11939,N_11100,N_11466);
nor U11940 (N_11940,N_11218,N_11013);
xor U11941 (N_11941,N_11026,N_11388);
xnor U11942 (N_11942,N_11249,N_11116);
and U11943 (N_11943,N_11046,N_11403);
or U11944 (N_11944,N_11053,N_11079);
and U11945 (N_11945,N_11050,N_11396);
and U11946 (N_11946,N_11191,N_11273);
or U11947 (N_11947,N_11399,N_11261);
nor U11948 (N_11948,N_11479,N_11220);
and U11949 (N_11949,N_11331,N_11220);
and U11950 (N_11950,N_11191,N_11437);
or U11951 (N_11951,N_11390,N_11289);
and U11952 (N_11952,N_11235,N_11061);
or U11953 (N_11953,N_11032,N_11173);
xnor U11954 (N_11954,N_11399,N_11180);
and U11955 (N_11955,N_11105,N_11223);
xnor U11956 (N_11956,N_11121,N_11033);
xnor U11957 (N_11957,N_11076,N_11156);
nor U11958 (N_11958,N_11361,N_11440);
nand U11959 (N_11959,N_11495,N_11052);
nor U11960 (N_11960,N_11319,N_11162);
nor U11961 (N_11961,N_11328,N_11376);
and U11962 (N_11962,N_11044,N_11078);
xor U11963 (N_11963,N_11253,N_11015);
xor U11964 (N_11964,N_11454,N_11455);
nor U11965 (N_11965,N_11228,N_11256);
and U11966 (N_11966,N_11080,N_11380);
or U11967 (N_11967,N_11062,N_11055);
nor U11968 (N_11968,N_11496,N_11459);
nand U11969 (N_11969,N_11272,N_11307);
xor U11970 (N_11970,N_11359,N_11322);
and U11971 (N_11971,N_11475,N_11296);
nor U11972 (N_11972,N_11407,N_11256);
nand U11973 (N_11973,N_11036,N_11333);
nor U11974 (N_11974,N_11263,N_11031);
or U11975 (N_11975,N_11393,N_11083);
nand U11976 (N_11976,N_11260,N_11220);
nor U11977 (N_11977,N_11360,N_11082);
xnor U11978 (N_11978,N_11423,N_11438);
or U11979 (N_11979,N_11045,N_11129);
xnor U11980 (N_11980,N_11091,N_11419);
xnor U11981 (N_11981,N_11430,N_11485);
and U11982 (N_11982,N_11429,N_11390);
or U11983 (N_11983,N_11236,N_11062);
xor U11984 (N_11984,N_11135,N_11298);
xnor U11985 (N_11985,N_11063,N_11291);
nor U11986 (N_11986,N_11422,N_11010);
nor U11987 (N_11987,N_11344,N_11025);
or U11988 (N_11988,N_11067,N_11217);
nand U11989 (N_11989,N_11083,N_11046);
or U11990 (N_11990,N_11290,N_11214);
xnor U11991 (N_11991,N_11235,N_11353);
xor U11992 (N_11992,N_11218,N_11487);
xnor U11993 (N_11993,N_11306,N_11202);
nand U11994 (N_11994,N_11414,N_11003);
and U11995 (N_11995,N_11445,N_11481);
nand U11996 (N_11996,N_11294,N_11260);
nor U11997 (N_11997,N_11474,N_11232);
nand U11998 (N_11998,N_11448,N_11451);
xor U11999 (N_11999,N_11160,N_11283);
nand U12000 (N_12000,N_11797,N_11624);
xor U12001 (N_12001,N_11800,N_11718);
nor U12002 (N_12002,N_11739,N_11985);
xnor U12003 (N_12003,N_11514,N_11935);
or U12004 (N_12004,N_11768,N_11654);
xor U12005 (N_12005,N_11970,N_11890);
nor U12006 (N_12006,N_11943,N_11773);
nor U12007 (N_12007,N_11877,N_11703);
nor U12008 (N_12008,N_11631,N_11893);
nor U12009 (N_12009,N_11861,N_11957);
nor U12010 (N_12010,N_11956,N_11963);
and U12011 (N_12011,N_11540,N_11645);
xor U12012 (N_12012,N_11700,N_11854);
nor U12013 (N_12013,N_11536,N_11999);
or U12014 (N_12014,N_11790,N_11586);
nand U12015 (N_12015,N_11682,N_11510);
nand U12016 (N_12016,N_11879,N_11575);
nor U12017 (N_12017,N_11753,N_11539);
xor U12018 (N_12018,N_11949,N_11961);
nor U12019 (N_12019,N_11728,N_11736);
nor U12020 (N_12020,N_11573,N_11746);
or U12021 (N_12021,N_11564,N_11931);
xnor U12022 (N_12022,N_11853,N_11844);
xnor U12023 (N_12023,N_11978,N_11636);
and U12024 (N_12024,N_11627,N_11785);
nand U12025 (N_12025,N_11997,N_11603);
nand U12026 (N_12026,N_11602,N_11686);
or U12027 (N_12027,N_11798,N_11755);
and U12028 (N_12028,N_11674,N_11707);
nor U12029 (N_12029,N_11621,N_11581);
or U12030 (N_12030,N_11634,N_11520);
xnor U12031 (N_12031,N_11538,N_11714);
and U12032 (N_12032,N_11860,N_11874);
and U12033 (N_12033,N_11817,N_11811);
nand U12034 (N_12034,N_11954,N_11926);
nand U12035 (N_12035,N_11919,N_11598);
nand U12036 (N_12036,N_11522,N_11834);
xnor U12037 (N_12037,N_11973,N_11620);
xor U12038 (N_12038,N_11565,N_11551);
nor U12039 (N_12039,N_11894,N_11613);
nand U12040 (N_12040,N_11868,N_11675);
nor U12041 (N_12041,N_11870,N_11717);
xor U12042 (N_12042,N_11698,N_11875);
and U12043 (N_12043,N_11866,N_11579);
xnor U12044 (N_12044,N_11976,N_11824);
and U12045 (N_12045,N_11867,N_11666);
xor U12046 (N_12046,N_11974,N_11643);
nor U12047 (N_12047,N_11914,N_11678);
xor U12048 (N_12048,N_11757,N_11938);
nor U12049 (N_12049,N_11726,N_11769);
xnor U12050 (N_12050,N_11826,N_11955);
nand U12051 (N_12051,N_11566,N_11715);
xor U12052 (N_12052,N_11735,N_11906);
xnor U12053 (N_12053,N_11713,N_11933);
nor U12054 (N_12054,N_11719,N_11502);
nor U12055 (N_12055,N_11544,N_11802);
and U12056 (N_12056,N_11990,N_11632);
and U12057 (N_12057,N_11756,N_11888);
nand U12058 (N_12058,N_11571,N_11737);
xnor U12059 (N_12059,N_11917,N_11887);
nor U12060 (N_12060,N_11821,N_11841);
xnor U12061 (N_12061,N_11695,N_11529);
or U12062 (N_12062,N_11863,N_11692);
or U12063 (N_12063,N_11837,N_11830);
xor U12064 (N_12064,N_11671,N_11886);
and U12065 (N_12065,N_11904,N_11584);
xor U12066 (N_12066,N_11663,N_11851);
and U12067 (N_12067,N_11848,N_11641);
and U12068 (N_12068,N_11688,N_11595);
nor U12069 (N_12069,N_11767,N_11977);
and U12070 (N_12070,N_11913,N_11947);
nand U12071 (N_12071,N_11774,N_11610);
xnor U12072 (N_12072,N_11659,N_11808);
nand U12073 (N_12073,N_11562,N_11941);
and U12074 (N_12074,N_11796,N_11582);
nor U12075 (N_12075,N_11795,N_11531);
xor U12076 (N_12076,N_11521,N_11537);
and U12077 (N_12077,N_11648,N_11911);
and U12078 (N_12078,N_11989,N_11747);
or U12079 (N_12079,N_11646,N_11852);
xor U12080 (N_12080,N_11743,N_11619);
xnor U12081 (N_12081,N_11618,N_11638);
nor U12082 (N_12082,N_11840,N_11683);
nand U12083 (N_12083,N_11762,N_11801);
and U12084 (N_12084,N_11778,N_11662);
xnor U12085 (N_12085,N_11548,N_11865);
nor U12086 (N_12086,N_11609,N_11936);
and U12087 (N_12087,N_11561,N_11816);
nand U12088 (N_12088,N_11898,N_11550);
and U12089 (N_12089,N_11667,N_11912);
and U12090 (N_12090,N_11950,N_11975);
or U12091 (N_12091,N_11818,N_11614);
and U12092 (N_12092,N_11526,N_11585);
and U12093 (N_12093,N_11501,N_11819);
and U12094 (N_12094,N_11729,N_11677);
or U12095 (N_12095,N_11690,N_11570);
or U12096 (N_12096,N_11708,N_11994);
nor U12097 (N_12097,N_11918,N_11611);
or U12098 (N_12098,N_11932,N_11846);
nor U12099 (N_12099,N_11823,N_11964);
or U12100 (N_12100,N_11925,N_11805);
and U12101 (N_12101,N_11828,N_11696);
nor U12102 (N_12102,N_11872,N_11992);
or U12103 (N_12103,N_11635,N_11549);
and U12104 (N_12104,N_11567,N_11916);
xnor U12105 (N_12105,N_11810,N_11530);
nor U12106 (N_12106,N_11754,N_11612);
or U12107 (N_12107,N_11554,N_11535);
nor U12108 (N_12108,N_11850,N_11901);
nor U12109 (N_12109,N_11759,N_11891);
or U12110 (N_12110,N_11655,N_11766);
xnor U12111 (N_12111,N_11574,N_11789);
xor U12112 (N_12112,N_11922,N_11684);
and U12113 (N_12113,N_11968,N_11959);
nor U12114 (N_12114,N_11711,N_11722);
and U12115 (N_12115,N_11515,N_11542);
and U12116 (N_12116,N_11902,N_11780);
or U12117 (N_12117,N_11556,N_11944);
or U12118 (N_12118,N_11709,N_11680);
nor U12119 (N_12119,N_11969,N_11665);
and U12120 (N_12120,N_11857,N_11706);
and U12121 (N_12121,N_11608,N_11721);
nor U12122 (N_12122,N_11731,N_11650);
nor U12123 (N_12123,N_11984,N_11734);
xnor U12124 (N_12124,N_11929,N_11583);
and U12125 (N_12125,N_11988,N_11664);
and U12126 (N_12126,N_11628,N_11604);
nor U12127 (N_12127,N_11601,N_11606);
and U12128 (N_12128,N_11849,N_11945);
and U12129 (N_12129,N_11694,N_11658);
and U12130 (N_12130,N_11783,N_11506);
nor U12131 (N_12131,N_11572,N_11878);
or U12132 (N_12132,N_11900,N_11587);
or U12133 (N_12133,N_11839,N_11884);
and U12134 (N_12134,N_11831,N_11668);
or U12135 (N_12135,N_11750,N_11749);
or U12136 (N_12136,N_11928,N_11647);
or U12137 (N_12137,N_11644,N_11740);
or U12138 (N_12138,N_11927,N_11725);
nand U12139 (N_12139,N_11651,N_11770);
nand U12140 (N_12140,N_11507,N_11794);
and U12141 (N_12141,N_11519,N_11503);
nor U12142 (N_12142,N_11909,N_11812);
and U12143 (N_12143,N_11880,N_11742);
nand U12144 (N_12144,N_11952,N_11560);
xnor U12145 (N_12145,N_11776,N_11862);
xor U12146 (N_12146,N_11751,N_11896);
and U12147 (N_12147,N_11764,N_11630);
nor U12148 (N_12148,N_11784,N_11642);
nor U12149 (N_12149,N_11799,N_11772);
or U12150 (N_12150,N_11845,N_11907);
xor U12151 (N_12151,N_11622,N_11516);
or U12152 (N_12152,N_11676,N_11793);
xnor U12153 (N_12153,N_11633,N_11553);
xnor U12154 (N_12154,N_11607,N_11993);
and U12155 (N_12155,N_11962,N_11822);
nor U12156 (N_12156,N_11543,N_11730);
xnor U12157 (N_12157,N_11983,N_11557);
xnor U12158 (N_12158,N_11827,N_11847);
and U12159 (N_12159,N_11649,N_11656);
nand U12160 (N_12160,N_11967,N_11527);
nand U12161 (N_12161,N_11741,N_11835);
nor U12162 (N_12162,N_11771,N_11889);
xnor U12163 (N_12163,N_11637,N_11563);
nand U12164 (N_12164,N_11777,N_11517);
or U12165 (N_12165,N_11547,N_11981);
and U12166 (N_12166,N_11758,N_11541);
xnor U12167 (N_12167,N_11524,N_11982);
nand U12168 (N_12168,N_11873,N_11825);
xnor U12169 (N_12169,N_11836,N_11804);
and U12170 (N_12170,N_11661,N_11672);
xnor U12171 (N_12171,N_11937,N_11761);
xnor U12172 (N_12172,N_11689,N_11939);
or U12173 (N_12173,N_11704,N_11552);
nor U12174 (N_12174,N_11966,N_11787);
and U12175 (N_12175,N_11528,N_11670);
nand U12176 (N_12176,N_11987,N_11723);
xor U12177 (N_12177,N_11523,N_11518);
or U12178 (N_12178,N_11720,N_11921);
nand U12179 (N_12179,N_11568,N_11685);
nand U12180 (N_12180,N_11669,N_11998);
xor U12181 (N_12181,N_11511,N_11681);
and U12182 (N_12182,N_11699,N_11915);
and U12183 (N_12183,N_11576,N_11905);
nand U12184 (N_12184,N_11829,N_11596);
xor U12185 (N_12185,N_11500,N_11732);
or U12186 (N_12186,N_11859,N_11979);
nand U12187 (N_12187,N_11814,N_11843);
and U12188 (N_12188,N_11727,N_11615);
or U12189 (N_12189,N_11972,N_11505);
nand U12190 (N_12190,N_11809,N_11640);
and U12191 (N_12191,N_11748,N_11705);
and U12192 (N_12192,N_11791,N_11593);
or U12193 (N_12193,N_11765,N_11555);
and U12194 (N_12194,N_11869,N_11948);
and U12195 (N_12195,N_11986,N_11693);
or U12196 (N_12196,N_11760,N_11991);
or U12197 (N_12197,N_11590,N_11558);
or U12198 (N_12198,N_11617,N_11792);
nand U12199 (N_12199,N_11920,N_11953);
or U12200 (N_12200,N_11856,N_11600);
or U12201 (N_12201,N_11813,N_11626);
nand U12202 (N_12202,N_11803,N_11958);
or U12203 (N_12203,N_11545,N_11965);
and U12204 (N_12204,N_11580,N_11702);
xor U12205 (N_12205,N_11577,N_11892);
nand U12206 (N_12206,N_11710,N_11591);
nand U12207 (N_12207,N_11930,N_11940);
nor U12208 (N_12208,N_11942,N_11908);
xor U12209 (N_12209,N_11652,N_11687);
and U12210 (N_12210,N_11995,N_11883);
xor U12211 (N_12211,N_11924,N_11980);
xnor U12212 (N_12212,N_11820,N_11605);
xnor U12213 (N_12213,N_11807,N_11569);
nand U12214 (N_12214,N_11513,N_11532);
and U12215 (N_12215,N_11960,N_11781);
nand U12216 (N_12216,N_11871,N_11855);
and U12217 (N_12217,N_11504,N_11733);
xnor U12218 (N_12218,N_11910,N_11763);
nand U12219 (N_12219,N_11625,N_11779);
xor U12220 (N_12220,N_11578,N_11934);
and U12221 (N_12221,N_11923,N_11903);
and U12222 (N_12222,N_11876,N_11508);
nand U12223 (N_12223,N_11895,N_11653);
xnor U12224 (N_12224,N_11864,N_11786);
nor U12225 (N_12225,N_11639,N_11782);
or U12226 (N_12226,N_11691,N_11716);
or U12227 (N_12227,N_11971,N_11673);
nor U12228 (N_12228,N_11697,N_11897);
nand U12229 (N_12229,N_11775,N_11599);
xor U12230 (N_12230,N_11712,N_11946);
or U12231 (N_12231,N_11592,N_11996);
or U12232 (N_12232,N_11546,N_11752);
nor U12233 (N_12233,N_11512,N_11588);
and U12234 (N_12234,N_11744,N_11594);
and U12235 (N_12235,N_11660,N_11838);
nand U12236 (N_12236,N_11701,N_11815);
or U12237 (N_12237,N_11899,N_11881);
xor U12238 (N_12238,N_11616,N_11629);
xnor U12239 (N_12239,N_11738,N_11788);
nand U12240 (N_12240,N_11623,N_11534);
and U12241 (N_12241,N_11533,N_11525);
or U12242 (N_12242,N_11882,N_11559);
or U12243 (N_12243,N_11833,N_11509);
nand U12244 (N_12244,N_11745,N_11657);
xnor U12245 (N_12245,N_11589,N_11806);
and U12246 (N_12246,N_11842,N_11597);
nand U12247 (N_12247,N_11885,N_11724);
nor U12248 (N_12248,N_11858,N_11679);
xor U12249 (N_12249,N_11951,N_11832);
or U12250 (N_12250,N_11792,N_11648);
xor U12251 (N_12251,N_11874,N_11510);
xnor U12252 (N_12252,N_11722,N_11778);
nor U12253 (N_12253,N_11758,N_11564);
xor U12254 (N_12254,N_11752,N_11600);
nor U12255 (N_12255,N_11600,N_11886);
and U12256 (N_12256,N_11907,N_11533);
or U12257 (N_12257,N_11553,N_11649);
xnor U12258 (N_12258,N_11748,N_11679);
and U12259 (N_12259,N_11770,N_11686);
or U12260 (N_12260,N_11538,N_11645);
or U12261 (N_12261,N_11571,N_11835);
and U12262 (N_12262,N_11688,N_11698);
or U12263 (N_12263,N_11720,N_11933);
or U12264 (N_12264,N_11612,N_11756);
and U12265 (N_12265,N_11757,N_11621);
nand U12266 (N_12266,N_11936,N_11754);
nand U12267 (N_12267,N_11766,N_11661);
or U12268 (N_12268,N_11619,N_11645);
nand U12269 (N_12269,N_11506,N_11533);
or U12270 (N_12270,N_11934,N_11738);
xor U12271 (N_12271,N_11670,N_11759);
xnor U12272 (N_12272,N_11524,N_11525);
nand U12273 (N_12273,N_11771,N_11618);
xor U12274 (N_12274,N_11970,N_11520);
nand U12275 (N_12275,N_11674,N_11961);
nand U12276 (N_12276,N_11733,N_11550);
nand U12277 (N_12277,N_11581,N_11606);
nand U12278 (N_12278,N_11595,N_11538);
xnor U12279 (N_12279,N_11924,N_11796);
nand U12280 (N_12280,N_11503,N_11990);
xnor U12281 (N_12281,N_11969,N_11978);
and U12282 (N_12282,N_11623,N_11973);
or U12283 (N_12283,N_11537,N_11737);
xor U12284 (N_12284,N_11634,N_11794);
or U12285 (N_12285,N_11824,N_11679);
and U12286 (N_12286,N_11639,N_11622);
or U12287 (N_12287,N_11666,N_11659);
or U12288 (N_12288,N_11943,N_11720);
nor U12289 (N_12289,N_11519,N_11920);
or U12290 (N_12290,N_11583,N_11533);
or U12291 (N_12291,N_11585,N_11904);
nand U12292 (N_12292,N_11701,N_11515);
nor U12293 (N_12293,N_11825,N_11844);
xnor U12294 (N_12294,N_11926,N_11918);
or U12295 (N_12295,N_11894,N_11827);
or U12296 (N_12296,N_11542,N_11530);
xor U12297 (N_12297,N_11649,N_11742);
nor U12298 (N_12298,N_11750,N_11801);
xor U12299 (N_12299,N_11807,N_11724);
and U12300 (N_12300,N_11908,N_11910);
xor U12301 (N_12301,N_11659,N_11615);
xor U12302 (N_12302,N_11677,N_11848);
and U12303 (N_12303,N_11691,N_11573);
nor U12304 (N_12304,N_11783,N_11558);
and U12305 (N_12305,N_11865,N_11758);
or U12306 (N_12306,N_11851,N_11725);
and U12307 (N_12307,N_11694,N_11602);
nand U12308 (N_12308,N_11661,N_11855);
nor U12309 (N_12309,N_11701,N_11555);
and U12310 (N_12310,N_11835,N_11734);
xor U12311 (N_12311,N_11832,N_11911);
and U12312 (N_12312,N_11605,N_11766);
nand U12313 (N_12313,N_11731,N_11539);
xor U12314 (N_12314,N_11751,N_11712);
nor U12315 (N_12315,N_11891,N_11503);
xnor U12316 (N_12316,N_11605,N_11803);
and U12317 (N_12317,N_11557,N_11688);
nand U12318 (N_12318,N_11859,N_11936);
nor U12319 (N_12319,N_11500,N_11680);
nor U12320 (N_12320,N_11518,N_11920);
and U12321 (N_12321,N_11588,N_11853);
nor U12322 (N_12322,N_11763,N_11631);
or U12323 (N_12323,N_11692,N_11669);
and U12324 (N_12324,N_11770,N_11683);
xnor U12325 (N_12325,N_11554,N_11962);
and U12326 (N_12326,N_11953,N_11734);
xor U12327 (N_12327,N_11869,N_11605);
nor U12328 (N_12328,N_11536,N_11688);
xor U12329 (N_12329,N_11912,N_11620);
xnor U12330 (N_12330,N_11890,N_11513);
nor U12331 (N_12331,N_11788,N_11902);
or U12332 (N_12332,N_11740,N_11862);
nand U12333 (N_12333,N_11598,N_11553);
nor U12334 (N_12334,N_11963,N_11955);
nand U12335 (N_12335,N_11840,N_11697);
or U12336 (N_12336,N_11530,N_11879);
nor U12337 (N_12337,N_11672,N_11570);
nor U12338 (N_12338,N_11828,N_11744);
and U12339 (N_12339,N_11931,N_11914);
xnor U12340 (N_12340,N_11683,N_11614);
xnor U12341 (N_12341,N_11731,N_11749);
xor U12342 (N_12342,N_11618,N_11528);
nor U12343 (N_12343,N_11512,N_11820);
xor U12344 (N_12344,N_11706,N_11949);
or U12345 (N_12345,N_11601,N_11702);
xor U12346 (N_12346,N_11936,N_11625);
or U12347 (N_12347,N_11562,N_11918);
or U12348 (N_12348,N_11506,N_11501);
nor U12349 (N_12349,N_11971,N_11995);
and U12350 (N_12350,N_11743,N_11800);
and U12351 (N_12351,N_11772,N_11656);
nor U12352 (N_12352,N_11727,N_11629);
nor U12353 (N_12353,N_11527,N_11594);
nor U12354 (N_12354,N_11657,N_11993);
nor U12355 (N_12355,N_11771,N_11755);
and U12356 (N_12356,N_11892,N_11651);
nand U12357 (N_12357,N_11518,N_11620);
or U12358 (N_12358,N_11889,N_11689);
and U12359 (N_12359,N_11871,N_11971);
or U12360 (N_12360,N_11549,N_11949);
nand U12361 (N_12361,N_11981,N_11548);
nor U12362 (N_12362,N_11936,N_11818);
xnor U12363 (N_12363,N_11958,N_11518);
xnor U12364 (N_12364,N_11583,N_11855);
nand U12365 (N_12365,N_11680,N_11510);
nor U12366 (N_12366,N_11678,N_11721);
nor U12367 (N_12367,N_11520,N_11978);
nand U12368 (N_12368,N_11681,N_11521);
xnor U12369 (N_12369,N_11516,N_11793);
or U12370 (N_12370,N_11728,N_11670);
xnor U12371 (N_12371,N_11721,N_11586);
nand U12372 (N_12372,N_11597,N_11985);
and U12373 (N_12373,N_11500,N_11648);
or U12374 (N_12374,N_11641,N_11650);
and U12375 (N_12375,N_11775,N_11850);
and U12376 (N_12376,N_11708,N_11710);
nor U12377 (N_12377,N_11939,N_11662);
nand U12378 (N_12378,N_11662,N_11931);
or U12379 (N_12379,N_11875,N_11526);
xnor U12380 (N_12380,N_11536,N_11828);
or U12381 (N_12381,N_11980,N_11638);
nand U12382 (N_12382,N_11608,N_11809);
nor U12383 (N_12383,N_11816,N_11635);
nand U12384 (N_12384,N_11739,N_11832);
nand U12385 (N_12385,N_11879,N_11924);
or U12386 (N_12386,N_11654,N_11535);
or U12387 (N_12387,N_11831,N_11948);
nor U12388 (N_12388,N_11742,N_11796);
or U12389 (N_12389,N_11606,N_11584);
nor U12390 (N_12390,N_11675,N_11679);
xnor U12391 (N_12391,N_11998,N_11547);
nor U12392 (N_12392,N_11707,N_11870);
xnor U12393 (N_12393,N_11587,N_11677);
xnor U12394 (N_12394,N_11863,N_11516);
or U12395 (N_12395,N_11739,N_11708);
and U12396 (N_12396,N_11790,N_11889);
and U12397 (N_12397,N_11576,N_11508);
and U12398 (N_12398,N_11940,N_11579);
nor U12399 (N_12399,N_11699,N_11731);
nor U12400 (N_12400,N_11711,N_11702);
and U12401 (N_12401,N_11678,N_11507);
nor U12402 (N_12402,N_11513,N_11602);
nand U12403 (N_12403,N_11742,N_11758);
and U12404 (N_12404,N_11977,N_11799);
and U12405 (N_12405,N_11725,N_11702);
xor U12406 (N_12406,N_11927,N_11612);
xnor U12407 (N_12407,N_11727,N_11779);
or U12408 (N_12408,N_11941,N_11940);
or U12409 (N_12409,N_11568,N_11992);
and U12410 (N_12410,N_11549,N_11681);
nor U12411 (N_12411,N_11852,N_11792);
or U12412 (N_12412,N_11847,N_11981);
xnor U12413 (N_12413,N_11509,N_11815);
nor U12414 (N_12414,N_11769,N_11958);
nand U12415 (N_12415,N_11562,N_11646);
xor U12416 (N_12416,N_11780,N_11598);
nor U12417 (N_12417,N_11925,N_11897);
xor U12418 (N_12418,N_11954,N_11516);
and U12419 (N_12419,N_11789,N_11983);
xor U12420 (N_12420,N_11506,N_11508);
and U12421 (N_12421,N_11607,N_11600);
xor U12422 (N_12422,N_11893,N_11603);
or U12423 (N_12423,N_11805,N_11996);
nor U12424 (N_12424,N_11727,N_11715);
nor U12425 (N_12425,N_11577,N_11527);
or U12426 (N_12426,N_11606,N_11769);
or U12427 (N_12427,N_11938,N_11743);
or U12428 (N_12428,N_11637,N_11972);
nand U12429 (N_12429,N_11901,N_11957);
nor U12430 (N_12430,N_11593,N_11646);
or U12431 (N_12431,N_11797,N_11770);
xor U12432 (N_12432,N_11779,N_11651);
or U12433 (N_12433,N_11552,N_11912);
xnor U12434 (N_12434,N_11885,N_11526);
nor U12435 (N_12435,N_11904,N_11669);
nand U12436 (N_12436,N_11681,N_11764);
xnor U12437 (N_12437,N_11521,N_11968);
nor U12438 (N_12438,N_11541,N_11542);
and U12439 (N_12439,N_11916,N_11999);
nor U12440 (N_12440,N_11739,N_11780);
nand U12441 (N_12441,N_11601,N_11854);
and U12442 (N_12442,N_11933,N_11751);
and U12443 (N_12443,N_11885,N_11720);
nor U12444 (N_12444,N_11589,N_11894);
xor U12445 (N_12445,N_11697,N_11866);
and U12446 (N_12446,N_11562,N_11773);
and U12447 (N_12447,N_11840,N_11740);
nor U12448 (N_12448,N_11879,N_11521);
and U12449 (N_12449,N_11728,N_11683);
nor U12450 (N_12450,N_11850,N_11645);
and U12451 (N_12451,N_11608,N_11569);
and U12452 (N_12452,N_11758,N_11955);
nor U12453 (N_12453,N_11971,N_11988);
nand U12454 (N_12454,N_11502,N_11635);
xnor U12455 (N_12455,N_11862,N_11764);
xor U12456 (N_12456,N_11990,N_11755);
nor U12457 (N_12457,N_11921,N_11589);
xor U12458 (N_12458,N_11537,N_11637);
and U12459 (N_12459,N_11766,N_11778);
xnor U12460 (N_12460,N_11585,N_11885);
nand U12461 (N_12461,N_11583,N_11883);
xor U12462 (N_12462,N_11787,N_11805);
and U12463 (N_12463,N_11878,N_11757);
xnor U12464 (N_12464,N_11802,N_11949);
and U12465 (N_12465,N_11660,N_11873);
xor U12466 (N_12466,N_11739,N_11639);
and U12467 (N_12467,N_11879,N_11947);
and U12468 (N_12468,N_11884,N_11968);
and U12469 (N_12469,N_11764,N_11903);
or U12470 (N_12470,N_11691,N_11698);
xnor U12471 (N_12471,N_11751,N_11936);
nor U12472 (N_12472,N_11616,N_11748);
or U12473 (N_12473,N_11816,N_11644);
or U12474 (N_12474,N_11548,N_11753);
and U12475 (N_12475,N_11956,N_11763);
and U12476 (N_12476,N_11791,N_11848);
or U12477 (N_12477,N_11880,N_11610);
nand U12478 (N_12478,N_11950,N_11744);
nor U12479 (N_12479,N_11623,N_11913);
xor U12480 (N_12480,N_11750,N_11528);
or U12481 (N_12481,N_11934,N_11588);
nand U12482 (N_12482,N_11828,N_11658);
xnor U12483 (N_12483,N_11923,N_11966);
and U12484 (N_12484,N_11538,N_11592);
or U12485 (N_12485,N_11697,N_11595);
or U12486 (N_12486,N_11940,N_11796);
or U12487 (N_12487,N_11618,N_11915);
nor U12488 (N_12488,N_11880,N_11579);
nand U12489 (N_12489,N_11768,N_11795);
or U12490 (N_12490,N_11720,N_11646);
nand U12491 (N_12491,N_11717,N_11791);
and U12492 (N_12492,N_11716,N_11986);
nor U12493 (N_12493,N_11988,N_11653);
and U12494 (N_12494,N_11737,N_11863);
xnor U12495 (N_12495,N_11665,N_11712);
nand U12496 (N_12496,N_11955,N_11594);
xnor U12497 (N_12497,N_11914,N_11883);
or U12498 (N_12498,N_11946,N_11661);
xnor U12499 (N_12499,N_11522,N_11959);
xor U12500 (N_12500,N_12311,N_12237);
nand U12501 (N_12501,N_12138,N_12422);
or U12502 (N_12502,N_12037,N_12192);
nor U12503 (N_12503,N_12174,N_12163);
and U12504 (N_12504,N_12032,N_12049);
nand U12505 (N_12505,N_12470,N_12019);
and U12506 (N_12506,N_12246,N_12279);
xnor U12507 (N_12507,N_12258,N_12053);
nand U12508 (N_12508,N_12484,N_12418);
or U12509 (N_12509,N_12287,N_12188);
nor U12510 (N_12510,N_12487,N_12055);
and U12511 (N_12511,N_12288,N_12227);
or U12512 (N_12512,N_12084,N_12464);
nand U12513 (N_12513,N_12369,N_12075);
and U12514 (N_12514,N_12080,N_12494);
xor U12515 (N_12515,N_12231,N_12147);
nor U12516 (N_12516,N_12426,N_12177);
or U12517 (N_12517,N_12186,N_12420);
xor U12518 (N_12518,N_12193,N_12078);
or U12519 (N_12519,N_12408,N_12136);
nand U12520 (N_12520,N_12140,N_12382);
or U12521 (N_12521,N_12180,N_12356);
nor U12522 (N_12522,N_12236,N_12299);
xnor U12523 (N_12523,N_12030,N_12085);
nor U12524 (N_12524,N_12374,N_12417);
and U12525 (N_12525,N_12387,N_12449);
and U12526 (N_12526,N_12437,N_12000);
nand U12527 (N_12527,N_12312,N_12359);
xnor U12528 (N_12528,N_12038,N_12284);
or U12529 (N_12529,N_12393,N_12006);
nor U12530 (N_12530,N_12152,N_12238);
or U12531 (N_12531,N_12275,N_12014);
or U12532 (N_12532,N_12303,N_12114);
and U12533 (N_12533,N_12282,N_12172);
and U12534 (N_12534,N_12414,N_12306);
or U12535 (N_12535,N_12293,N_12065);
nor U12536 (N_12536,N_12101,N_12241);
nor U12537 (N_12537,N_12212,N_12351);
or U12538 (N_12538,N_12024,N_12254);
and U12539 (N_12539,N_12283,N_12402);
or U12540 (N_12540,N_12358,N_12371);
nand U12541 (N_12541,N_12438,N_12433);
and U12542 (N_12542,N_12073,N_12416);
xor U12543 (N_12543,N_12201,N_12466);
nand U12544 (N_12544,N_12357,N_12045);
or U12545 (N_12545,N_12394,N_12345);
nand U12546 (N_12546,N_12327,N_12329);
and U12547 (N_12547,N_12046,N_12107);
or U12548 (N_12548,N_12074,N_12267);
and U12549 (N_12549,N_12217,N_12453);
nand U12550 (N_12550,N_12009,N_12111);
nor U12551 (N_12551,N_12167,N_12131);
nor U12552 (N_12552,N_12214,N_12054);
or U12553 (N_12553,N_12092,N_12368);
or U12554 (N_12554,N_12292,N_12025);
xnor U12555 (N_12555,N_12332,N_12120);
nor U12556 (N_12556,N_12134,N_12017);
nand U12557 (N_12557,N_12335,N_12353);
nand U12558 (N_12558,N_12277,N_12404);
xor U12559 (N_12559,N_12226,N_12289);
or U12560 (N_12560,N_12137,N_12033);
and U12561 (N_12561,N_12328,N_12251);
nor U12562 (N_12562,N_12469,N_12446);
xnor U12563 (N_12563,N_12386,N_12350);
xnor U12564 (N_12564,N_12118,N_12452);
or U12565 (N_12565,N_12139,N_12223);
nand U12566 (N_12566,N_12082,N_12077);
or U12567 (N_12567,N_12268,N_12336);
or U12568 (N_12568,N_12243,N_12304);
xor U12569 (N_12569,N_12108,N_12124);
and U12570 (N_12570,N_12203,N_12381);
or U12571 (N_12571,N_12432,N_12298);
nand U12572 (N_12572,N_12479,N_12086);
nand U12573 (N_12573,N_12185,N_12153);
or U12574 (N_12574,N_12112,N_12070);
nand U12575 (N_12575,N_12383,N_12321);
nor U12576 (N_12576,N_12181,N_12158);
nor U12577 (N_12577,N_12228,N_12144);
and U12578 (N_12578,N_12061,N_12057);
or U12579 (N_12579,N_12388,N_12488);
nor U12580 (N_12580,N_12104,N_12278);
nor U12581 (N_12581,N_12233,N_12378);
nor U12582 (N_12582,N_12151,N_12483);
or U12583 (N_12583,N_12271,N_12083);
or U12584 (N_12584,N_12413,N_12333);
nand U12585 (N_12585,N_12425,N_12302);
or U12586 (N_12586,N_12015,N_12314);
xnor U12587 (N_12587,N_12410,N_12389);
xnor U12588 (N_12588,N_12317,N_12175);
xor U12589 (N_12589,N_12361,N_12334);
or U12590 (N_12590,N_12263,N_12403);
nor U12591 (N_12591,N_12097,N_12339);
nor U12592 (N_12592,N_12016,N_12222);
or U12593 (N_12593,N_12265,N_12255);
nor U12594 (N_12594,N_12338,N_12225);
nor U12595 (N_12595,N_12309,N_12471);
nand U12596 (N_12596,N_12218,N_12341);
or U12597 (N_12597,N_12149,N_12459);
nand U12598 (N_12598,N_12297,N_12021);
xor U12599 (N_12599,N_12373,N_12044);
and U12600 (N_12600,N_12444,N_12322);
xor U12601 (N_12601,N_12472,N_12012);
nand U12602 (N_12602,N_12011,N_12262);
nand U12603 (N_12603,N_12160,N_12123);
nand U12604 (N_12604,N_12455,N_12477);
xnor U12605 (N_12605,N_12428,N_12161);
nor U12606 (N_12606,N_12220,N_12276);
nor U12607 (N_12607,N_12330,N_12463);
nor U12608 (N_12608,N_12247,N_12252);
or U12609 (N_12609,N_12056,N_12031);
and U12610 (N_12610,N_12081,N_12424);
xnor U12611 (N_12611,N_12029,N_12407);
nand U12612 (N_12612,N_12259,N_12480);
and U12613 (N_12613,N_12261,N_12363);
xor U12614 (N_12614,N_12191,N_12256);
nor U12615 (N_12615,N_12397,N_12244);
and U12616 (N_12616,N_12266,N_12089);
nand U12617 (N_12617,N_12187,N_12143);
nand U12618 (N_12618,N_12476,N_12431);
nand U12619 (N_12619,N_12051,N_12286);
or U12620 (N_12620,N_12159,N_12064);
nor U12621 (N_12621,N_12179,N_12347);
nor U12622 (N_12622,N_12039,N_12168);
and U12623 (N_12623,N_12170,N_12202);
nand U12624 (N_12624,N_12491,N_12035);
xnor U12625 (N_12625,N_12221,N_12496);
or U12626 (N_12626,N_12028,N_12235);
and U12627 (N_12627,N_12430,N_12337);
and U12628 (N_12628,N_12154,N_12385);
or U12629 (N_12629,N_12047,N_12142);
nor U12630 (N_12630,N_12490,N_12069);
xnor U12631 (N_12631,N_12224,N_12245);
nor U12632 (N_12632,N_12117,N_12189);
or U12633 (N_12633,N_12421,N_12102);
nor U12634 (N_12634,N_12380,N_12248);
nand U12635 (N_12635,N_12088,N_12105);
xnor U12636 (N_12636,N_12099,N_12364);
and U12637 (N_12637,N_12473,N_12023);
or U12638 (N_12638,N_12405,N_12448);
or U12639 (N_12639,N_12443,N_12209);
nand U12640 (N_12640,N_12468,N_12100);
xnor U12641 (N_12641,N_12270,N_12348);
or U12642 (N_12642,N_12458,N_12076);
nand U12643 (N_12643,N_12384,N_12213);
and U12644 (N_12644,N_12207,N_12122);
xnor U12645 (N_12645,N_12253,N_12162);
nor U12646 (N_12646,N_12127,N_12194);
and U12647 (N_12647,N_12157,N_12485);
or U12648 (N_12648,N_12445,N_12022);
and U12649 (N_12649,N_12280,N_12467);
and U12650 (N_12650,N_12439,N_12215);
nor U12651 (N_12651,N_12001,N_12310);
xnor U12652 (N_12652,N_12447,N_12242);
and U12653 (N_12653,N_12323,N_12027);
and U12654 (N_12654,N_12205,N_12096);
nor U12655 (N_12655,N_12273,N_12199);
nand U12656 (N_12656,N_12498,N_12190);
xnor U12657 (N_12657,N_12481,N_12379);
xor U12658 (N_12658,N_12367,N_12493);
xnor U12659 (N_12659,N_12419,N_12132);
xnor U12660 (N_12660,N_12034,N_12206);
nor U12661 (N_12661,N_12440,N_12020);
nand U12662 (N_12662,N_12435,N_12366);
nand U12663 (N_12663,N_12489,N_12094);
nand U12664 (N_12664,N_12307,N_12198);
and U12665 (N_12665,N_12274,N_12173);
or U12666 (N_12666,N_12450,N_12063);
nor U12667 (N_12667,N_12135,N_12121);
and U12668 (N_12668,N_12462,N_12036);
nor U12669 (N_12669,N_12331,N_12040);
and U12670 (N_12670,N_12294,N_12442);
nor U12671 (N_12671,N_12395,N_12377);
or U12672 (N_12672,N_12360,N_12058);
xor U12673 (N_12673,N_12349,N_12184);
xor U12674 (N_12674,N_12146,N_12013);
nor U12675 (N_12675,N_12313,N_12090);
xnor U12676 (N_12676,N_12316,N_12461);
nand U12677 (N_12677,N_12296,N_12196);
nand U12678 (N_12678,N_12067,N_12370);
nand U12679 (N_12679,N_12007,N_12043);
or U12680 (N_12680,N_12026,N_12399);
xor U12681 (N_12681,N_12457,N_12400);
and U12682 (N_12682,N_12326,N_12178);
nand U12683 (N_12683,N_12062,N_12441);
and U12684 (N_12684,N_12346,N_12355);
and U12685 (N_12685,N_12318,N_12176);
and U12686 (N_12686,N_12492,N_12269);
xnor U12687 (N_12687,N_12018,N_12182);
nand U12688 (N_12688,N_12210,N_12465);
xor U12689 (N_12689,N_12169,N_12008);
nor U12690 (N_12690,N_12362,N_12406);
nor U12691 (N_12691,N_12133,N_12423);
nand U12692 (N_12692,N_12125,N_12415);
and U12693 (N_12693,N_12434,N_12300);
nand U12694 (N_12694,N_12071,N_12052);
and U12695 (N_12695,N_12087,N_12150);
xor U12696 (N_12696,N_12281,N_12059);
and U12697 (N_12697,N_12372,N_12454);
nand U12698 (N_12698,N_12079,N_12340);
nand U12699 (N_12699,N_12155,N_12165);
nor U12700 (N_12700,N_12230,N_12392);
nand U12701 (N_12701,N_12456,N_12482);
or U12702 (N_12702,N_12436,N_12126);
and U12703 (N_12703,N_12048,N_12451);
or U12704 (N_12704,N_12145,N_12325);
xor U12705 (N_12705,N_12103,N_12042);
xnor U12706 (N_12706,N_12156,N_12211);
xnor U12707 (N_12707,N_12290,N_12344);
and U12708 (N_12708,N_12411,N_12401);
nor U12709 (N_12709,N_12010,N_12116);
and U12710 (N_12710,N_12308,N_12072);
nand U12711 (N_12711,N_12365,N_12249);
or U12712 (N_12712,N_12115,N_12319);
nor U12713 (N_12713,N_12301,N_12068);
nor U12714 (N_12714,N_12128,N_12352);
or U12715 (N_12715,N_12091,N_12095);
xor U12716 (N_12716,N_12171,N_12412);
nand U12717 (N_12717,N_12342,N_12396);
and U12718 (N_12718,N_12390,N_12129);
or U12719 (N_12719,N_12130,N_12315);
nand U12720 (N_12720,N_12429,N_12183);
nor U12721 (N_12721,N_12106,N_12041);
nand U12722 (N_12722,N_12200,N_12208);
or U12723 (N_12723,N_12272,N_12164);
xor U12724 (N_12724,N_12295,N_12232);
nor U12725 (N_12725,N_12305,N_12148);
or U12726 (N_12726,N_12197,N_12005);
nor U12727 (N_12727,N_12166,N_12427);
nand U12728 (N_12728,N_12003,N_12285);
or U12729 (N_12729,N_12050,N_12478);
nor U12730 (N_12730,N_12219,N_12320);
and U12731 (N_12731,N_12098,N_12240);
xnor U12732 (N_12732,N_12002,N_12474);
xor U12733 (N_12733,N_12324,N_12460);
or U12734 (N_12734,N_12497,N_12113);
nor U12735 (N_12735,N_12495,N_12234);
nor U12736 (N_12736,N_12376,N_12093);
xnor U12737 (N_12737,N_12260,N_12004);
and U12738 (N_12738,N_12216,N_12486);
and U12739 (N_12739,N_12391,N_12264);
and U12740 (N_12740,N_12250,N_12060);
and U12741 (N_12741,N_12119,N_12110);
nor U12742 (N_12742,N_12109,N_12239);
and U12743 (N_12743,N_12066,N_12343);
xor U12744 (N_12744,N_12141,N_12354);
or U12745 (N_12745,N_12499,N_12398);
or U12746 (N_12746,N_12195,N_12475);
or U12747 (N_12747,N_12409,N_12375);
nand U12748 (N_12748,N_12257,N_12229);
or U12749 (N_12749,N_12204,N_12291);
and U12750 (N_12750,N_12132,N_12480);
nand U12751 (N_12751,N_12031,N_12484);
nand U12752 (N_12752,N_12046,N_12088);
or U12753 (N_12753,N_12021,N_12012);
nand U12754 (N_12754,N_12373,N_12021);
xnor U12755 (N_12755,N_12264,N_12080);
and U12756 (N_12756,N_12094,N_12230);
and U12757 (N_12757,N_12037,N_12165);
or U12758 (N_12758,N_12305,N_12226);
nor U12759 (N_12759,N_12265,N_12115);
nand U12760 (N_12760,N_12465,N_12411);
or U12761 (N_12761,N_12206,N_12143);
nor U12762 (N_12762,N_12235,N_12365);
nor U12763 (N_12763,N_12395,N_12126);
nand U12764 (N_12764,N_12345,N_12443);
and U12765 (N_12765,N_12048,N_12342);
xnor U12766 (N_12766,N_12174,N_12252);
and U12767 (N_12767,N_12211,N_12019);
nor U12768 (N_12768,N_12337,N_12051);
nand U12769 (N_12769,N_12056,N_12151);
nor U12770 (N_12770,N_12220,N_12080);
xor U12771 (N_12771,N_12030,N_12273);
nor U12772 (N_12772,N_12294,N_12093);
nor U12773 (N_12773,N_12175,N_12133);
nor U12774 (N_12774,N_12454,N_12416);
xnor U12775 (N_12775,N_12322,N_12244);
and U12776 (N_12776,N_12131,N_12130);
and U12777 (N_12777,N_12359,N_12206);
and U12778 (N_12778,N_12493,N_12019);
and U12779 (N_12779,N_12361,N_12019);
nand U12780 (N_12780,N_12403,N_12286);
and U12781 (N_12781,N_12370,N_12007);
or U12782 (N_12782,N_12382,N_12116);
or U12783 (N_12783,N_12268,N_12389);
and U12784 (N_12784,N_12397,N_12084);
nand U12785 (N_12785,N_12239,N_12448);
or U12786 (N_12786,N_12493,N_12000);
and U12787 (N_12787,N_12159,N_12343);
nor U12788 (N_12788,N_12374,N_12461);
nor U12789 (N_12789,N_12237,N_12352);
or U12790 (N_12790,N_12492,N_12026);
xnor U12791 (N_12791,N_12418,N_12366);
xnor U12792 (N_12792,N_12493,N_12246);
nor U12793 (N_12793,N_12391,N_12135);
nand U12794 (N_12794,N_12432,N_12299);
nand U12795 (N_12795,N_12346,N_12038);
xor U12796 (N_12796,N_12081,N_12005);
nor U12797 (N_12797,N_12298,N_12389);
nor U12798 (N_12798,N_12474,N_12091);
nor U12799 (N_12799,N_12040,N_12377);
or U12800 (N_12800,N_12196,N_12217);
and U12801 (N_12801,N_12249,N_12360);
or U12802 (N_12802,N_12368,N_12072);
nand U12803 (N_12803,N_12416,N_12450);
nand U12804 (N_12804,N_12318,N_12144);
or U12805 (N_12805,N_12368,N_12022);
nor U12806 (N_12806,N_12297,N_12286);
nor U12807 (N_12807,N_12059,N_12421);
nand U12808 (N_12808,N_12221,N_12311);
nor U12809 (N_12809,N_12263,N_12179);
or U12810 (N_12810,N_12264,N_12289);
nand U12811 (N_12811,N_12135,N_12126);
nor U12812 (N_12812,N_12069,N_12292);
nand U12813 (N_12813,N_12339,N_12382);
and U12814 (N_12814,N_12319,N_12302);
nor U12815 (N_12815,N_12327,N_12266);
or U12816 (N_12816,N_12286,N_12339);
and U12817 (N_12817,N_12309,N_12132);
nor U12818 (N_12818,N_12062,N_12423);
or U12819 (N_12819,N_12472,N_12294);
and U12820 (N_12820,N_12214,N_12453);
nand U12821 (N_12821,N_12405,N_12463);
or U12822 (N_12822,N_12409,N_12221);
nand U12823 (N_12823,N_12038,N_12106);
and U12824 (N_12824,N_12418,N_12241);
nor U12825 (N_12825,N_12245,N_12422);
and U12826 (N_12826,N_12488,N_12357);
nor U12827 (N_12827,N_12414,N_12423);
and U12828 (N_12828,N_12181,N_12236);
and U12829 (N_12829,N_12171,N_12161);
or U12830 (N_12830,N_12009,N_12317);
xor U12831 (N_12831,N_12352,N_12365);
nand U12832 (N_12832,N_12066,N_12048);
nor U12833 (N_12833,N_12322,N_12251);
and U12834 (N_12834,N_12276,N_12024);
or U12835 (N_12835,N_12207,N_12202);
and U12836 (N_12836,N_12345,N_12075);
or U12837 (N_12837,N_12291,N_12159);
nand U12838 (N_12838,N_12351,N_12060);
nand U12839 (N_12839,N_12225,N_12040);
and U12840 (N_12840,N_12246,N_12093);
xnor U12841 (N_12841,N_12285,N_12220);
and U12842 (N_12842,N_12377,N_12437);
xnor U12843 (N_12843,N_12179,N_12498);
nor U12844 (N_12844,N_12343,N_12262);
xor U12845 (N_12845,N_12142,N_12366);
xnor U12846 (N_12846,N_12448,N_12197);
xor U12847 (N_12847,N_12015,N_12242);
nor U12848 (N_12848,N_12312,N_12147);
xnor U12849 (N_12849,N_12394,N_12032);
nand U12850 (N_12850,N_12471,N_12259);
nand U12851 (N_12851,N_12196,N_12346);
nor U12852 (N_12852,N_12189,N_12106);
or U12853 (N_12853,N_12326,N_12004);
nor U12854 (N_12854,N_12489,N_12130);
or U12855 (N_12855,N_12407,N_12030);
nor U12856 (N_12856,N_12052,N_12462);
xor U12857 (N_12857,N_12078,N_12158);
xnor U12858 (N_12858,N_12144,N_12158);
and U12859 (N_12859,N_12396,N_12442);
and U12860 (N_12860,N_12389,N_12222);
nor U12861 (N_12861,N_12078,N_12368);
and U12862 (N_12862,N_12119,N_12239);
and U12863 (N_12863,N_12064,N_12405);
and U12864 (N_12864,N_12270,N_12356);
and U12865 (N_12865,N_12296,N_12470);
xor U12866 (N_12866,N_12231,N_12150);
or U12867 (N_12867,N_12025,N_12082);
and U12868 (N_12868,N_12367,N_12408);
or U12869 (N_12869,N_12305,N_12278);
xor U12870 (N_12870,N_12077,N_12089);
xor U12871 (N_12871,N_12292,N_12229);
xnor U12872 (N_12872,N_12437,N_12021);
nand U12873 (N_12873,N_12168,N_12161);
xnor U12874 (N_12874,N_12009,N_12052);
nand U12875 (N_12875,N_12354,N_12427);
nand U12876 (N_12876,N_12093,N_12156);
and U12877 (N_12877,N_12045,N_12054);
nand U12878 (N_12878,N_12212,N_12285);
xor U12879 (N_12879,N_12133,N_12293);
xnor U12880 (N_12880,N_12132,N_12161);
nand U12881 (N_12881,N_12447,N_12002);
nor U12882 (N_12882,N_12189,N_12482);
xnor U12883 (N_12883,N_12420,N_12298);
or U12884 (N_12884,N_12383,N_12384);
xnor U12885 (N_12885,N_12042,N_12040);
and U12886 (N_12886,N_12224,N_12403);
nor U12887 (N_12887,N_12260,N_12171);
xor U12888 (N_12888,N_12026,N_12483);
or U12889 (N_12889,N_12390,N_12242);
and U12890 (N_12890,N_12179,N_12458);
nor U12891 (N_12891,N_12239,N_12026);
nand U12892 (N_12892,N_12329,N_12155);
xnor U12893 (N_12893,N_12151,N_12475);
and U12894 (N_12894,N_12436,N_12238);
nand U12895 (N_12895,N_12157,N_12436);
and U12896 (N_12896,N_12224,N_12213);
and U12897 (N_12897,N_12284,N_12491);
or U12898 (N_12898,N_12032,N_12171);
and U12899 (N_12899,N_12209,N_12163);
nor U12900 (N_12900,N_12469,N_12103);
or U12901 (N_12901,N_12400,N_12420);
and U12902 (N_12902,N_12029,N_12062);
nand U12903 (N_12903,N_12196,N_12429);
or U12904 (N_12904,N_12146,N_12316);
nand U12905 (N_12905,N_12300,N_12438);
nand U12906 (N_12906,N_12370,N_12099);
or U12907 (N_12907,N_12462,N_12210);
or U12908 (N_12908,N_12056,N_12350);
and U12909 (N_12909,N_12047,N_12038);
and U12910 (N_12910,N_12005,N_12107);
xor U12911 (N_12911,N_12222,N_12057);
and U12912 (N_12912,N_12312,N_12156);
and U12913 (N_12913,N_12499,N_12381);
xnor U12914 (N_12914,N_12065,N_12260);
and U12915 (N_12915,N_12258,N_12288);
and U12916 (N_12916,N_12041,N_12214);
and U12917 (N_12917,N_12072,N_12065);
nand U12918 (N_12918,N_12000,N_12400);
nor U12919 (N_12919,N_12085,N_12202);
nand U12920 (N_12920,N_12006,N_12190);
xnor U12921 (N_12921,N_12418,N_12444);
nor U12922 (N_12922,N_12476,N_12156);
xor U12923 (N_12923,N_12315,N_12465);
nor U12924 (N_12924,N_12470,N_12267);
and U12925 (N_12925,N_12368,N_12087);
or U12926 (N_12926,N_12289,N_12182);
and U12927 (N_12927,N_12399,N_12069);
nand U12928 (N_12928,N_12486,N_12326);
xor U12929 (N_12929,N_12042,N_12241);
nor U12930 (N_12930,N_12181,N_12329);
nand U12931 (N_12931,N_12317,N_12179);
nand U12932 (N_12932,N_12201,N_12181);
xnor U12933 (N_12933,N_12496,N_12290);
or U12934 (N_12934,N_12181,N_12426);
nor U12935 (N_12935,N_12423,N_12446);
nand U12936 (N_12936,N_12345,N_12248);
or U12937 (N_12937,N_12159,N_12120);
nor U12938 (N_12938,N_12048,N_12133);
nor U12939 (N_12939,N_12264,N_12208);
or U12940 (N_12940,N_12459,N_12439);
nor U12941 (N_12941,N_12127,N_12284);
nor U12942 (N_12942,N_12197,N_12371);
or U12943 (N_12943,N_12355,N_12056);
nand U12944 (N_12944,N_12100,N_12312);
nor U12945 (N_12945,N_12201,N_12125);
or U12946 (N_12946,N_12484,N_12245);
and U12947 (N_12947,N_12356,N_12396);
and U12948 (N_12948,N_12416,N_12077);
xnor U12949 (N_12949,N_12164,N_12479);
nand U12950 (N_12950,N_12190,N_12301);
nor U12951 (N_12951,N_12159,N_12233);
nand U12952 (N_12952,N_12052,N_12162);
or U12953 (N_12953,N_12269,N_12464);
or U12954 (N_12954,N_12150,N_12102);
xor U12955 (N_12955,N_12454,N_12487);
xnor U12956 (N_12956,N_12125,N_12357);
and U12957 (N_12957,N_12000,N_12019);
nor U12958 (N_12958,N_12359,N_12069);
nand U12959 (N_12959,N_12099,N_12098);
and U12960 (N_12960,N_12319,N_12409);
or U12961 (N_12961,N_12278,N_12413);
nor U12962 (N_12962,N_12462,N_12109);
xor U12963 (N_12963,N_12129,N_12114);
or U12964 (N_12964,N_12061,N_12173);
or U12965 (N_12965,N_12288,N_12247);
nand U12966 (N_12966,N_12450,N_12028);
and U12967 (N_12967,N_12336,N_12385);
xnor U12968 (N_12968,N_12215,N_12426);
xnor U12969 (N_12969,N_12455,N_12183);
or U12970 (N_12970,N_12185,N_12028);
nand U12971 (N_12971,N_12067,N_12071);
or U12972 (N_12972,N_12153,N_12494);
and U12973 (N_12973,N_12341,N_12068);
or U12974 (N_12974,N_12302,N_12260);
nand U12975 (N_12975,N_12468,N_12062);
xor U12976 (N_12976,N_12216,N_12186);
nor U12977 (N_12977,N_12143,N_12152);
nand U12978 (N_12978,N_12427,N_12095);
or U12979 (N_12979,N_12278,N_12009);
nand U12980 (N_12980,N_12206,N_12337);
nor U12981 (N_12981,N_12283,N_12329);
and U12982 (N_12982,N_12222,N_12118);
nand U12983 (N_12983,N_12197,N_12166);
nand U12984 (N_12984,N_12480,N_12179);
xor U12985 (N_12985,N_12065,N_12305);
nand U12986 (N_12986,N_12160,N_12353);
xnor U12987 (N_12987,N_12304,N_12184);
nand U12988 (N_12988,N_12366,N_12362);
or U12989 (N_12989,N_12269,N_12461);
xnor U12990 (N_12990,N_12060,N_12488);
and U12991 (N_12991,N_12182,N_12016);
nor U12992 (N_12992,N_12243,N_12221);
and U12993 (N_12993,N_12053,N_12072);
and U12994 (N_12994,N_12434,N_12138);
or U12995 (N_12995,N_12146,N_12492);
nand U12996 (N_12996,N_12241,N_12108);
and U12997 (N_12997,N_12146,N_12290);
xor U12998 (N_12998,N_12464,N_12454);
and U12999 (N_12999,N_12266,N_12445);
nor U13000 (N_13000,N_12801,N_12934);
xor U13001 (N_13001,N_12969,N_12998);
nand U13002 (N_13002,N_12936,N_12868);
and U13003 (N_13003,N_12614,N_12895);
nand U13004 (N_13004,N_12797,N_12566);
nand U13005 (N_13005,N_12767,N_12911);
nand U13006 (N_13006,N_12514,N_12510);
or U13007 (N_13007,N_12594,N_12737);
nand U13008 (N_13008,N_12757,N_12610);
and U13009 (N_13009,N_12677,N_12504);
nor U13010 (N_13010,N_12662,N_12974);
nand U13011 (N_13011,N_12512,N_12517);
xor U13012 (N_13012,N_12861,N_12946);
and U13013 (N_13013,N_12620,N_12845);
or U13014 (N_13014,N_12597,N_12756);
and U13015 (N_13015,N_12755,N_12778);
nand U13016 (N_13016,N_12670,N_12844);
or U13017 (N_13017,N_12718,N_12678);
nor U13018 (N_13018,N_12912,N_12683);
nand U13019 (N_13019,N_12838,N_12686);
and U13020 (N_13020,N_12891,N_12884);
and U13021 (N_13021,N_12712,N_12704);
xor U13022 (N_13022,N_12954,N_12656);
nand U13023 (N_13023,N_12876,N_12859);
xnor U13024 (N_13024,N_12506,N_12933);
xor U13025 (N_13025,N_12693,N_12994);
or U13026 (N_13026,N_12643,N_12765);
and U13027 (N_13027,N_12802,N_12703);
or U13028 (N_13028,N_12874,N_12654);
xnor U13029 (N_13029,N_12511,N_12720);
nand U13030 (N_13030,N_12746,N_12803);
nand U13031 (N_13031,N_12525,N_12878);
or U13032 (N_13032,N_12988,N_12665);
or U13033 (N_13033,N_12534,N_12873);
nor U13034 (N_13034,N_12660,N_12653);
and U13035 (N_13035,N_12667,N_12918);
nand U13036 (N_13036,N_12550,N_12531);
or U13037 (N_13037,N_12714,N_12707);
xor U13038 (N_13038,N_12561,N_12927);
and U13039 (N_13039,N_12948,N_12817);
xor U13040 (N_13040,N_12735,N_12505);
nor U13041 (N_13041,N_12698,N_12930);
xor U13042 (N_13042,N_12513,N_12533);
or U13043 (N_13043,N_12983,N_12588);
and U13044 (N_13044,N_12527,N_12890);
nand U13045 (N_13045,N_12907,N_12734);
nand U13046 (N_13046,N_12780,N_12771);
xor U13047 (N_13047,N_12701,N_12999);
nand U13048 (N_13048,N_12809,N_12582);
or U13049 (N_13049,N_12556,N_12549);
nor U13050 (N_13050,N_12799,N_12949);
nand U13051 (N_13051,N_12975,N_12553);
nor U13052 (N_13052,N_12924,N_12840);
xor U13053 (N_13053,N_12634,N_12896);
xor U13054 (N_13054,N_12617,N_12547);
or U13055 (N_13055,N_12788,N_12708);
nand U13056 (N_13056,N_12627,N_12622);
xor U13057 (N_13057,N_12978,N_12850);
xor U13058 (N_13058,N_12903,N_12623);
and U13059 (N_13059,N_12702,N_12601);
nor U13060 (N_13060,N_12650,N_12926);
nor U13061 (N_13061,N_12851,N_12532);
xor U13062 (N_13062,N_12747,N_12633);
or U13063 (N_13063,N_12822,N_12996);
nor U13064 (N_13064,N_12958,N_12543);
xnor U13065 (N_13065,N_12570,N_12986);
nand U13066 (N_13066,N_12618,N_12729);
nor U13067 (N_13067,N_12834,N_12919);
xnor U13068 (N_13068,N_12824,N_12640);
and U13069 (N_13069,N_12880,N_12877);
xnor U13070 (N_13070,N_12571,N_12843);
xnor U13071 (N_13071,N_12738,N_12816);
nor U13072 (N_13072,N_12631,N_12544);
xor U13073 (N_13073,N_12967,N_12515);
nand U13074 (N_13074,N_12624,N_12675);
and U13075 (N_13075,N_12836,N_12914);
nor U13076 (N_13076,N_12984,N_12893);
xor U13077 (N_13077,N_12774,N_12727);
or U13078 (N_13078,N_12555,N_12962);
nand U13079 (N_13079,N_12917,N_12853);
nor U13080 (N_13080,N_12621,N_12945);
or U13081 (N_13081,N_12760,N_12639);
nor U13082 (N_13082,N_12754,N_12689);
nand U13083 (N_13083,N_12635,N_12957);
and U13084 (N_13084,N_12781,N_12856);
and U13085 (N_13085,N_12661,N_12966);
or U13086 (N_13086,N_12598,N_12637);
xnor U13087 (N_13087,N_12813,N_12695);
nand U13088 (N_13088,N_12832,N_12937);
nand U13089 (N_13089,N_12723,N_12811);
or U13090 (N_13090,N_12779,N_12894);
nor U13091 (N_13091,N_12666,N_12649);
or U13092 (N_13092,N_12605,N_12535);
xor U13093 (N_13093,N_12697,N_12971);
nand U13094 (N_13094,N_12943,N_12915);
and U13095 (N_13095,N_12955,N_12795);
xor U13096 (N_13096,N_12992,N_12730);
and U13097 (N_13097,N_12710,N_12787);
xnor U13098 (N_13098,N_12608,N_12910);
xnor U13099 (N_13099,N_12941,N_12833);
and U13100 (N_13100,N_12920,N_12560);
xnor U13101 (N_13101,N_12672,N_12800);
nor U13102 (N_13102,N_12961,N_12573);
or U13103 (N_13103,N_12987,N_12558);
nand U13104 (N_13104,N_12596,N_12794);
nor U13105 (N_13105,N_12763,N_12518);
or U13106 (N_13106,N_12806,N_12991);
nand U13107 (N_13107,N_12509,N_12959);
xor U13108 (N_13108,N_12557,N_12897);
and U13109 (N_13109,N_12883,N_12977);
or U13110 (N_13110,N_12798,N_12644);
nand U13111 (N_13111,N_12785,N_12725);
or U13112 (N_13112,N_12839,N_12860);
nand U13113 (N_13113,N_12748,N_12939);
xnor U13114 (N_13114,N_12989,N_12953);
or U13115 (N_13115,N_12786,N_12516);
nor U13116 (N_13116,N_12659,N_12993);
nand U13117 (N_13117,N_12849,N_12715);
or U13118 (N_13118,N_12902,N_12674);
nand U13119 (N_13119,N_12805,N_12777);
and U13120 (N_13120,N_12673,N_12972);
nor U13121 (N_13121,N_12886,N_12562);
and U13122 (N_13122,N_12584,N_12600);
nand U13123 (N_13123,N_12854,N_12935);
and U13124 (N_13124,N_12576,N_12846);
nor U13125 (N_13125,N_12680,N_12830);
xor U13126 (N_13126,N_12864,N_12690);
or U13127 (N_13127,N_12810,N_12572);
or U13128 (N_13128,N_12647,N_12990);
nor U13129 (N_13129,N_12537,N_12828);
xor U13130 (N_13130,N_12554,N_12520);
nand U13131 (N_13131,N_12741,N_12539);
xnor U13132 (N_13132,N_12646,N_12595);
nand U13133 (N_13133,N_12500,N_12751);
xnor U13134 (N_13134,N_12913,N_12835);
and U13135 (N_13135,N_12808,N_12724);
xnor U13136 (N_13136,N_12812,N_12616);
xor U13137 (N_13137,N_12916,N_12540);
and U13138 (N_13138,N_12932,N_12743);
nand U13139 (N_13139,N_12577,N_12638);
or U13140 (N_13140,N_12973,N_12669);
nor U13141 (N_13141,N_12931,N_12521);
nor U13142 (N_13142,N_12681,N_12736);
nor U13143 (N_13143,N_12745,N_12970);
and U13144 (N_13144,N_12776,N_12579);
nor U13145 (N_13145,N_12688,N_12591);
nor U13146 (N_13146,N_12732,N_12648);
nand U13147 (N_13147,N_12565,N_12968);
nor U13148 (N_13148,N_12821,N_12586);
nand U13149 (N_13149,N_12872,N_12536);
xnor U13150 (N_13150,N_12726,N_12524);
and U13151 (N_13151,N_12879,N_12921);
and U13152 (N_13152,N_12892,N_12869);
or U13153 (N_13153,N_12789,N_12578);
nand U13154 (N_13154,N_12522,N_12655);
nor U13155 (N_13155,N_12641,N_12530);
or U13156 (N_13156,N_12719,N_12875);
nand U13157 (N_13157,N_12923,N_12705);
xnor U13158 (N_13158,N_12906,N_12713);
xor U13159 (N_13159,N_12548,N_12749);
nor U13160 (N_13160,N_12752,N_12717);
and U13161 (N_13161,N_12866,N_12908);
xor U13162 (N_13162,N_12568,N_12676);
nand U13163 (N_13163,N_12758,N_12694);
or U13164 (N_13164,N_12569,N_12528);
xor U13165 (N_13165,N_12855,N_12825);
nand U13166 (N_13166,N_12657,N_12602);
or U13167 (N_13167,N_12862,N_12699);
nand U13168 (N_13168,N_12503,N_12619);
and U13169 (N_13169,N_12700,N_12909);
nand U13170 (N_13170,N_12750,N_12881);
and U13171 (N_13171,N_12938,N_12922);
nor U13172 (N_13172,N_12963,N_12819);
and U13173 (N_13173,N_12564,N_12629);
nand U13174 (N_13174,N_12904,N_12739);
nand U13175 (N_13175,N_12815,N_12740);
xnor U13176 (N_13176,N_12615,N_12706);
nand U13177 (N_13177,N_12529,N_12563);
nor U13178 (N_13178,N_12867,N_12980);
nand U13179 (N_13179,N_12545,N_12642);
or U13180 (N_13180,N_12956,N_12508);
nand U13181 (N_13181,N_12589,N_12679);
and U13182 (N_13182,N_12841,N_12901);
or U13183 (N_13183,N_12784,N_12685);
nand U13184 (N_13184,N_12769,N_12728);
xor U13185 (N_13185,N_12722,N_12606);
or U13186 (N_13186,N_12898,N_12796);
xor U13187 (N_13187,N_12603,N_12753);
and U13188 (N_13188,N_12772,N_12976);
xor U13189 (N_13189,N_12590,N_12742);
xor U13190 (N_13190,N_12551,N_12546);
or U13191 (N_13191,N_12538,N_12950);
nor U13192 (N_13192,N_12501,N_12768);
xor U13193 (N_13193,N_12721,N_12733);
or U13194 (N_13194,N_12965,N_12502);
nor U13195 (N_13195,N_12609,N_12814);
nand U13196 (N_13196,N_12793,N_12611);
and U13197 (N_13197,N_12773,N_12942);
nor U13198 (N_13198,N_12684,N_12592);
and U13199 (N_13199,N_12507,N_12857);
nand U13200 (N_13200,N_12865,N_12671);
and U13201 (N_13201,N_12587,N_12552);
nor U13202 (N_13202,N_12925,N_12762);
and U13203 (N_13203,N_12766,N_12652);
nand U13204 (N_13204,N_12632,N_12870);
nor U13205 (N_13205,N_12775,N_12628);
or U13206 (N_13206,N_12668,N_12663);
and U13207 (N_13207,N_12636,N_12790);
nand U13208 (N_13208,N_12613,N_12519);
or U13209 (N_13209,N_12687,N_12574);
and U13210 (N_13210,N_12691,N_12709);
nand U13211 (N_13211,N_12651,N_12964);
xor U13212 (N_13212,N_12630,N_12607);
or U13213 (N_13213,N_12940,N_12744);
xnor U13214 (N_13214,N_12583,N_12848);
nand U13215 (N_13215,N_12682,N_12782);
xor U13216 (N_13216,N_12542,N_12858);
nand U13217 (N_13217,N_12826,N_12696);
nor U13218 (N_13218,N_12541,N_12951);
nand U13219 (N_13219,N_12559,N_12581);
nand U13220 (N_13220,N_12580,N_12887);
nand U13221 (N_13221,N_12626,N_12842);
nor U13222 (N_13222,N_12820,N_12585);
xor U13223 (N_13223,N_12567,N_12612);
xnor U13224 (N_13224,N_12863,N_12625);
nand U13225 (N_13225,N_12731,N_12952);
and U13226 (N_13226,N_12900,N_12905);
xnor U13227 (N_13227,N_12761,N_12960);
nand U13228 (N_13228,N_12783,N_12716);
or U13229 (N_13229,N_12827,N_12791);
nand U13230 (N_13230,N_12829,N_12985);
nand U13231 (N_13231,N_12979,N_12889);
or U13232 (N_13232,N_12947,N_12852);
nor U13233 (N_13233,N_12804,N_12692);
or U13234 (N_13234,N_12837,N_12645);
nor U13235 (N_13235,N_12831,N_12885);
xnor U13236 (N_13236,N_12818,N_12604);
and U13237 (N_13237,N_12929,N_12770);
or U13238 (N_13238,N_12658,N_12888);
or U13239 (N_13239,N_12523,N_12944);
nand U13240 (N_13240,N_12575,N_12764);
nor U13241 (N_13241,N_12871,N_12981);
xor U13242 (N_13242,N_12792,N_12711);
xnor U13243 (N_13243,N_12599,N_12664);
nand U13244 (N_13244,N_12823,N_12759);
nor U13245 (N_13245,N_12995,N_12997);
nor U13246 (N_13246,N_12899,N_12982);
and U13247 (N_13247,N_12807,N_12526);
nor U13248 (N_13248,N_12882,N_12847);
xnor U13249 (N_13249,N_12593,N_12928);
xor U13250 (N_13250,N_12678,N_12668);
and U13251 (N_13251,N_12880,N_12760);
xnor U13252 (N_13252,N_12755,N_12941);
or U13253 (N_13253,N_12684,N_12876);
nor U13254 (N_13254,N_12606,N_12623);
nor U13255 (N_13255,N_12746,N_12686);
and U13256 (N_13256,N_12637,N_12992);
nor U13257 (N_13257,N_12907,N_12582);
nor U13258 (N_13258,N_12542,N_12518);
or U13259 (N_13259,N_12816,N_12672);
or U13260 (N_13260,N_12787,N_12827);
xor U13261 (N_13261,N_12776,N_12699);
nand U13262 (N_13262,N_12552,N_12941);
xnor U13263 (N_13263,N_12927,N_12799);
xor U13264 (N_13264,N_12959,N_12543);
and U13265 (N_13265,N_12604,N_12971);
xor U13266 (N_13266,N_12623,N_12799);
xor U13267 (N_13267,N_12738,N_12610);
or U13268 (N_13268,N_12767,N_12895);
or U13269 (N_13269,N_12904,N_12529);
or U13270 (N_13270,N_12780,N_12876);
nand U13271 (N_13271,N_12773,N_12703);
and U13272 (N_13272,N_12547,N_12576);
nand U13273 (N_13273,N_12998,N_12995);
and U13274 (N_13274,N_12764,N_12622);
and U13275 (N_13275,N_12780,N_12593);
or U13276 (N_13276,N_12867,N_12709);
nand U13277 (N_13277,N_12967,N_12832);
nand U13278 (N_13278,N_12989,N_12757);
and U13279 (N_13279,N_12920,N_12827);
nand U13280 (N_13280,N_12783,N_12526);
or U13281 (N_13281,N_12681,N_12873);
xnor U13282 (N_13282,N_12855,N_12699);
nor U13283 (N_13283,N_12537,N_12763);
or U13284 (N_13284,N_12571,N_12848);
nand U13285 (N_13285,N_12793,N_12698);
xor U13286 (N_13286,N_12995,N_12746);
and U13287 (N_13287,N_12859,N_12916);
and U13288 (N_13288,N_12861,N_12798);
nand U13289 (N_13289,N_12648,N_12843);
nor U13290 (N_13290,N_12919,N_12518);
and U13291 (N_13291,N_12817,N_12500);
xor U13292 (N_13292,N_12539,N_12788);
or U13293 (N_13293,N_12858,N_12532);
nand U13294 (N_13294,N_12617,N_12722);
and U13295 (N_13295,N_12651,N_12617);
or U13296 (N_13296,N_12980,N_12845);
and U13297 (N_13297,N_12785,N_12513);
or U13298 (N_13298,N_12631,N_12832);
nand U13299 (N_13299,N_12958,N_12832);
or U13300 (N_13300,N_12609,N_12936);
nor U13301 (N_13301,N_12530,N_12925);
nor U13302 (N_13302,N_12511,N_12679);
nand U13303 (N_13303,N_12930,N_12929);
nand U13304 (N_13304,N_12702,N_12916);
nor U13305 (N_13305,N_12657,N_12662);
xnor U13306 (N_13306,N_12921,N_12996);
xor U13307 (N_13307,N_12819,N_12798);
nand U13308 (N_13308,N_12523,N_12981);
or U13309 (N_13309,N_12576,N_12758);
xnor U13310 (N_13310,N_12865,N_12979);
xor U13311 (N_13311,N_12787,N_12846);
or U13312 (N_13312,N_12600,N_12616);
nand U13313 (N_13313,N_12605,N_12610);
nand U13314 (N_13314,N_12550,N_12744);
and U13315 (N_13315,N_12808,N_12874);
or U13316 (N_13316,N_12988,N_12898);
nand U13317 (N_13317,N_12724,N_12729);
xnor U13318 (N_13318,N_12581,N_12743);
xor U13319 (N_13319,N_12843,N_12530);
xnor U13320 (N_13320,N_12767,N_12816);
xor U13321 (N_13321,N_12521,N_12765);
or U13322 (N_13322,N_12879,N_12896);
and U13323 (N_13323,N_12726,N_12571);
nand U13324 (N_13324,N_12654,N_12899);
xnor U13325 (N_13325,N_12770,N_12504);
xnor U13326 (N_13326,N_12506,N_12771);
and U13327 (N_13327,N_12935,N_12916);
nor U13328 (N_13328,N_12694,N_12568);
or U13329 (N_13329,N_12593,N_12879);
xor U13330 (N_13330,N_12584,N_12572);
and U13331 (N_13331,N_12840,N_12691);
and U13332 (N_13332,N_12579,N_12878);
or U13333 (N_13333,N_12671,N_12872);
nand U13334 (N_13334,N_12669,N_12792);
xnor U13335 (N_13335,N_12652,N_12859);
xor U13336 (N_13336,N_12560,N_12637);
xor U13337 (N_13337,N_12830,N_12526);
nor U13338 (N_13338,N_12738,N_12647);
nor U13339 (N_13339,N_12596,N_12921);
or U13340 (N_13340,N_12806,N_12843);
or U13341 (N_13341,N_12997,N_12594);
nor U13342 (N_13342,N_12781,N_12860);
nor U13343 (N_13343,N_12688,N_12657);
nand U13344 (N_13344,N_12946,N_12716);
nand U13345 (N_13345,N_12517,N_12936);
xnor U13346 (N_13346,N_12519,N_12753);
or U13347 (N_13347,N_12566,N_12697);
or U13348 (N_13348,N_12993,N_12925);
nor U13349 (N_13349,N_12684,N_12808);
xnor U13350 (N_13350,N_12919,N_12605);
nor U13351 (N_13351,N_12695,N_12550);
and U13352 (N_13352,N_12873,N_12657);
or U13353 (N_13353,N_12688,N_12735);
xor U13354 (N_13354,N_12714,N_12541);
or U13355 (N_13355,N_12929,N_12780);
or U13356 (N_13356,N_12737,N_12938);
or U13357 (N_13357,N_12729,N_12680);
xnor U13358 (N_13358,N_12621,N_12661);
xnor U13359 (N_13359,N_12809,N_12782);
nand U13360 (N_13360,N_12978,N_12826);
or U13361 (N_13361,N_12940,N_12585);
or U13362 (N_13362,N_12889,N_12544);
nor U13363 (N_13363,N_12933,N_12776);
or U13364 (N_13364,N_12649,N_12792);
nor U13365 (N_13365,N_12858,N_12752);
or U13366 (N_13366,N_12521,N_12692);
or U13367 (N_13367,N_12905,N_12756);
nor U13368 (N_13368,N_12691,N_12898);
and U13369 (N_13369,N_12699,N_12695);
or U13370 (N_13370,N_12583,N_12982);
nor U13371 (N_13371,N_12690,N_12522);
xnor U13372 (N_13372,N_12713,N_12652);
and U13373 (N_13373,N_12619,N_12775);
nor U13374 (N_13374,N_12624,N_12746);
nor U13375 (N_13375,N_12623,N_12994);
xor U13376 (N_13376,N_12663,N_12889);
nand U13377 (N_13377,N_12957,N_12970);
xnor U13378 (N_13378,N_12537,N_12699);
or U13379 (N_13379,N_12824,N_12706);
xor U13380 (N_13380,N_12511,N_12626);
or U13381 (N_13381,N_12988,N_12735);
or U13382 (N_13382,N_12783,N_12877);
xnor U13383 (N_13383,N_12852,N_12562);
xnor U13384 (N_13384,N_12842,N_12908);
nor U13385 (N_13385,N_12586,N_12514);
xor U13386 (N_13386,N_12961,N_12500);
xor U13387 (N_13387,N_12588,N_12522);
nand U13388 (N_13388,N_12928,N_12793);
nand U13389 (N_13389,N_12542,N_12952);
or U13390 (N_13390,N_12604,N_12607);
and U13391 (N_13391,N_12543,N_12818);
nor U13392 (N_13392,N_12664,N_12730);
or U13393 (N_13393,N_12755,N_12796);
nor U13394 (N_13394,N_12837,N_12506);
xnor U13395 (N_13395,N_12892,N_12502);
nor U13396 (N_13396,N_12697,N_12745);
and U13397 (N_13397,N_12929,N_12527);
or U13398 (N_13398,N_12814,N_12648);
or U13399 (N_13399,N_12894,N_12516);
nand U13400 (N_13400,N_12869,N_12804);
or U13401 (N_13401,N_12837,N_12919);
nand U13402 (N_13402,N_12827,N_12708);
nand U13403 (N_13403,N_12988,N_12635);
xor U13404 (N_13404,N_12651,N_12509);
nand U13405 (N_13405,N_12899,N_12636);
or U13406 (N_13406,N_12785,N_12930);
and U13407 (N_13407,N_12987,N_12859);
nand U13408 (N_13408,N_12785,N_12698);
nor U13409 (N_13409,N_12631,N_12728);
xor U13410 (N_13410,N_12708,N_12779);
xnor U13411 (N_13411,N_12509,N_12582);
xnor U13412 (N_13412,N_12731,N_12797);
nand U13413 (N_13413,N_12939,N_12888);
or U13414 (N_13414,N_12987,N_12649);
xor U13415 (N_13415,N_12579,N_12684);
or U13416 (N_13416,N_12646,N_12759);
and U13417 (N_13417,N_12779,N_12525);
and U13418 (N_13418,N_12939,N_12771);
or U13419 (N_13419,N_12745,N_12849);
nand U13420 (N_13420,N_12876,N_12662);
or U13421 (N_13421,N_12985,N_12629);
and U13422 (N_13422,N_12890,N_12773);
xor U13423 (N_13423,N_12706,N_12797);
or U13424 (N_13424,N_12545,N_12935);
and U13425 (N_13425,N_12762,N_12849);
nor U13426 (N_13426,N_12983,N_12982);
or U13427 (N_13427,N_12975,N_12796);
and U13428 (N_13428,N_12753,N_12646);
xnor U13429 (N_13429,N_12537,N_12847);
and U13430 (N_13430,N_12977,N_12708);
nand U13431 (N_13431,N_12859,N_12815);
nor U13432 (N_13432,N_12536,N_12807);
or U13433 (N_13433,N_12986,N_12898);
xor U13434 (N_13434,N_12980,N_12549);
xor U13435 (N_13435,N_12552,N_12734);
nand U13436 (N_13436,N_12799,N_12585);
nor U13437 (N_13437,N_12627,N_12681);
xnor U13438 (N_13438,N_12539,N_12508);
nor U13439 (N_13439,N_12750,N_12679);
and U13440 (N_13440,N_12650,N_12503);
nand U13441 (N_13441,N_12909,N_12530);
nand U13442 (N_13442,N_12888,N_12559);
xnor U13443 (N_13443,N_12846,N_12877);
and U13444 (N_13444,N_12642,N_12842);
and U13445 (N_13445,N_12582,N_12610);
xnor U13446 (N_13446,N_12911,N_12636);
or U13447 (N_13447,N_12966,N_12939);
and U13448 (N_13448,N_12923,N_12875);
and U13449 (N_13449,N_12724,N_12772);
xnor U13450 (N_13450,N_12991,N_12742);
nand U13451 (N_13451,N_12726,N_12588);
nand U13452 (N_13452,N_12775,N_12575);
nand U13453 (N_13453,N_12728,N_12990);
xor U13454 (N_13454,N_12685,N_12545);
or U13455 (N_13455,N_12918,N_12549);
xnor U13456 (N_13456,N_12875,N_12570);
xnor U13457 (N_13457,N_12898,N_12794);
xnor U13458 (N_13458,N_12786,N_12526);
xnor U13459 (N_13459,N_12700,N_12704);
or U13460 (N_13460,N_12634,N_12724);
and U13461 (N_13461,N_12663,N_12807);
nand U13462 (N_13462,N_12654,N_12979);
or U13463 (N_13463,N_12995,N_12931);
and U13464 (N_13464,N_12830,N_12977);
nand U13465 (N_13465,N_12591,N_12659);
nor U13466 (N_13466,N_12672,N_12984);
xnor U13467 (N_13467,N_12956,N_12980);
xor U13468 (N_13468,N_12758,N_12788);
xor U13469 (N_13469,N_12702,N_12597);
nor U13470 (N_13470,N_12922,N_12520);
nand U13471 (N_13471,N_12649,N_12816);
nor U13472 (N_13472,N_12954,N_12616);
and U13473 (N_13473,N_12542,N_12560);
or U13474 (N_13474,N_12900,N_12681);
nand U13475 (N_13475,N_12676,N_12528);
and U13476 (N_13476,N_12709,N_12974);
xnor U13477 (N_13477,N_12818,N_12643);
or U13478 (N_13478,N_12863,N_12590);
xor U13479 (N_13479,N_12515,N_12959);
and U13480 (N_13480,N_12522,N_12815);
and U13481 (N_13481,N_12876,N_12619);
xor U13482 (N_13482,N_12996,N_12529);
nand U13483 (N_13483,N_12949,N_12985);
or U13484 (N_13484,N_12687,N_12589);
nor U13485 (N_13485,N_12802,N_12882);
nor U13486 (N_13486,N_12652,N_12921);
and U13487 (N_13487,N_12599,N_12594);
and U13488 (N_13488,N_12734,N_12674);
or U13489 (N_13489,N_12535,N_12908);
or U13490 (N_13490,N_12928,N_12837);
or U13491 (N_13491,N_12580,N_12864);
and U13492 (N_13492,N_12515,N_12953);
nand U13493 (N_13493,N_12907,N_12776);
xnor U13494 (N_13494,N_12936,N_12550);
xnor U13495 (N_13495,N_12826,N_12609);
and U13496 (N_13496,N_12873,N_12976);
nand U13497 (N_13497,N_12789,N_12652);
xor U13498 (N_13498,N_12662,N_12916);
and U13499 (N_13499,N_12889,N_12634);
xnor U13500 (N_13500,N_13205,N_13480);
nor U13501 (N_13501,N_13276,N_13283);
or U13502 (N_13502,N_13377,N_13415);
nand U13503 (N_13503,N_13040,N_13340);
nand U13504 (N_13504,N_13211,N_13179);
or U13505 (N_13505,N_13168,N_13101);
nand U13506 (N_13506,N_13417,N_13486);
xnor U13507 (N_13507,N_13331,N_13430);
nor U13508 (N_13508,N_13212,N_13232);
and U13509 (N_13509,N_13127,N_13363);
or U13510 (N_13510,N_13344,N_13152);
and U13511 (N_13511,N_13467,N_13375);
or U13512 (N_13512,N_13056,N_13013);
or U13513 (N_13513,N_13139,N_13045);
and U13514 (N_13514,N_13450,N_13145);
nand U13515 (N_13515,N_13370,N_13449);
nand U13516 (N_13516,N_13104,N_13064);
nand U13517 (N_13517,N_13437,N_13435);
or U13518 (N_13518,N_13014,N_13030);
nor U13519 (N_13519,N_13359,N_13003);
nand U13520 (N_13520,N_13349,N_13452);
nand U13521 (N_13521,N_13345,N_13106);
nor U13522 (N_13522,N_13258,N_13111);
or U13523 (N_13523,N_13220,N_13381);
nor U13524 (N_13524,N_13095,N_13343);
nand U13525 (N_13525,N_13119,N_13260);
xor U13526 (N_13526,N_13376,N_13184);
nor U13527 (N_13527,N_13029,N_13275);
xnor U13528 (N_13528,N_13075,N_13138);
nor U13529 (N_13529,N_13112,N_13265);
and U13530 (N_13530,N_13102,N_13140);
nand U13531 (N_13531,N_13099,N_13218);
or U13532 (N_13532,N_13327,N_13170);
nand U13533 (N_13533,N_13188,N_13114);
xnor U13534 (N_13534,N_13100,N_13169);
nand U13535 (N_13535,N_13289,N_13433);
and U13536 (N_13536,N_13019,N_13317);
or U13537 (N_13537,N_13465,N_13154);
nor U13538 (N_13538,N_13118,N_13403);
nand U13539 (N_13539,N_13052,N_13354);
and U13540 (N_13540,N_13439,N_13028);
nand U13541 (N_13541,N_13132,N_13294);
xor U13542 (N_13542,N_13455,N_13459);
or U13543 (N_13543,N_13297,N_13053);
or U13544 (N_13544,N_13046,N_13478);
and U13545 (N_13545,N_13269,N_13057);
nand U13546 (N_13546,N_13235,N_13284);
nand U13547 (N_13547,N_13068,N_13213);
xor U13548 (N_13548,N_13307,N_13155);
nand U13549 (N_13549,N_13059,N_13316);
xor U13550 (N_13550,N_13157,N_13191);
nand U13551 (N_13551,N_13248,N_13308);
nand U13552 (N_13552,N_13388,N_13219);
xor U13553 (N_13553,N_13079,N_13458);
and U13554 (N_13554,N_13035,N_13183);
and U13555 (N_13555,N_13251,N_13339);
xnor U13556 (N_13556,N_13356,N_13051);
or U13557 (N_13557,N_13350,N_13087);
nand U13558 (N_13558,N_13399,N_13338);
or U13559 (N_13559,N_13278,N_13429);
and U13560 (N_13560,N_13049,N_13266);
nand U13561 (N_13561,N_13018,N_13025);
xnor U13562 (N_13562,N_13004,N_13328);
nor U13563 (N_13563,N_13368,N_13195);
and U13564 (N_13564,N_13481,N_13009);
and U13565 (N_13565,N_13136,N_13400);
nand U13566 (N_13566,N_13390,N_13158);
xnor U13567 (N_13567,N_13364,N_13162);
xor U13568 (N_13568,N_13134,N_13475);
xor U13569 (N_13569,N_13161,N_13373);
xnor U13570 (N_13570,N_13225,N_13245);
or U13571 (N_13571,N_13207,N_13182);
xnor U13572 (N_13572,N_13011,N_13393);
and U13573 (N_13573,N_13401,N_13330);
and U13574 (N_13574,N_13304,N_13063);
xnor U13575 (N_13575,N_13259,N_13187);
nand U13576 (N_13576,N_13228,N_13446);
xor U13577 (N_13577,N_13466,N_13074);
or U13578 (N_13578,N_13434,N_13443);
nand U13579 (N_13579,N_13082,N_13243);
or U13580 (N_13580,N_13312,N_13414);
and U13581 (N_13581,N_13410,N_13124);
and U13582 (N_13582,N_13357,N_13027);
nor U13583 (N_13583,N_13066,N_13423);
xor U13584 (N_13584,N_13402,N_13242);
nand U13585 (N_13585,N_13409,N_13424);
and U13586 (N_13586,N_13367,N_13285);
or U13587 (N_13587,N_13442,N_13073);
or U13588 (N_13588,N_13214,N_13165);
nand U13589 (N_13589,N_13016,N_13203);
and U13590 (N_13590,N_13432,N_13351);
nor U13591 (N_13591,N_13060,N_13230);
xnor U13592 (N_13592,N_13078,N_13039);
nor U13593 (N_13593,N_13389,N_13058);
or U13594 (N_13594,N_13324,N_13451);
nand U13595 (N_13595,N_13034,N_13148);
nand U13596 (N_13596,N_13067,N_13055);
xor U13597 (N_13597,N_13084,N_13318);
nand U13598 (N_13598,N_13361,N_13071);
xor U13599 (N_13599,N_13091,N_13426);
xor U13600 (N_13600,N_13301,N_13204);
and U13601 (N_13601,N_13453,N_13186);
nor U13602 (N_13602,N_13441,N_13386);
nor U13603 (N_13603,N_13236,N_13109);
nand U13604 (N_13604,N_13076,N_13135);
nor U13605 (N_13605,N_13210,N_13250);
or U13606 (N_13606,N_13180,N_13295);
xor U13607 (N_13607,N_13024,N_13116);
xor U13608 (N_13608,N_13348,N_13305);
or U13609 (N_13609,N_13280,N_13252);
xor U13610 (N_13610,N_13031,N_13302);
or U13611 (N_13611,N_13108,N_13226);
and U13612 (N_13612,N_13319,N_13037);
and U13613 (N_13613,N_13271,N_13394);
xor U13614 (N_13614,N_13476,N_13153);
xor U13615 (N_13615,N_13290,N_13227);
and U13616 (N_13616,N_13038,N_13143);
or U13617 (N_13617,N_13445,N_13436);
or U13618 (N_13618,N_13425,N_13048);
or U13619 (N_13619,N_13103,N_13181);
nand U13620 (N_13620,N_13217,N_13264);
or U13621 (N_13621,N_13342,N_13485);
or U13622 (N_13622,N_13257,N_13065);
xor U13623 (N_13623,N_13070,N_13144);
nand U13624 (N_13624,N_13096,N_13173);
or U13625 (N_13625,N_13496,N_13438);
and U13626 (N_13626,N_13199,N_13137);
and U13627 (N_13627,N_13223,N_13092);
xnor U13628 (N_13628,N_13147,N_13471);
nand U13629 (N_13629,N_13385,N_13042);
and U13630 (N_13630,N_13347,N_13404);
nand U13631 (N_13631,N_13279,N_13151);
or U13632 (N_13632,N_13020,N_13499);
nand U13633 (N_13633,N_13282,N_13296);
and U13634 (N_13634,N_13237,N_13202);
xor U13635 (N_13635,N_13081,N_13416);
and U13636 (N_13636,N_13088,N_13315);
nor U13637 (N_13637,N_13298,N_13130);
nand U13638 (N_13638,N_13120,N_13474);
or U13639 (N_13639,N_13365,N_13291);
or U13640 (N_13640,N_13167,N_13050);
nand U13641 (N_13641,N_13387,N_13461);
and U13642 (N_13642,N_13456,N_13083);
xnor U13643 (N_13643,N_13352,N_13177);
or U13644 (N_13644,N_13372,N_13469);
nand U13645 (N_13645,N_13125,N_13273);
and U13646 (N_13646,N_13470,N_13497);
nand U13647 (N_13647,N_13277,N_13335);
xor U13648 (N_13648,N_13263,N_13208);
or U13649 (N_13649,N_13371,N_13159);
nand U13650 (N_13650,N_13249,N_13491);
and U13651 (N_13651,N_13479,N_13326);
xor U13652 (N_13652,N_13054,N_13353);
xnor U13653 (N_13653,N_13128,N_13041);
xnor U13654 (N_13654,N_13380,N_13336);
or U13655 (N_13655,N_13231,N_13200);
xnor U13656 (N_13656,N_13411,N_13008);
xnor U13657 (N_13657,N_13369,N_13407);
nor U13658 (N_13658,N_13396,N_13010);
or U13659 (N_13659,N_13239,N_13460);
xor U13660 (N_13660,N_13493,N_13093);
or U13661 (N_13661,N_13448,N_13012);
xor U13662 (N_13662,N_13314,N_13378);
or U13663 (N_13663,N_13309,N_13192);
and U13664 (N_13664,N_13440,N_13420);
and U13665 (N_13665,N_13172,N_13487);
or U13666 (N_13666,N_13062,N_13254);
or U13667 (N_13667,N_13146,N_13270);
xor U13668 (N_13668,N_13141,N_13366);
nor U13669 (N_13669,N_13406,N_13215);
and U13670 (N_13670,N_13043,N_13001);
nor U13671 (N_13671,N_13241,N_13412);
and U13672 (N_13672,N_13395,N_13150);
xor U13673 (N_13673,N_13117,N_13121);
xor U13674 (N_13674,N_13299,N_13334);
nor U13675 (N_13675,N_13176,N_13189);
nand U13676 (N_13676,N_13198,N_13490);
nand U13677 (N_13677,N_13178,N_13321);
nor U13678 (N_13678,N_13457,N_13379);
or U13679 (N_13679,N_13268,N_13427);
and U13680 (N_13680,N_13171,N_13454);
nand U13681 (N_13681,N_13355,N_13281);
or U13682 (N_13682,N_13149,N_13222);
xor U13683 (N_13683,N_13422,N_13122);
nand U13684 (N_13684,N_13287,N_13293);
nor U13685 (N_13685,N_13240,N_13384);
xnor U13686 (N_13686,N_13383,N_13494);
nor U13687 (N_13687,N_13473,N_13026);
xor U13688 (N_13688,N_13462,N_13126);
nand U13689 (N_13689,N_13175,N_13300);
or U13690 (N_13690,N_13392,N_13320);
xor U13691 (N_13691,N_13274,N_13272);
nand U13692 (N_13692,N_13174,N_13129);
or U13693 (N_13693,N_13061,N_13498);
nor U13694 (N_13694,N_13123,N_13142);
or U13695 (N_13695,N_13492,N_13488);
and U13696 (N_13696,N_13197,N_13472);
nand U13697 (N_13697,N_13089,N_13005);
or U13698 (N_13698,N_13382,N_13164);
and U13699 (N_13699,N_13463,N_13397);
nand U13700 (N_13700,N_13329,N_13015);
nand U13701 (N_13701,N_13358,N_13253);
nor U13702 (N_13702,N_13484,N_13224);
or U13703 (N_13703,N_13477,N_13482);
nand U13704 (N_13704,N_13190,N_13021);
and U13705 (N_13705,N_13072,N_13085);
xor U13706 (N_13706,N_13194,N_13238);
and U13707 (N_13707,N_13495,N_13292);
nand U13708 (N_13708,N_13206,N_13080);
or U13709 (N_13709,N_13323,N_13255);
nor U13710 (N_13710,N_13261,N_13325);
nand U13711 (N_13711,N_13047,N_13032);
and U13712 (N_13712,N_13362,N_13247);
xor U13713 (N_13713,N_13110,N_13086);
or U13714 (N_13714,N_13007,N_13000);
or U13715 (N_13715,N_13421,N_13303);
or U13716 (N_13716,N_13069,N_13131);
nor U13717 (N_13717,N_13017,N_13023);
xnor U13718 (N_13718,N_13156,N_13288);
or U13719 (N_13719,N_13209,N_13405);
xor U13720 (N_13720,N_13036,N_13160);
xor U13721 (N_13721,N_13374,N_13105);
or U13722 (N_13722,N_13113,N_13094);
xor U13723 (N_13723,N_13002,N_13185);
nor U13724 (N_13724,N_13332,N_13391);
nand U13725 (N_13725,N_13166,N_13107);
or U13726 (N_13726,N_13246,N_13115);
nor U13727 (N_13727,N_13464,N_13090);
nor U13728 (N_13728,N_13311,N_13483);
and U13729 (N_13729,N_13337,N_13077);
or U13730 (N_13730,N_13444,N_13333);
and U13731 (N_13731,N_13408,N_13163);
xor U13732 (N_13732,N_13098,N_13256);
nor U13733 (N_13733,N_13413,N_13286);
or U13734 (N_13734,N_13196,N_13419);
nor U13735 (N_13735,N_13346,N_13360);
nand U13736 (N_13736,N_13044,N_13097);
xor U13737 (N_13737,N_13033,N_13428);
nand U13738 (N_13738,N_13313,N_13322);
or U13739 (N_13739,N_13489,N_13234);
or U13740 (N_13740,N_13262,N_13306);
xor U13741 (N_13741,N_13310,N_13006);
or U13742 (N_13742,N_13244,N_13233);
nand U13743 (N_13743,N_13229,N_13216);
or U13744 (N_13744,N_13193,N_13431);
and U13745 (N_13745,N_13398,N_13201);
and U13746 (N_13746,N_13221,N_13133);
xnor U13747 (N_13747,N_13022,N_13267);
or U13748 (N_13748,N_13341,N_13447);
or U13749 (N_13749,N_13418,N_13468);
xnor U13750 (N_13750,N_13266,N_13240);
or U13751 (N_13751,N_13490,N_13390);
nand U13752 (N_13752,N_13346,N_13344);
and U13753 (N_13753,N_13492,N_13236);
nand U13754 (N_13754,N_13277,N_13230);
nand U13755 (N_13755,N_13198,N_13491);
or U13756 (N_13756,N_13026,N_13402);
nand U13757 (N_13757,N_13486,N_13092);
and U13758 (N_13758,N_13491,N_13373);
and U13759 (N_13759,N_13271,N_13257);
nor U13760 (N_13760,N_13232,N_13145);
nor U13761 (N_13761,N_13005,N_13213);
nand U13762 (N_13762,N_13010,N_13431);
xor U13763 (N_13763,N_13173,N_13175);
nor U13764 (N_13764,N_13024,N_13336);
xnor U13765 (N_13765,N_13356,N_13111);
xor U13766 (N_13766,N_13057,N_13415);
and U13767 (N_13767,N_13058,N_13129);
nor U13768 (N_13768,N_13168,N_13154);
nor U13769 (N_13769,N_13316,N_13071);
and U13770 (N_13770,N_13125,N_13025);
or U13771 (N_13771,N_13313,N_13393);
or U13772 (N_13772,N_13194,N_13497);
and U13773 (N_13773,N_13412,N_13116);
or U13774 (N_13774,N_13429,N_13105);
or U13775 (N_13775,N_13144,N_13013);
and U13776 (N_13776,N_13323,N_13049);
nor U13777 (N_13777,N_13479,N_13341);
or U13778 (N_13778,N_13447,N_13252);
xnor U13779 (N_13779,N_13246,N_13251);
xnor U13780 (N_13780,N_13248,N_13162);
xnor U13781 (N_13781,N_13325,N_13276);
xnor U13782 (N_13782,N_13251,N_13119);
nor U13783 (N_13783,N_13464,N_13022);
nor U13784 (N_13784,N_13176,N_13152);
nand U13785 (N_13785,N_13206,N_13454);
nand U13786 (N_13786,N_13105,N_13446);
nand U13787 (N_13787,N_13365,N_13342);
xor U13788 (N_13788,N_13472,N_13296);
and U13789 (N_13789,N_13252,N_13291);
nand U13790 (N_13790,N_13209,N_13292);
xnor U13791 (N_13791,N_13362,N_13344);
or U13792 (N_13792,N_13010,N_13341);
or U13793 (N_13793,N_13136,N_13046);
nor U13794 (N_13794,N_13023,N_13239);
and U13795 (N_13795,N_13045,N_13407);
nor U13796 (N_13796,N_13058,N_13423);
or U13797 (N_13797,N_13036,N_13019);
xor U13798 (N_13798,N_13023,N_13356);
nor U13799 (N_13799,N_13366,N_13100);
nor U13800 (N_13800,N_13117,N_13194);
and U13801 (N_13801,N_13372,N_13438);
nor U13802 (N_13802,N_13029,N_13136);
nor U13803 (N_13803,N_13091,N_13071);
or U13804 (N_13804,N_13439,N_13280);
and U13805 (N_13805,N_13294,N_13166);
nor U13806 (N_13806,N_13251,N_13384);
nand U13807 (N_13807,N_13422,N_13214);
and U13808 (N_13808,N_13313,N_13287);
or U13809 (N_13809,N_13403,N_13265);
and U13810 (N_13810,N_13077,N_13446);
xor U13811 (N_13811,N_13050,N_13424);
or U13812 (N_13812,N_13418,N_13004);
xnor U13813 (N_13813,N_13363,N_13068);
or U13814 (N_13814,N_13061,N_13065);
or U13815 (N_13815,N_13124,N_13054);
xor U13816 (N_13816,N_13287,N_13107);
nand U13817 (N_13817,N_13272,N_13408);
and U13818 (N_13818,N_13474,N_13183);
xor U13819 (N_13819,N_13081,N_13402);
nor U13820 (N_13820,N_13120,N_13428);
or U13821 (N_13821,N_13136,N_13211);
nand U13822 (N_13822,N_13435,N_13387);
nor U13823 (N_13823,N_13141,N_13055);
or U13824 (N_13824,N_13372,N_13308);
and U13825 (N_13825,N_13019,N_13292);
xnor U13826 (N_13826,N_13183,N_13216);
and U13827 (N_13827,N_13407,N_13324);
xor U13828 (N_13828,N_13450,N_13132);
nor U13829 (N_13829,N_13101,N_13023);
nor U13830 (N_13830,N_13018,N_13002);
nor U13831 (N_13831,N_13039,N_13217);
xnor U13832 (N_13832,N_13295,N_13479);
nor U13833 (N_13833,N_13392,N_13081);
and U13834 (N_13834,N_13016,N_13032);
and U13835 (N_13835,N_13440,N_13180);
nand U13836 (N_13836,N_13068,N_13029);
or U13837 (N_13837,N_13039,N_13124);
xor U13838 (N_13838,N_13267,N_13290);
nand U13839 (N_13839,N_13174,N_13456);
nand U13840 (N_13840,N_13250,N_13311);
nand U13841 (N_13841,N_13256,N_13169);
xor U13842 (N_13842,N_13277,N_13002);
and U13843 (N_13843,N_13233,N_13372);
xor U13844 (N_13844,N_13198,N_13178);
and U13845 (N_13845,N_13172,N_13221);
nor U13846 (N_13846,N_13258,N_13195);
nor U13847 (N_13847,N_13216,N_13303);
nor U13848 (N_13848,N_13365,N_13429);
xnor U13849 (N_13849,N_13268,N_13279);
xor U13850 (N_13850,N_13293,N_13402);
and U13851 (N_13851,N_13304,N_13412);
or U13852 (N_13852,N_13359,N_13252);
nand U13853 (N_13853,N_13077,N_13280);
xor U13854 (N_13854,N_13112,N_13340);
nand U13855 (N_13855,N_13243,N_13284);
and U13856 (N_13856,N_13426,N_13153);
xnor U13857 (N_13857,N_13240,N_13391);
nor U13858 (N_13858,N_13474,N_13171);
nor U13859 (N_13859,N_13140,N_13291);
or U13860 (N_13860,N_13405,N_13023);
and U13861 (N_13861,N_13398,N_13229);
nor U13862 (N_13862,N_13390,N_13423);
xnor U13863 (N_13863,N_13093,N_13016);
and U13864 (N_13864,N_13284,N_13391);
xnor U13865 (N_13865,N_13312,N_13140);
and U13866 (N_13866,N_13075,N_13340);
or U13867 (N_13867,N_13018,N_13001);
nand U13868 (N_13868,N_13303,N_13178);
nor U13869 (N_13869,N_13372,N_13217);
nor U13870 (N_13870,N_13401,N_13131);
nand U13871 (N_13871,N_13330,N_13059);
or U13872 (N_13872,N_13375,N_13324);
nand U13873 (N_13873,N_13486,N_13238);
or U13874 (N_13874,N_13071,N_13428);
and U13875 (N_13875,N_13055,N_13015);
nor U13876 (N_13876,N_13227,N_13368);
nor U13877 (N_13877,N_13158,N_13254);
nand U13878 (N_13878,N_13179,N_13445);
nand U13879 (N_13879,N_13499,N_13247);
nand U13880 (N_13880,N_13401,N_13495);
or U13881 (N_13881,N_13092,N_13226);
nand U13882 (N_13882,N_13380,N_13243);
xor U13883 (N_13883,N_13054,N_13310);
xor U13884 (N_13884,N_13186,N_13020);
nand U13885 (N_13885,N_13320,N_13208);
or U13886 (N_13886,N_13381,N_13087);
nor U13887 (N_13887,N_13010,N_13452);
nand U13888 (N_13888,N_13492,N_13341);
nor U13889 (N_13889,N_13394,N_13230);
nand U13890 (N_13890,N_13175,N_13397);
nor U13891 (N_13891,N_13321,N_13370);
nand U13892 (N_13892,N_13026,N_13421);
nand U13893 (N_13893,N_13407,N_13235);
xor U13894 (N_13894,N_13240,N_13261);
nor U13895 (N_13895,N_13295,N_13422);
xnor U13896 (N_13896,N_13242,N_13321);
and U13897 (N_13897,N_13093,N_13090);
nand U13898 (N_13898,N_13273,N_13165);
or U13899 (N_13899,N_13013,N_13499);
nand U13900 (N_13900,N_13344,N_13123);
nor U13901 (N_13901,N_13347,N_13117);
nand U13902 (N_13902,N_13412,N_13118);
and U13903 (N_13903,N_13196,N_13036);
nor U13904 (N_13904,N_13331,N_13043);
and U13905 (N_13905,N_13023,N_13316);
xor U13906 (N_13906,N_13404,N_13167);
or U13907 (N_13907,N_13350,N_13251);
xnor U13908 (N_13908,N_13377,N_13291);
xor U13909 (N_13909,N_13464,N_13232);
nand U13910 (N_13910,N_13004,N_13445);
or U13911 (N_13911,N_13155,N_13011);
nand U13912 (N_13912,N_13427,N_13318);
or U13913 (N_13913,N_13319,N_13428);
xor U13914 (N_13914,N_13382,N_13051);
or U13915 (N_13915,N_13136,N_13397);
and U13916 (N_13916,N_13007,N_13190);
or U13917 (N_13917,N_13106,N_13038);
or U13918 (N_13918,N_13361,N_13375);
xor U13919 (N_13919,N_13225,N_13002);
xnor U13920 (N_13920,N_13393,N_13316);
or U13921 (N_13921,N_13194,N_13147);
nor U13922 (N_13922,N_13252,N_13256);
nor U13923 (N_13923,N_13443,N_13473);
nor U13924 (N_13924,N_13204,N_13131);
or U13925 (N_13925,N_13411,N_13391);
and U13926 (N_13926,N_13037,N_13303);
xnor U13927 (N_13927,N_13086,N_13361);
nor U13928 (N_13928,N_13224,N_13086);
and U13929 (N_13929,N_13175,N_13197);
and U13930 (N_13930,N_13181,N_13190);
xor U13931 (N_13931,N_13054,N_13414);
nand U13932 (N_13932,N_13101,N_13404);
and U13933 (N_13933,N_13124,N_13268);
and U13934 (N_13934,N_13224,N_13178);
nand U13935 (N_13935,N_13349,N_13473);
and U13936 (N_13936,N_13211,N_13026);
nand U13937 (N_13937,N_13103,N_13320);
and U13938 (N_13938,N_13302,N_13464);
nand U13939 (N_13939,N_13143,N_13257);
xor U13940 (N_13940,N_13108,N_13203);
nor U13941 (N_13941,N_13246,N_13320);
nor U13942 (N_13942,N_13280,N_13090);
and U13943 (N_13943,N_13305,N_13105);
or U13944 (N_13944,N_13477,N_13064);
nand U13945 (N_13945,N_13105,N_13017);
and U13946 (N_13946,N_13428,N_13301);
nand U13947 (N_13947,N_13466,N_13327);
or U13948 (N_13948,N_13367,N_13397);
nand U13949 (N_13949,N_13351,N_13264);
nand U13950 (N_13950,N_13189,N_13204);
nand U13951 (N_13951,N_13386,N_13382);
nand U13952 (N_13952,N_13188,N_13264);
xor U13953 (N_13953,N_13234,N_13367);
nor U13954 (N_13954,N_13247,N_13386);
xor U13955 (N_13955,N_13391,N_13131);
xor U13956 (N_13956,N_13196,N_13475);
xor U13957 (N_13957,N_13030,N_13117);
nand U13958 (N_13958,N_13206,N_13271);
nor U13959 (N_13959,N_13208,N_13118);
nand U13960 (N_13960,N_13017,N_13039);
nor U13961 (N_13961,N_13364,N_13400);
and U13962 (N_13962,N_13311,N_13027);
nand U13963 (N_13963,N_13077,N_13318);
or U13964 (N_13964,N_13480,N_13272);
or U13965 (N_13965,N_13258,N_13468);
nand U13966 (N_13966,N_13439,N_13139);
and U13967 (N_13967,N_13430,N_13090);
or U13968 (N_13968,N_13442,N_13207);
or U13969 (N_13969,N_13169,N_13128);
nand U13970 (N_13970,N_13087,N_13201);
xnor U13971 (N_13971,N_13428,N_13365);
nor U13972 (N_13972,N_13247,N_13489);
or U13973 (N_13973,N_13367,N_13100);
nand U13974 (N_13974,N_13162,N_13040);
nand U13975 (N_13975,N_13274,N_13458);
and U13976 (N_13976,N_13136,N_13155);
nand U13977 (N_13977,N_13051,N_13178);
nor U13978 (N_13978,N_13244,N_13089);
or U13979 (N_13979,N_13274,N_13208);
nor U13980 (N_13980,N_13092,N_13068);
or U13981 (N_13981,N_13273,N_13190);
xor U13982 (N_13982,N_13314,N_13170);
or U13983 (N_13983,N_13451,N_13222);
xor U13984 (N_13984,N_13000,N_13114);
nand U13985 (N_13985,N_13068,N_13462);
xor U13986 (N_13986,N_13499,N_13156);
and U13987 (N_13987,N_13231,N_13334);
xor U13988 (N_13988,N_13031,N_13076);
xnor U13989 (N_13989,N_13290,N_13498);
nand U13990 (N_13990,N_13348,N_13451);
or U13991 (N_13991,N_13226,N_13029);
or U13992 (N_13992,N_13153,N_13129);
and U13993 (N_13993,N_13395,N_13128);
nand U13994 (N_13994,N_13225,N_13350);
xor U13995 (N_13995,N_13142,N_13278);
nand U13996 (N_13996,N_13448,N_13259);
nand U13997 (N_13997,N_13229,N_13377);
nand U13998 (N_13998,N_13129,N_13266);
or U13999 (N_13999,N_13224,N_13284);
and U14000 (N_14000,N_13518,N_13898);
nor U14001 (N_14001,N_13923,N_13896);
and U14002 (N_14002,N_13734,N_13796);
xnor U14003 (N_14003,N_13968,N_13885);
nand U14004 (N_14004,N_13823,N_13826);
nor U14005 (N_14005,N_13756,N_13805);
or U14006 (N_14006,N_13612,N_13937);
and U14007 (N_14007,N_13830,N_13754);
nand U14008 (N_14008,N_13800,N_13666);
nor U14009 (N_14009,N_13525,N_13955);
and U14010 (N_14010,N_13960,N_13654);
and U14011 (N_14011,N_13752,N_13635);
or U14012 (N_14012,N_13982,N_13636);
and U14013 (N_14013,N_13711,N_13630);
xor U14014 (N_14014,N_13869,N_13907);
xnor U14015 (N_14015,N_13879,N_13639);
nand U14016 (N_14016,N_13777,N_13884);
xnor U14017 (N_14017,N_13638,N_13994);
nand U14018 (N_14018,N_13645,N_13615);
nor U14019 (N_14019,N_13978,N_13716);
nand U14020 (N_14020,N_13552,N_13780);
or U14021 (N_14021,N_13958,N_13748);
nor U14022 (N_14022,N_13905,N_13784);
or U14023 (N_14023,N_13587,N_13585);
nor U14024 (N_14024,N_13562,N_13741);
xnor U14025 (N_14025,N_13505,N_13837);
and U14026 (N_14026,N_13701,N_13914);
nor U14027 (N_14027,N_13875,N_13502);
xnor U14028 (N_14028,N_13992,N_13738);
or U14029 (N_14029,N_13825,N_13529);
or U14030 (N_14030,N_13678,N_13928);
nor U14031 (N_14031,N_13922,N_13693);
xor U14032 (N_14032,N_13990,N_13582);
nor U14033 (N_14033,N_13974,N_13783);
xnor U14034 (N_14034,N_13705,N_13713);
or U14035 (N_14035,N_13633,N_13593);
or U14036 (N_14036,N_13927,N_13657);
nor U14037 (N_14037,N_13785,N_13662);
xor U14038 (N_14038,N_13653,N_13604);
or U14039 (N_14039,N_13833,N_13983);
or U14040 (N_14040,N_13817,N_13915);
nor U14041 (N_14041,N_13570,N_13806);
or U14042 (N_14042,N_13808,N_13700);
xor U14043 (N_14043,N_13999,N_13569);
nor U14044 (N_14044,N_13803,N_13841);
nor U14045 (N_14045,N_13829,N_13963);
nor U14046 (N_14046,N_13913,N_13849);
nor U14047 (N_14047,N_13957,N_13682);
or U14048 (N_14048,N_13984,N_13945);
nand U14049 (N_14049,N_13961,N_13673);
nand U14050 (N_14050,N_13820,N_13627);
nand U14051 (N_14051,N_13846,N_13672);
or U14052 (N_14052,N_13522,N_13563);
nand U14053 (N_14053,N_13819,N_13669);
or U14054 (N_14054,N_13768,N_13954);
nor U14055 (N_14055,N_13942,N_13643);
nor U14056 (N_14056,N_13815,N_13707);
xor U14057 (N_14057,N_13576,N_13967);
nand U14058 (N_14058,N_13509,N_13719);
and U14059 (N_14059,N_13772,N_13890);
nand U14060 (N_14060,N_13517,N_13532);
or U14061 (N_14061,N_13684,N_13926);
xnor U14062 (N_14062,N_13641,N_13521);
or U14063 (N_14063,N_13583,N_13610);
xor U14064 (N_14064,N_13949,N_13544);
nand U14065 (N_14065,N_13631,N_13918);
and U14066 (N_14066,N_13564,N_13753);
or U14067 (N_14067,N_13924,N_13989);
and U14068 (N_14068,N_13947,N_13845);
xor U14069 (N_14069,N_13658,N_13725);
nor U14070 (N_14070,N_13867,N_13606);
or U14071 (N_14071,N_13788,N_13721);
and U14072 (N_14072,N_13795,N_13647);
or U14073 (N_14073,N_13834,N_13870);
and U14074 (N_14074,N_13577,N_13733);
nor U14075 (N_14075,N_13860,N_13740);
or U14076 (N_14076,N_13852,N_13911);
xnor U14077 (N_14077,N_13687,N_13547);
and U14078 (N_14078,N_13728,N_13650);
and U14079 (N_14079,N_13797,N_13746);
nor U14080 (N_14080,N_13702,N_13977);
and U14081 (N_14081,N_13871,N_13973);
nor U14082 (N_14082,N_13946,N_13995);
and U14083 (N_14083,N_13765,N_13644);
nor U14084 (N_14084,N_13932,N_13877);
nor U14085 (N_14085,N_13730,N_13514);
or U14086 (N_14086,N_13718,N_13536);
nand U14087 (N_14087,N_13934,N_13873);
nor U14088 (N_14088,N_13757,N_13512);
nor U14089 (N_14089,N_13603,N_13715);
nand U14090 (N_14090,N_13726,N_13588);
nand U14091 (N_14091,N_13900,N_13520);
xor U14092 (N_14092,N_13590,N_13787);
or U14093 (N_14093,N_13646,N_13649);
nor U14094 (N_14094,N_13882,N_13773);
xor U14095 (N_14095,N_13936,N_13868);
xor U14096 (N_14096,N_13809,N_13920);
nor U14097 (N_14097,N_13642,N_13824);
nor U14098 (N_14098,N_13952,N_13943);
xor U14099 (N_14099,N_13939,N_13774);
nor U14100 (N_14100,N_13901,N_13565);
and U14101 (N_14101,N_13617,N_13921);
nand U14102 (N_14102,N_13962,N_13656);
nor U14103 (N_14103,N_13729,N_13699);
or U14104 (N_14104,N_13807,N_13696);
or U14105 (N_14105,N_13661,N_13866);
nand U14106 (N_14106,N_13747,N_13616);
xnor U14107 (N_14107,N_13762,N_13766);
nor U14108 (N_14108,N_13695,N_13601);
nor U14109 (N_14109,N_13976,N_13948);
nand U14110 (N_14110,N_13531,N_13703);
nand U14111 (N_14111,N_13909,N_13572);
and U14112 (N_14112,N_13567,N_13580);
or U14113 (N_14113,N_13902,N_13811);
xnor U14114 (N_14114,N_13670,N_13743);
nor U14115 (N_14115,N_13692,N_13523);
and U14116 (N_14116,N_13789,N_13640);
and U14117 (N_14117,N_13542,N_13761);
and U14118 (N_14118,N_13651,N_13732);
or U14119 (N_14119,N_13775,N_13941);
nand U14120 (N_14120,N_13595,N_13810);
and U14121 (N_14121,N_13916,N_13883);
or U14122 (N_14122,N_13735,N_13889);
and U14123 (N_14123,N_13737,N_13767);
and U14124 (N_14124,N_13938,N_13979);
and U14125 (N_14125,N_13663,N_13888);
or U14126 (N_14126,N_13683,N_13814);
xnor U14127 (N_14127,N_13589,N_13623);
nand U14128 (N_14128,N_13782,N_13998);
or U14129 (N_14129,N_13929,N_13770);
nand U14130 (N_14130,N_13812,N_13951);
xor U14131 (N_14131,N_13930,N_13804);
and U14132 (N_14132,N_13686,N_13854);
xnor U14133 (N_14133,N_13620,N_13530);
nand U14134 (N_14134,N_13550,N_13848);
and U14135 (N_14135,N_13515,N_13608);
xnor U14136 (N_14136,N_13690,N_13791);
and U14137 (N_14137,N_13828,N_13971);
or U14138 (N_14138,N_13553,N_13910);
and U14139 (N_14139,N_13560,N_13584);
xnor U14140 (N_14140,N_13573,N_13539);
or U14141 (N_14141,N_13827,N_13844);
nand U14142 (N_14142,N_13778,N_13821);
nor U14143 (N_14143,N_13533,N_13894);
or U14144 (N_14144,N_13925,N_13917);
xor U14145 (N_14145,N_13543,N_13581);
and U14146 (N_14146,N_13600,N_13674);
or U14147 (N_14147,N_13818,N_13609);
and U14148 (N_14148,N_13549,N_13986);
nand U14149 (N_14149,N_13832,N_13759);
nand U14150 (N_14150,N_13763,N_13853);
nand U14151 (N_14151,N_13836,N_13959);
nor U14152 (N_14152,N_13628,N_13507);
and U14153 (N_14153,N_13972,N_13802);
nand U14154 (N_14154,N_13680,N_13771);
and U14155 (N_14155,N_13997,N_13751);
nor U14156 (N_14156,N_13838,N_13534);
nor U14157 (N_14157,N_13632,N_13671);
nand U14158 (N_14158,N_13822,N_13776);
nand U14159 (N_14159,N_13545,N_13559);
and U14160 (N_14160,N_13876,N_13602);
nor U14161 (N_14161,N_13769,N_13893);
nor U14162 (N_14162,N_13906,N_13935);
or U14163 (N_14163,N_13704,N_13862);
and U14164 (N_14164,N_13835,N_13712);
and U14165 (N_14165,N_13622,N_13933);
nor U14166 (N_14166,N_13537,N_13966);
nor U14167 (N_14167,N_13503,N_13981);
xor U14168 (N_14168,N_13742,N_13506);
nor U14169 (N_14169,N_13739,N_13919);
or U14170 (N_14170,N_13895,N_13750);
nand U14171 (N_14171,N_13504,N_13685);
xor U14172 (N_14172,N_13886,N_13764);
or U14173 (N_14173,N_13664,N_13799);
nor U14174 (N_14174,N_13681,N_13991);
nor U14175 (N_14175,N_13781,N_13798);
nor U14176 (N_14176,N_13665,N_13864);
xnor U14177 (N_14177,N_13511,N_13586);
nand U14178 (N_14178,N_13731,N_13874);
or U14179 (N_14179,N_13985,N_13760);
nor U14180 (N_14180,N_13790,N_13655);
or U14181 (N_14181,N_13677,N_13648);
xor U14182 (N_14182,N_13596,N_13574);
nor U14183 (N_14183,N_13912,N_13708);
and U14184 (N_14184,N_13840,N_13566);
xor U14185 (N_14185,N_13993,N_13720);
and U14186 (N_14186,N_13568,N_13859);
nor U14187 (N_14187,N_13891,N_13987);
and U14188 (N_14188,N_13541,N_13527);
or U14189 (N_14189,N_13652,N_13839);
nand U14190 (N_14190,N_13897,N_13717);
and U14191 (N_14191,N_13667,N_13558);
nor U14192 (N_14192,N_13956,N_13709);
nor U14193 (N_14193,N_13689,N_13755);
nand U14194 (N_14194,N_13579,N_13621);
or U14195 (N_14195,N_13843,N_13749);
nor U14196 (N_14196,N_13598,N_13940);
and U14197 (N_14197,N_13613,N_13551);
or U14198 (N_14198,N_13816,N_13851);
or U14199 (N_14199,N_13519,N_13758);
or U14200 (N_14200,N_13634,N_13524);
nor U14201 (N_14201,N_13881,N_13980);
nor U14202 (N_14202,N_13697,N_13500);
xnor U14203 (N_14203,N_13614,N_13675);
or U14204 (N_14204,N_13831,N_13607);
nor U14205 (N_14205,N_13944,N_13528);
xor U14206 (N_14206,N_13969,N_13599);
and U14207 (N_14207,N_13710,N_13745);
xor U14208 (N_14208,N_13724,N_13548);
and U14209 (N_14209,N_13988,N_13611);
nor U14210 (N_14210,N_13660,N_13801);
and U14211 (N_14211,N_13694,N_13950);
nand U14212 (N_14212,N_13501,N_13736);
nand U14213 (N_14213,N_13668,N_13793);
nand U14214 (N_14214,N_13540,N_13706);
nor U14215 (N_14215,N_13676,N_13723);
and U14216 (N_14216,N_13850,N_13953);
xor U14217 (N_14217,N_13727,N_13624);
or U14218 (N_14218,N_13629,N_13637);
or U14219 (N_14219,N_13899,N_13555);
nand U14220 (N_14220,N_13578,N_13813);
and U14221 (N_14221,N_13904,N_13903);
or U14222 (N_14222,N_13526,N_13965);
and U14223 (N_14223,N_13508,N_13691);
or U14224 (N_14224,N_13554,N_13513);
and U14225 (N_14225,N_13779,N_13878);
nor U14226 (N_14226,N_13575,N_13892);
or U14227 (N_14227,N_13557,N_13679);
and U14228 (N_14228,N_13970,N_13714);
xor U14229 (N_14229,N_13516,N_13887);
xor U14230 (N_14230,N_13880,N_13872);
or U14231 (N_14231,N_13722,N_13847);
nor U14232 (N_14232,N_13626,N_13535);
or U14233 (N_14233,N_13858,N_13861);
nor U14234 (N_14234,N_13619,N_13546);
or U14235 (N_14235,N_13698,N_13688);
nor U14236 (N_14236,N_13908,N_13792);
or U14237 (N_14237,N_13856,N_13842);
and U14238 (N_14238,N_13996,N_13931);
or U14239 (N_14239,N_13786,N_13744);
nor U14240 (N_14240,N_13975,N_13510);
or U14241 (N_14241,N_13538,N_13964);
or U14242 (N_14242,N_13855,N_13561);
nor U14243 (N_14243,N_13597,N_13794);
nand U14244 (N_14244,N_13556,N_13605);
nand U14245 (N_14245,N_13618,N_13659);
nand U14246 (N_14246,N_13571,N_13863);
nor U14247 (N_14247,N_13857,N_13865);
nand U14248 (N_14248,N_13592,N_13625);
xnor U14249 (N_14249,N_13591,N_13594);
xnor U14250 (N_14250,N_13928,N_13749);
nand U14251 (N_14251,N_13902,N_13652);
and U14252 (N_14252,N_13790,N_13521);
nor U14253 (N_14253,N_13502,N_13526);
nor U14254 (N_14254,N_13509,N_13707);
nor U14255 (N_14255,N_13731,N_13845);
and U14256 (N_14256,N_13685,N_13991);
or U14257 (N_14257,N_13936,N_13876);
or U14258 (N_14258,N_13712,N_13820);
xor U14259 (N_14259,N_13564,N_13526);
and U14260 (N_14260,N_13673,N_13956);
and U14261 (N_14261,N_13575,N_13555);
or U14262 (N_14262,N_13864,N_13936);
and U14263 (N_14263,N_13719,N_13819);
xnor U14264 (N_14264,N_13555,N_13707);
and U14265 (N_14265,N_13841,N_13734);
and U14266 (N_14266,N_13563,N_13613);
nand U14267 (N_14267,N_13894,N_13563);
nor U14268 (N_14268,N_13666,N_13526);
and U14269 (N_14269,N_13785,N_13886);
nand U14270 (N_14270,N_13848,N_13630);
or U14271 (N_14271,N_13976,N_13909);
or U14272 (N_14272,N_13746,N_13705);
nand U14273 (N_14273,N_13988,N_13839);
xnor U14274 (N_14274,N_13826,N_13864);
xor U14275 (N_14275,N_13834,N_13632);
and U14276 (N_14276,N_13849,N_13560);
and U14277 (N_14277,N_13751,N_13736);
or U14278 (N_14278,N_13812,N_13862);
xnor U14279 (N_14279,N_13643,N_13974);
or U14280 (N_14280,N_13729,N_13826);
nor U14281 (N_14281,N_13522,N_13699);
nand U14282 (N_14282,N_13588,N_13561);
nand U14283 (N_14283,N_13842,N_13804);
or U14284 (N_14284,N_13681,N_13746);
or U14285 (N_14285,N_13509,N_13526);
nand U14286 (N_14286,N_13861,N_13900);
nor U14287 (N_14287,N_13986,N_13535);
nand U14288 (N_14288,N_13640,N_13993);
nor U14289 (N_14289,N_13929,N_13734);
or U14290 (N_14290,N_13813,N_13600);
and U14291 (N_14291,N_13868,N_13951);
xnor U14292 (N_14292,N_13613,N_13843);
nand U14293 (N_14293,N_13802,N_13900);
or U14294 (N_14294,N_13854,N_13682);
and U14295 (N_14295,N_13991,N_13558);
xnor U14296 (N_14296,N_13779,N_13732);
or U14297 (N_14297,N_13873,N_13940);
nor U14298 (N_14298,N_13944,N_13687);
or U14299 (N_14299,N_13555,N_13827);
and U14300 (N_14300,N_13679,N_13895);
nor U14301 (N_14301,N_13553,N_13551);
or U14302 (N_14302,N_13809,N_13774);
xor U14303 (N_14303,N_13709,N_13528);
nor U14304 (N_14304,N_13574,N_13882);
and U14305 (N_14305,N_13826,N_13649);
xor U14306 (N_14306,N_13515,N_13948);
or U14307 (N_14307,N_13560,N_13986);
nand U14308 (N_14308,N_13859,N_13937);
xnor U14309 (N_14309,N_13614,N_13663);
nand U14310 (N_14310,N_13736,N_13733);
and U14311 (N_14311,N_13538,N_13512);
and U14312 (N_14312,N_13824,N_13580);
nand U14313 (N_14313,N_13851,N_13942);
xor U14314 (N_14314,N_13672,N_13676);
xnor U14315 (N_14315,N_13642,N_13968);
or U14316 (N_14316,N_13746,N_13908);
nor U14317 (N_14317,N_13870,N_13556);
xnor U14318 (N_14318,N_13780,N_13577);
or U14319 (N_14319,N_13603,N_13685);
nor U14320 (N_14320,N_13906,N_13712);
nand U14321 (N_14321,N_13605,N_13559);
nand U14322 (N_14322,N_13721,N_13688);
or U14323 (N_14323,N_13786,N_13647);
nand U14324 (N_14324,N_13876,N_13560);
nand U14325 (N_14325,N_13762,N_13692);
nor U14326 (N_14326,N_13716,N_13888);
and U14327 (N_14327,N_13898,N_13848);
xnor U14328 (N_14328,N_13792,N_13550);
nand U14329 (N_14329,N_13743,N_13992);
nor U14330 (N_14330,N_13674,N_13976);
nor U14331 (N_14331,N_13741,N_13678);
nand U14332 (N_14332,N_13908,N_13719);
nand U14333 (N_14333,N_13557,N_13776);
and U14334 (N_14334,N_13988,N_13533);
and U14335 (N_14335,N_13555,N_13673);
nand U14336 (N_14336,N_13960,N_13893);
nand U14337 (N_14337,N_13877,N_13959);
or U14338 (N_14338,N_13528,N_13663);
nor U14339 (N_14339,N_13595,N_13548);
nand U14340 (N_14340,N_13932,N_13748);
nor U14341 (N_14341,N_13541,N_13613);
nand U14342 (N_14342,N_13566,N_13512);
or U14343 (N_14343,N_13759,N_13762);
nor U14344 (N_14344,N_13937,N_13671);
nor U14345 (N_14345,N_13881,N_13943);
and U14346 (N_14346,N_13782,N_13539);
or U14347 (N_14347,N_13652,N_13519);
nand U14348 (N_14348,N_13936,N_13551);
nand U14349 (N_14349,N_13874,N_13678);
xor U14350 (N_14350,N_13848,N_13922);
nand U14351 (N_14351,N_13676,N_13927);
xnor U14352 (N_14352,N_13505,N_13887);
and U14353 (N_14353,N_13700,N_13716);
nand U14354 (N_14354,N_13933,N_13825);
xor U14355 (N_14355,N_13967,N_13859);
xor U14356 (N_14356,N_13602,N_13737);
xnor U14357 (N_14357,N_13832,N_13993);
nand U14358 (N_14358,N_13531,N_13665);
nand U14359 (N_14359,N_13633,N_13675);
and U14360 (N_14360,N_13544,N_13689);
nor U14361 (N_14361,N_13631,N_13501);
xor U14362 (N_14362,N_13787,N_13880);
nand U14363 (N_14363,N_13586,N_13680);
and U14364 (N_14364,N_13940,N_13986);
nor U14365 (N_14365,N_13791,N_13785);
nor U14366 (N_14366,N_13831,N_13871);
and U14367 (N_14367,N_13979,N_13602);
xor U14368 (N_14368,N_13597,N_13920);
or U14369 (N_14369,N_13602,N_13971);
or U14370 (N_14370,N_13861,N_13813);
nand U14371 (N_14371,N_13839,N_13821);
nand U14372 (N_14372,N_13627,N_13833);
nor U14373 (N_14373,N_13790,N_13552);
and U14374 (N_14374,N_13752,N_13972);
and U14375 (N_14375,N_13650,N_13845);
and U14376 (N_14376,N_13939,N_13752);
or U14377 (N_14377,N_13949,N_13510);
and U14378 (N_14378,N_13642,N_13567);
nor U14379 (N_14379,N_13677,N_13617);
or U14380 (N_14380,N_13962,N_13950);
and U14381 (N_14381,N_13679,N_13689);
xnor U14382 (N_14382,N_13543,N_13777);
and U14383 (N_14383,N_13532,N_13657);
or U14384 (N_14384,N_13777,N_13688);
and U14385 (N_14385,N_13928,N_13563);
or U14386 (N_14386,N_13744,N_13516);
or U14387 (N_14387,N_13606,N_13624);
xnor U14388 (N_14388,N_13594,N_13773);
nand U14389 (N_14389,N_13928,N_13934);
nand U14390 (N_14390,N_13952,N_13607);
or U14391 (N_14391,N_13785,N_13735);
nor U14392 (N_14392,N_13781,N_13903);
xnor U14393 (N_14393,N_13571,N_13701);
or U14394 (N_14394,N_13729,N_13632);
or U14395 (N_14395,N_13539,N_13547);
or U14396 (N_14396,N_13541,N_13848);
nor U14397 (N_14397,N_13630,N_13689);
nor U14398 (N_14398,N_13680,N_13584);
nand U14399 (N_14399,N_13981,N_13613);
xnor U14400 (N_14400,N_13791,N_13547);
nand U14401 (N_14401,N_13520,N_13747);
xor U14402 (N_14402,N_13683,N_13927);
or U14403 (N_14403,N_13994,N_13887);
or U14404 (N_14404,N_13922,N_13784);
nand U14405 (N_14405,N_13684,N_13549);
xnor U14406 (N_14406,N_13632,N_13653);
nor U14407 (N_14407,N_13600,N_13824);
or U14408 (N_14408,N_13589,N_13706);
or U14409 (N_14409,N_13657,N_13632);
or U14410 (N_14410,N_13607,N_13962);
or U14411 (N_14411,N_13894,N_13584);
and U14412 (N_14412,N_13946,N_13672);
xor U14413 (N_14413,N_13637,N_13985);
and U14414 (N_14414,N_13796,N_13812);
nor U14415 (N_14415,N_13609,N_13863);
or U14416 (N_14416,N_13984,N_13914);
xnor U14417 (N_14417,N_13617,N_13531);
xnor U14418 (N_14418,N_13914,N_13614);
xor U14419 (N_14419,N_13839,N_13658);
and U14420 (N_14420,N_13878,N_13552);
nor U14421 (N_14421,N_13606,N_13779);
nor U14422 (N_14422,N_13650,N_13641);
nor U14423 (N_14423,N_13816,N_13754);
xor U14424 (N_14424,N_13984,N_13837);
xnor U14425 (N_14425,N_13960,N_13605);
xnor U14426 (N_14426,N_13549,N_13720);
nand U14427 (N_14427,N_13755,N_13614);
and U14428 (N_14428,N_13994,N_13957);
nor U14429 (N_14429,N_13836,N_13550);
xor U14430 (N_14430,N_13911,N_13949);
xor U14431 (N_14431,N_13802,N_13626);
xnor U14432 (N_14432,N_13859,N_13775);
and U14433 (N_14433,N_13761,N_13916);
and U14434 (N_14434,N_13531,N_13671);
nand U14435 (N_14435,N_13718,N_13619);
or U14436 (N_14436,N_13546,N_13736);
xnor U14437 (N_14437,N_13908,N_13714);
xnor U14438 (N_14438,N_13954,N_13977);
xnor U14439 (N_14439,N_13989,N_13558);
and U14440 (N_14440,N_13683,N_13714);
and U14441 (N_14441,N_13876,N_13739);
nand U14442 (N_14442,N_13623,N_13572);
nand U14443 (N_14443,N_13643,N_13911);
or U14444 (N_14444,N_13921,N_13781);
or U14445 (N_14445,N_13970,N_13786);
nor U14446 (N_14446,N_13632,N_13873);
nor U14447 (N_14447,N_13774,N_13662);
and U14448 (N_14448,N_13554,N_13972);
nor U14449 (N_14449,N_13911,N_13598);
xor U14450 (N_14450,N_13939,N_13671);
or U14451 (N_14451,N_13717,N_13887);
xor U14452 (N_14452,N_13908,N_13763);
nor U14453 (N_14453,N_13881,N_13777);
nor U14454 (N_14454,N_13647,N_13715);
nor U14455 (N_14455,N_13588,N_13940);
nor U14456 (N_14456,N_13842,N_13664);
and U14457 (N_14457,N_13782,N_13641);
nand U14458 (N_14458,N_13961,N_13888);
and U14459 (N_14459,N_13957,N_13972);
xor U14460 (N_14460,N_13680,N_13835);
nand U14461 (N_14461,N_13729,N_13595);
or U14462 (N_14462,N_13646,N_13531);
xnor U14463 (N_14463,N_13844,N_13606);
nor U14464 (N_14464,N_13855,N_13757);
xor U14465 (N_14465,N_13651,N_13832);
nor U14466 (N_14466,N_13916,N_13998);
or U14467 (N_14467,N_13924,N_13630);
xnor U14468 (N_14468,N_13698,N_13551);
nand U14469 (N_14469,N_13604,N_13877);
and U14470 (N_14470,N_13628,N_13583);
and U14471 (N_14471,N_13872,N_13516);
and U14472 (N_14472,N_13914,N_13735);
and U14473 (N_14473,N_13613,N_13923);
nand U14474 (N_14474,N_13717,N_13744);
or U14475 (N_14475,N_13552,N_13999);
and U14476 (N_14476,N_13692,N_13764);
or U14477 (N_14477,N_13983,N_13769);
and U14478 (N_14478,N_13733,N_13642);
or U14479 (N_14479,N_13914,N_13603);
xor U14480 (N_14480,N_13527,N_13755);
and U14481 (N_14481,N_13974,N_13700);
or U14482 (N_14482,N_13616,N_13523);
or U14483 (N_14483,N_13618,N_13750);
nand U14484 (N_14484,N_13643,N_13699);
nor U14485 (N_14485,N_13582,N_13750);
and U14486 (N_14486,N_13776,N_13892);
and U14487 (N_14487,N_13527,N_13552);
and U14488 (N_14488,N_13502,N_13514);
nand U14489 (N_14489,N_13637,N_13937);
nand U14490 (N_14490,N_13579,N_13581);
nand U14491 (N_14491,N_13749,N_13613);
nand U14492 (N_14492,N_13861,N_13529);
xnor U14493 (N_14493,N_13534,N_13703);
or U14494 (N_14494,N_13510,N_13914);
and U14495 (N_14495,N_13963,N_13824);
nor U14496 (N_14496,N_13635,N_13780);
nor U14497 (N_14497,N_13553,N_13620);
and U14498 (N_14498,N_13726,N_13814);
or U14499 (N_14499,N_13987,N_13520);
nand U14500 (N_14500,N_14388,N_14126);
and U14501 (N_14501,N_14033,N_14403);
nand U14502 (N_14502,N_14378,N_14384);
nor U14503 (N_14503,N_14032,N_14373);
nor U14504 (N_14504,N_14105,N_14390);
or U14505 (N_14505,N_14211,N_14432);
and U14506 (N_14506,N_14053,N_14216);
xor U14507 (N_14507,N_14336,N_14149);
nand U14508 (N_14508,N_14480,N_14293);
xnor U14509 (N_14509,N_14494,N_14009);
or U14510 (N_14510,N_14072,N_14365);
and U14511 (N_14511,N_14044,N_14245);
and U14512 (N_14512,N_14212,N_14435);
nor U14513 (N_14513,N_14246,N_14055);
nand U14514 (N_14514,N_14230,N_14300);
or U14515 (N_14515,N_14454,N_14027);
nand U14516 (N_14516,N_14345,N_14304);
nand U14517 (N_14517,N_14376,N_14213);
nand U14518 (N_14518,N_14007,N_14228);
xor U14519 (N_14519,N_14325,N_14363);
nor U14520 (N_14520,N_14205,N_14194);
xnor U14521 (N_14521,N_14364,N_14477);
or U14522 (N_14522,N_14100,N_14183);
nand U14523 (N_14523,N_14050,N_14111);
xnor U14524 (N_14524,N_14433,N_14485);
and U14525 (N_14525,N_14052,N_14233);
and U14526 (N_14526,N_14441,N_14056);
or U14527 (N_14527,N_14393,N_14356);
or U14528 (N_14528,N_14201,N_14457);
and U14529 (N_14529,N_14179,N_14078);
or U14530 (N_14530,N_14051,N_14286);
and U14531 (N_14531,N_14115,N_14085);
nand U14532 (N_14532,N_14215,N_14317);
or U14533 (N_14533,N_14147,N_14295);
nand U14534 (N_14534,N_14255,N_14483);
and U14535 (N_14535,N_14283,N_14349);
or U14536 (N_14536,N_14272,N_14309);
and U14537 (N_14537,N_14497,N_14342);
or U14538 (N_14538,N_14186,N_14297);
and U14539 (N_14539,N_14326,N_14404);
nand U14540 (N_14540,N_14067,N_14410);
nand U14541 (N_14541,N_14308,N_14202);
or U14542 (N_14542,N_14266,N_14341);
nand U14543 (N_14543,N_14134,N_14427);
nand U14544 (N_14544,N_14118,N_14425);
nand U14545 (N_14545,N_14301,N_14486);
nor U14546 (N_14546,N_14362,N_14018);
nand U14547 (N_14547,N_14139,N_14200);
xor U14548 (N_14548,N_14145,N_14076);
nor U14549 (N_14549,N_14185,N_14413);
xor U14550 (N_14550,N_14140,N_14204);
and U14551 (N_14551,N_14237,N_14334);
xor U14552 (N_14552,N_14244,N_14288);
and U14553 (N_14553,N_14263,N_14088);
or U14554 (N_14554,N_14419,N_14068);
nand U14555 (N_14555,N_14241,N_14192);
and U14556 (N_14556,N_14357,N_14040);
xor U14557 (N_14557,N_14273,N_14226);
or U14558 (N_14558,N_14391,N_14096);
xor U14559 (N_14559,N_14375,N_14157);
and U14560 (N_14560,N_14093,N_14382);
and U14561 (N_14561,N_14089,N_14219);
or U14562 (N_14562,N_14343,N_14409);
nor U14563 (N_14563,N_14170,N_14478);
and U14564 (N_14564,N_14449,N_14469);
and U14565 (N_14565,N_14476,N_14337);
or U14566 (N_14566,N_14499,N_14119);
and U14567 (N_14567,N_14164,N_14199);
xor U14568 (N_14568,N_14066,N_14493);
xor U14569 (N_14569,N_14101,N_14247);
or U14570 (N_14570,N_14175,N_14374);
and U14571 (N_14571,N_14191,N_14043);
nor U14572 (N_14572,N_14097,N_14198);
nor U14573 (N_14573,N_14242,N_14369);
or U14574 (N_14574,N_14367,N_14468);
or U14575 (N_14575,N_14239,N_14253);
xnor U14576 (N_14576,N_14495,N_14073);
nand U14577 (N_14577,N_14269,N_14182);
or U14578 (N_14578,N_14310,N_14133);
xnor U14579 (N_14579,N_14046,N_14277);
and U14580 (N_14580,N_14082,N_14303);
and U14581 (N_14581,N_14138,N_14117);
nor U14582 (N_14582,N_14030,N_14487);
xnor U14583 (N_14583,N_14172,N_14002);
xnor U14584 (N_14584,N_14284,N_14077);
xor U14585 (N_14585,N_14123,N_14292);
xor U14586 (N_14586,N_14346,N_14445);
nand U14587 (N_14587,N_14348,N_14017);
nand U14588 (N_14588,N_14271,N_14421);
and U14589 (N_14589,N_14232,N_14305);
xor U14590 (N_14590,N_14360,N_14312);
nor U14591 (N_14591,N_14095,N_14423);
nor U14592 (N_14592,N_14158,N_14322);
nand U14593 (N_14593,N_14354,N_14315);
xnor U14594 (N_14594,N_14108,N_14311);
or U14595 (N_14595,N_14352,N_14406);
or U14596 (N_14596,N_14127,N_14021);
and U14597 (N_14597,N_14006,N_14025);
nand U14598 (N_14598,N_14217,N_14104);
nor U14599 (N_14599,N_14261,N_14162);
and U14600 (N_14600,N_14203,N_14439);
and U14601 (N_14601,N_14330,N_14022);
xnor U14602 (N_14602,N_14110,N_14426);
nand U14603 (N_14603,N_14359,N_14069);
or U14604 (N_14604,N_14103,N_14287);
nand U14605 (N_14605,N_14159,N_14278);
nor U14606 (N_14606,N_14235,N_14451);
or U14607 (N_14607,N_14090,N_14178);
nand U14608 (N_14608,N_14383,N_14148);
xnor U14609 (N_14609,N_14173,N_14321);
nor U14610 (N_14610,N_14234,N_14092);
and U14611 (N_14611,N_14328,N_14381);
nand U14612 (N_14612,N_14080,N_14222);
or U14613 (N_14613,N_14465,N_14169);
nand U14614 (N_14614,N_14231,N_14256);
xor U14615 (N_14615,N_14070,N_14129);
or U14616 (N_14616,N_14141,N_14026);
nand U14617 (N_14617,N_14320,N_14464);
nor U14618 (N_14618,N_14387,N_14282);
or U14619 (N_14619,N_14307,N_14001);
and U14620 (N_14620,N_14392,N_14063);
xor U14621 (N_14621,N_14177,N_14482);
nand U14622 (N_14622,N_14071,N_14397);
or U14623 (N_14623,N_14210,N_14339);
nand U14624 (N_14624,N_14340,N_14035);
and U14625 (N_14625,N_14227,N_14130);
or U14626 (N_14626,N_14492,N_14412);
or U14627 (N_14627,N_14415,N_14031);
xor U14628 (N_14628,N_14181,N_14087);
xor U14629 (N_14629,N_14190,N_14324);
or U14630 (N_14630,N_14098,N_14466);
nor U14631 (N_14631,N_14417,N_14298);
nand U14632 (N_14632,N_14459,N_14472);
or U14633 (N_14633,N_14012,N_14316);
or U14634 (N_14634,N_14251,N_14450);
xnor U14635 (N_14635,N_14489,N_14456);
xnor U14636 (N_14636,N_14106,N_14274);
and U14637 (N_14637,N_14121,N_14120);
and U14638 (N_14638,N_14418,N_14453);
or U14639 (N_14639,N_14462,N_14491);
nand U14640 (N_14640,N_14019,N_14084);
xor U14641 (N_14641,N_14248,N_14395);
nor U14642 (N_14642,N_14313,N_14028);
nor U14643 (N_14643,N_14344,N_14276);
or U14644 (N_14644,N_14153,N_14306);
or U14645 (N_14645,N_14408,N_14353);
nand U14646 (N_14646,N_14240,N_14029);
nand U14647 (N_14647,N_14180,N_14010);
and U14648 (N_14648,N_14401,N_14490);
or U14649 (N_14649,N_14064,N_14386);
nand U14650 (N_14650,N_14000,N_14350);
nand U14651 (N_14651,N_14150,N_14275);
nor U14652 (N_14652,N_14137,N_14446);
or U14653 (N_14653,N_14368,N_14124);
or U14654 (N_14654,N_14249,N_14079);
and U14655 (N_14655,N_14143,N_14498);
and U14656 (N_14656,N_14132,N_14188);
or U14657 (N_14657,N_14004,N_14038);
or U14658 (N_14658,N_14224,N_14122);
nor U14659 (N_14659,N_14061,N_14400);
or U14660 (N_14660,N_14291,N_14396);
xor U14661 (N_14661,N_14189,N_14016);
nand U14662 (N_14662,N_14264,N_14081);
nand U14663 (N_14663,N_14280,N_14474);
xor U14664 (N_14664,N_14014,N_14463);
or U14665 (N_14665,N_14428,N_14430);
nor U14666 (N_14666,N_14333,N_14060);
xor U14667 (N_14667,N_14460,N_14323);
nand U14668 (N_14668,N_14452,N_14218);
and U14669 (N_14669,N_14370,N_14161);
or U14670 (N_14670,N_14065,N_14358);
and U14671 (N_14671,N_14429,N_14023);
or U14672 (N_14672,N_14057,N_14059);
xnor U14673 (N_14673,N_14146,N_14444);
nor U14674 (N_14674,N_14163,N_14385);
and U14675 (N_14675,N_14112,N_14434);
and U14676 (N_14676,N_14260,N_14473);
and U14677 (N_14677,N_14207,N_14187);
xor U14678 (N_14678,N_14225,N_14042);
and U14679 (N_14679,N_14135,N_14389);
nand U14680 (N_14680,N_14037,N_14318);
or U14681 (N_14681,N_14281,N_14047);
nand U14682 (N_14682,N_14327,N_14236);
nor U14683 (N_14683,N_14167,N_14171);
nor U14684 (N_14684,N_14458,N_14144);
or U14685 (N_14685,N_14270,N_14195);
xor U14686 (N_14686,N_14262,N_14223);
or U14687 (N_14687,N_14160,N_14351);
or U14688 (N_14688,N_14074,N_14214);
nor U14689 (N_14689,N_14285,N_14398);
nor U14690 (N_14690,N_14099,N_14443);
and U14691 (N_14691,N_14184,N_14402);
and U14692 (N_14692,N_14411,N_14447);
xor U14693 (N_14693,N_14405,N_14128);
nand U14694 (N_14694,N_14252,N_14366);
or U14695 (N_14695,N_14335,N_14156);
xnor U14696 (N_14696,N_14048,N_14086);
and U14697 (N_14697,N_14221,N_14475);
and U14698 (N_14698,N_14414,N_14289);
xnor U14699 (N_14699,N_14174,N_14470);
and U14700 (N_14700,N_14267,N_14039);
or U14701 (N_14701,N_14015,N_14008);
nand U14702 (N_14702,N_14455,N_14259);
nor U14703 (N_14703,N_14416,N_14440);
and U14704 (N_14704,N_14250,N_14054);
and U14705 (N_14705,N_14116,N_14003);
or U14706 (N_14706,N_14020,N_14290);
nand U14707 (N_14707,N_14302,N_14329);
and U14708 (N_14708,N_14131,N_14347);
xnor U14709 (N_14709,N_14151,N_14107);
and U14710 (N_14710,N_14265,N_14091);
xor U14711 (N_14711,N_14407,N_14005);
and U14712 (N_14712,N_14257,N_14154);
and U14713 (N_14713,N_14377,N_14319);
nor U14714 (N_14714,N_14243,N_14299);
nor U14715 (N_14715,N_14294,N_14206);
and U14716 (N_14716,N_14279,N_14371);
nand U14717 (N_14717,N_14484,N_14422);
or U14718 (N_14718,N_14361,N_14471);
or U14719 (N_14719,N_14049,N_14166);
or U14720 (N_14720,N_14034,N_14220);
xnor U14721 (N_14721,N_14045,N_14196);
and U14722 (N_14722,N_14296,N_14461);
nor U14723 (N_14723,N_14436,N_14152);
and U14724 (N_14724,N_14399,N_14420);
nand U14725 (N_14725,N_14332,N_14431);
or U14726 (N_14726,N_14102,N_14125);
or U14727 (N_14727,N_14467,N_14041);
and U14728 (N_14728,N_14136,N_14379);
nand U14729 (N_14729,N_14238,N_14155);
xnor U14730 (N_14730,N_14024,N_14165);
nand U14731 (N_14731,N_14209,N_14083);
nor U14732 (N_14732,N_14448,N_14488);
nor U14733 (N_14733,N_14481,N_14193);
and U14734 (N_14734,N_14109,N_14062);
or U14735 (N_14735,N_14442,N_14331);
xor U14736 (N_14736,N_14268,N_14380);
or U14737 (N_14737,N_14355,N_14394);
and U14738 (N_14738,N_14094,N_14479);
or U14739 (N_14739,N_14496,N_14114);
nand U14740 (N_14740,N_14208,N_14113);
nand U14741 (N_14741,N_14075,N_14176);
nand U14742 (N_14742,N_14011,N_14372);
and U14743 (N_14743,N_14229,N_14437);
nand U14744 (N_14744,N_14142,N_14314);
nor U14745 (N_14745,N_14424,N_14036);
and U14746 (N_14746,N_14258,N_14168);
and U14747 (N_14747,N_14058,N_14438);
xnor U14748 (N_14748,N_14197,N_14338);
and U14749 (N_14749,N_14254,N_14013);
or U14750 (N_14750,N_14051,N_14291);
and U14751 (N_14751,N_14207,N_14427);
xor U14752 (N_14752,N_14499,N_14114);
nand U14753 (N_14753,N_14022,N_14449);
or U14754 (N_14754,N_14264,N_14371);
nand U14755 (N_14755,N_14133,N_14393);
nor U14756 (N_14756,N_14155,N_14318);
or U14757 (N_14757,N_14002,N_14144);
and U14758 (N_14758,N_14137,N_14263);
and U14759 (N_14759,N_14311,N_14343);
nand U14760 (N_14760,N_14317,N_14194);
nor U14761 (N_14761,N_14057,N_14379);
nor U14762 (N_14762,N_14193,N_14045);
xor U14763 (N_14763,N_14463,N_14409);
nor U14764 (N_14764,N_14490,N_14038);
nor U14765 (N_14765,N_14246,N_14182);
and U14766 (N_14766,N_14290,N_14328);
nor U14767 (N_14767,N_14249,N_14343);
or U14768 (N_14768,N_14170,N_14025);
nand U14769 (N_14769,N_14020,N_14404);
or U14770 (N_14770,N_14164,N_14107);
nand U14771 (N_14771,N_14354,N_14112);
xor U14772 (N_14772,N_14446,N_14079);
nand U14773 (N_14773,N_14196,N_14338);
nor U14774 (N_14774,N_14160,N_14326);
nand U14775 (N_14775,N_14248,N_14116);
or U14776 (N_14776,N_14096,N_14293);
nand U14777 (N_14777,N_14204,N_14231);
nor U14778 (N_14778,N_14196,N_14089);
nand U14779 (N_14779,N_14447,N_14499);
nor U14780 (N_14780,N_14313,N_14439);
nand U14781 (N_14781,N_14303,N_14346);
nand U14782 (N_14782,N_14148,N_14179);
xor U14783 (N_14783,N_14102,N_14259);
and U14784 (N_14784,N_14395,N_14154);
nor U14785 (N_14785,N_14031,N_14356);
xor U14786 (N_14786,N_14454,N_14243);
nand U14787 (N_14787,N_14121,N_14367);
xor U14788 (N_14788,N_14069,N_14135);
and U14789 (N_14789,N_14313,N_14365);
xor U14790 (N_14790,N_14137,N_14485);
or U14791 (N_14791,N_14032,N_14497);
xor U14792 (N_14792,N_14394,N_14445);
or U14793 (N_14793,N_14361,N_14118);
nor U14794 (N_14794,N_14391,N_14429);
or U14795 (N_14795,N_14259,N_14463);
xor U14796 (N_14796,N_14199,N_14190);
or U14797 (N_14797,N_14245,N_14069);
or U14798 (N_14798,N_14417,N_14025);
nor U14799 (N_14799,N_14497,N_14217);
or U14800 (N_14800,N_14107,N_14322);
or U14801 (N_14801,N_14285,N_14277);
xor U14802 (N_14802,N_14264,N_14338);
nor U14803 (N_14803,N_14476,N_14297);
and U14804 (N_14804,N_14184,N_14248);
xnor U14805 (N_14805,N_14391,N_14146);
and U14806 (N_14806,N_14241,N_14397);
nor U14807 (N_14807,N_14419,N_14087);
or U14808 (N_14808,N_14002,N_14091);
nand U14809 (N_14809,N_14197,N_14318);
and U14810 (N_14810,N_14477,N_14173);
nor U14811 (N_14811,N_14424,N_14190);
nand U14812 (N_14812,N_14432,N_14353);
nand U14813 (N_14813,N_14105,N_14328);
nand U14814 (N_14814,N_14196,N_14246);
nor U14815 (N_14815,N_14396,N_14494);
and U14816 (N_14816,N_14024,N_14447);
nor U14817 (N_14817,N_14165,N_14218);
xor U14818 (N_14818,N_14300,N_14457);
and U14819 (N_14819,N_14096,N_14133);
nor U14820 (N_14820,N_14092,N_14110);
xor U14821 (N_14821,N_14464,N_14066);
nor U14822 (N_14822,N_14050,N_14261);
or U14823 (N_14823,N_14204,N_14130);
xor U14824 (N_14824,N_14345,N_14123);
nand U14825 (N_14825,N_14031,N_14155);
xor U14826 (N_14826,N_14041,N_14428);
and U14827 (N_14827,N_14271,N_14034);
nor U14828 (N_14828,N_14136,N_14401);
nor U14829 (N_14829,N_14496,N_14420);
nand U14830 (N_14830,N_14400,N_14439);
xor U14831 (N_14831,N_14403,N_14162);
xnor U14832 (N_14832,N_14347,N_14059);
xor U14833 (N_14833,N_14076,N_14049);
nor U14834 (N_14834,N_14282,N_14174);
nor U14835 (N_14835,N_14230,N_14167);
nor U14836 (N_14836,N_14348,N_14001);
and U14837 (N_14837,N_14283,N_14144);
nand U14838 (N_14838,N_14395,N_14160);
or U14839 (N_14839,N_14277,N_14486);
xnor U14840 (N_14840,N_14474,N_14104);
xor U14841 (N_14841,N_14419,N_14091);
or U14842 (N_14842,N_14191,N_14274);
nor U14843 (N_14843,N_14460,N_14107);
xor U14844 (N_14844,N_14190,N_14253);
nor U14845 (N_14845,N_14024,N_14396);
nand U14846 (N_14846,N_14183,N_14287);
or U14847 (N_14847,N_14421,N_14232);
nor U14848 (N_14848,N_14334,N_14074);
nor U14849 (N_14849,N_14100,N_14286);
or U14850 (N_14850,N_14049,N_14384);
and U14851 (N_14851,N_14392,N_14231);
nor U14852 (N_14852,N_14019,N_14456);
and U14853 (N_14853,N_14023,N_14409);
nor U14854 (N_14854,N_14047,N_14489);
and U14855 (N_14855,N_14371,N_14461);
xor U14856 (N_14856,N_14370,N_14214);
nor U14857 (N_14857,N_14171,N_14473);
nand U14858 (N_14858,N_14423,N_14278);
and U14859 (N_14859,N_14274,N_14196);
nor U14860 (N_14860,N_14144,N_14499);
and U14861 (N_14861,N_14397,N_14086);
or U14862 (N_14862,N_14324,N_14145);
nand U14863 (N_14863,N_14103,N_14260);
nor U14864 (N_14864,N_14141,N_14114);
and U14865 (N_14865,N_14220,N_14459);
or U14866 (N_14866,N_14304,N_14228);
or U14867 (N_14867,N_14358,N_14437);
nand U14868 (N_14868,N_14329,N_14489);
nor U14869 (N_14869,N_14376,N_14400);
or U14870 (N_14870,N_14469,N_14450);
and U14871 (N_14871,N_14183,N_14369);
and U14872 (N_14872,N_14494,N_14168);
nor U14873 (N_14873,N_14089,N_14107);
nand U14874 (N_14874,N_14199,N_14320);
nand U14875 (N_14875,N_14174,N_14298);
nand U14876 (N_14876,N_14344,N_14301);
nand U14877 (N_14877,N_14324,N_14353);
nor U14878 (N_14878,N_14212,N_14051);
and U14879 (N_14879,N_14463,N_14430);
or U14880 (N_14880,N_14036,N_14223);
nand U14881 (N_14881,N_14181,N_14261);
and U14882 (N_14882,N_14343,N_14266);
and U14883 (N_14883,N_14064,N_14089);
nand U14884 (N_14884,N_14133,N_14448);
or U14885 (N_14885,N_14304,N_14222);
or U14886 (N_14886,N_14036,N_14124);
nand U14887 (N_14887,N_14298,N_14196);
nand U14888 (N_14888,N_14461,N_14349);
xor U14889 (N_14889,N_14479,N_14280);
and U14890 (N_14890,N_14474,N_14160);
nor U14891 (N_14891,N_14129,N_14227);
nand U14892 (N_14892,N_14266,N_14481);
or U14893 (N_14893,N_14053,N_14402);
and U14894 (N_14894,N_14286,N_14211);
nand U14895 (N_14895,N_14333,N_14415);
or U14896 (N_14896,N_14029,N_14044);
nand U14897 (N_14897,N_14115,N_14465);
or U14898 (N_14898,N_14422,N_14098);
or U14899 (N_14899,N_14004,N_14251);
nand U14900 (N_14900,N_14004,N_14210);
nor U14901 (N_14901,N_14271,N_14089);
xnor U14902 (N_14902,N_14205,N_14259);
nand U14903 (N_14903,N_14060,N_14195);
xnor U14904 (N_14904,N_14369,N_14238);
nor U14905 (N_14905,N_14465,N_14451);
nand U14906 (N_14906,N_14115,N_14469);
nor U14907 (N_14907,N_14428,N_14409);
and U14908 (N_14908,N_14067,N_14119);
nor U14909 (N_14909,N_14496,N_14498);
nor U14910 (N_14910,N_14111,N_14454);
and U14911 (N_14911,N_14379,N_14496);
nand U14912 (N_14912,N_14488,N_14442);
and U14913 (N_14913,N_14268,N_14095);
and U14914 (N_14914,N_14489,N_14111);
or U14915 (N_14915,N_14256,N_14102);
xnor U14916 (N_14916,N_14069,N_14318);
nand U14917 (N_14917,N_14065,N_14428);
and U14918 (N_14918,N_14043,N_14495);
and U14919 (N_14919,N_14474,N_14266);
or U14920 (N_14920,N_14218,N_14441);
or U14921 (N_14921,N_14356,N_14233);
nor U14922 (N_14922,N_14379,N_14048);
and U14923 (N_14923,N_14177,N_14470);
nand U14924 (N_14924,N_14216,N_14424);
or U14925 (N_14925,N_14216,N_14290);
and U14926 (N_14926,N_14441,N_14376);
nand U14927 (N_14927,N_14079,N_14108);
nand U14928 (N_14928,N_14288,N_14128);
and U14929 (N_14929,N_14379,N_14132);
nor U14930 (N_14930,N_14158,N_14186);
or U14931 (N_14931,N_14257,N_14488);
and U14932 (N_14932,N_14364,N_14097);
xor U14933 (N_14933,N_14152,N_14138);
xnor U14934 (N_14934,N_14024,N_14145);
and U14935 (N_14935,N_14129,N_14255);
and U14936 (N_14936,N_14337,N_14165);
or U14937 (N_14937,N_14199,N_14463);
nand U14938 (N_14938,N_14257,N_14404);
nand U14939 (N_14939,N_14209,N_14313);
nor U14940 (N_14940,N_14150,N_14295);
or U14941 (N_14941,N_14222,N_14030);
and U14942 (N_14942,N_14187,N_14066);
nand U14943 (N_14943,N_14374,N_14006);
nand U14944 (N_14944,N_14130,N_14132);
nand U14945 (N_14945,N_14374,N_14046);
nor U14946 (N_14946,N_14314,N_14430);
or U14947 (N_14947,N_14438,N_14499);
or U14948 (N_14948,N_14295,N_14356);
and U14949 (N_14949,N_14228,N_14158);
or U14950 (N_14950,N_14381,N_14156);
or U14951 (N_14951,N_14395,N_14071);
xnor U14952 (N_14952,N_14058,N_14378);
or U14953 (N_14953,N_14440,N_14181);
xor U14954 (N_14954,N_14119,N_14312);
and U14955 (N_14955,N_14165,N_14399);
nor U14956 (N_14956,N_14035,N_14385);
xnor U14957 (N_14957,N_14267,N_14103);
and U14958 (N_14958,N_14207,N_14156);
nor U14959 (N_14959,N_14017,N_14339);
nand U14960 (N_14960,N_14257,N_14011);
xor U14961 (N_14961,N_14237,N_14046);
or U14962 (N_14962,N_14399,N_14236);
or U14963 (N_14963,N_14210,N_14103);
and U14964 (N_14964,N_14077,N_14097);
and U14965 (N_14965,N_14469,N_14090);
nand U14966 (N_14966,N_14358,N_14401);
nor U14967 (N_14967,N_14003,N_14412);
or U14968 (N_14968,N_14393,N_14192);
nand U14969 (N_14969,N_14136,N_14190);
or U14970 (N_14970,N_14121,N_14317);
nand U14971 (N_14971,N_14179,N_14118);
xor U14972 (N_14972,N_14003,N_14089);
nor U14973 (N_14973,N_14320,N_14287);
or U14974 (N_14974,N_14473,N_14067);
and U14975 (N_14975,N_14367,N_14321);
and U14976 (N_14976,N_14214,N_14167);
nand U14977 (N_14977,N_14067,N_14348);
and U14978 (N_14978,N_14231,N_14492);
nand U14979 (N_14979,N_14350,N_14080);
nor U14980 (N_14980,N_14304,N_14086);
or U14981 (N_14981,N_14059,N_14215);
or U14982 (N_14982,N_14310,N_14258);
or U14983 (N_14983,N_14114,N_14360);
and U14984 (N_14984,N_14325,N_14357);
xnor U14985 (N_14985,N_14130,N_14353);
nor U14986 (N_14986,N_14149,N_14179);
or U14987 (N_14987,N_14016,N_14105);
nand U14988 (N_14988,N_14434,N_14090);
and U14989 (N_14989,N_14411,N_14166);
xor U14990 (N_14990,N_14040,N_14478);
and U14991 (N_14991,N_14431,N_14050);
xor U14992 (N_14992,N_14270,N_14043);
nand U14993 (N_14993,N_14024,N_14185);
xnor U14994 (N_14994,N_14161,N_14409);
and U14995 (N_14995,N_14150,N_14459);
nor U14996 (N_14996,N_14077,N_14289);
xnor U14997 (N_14997,N_14344,N_14078);
or U14998 (N_14998,N_14026,N_14174);
nor U14999 (N_14999,N_14373,N_14114);
nand U15000 (N_15000,N_14620,N_14577);
nor U15001 (N_15001,N_14957,N_14507);
and U15002 (N_15002,N_14615,N_14902);
xor U15003 (N_15003,N_14686,N_14523);
and U15004 (N_15004,N_14500,N_14881);
or U15005 (N_15005,N_14808,N_14602);
or U15006 (N_15006,N_14767,N_14742);
xnor U15007 (N_15007,N_14780,N_14914);
xor U15008 (N_15008,N_14975,N_14913);
nor U15009 (N_15009,N_14885,N_14586);
xor U15010 (N_15010,N_14922,N_14786);
nor U15011 (N_15011,N_14709,N_14833);
nand U15012 (N_15012,N_14992,N_14530);
or U15013 (N_15013,N_14733,N_14774);
nor U15014 (N_15014,N_14809,N_14525);
or U15015 (N_15015,N_14793,N_14639);
and U15016 (N_15016,N_14983,N_14510);
nor U15017 (N_15017,N_14839,N_14832);
or U15018 (N_15018,N_14807,N_14726);
nor U15019 (N_15019,N_14869,N_14846);
nand U15020 (N_15020,N_14712,N_14916);
xor U15021 (N_15021,N_14685,N_14900);
nor U15022 (N_15022,N_14835,N_14876);
or U15023 (N_15023,N_14631,N_14782);
nand U15024 (N_15024,N_14581,N_14958);
or U15025 (N_15025,N_14842,N_14871);
or U15026 (N_15026,N_14562,N_14788);
and U15027 (N_15027,N_14528,N_14805);
and U15028 (N_15028,N_14859,N_14536);
and U15029 (N_15029,N_14821,N_14830);
nor U15030 (N_15030,N_14894,N_14598);
nor U15031 (N_15031,N_14647,N_14641);
and U15032 (N_15032,N_14897,N_14745);
nor U15033 (N_15033,N_14918,N_14648);
xor U15034 (N_15034,N_14718,N_14969);
xor U15035 (N_15035,N_14880,N_14725);
nor U15036 (N_15036,N_14700,N_14820);
and U15037 (N_15037,N_14795,N_14844);
and U15038 (N_15038,N_14868,N_14759);
and U15039 (N_15039,N_14961,N_14657);
xor U15040 (N_15040,N_14890,N_14948);
nor U15041 (N_15041,N_14758,N_14895);
nor U15042 (N_15042,N_14937,N_14978);
or U15043 (N_15043,N_14804,N_14790);
and U15044 (N_15044,N_14595,N_14582);
and U15045 (N_15045,N_14789,N_14703);
nand U15046 (N_15046,N_14662,N_14870);
nor U15047 (N_15047,N_14716,N_14651);
or U15048 (N_15048,N_14908,N_14889);
xnor U15049 (N_15049,N_14738,N_14732);
nor U15050 (N_15050,N_14650,N_14968);
and U15051 (N_15051,N_14588,N_14971);
or U15052 (N_15052,N_14683,N_14678);
and U15053 (N_15053,N_14719,N_14556);
nor U15054 (N_15054,N_14501,N_14864);
nand U15055 (N_15055,N_14765,N_14569);
nor U15056 (N_15056,N_14543,N_14625);
and U15057 (N_15057,N_14851,N_14772);
or U15058 (N_15058,N_14552,N_14954);
nand U15059 (N_15059,N_14611,N_14862);
xnor U15060 (N_15060,N_14850,N_14981);
nor U15061 (N_15061,N_14551,N_14997);
or U15062 (N_15062,N_14592,N_14730);
or U15063 (N_15063,N_14801,N_14663);
nand U15064 (N_15064,N_14816,N_14548);
nand U15065 (N_15065,N_14882,N_14875);
nand U15066 (N_15066,N_14815,N_14570);
or U15067 (N_15067,N_14672,N_14915);
and U15068 (N_15068,N_14729,N_14585);
and U15069 (N_15069,N_14603,N_14559);
nor U15070 (N_15070,N_14898,N_14563);
nand U15071 (N_15071,N_14993,N_14931);
or U15072 (N_15072,N_14995,N_14896);
nor U15073 (N_15073,N_14658,N_14814);
nand U15074 (N_15074,N_14887,N_14760);
xnor U15075 (N_15075,N_14917,N_14787);
nand U15076 (N_15076,N_14813,N_14679);
or U15077 (N_15077,N_14610,N_14688);
nand U15078 (N_15078,N_14819,N_14622);
nor U15079 (N_15079,N_14989,N_14566);
nand U15080 (N_15080,N_14963,N_14901);
xor U15081 (N_15081,N_14825,N_14812);
nand U15082 (N_15082,N_14985,N_14926);
nor U15083 (N_15083,N_14539,N_14628);
or U15084 (N_15084,N_14635,N_14853);
nor U15085 (N_15085,N_14560,N_14692);
or U15086 (N_15086,N_14634,N_14544);
and U15087 (N_15087,N_14721,N_14823);
nor U15088 (N_15088,N_14506,N_14601);
xor U15089 (N_15089,N_14763,N_14964);
xor U15090 (N_15090,N_14514,N_14687);
and U15091 (N_15091,N_14966,N_14843);
xnor U15092 (N_15092,N_14715,N_14521);
and U15093 (N_15093,N_14974,N_14681);
nor U15094 (N_15094,N_14670,N_14652);
or U15095 (N_15095,N_14865,N_14699);
and U15096 (N_15096,N_14669,N_14932);
xor U15097 (N_15097,N_14925,N_14845);
and U15098 (N_15098,N_14527,N_14590);
nand U15099 (N_15099,N_14959,N_14504);
and U15100 (N_15100,N_14910,N_14661);
nor U15101 (N_15101,N_14701,N_14751);
xnor U15102 (N_15102,N_14659,N_14867);
nor U15103 (N_15103,N_14747,N_14637);
nand U15104 (N_15104,N_14860,N_14776);
nand U15105 (N_15105,N_14677,N_14855);
and U15106 (N_15106,N_14660,N_14710);
xor U15107 (N_15107,N_14877,N_14704);
and U15108 (N_15108,N_14593,N_14938);
xor U15109 (N_15109,N_14942,N_14972);
nand U15110 (N_15110,N_14568,N_14583);
nor U15111 (N_15111,N_14542,N_14798);
and U15112 (N_15112,N_14769,N_14824);
and U15113 (N_15113,N_14884,N_14723);
xnor U15114 (N_15114,N_14731,N_14785);
and U15115 (N_15115,N_14575,N_14535);
nand U15116 (N_15116,N_14606,N_14711);
or U15117 (N_15117,N_14676,N_14573);
xor U15118 (N_15118,N_14891,N_14698);
and U15119 (N_15119,N_14779,N_14511);
nor U15120 (N_15120,N_14892,N_14690);
nand U15121 (N_15121,N_14567,N_14649);
xor U15122 (N_15122,N_14965,N_14984);
xor U15123 (N_15123,N_14572,N_14854);
nand U15124 (N_15124,N_14671,N_14520);
xor U15125 (N_15125,N_14534,N_14643);
or U15126 (N_15126,N_14803,N_14944);
nand U15127 (N_15127,N_14802,N_14717);
nor U15128 (N_15128,N_14666,N_14754);
or U15129 (N_15129,N_14656,N_14653);
nand U15130 (N_15130,N_14513,N_14980);
nor U15131 (N_15131,N_14927,N_14952);
xnor U15132 (N_15132,N_14951,N_14970);
or U15133 (N_15133,N_14783,N_14674);
nor U15134 (N_15134,N_14904,N_14773);
and U15135 (N_15135,N_14784,N_14982);
and U15136 (N_15136,N_14722,N_14811);
nor U15137 (N_15137,N_14939,N_14858);
and U15138 (N_15138,N_14537,N_14998);
nor U15139 (N_15139,N_14591,N_14841);
or U15140 (N_15140,N_14667,N_14578);
xnor U15141 (N_15141,N_14720,N_14574);
nand U15142 (N_15142,N_14940,N_14605);
nor U15143 (N_15143,N_14553,N_14621);
nand U15144 (N_15144,N_14827,N_14757);
nor U15145 (N_15145,N_14706,N_14579);
or U15146 (N_15146,N_14693,N_14792);
nor U15147 (N_15147,N_14714,N_14818);
and U15148 (N_15148,N_14599,N_14909);
and U15149 (N_15149,N_14684,N_14538);
and U15150 (N_15150,N_14626,N_14771);
xnor U15151 (N_15151,N_14987,N_14873);
nand U15152 (N_15152,N_14531,N_14999);
or U15153 (N_15153,N_14800,N_14848);
or U15154 (N_15154,N_14967,N_14755);
xnor U15155 (N_15155,N_14929,N_14608);
or U15156 (N_15156,N_14517,N_14673);
and U15157 (N_15157,N_14616,N_14600);
or U15158 (N_15158,N_14636,N_14632);
or U15159 (N_15159,N_14797,N_14629);
nor U15160 (N_15160,N_14863,N_14597);
xnor U15161 (N_15161,N_14654,N_14878);
xnor U15162 (N_15162,N_14990,N_14645);
and U15163 (N_15163,N_14935,N_14613);
nand U15164 (N_15164,N_14509,N_14956);
and U15165 (N_15165,N_14565,N_14630);
nand U15166 (N_15166,N_14766,N_14644);
xnor U15167 (N_15167,N_14837,N_14829);
nand U15168 (N_15168,N_14576,N_14852);
nor U15169 (N_15169,N_14541,N_14886);
or U15170 (N_15170,N_14768,N_14883);
nand U15171 (N_15171,N_14532,N_14976);
nand U15172 (N_15172,N_14695,N_14612);
nor U15173 (N_15173,N_14508,N_14986);
and U15174 (N_15174,N_14596,N_14737);
nand U15175 (N_15175,N_14906,N_14817);
nor U15176 (N_15176,N_14555,N_14946);
nand U15177 (N_15177,N_14919,N_14540);
or U15178 (N_15178,N_14941,N_14584);
xnor U15179 (N_15179,N_14750,N_14840);
and U15180 (N_15180,N_14694,N_14557);
xnor U15181 (N_15181,N_14638,N_14713);
or U15182 (N_15182,N_14587,N_14761);
xor U15183 (N_15183,N_14955,N_14623);
and U15184 (N_15184,N_14943,N_14907);
xor U15185 (N_15185,N_14728,N_14911);
xnor U15186 (N_15186,N_14502,N_14834);
or U15187 (N_15187,N_14594,N_14522);
nor U15188 (N_15188,N_14627,N_14791);
and U15189 (N_15189,N_14736,N_14794);
or U15190 (N_15190,N_14614,N_14775);
and U15191 (N_15191,N_14561,N_14705);
or U15192 (N_15192,N_14633,N_14697);
or U15193 (N_15193,N_14903,N_14962);
xnor U15194 (N_15194,N_14624,N_14640);
or U15195 (N_15195,N_14826,N_14988);
and U15196 (N_15196,N_14960,N_14533);
nand U15197 (N_15197,N_14740,N_14580);
xnor U15198 (N_15198,N_14753,N_14949);
nand U15199 (N_15199,N_14756,N_14642);
and U15200 (N_15200,N_14899,N_14879);
or U15201 (N_15201,N_14836,N_14828);
and U15202 (N_15202,N_14778,N_14810);
nor U15203 (N_15203,N_14519,N_14646);
xnor U15204 (N_15204,N_14668,N_14696);
nor U15205 (N_15205,N_14609,N_14905);
xor U15206 (N_15206,N_14856,N_14739);
xor U15207 (N_15207,N_14743,N_14589);
nand U15208 (N_15208,N_14973,N_14545);
and U15209 (N_15209,N_14746,N_14764);
or U15210 (N_15210,N_14618,N_14707);
nor U15211 (N_15211,N_14912,N_14977);
or U15212 (N_15212,N_14607,N_14680);
xnor U15213 (N_15213,N_14702,N_14546);
nor U15214 (N_15214,N_14799,N_14518);
xor U15215 (N_15215,N_14777,N_14617);
nand U15216 (N_15216,N_14547,N_14920);
nand U15217 (N_15217,N_14770,N_14921);
or U15218 (N_15218,N_14874,N_14564);
or U15219 (N_15219,N_14708,N_14930);
or U15220 (N_15220,N_14619,N_14516);
nand U15221 (N_15221,N_14861,N_14675);
xnor U15222 (N_15222,N_14950,N_14554);
nor U15223 (N_15223,N_14505,N_14665);
nor U15224 (N_15224,N_14847,N_14604);
nand U15225 (N_15225,N_14734,N_14558);
or U15226 (N_15226,N_14831,N_14748);
nand U15227 (N_15227,N_14664,N_14953);
nand U15228 (N_15228,N_14934,N_14849);
nor U15229 (N_15229,N_14945,N_14524);
nand U15230 (N_15230,N_14724,N_14857);
nor U15231 (N_15231,N_14893,N_14571);
xnor U15232 (N_15232,N_14503,N_14727);
nor U15233 (N_15233,N_14822,N_14655);
xnor U15234 (N_15234,N_14735,N_14526);
nor U15235 (N_15235,N_14752,N_14682);
nand U15236 (N_15236,N_14872,N_14996);
nand U15237 (N_15237,N_14923,N_14781);
and U15238 (N_15238,N_14928,N_14806);
xor U15239 (N_15239,N_14512,N_14741);
xnor U15240 (N_15240,N_14762,N_14994);
and U15241 (N_15241,N_14888,N_14924);
xnor U15242 (N_15242,N_14979,N_14515);
or U15243 (N_15243,N_14744,N_14549);
nand U15244 (N_15244,N_14866,N_14936);
or U15245 (N_15245,N_14691,N_14947);
or U15246 (N_15246,N_14991,N_14838);
or U15247 (N_15247,N_14749,N_14933);
xor U15248 (N_15248,N_14796,N_14529);
xor U15249 (N_15249,N_14550,N_14689);
xor U15250 (N_15250,N_14705,N_14734);
and U15251 (N_15251,N_14545,N_14908);
nand U15252 (N_15252,N_14606,N_14645);
nand U15253 (N_15253,N_14924,N_14928);
xor U15254 (N_15254,N_14914,N_14739);
or U15255 (N_15255,N_14988,N_14944);
xnor U15256 (N_15256,N_14619,N_14853);
nand U15257 (N_15257,N_14678,N_14650);
nand U15258 (N_15258,N_14957,N_14606);
xor U15259 (N_15259,N_14913,N_14926);
and U15260 (N_15260,N_14897,N_14550);
nand U15261 (N_15261,N_14835,N_14757);
xnor U15262 (N_15262,N_14544,N_14593);
or U15263 (N_15263,N_14724,N_14909);
and U15264 (N_15264,N_14797,N_14618);
nor U15265 (N_15265,N_14799,N_14889);
xor U15266 (N_15266,N_14616,N_14542);
xor U15267 (N_15267,N_14966,N_14614);
or U15268 (N_15268,N_14723,N_14826);
nand U15269 (N_15269,N_14569,N_14940);
nor U15270 (N_15270,N_14915,N_14558);
or U15271 (N_15271,N_14967,N_14578);
or U15272 (N_15272,N_14893,N_14538);
or U15273 (N_15273,N_14634,N_14972);
nand U15274 (N_15274,N_14512,N_14902);
xor U15275 (N_15275,N_14762,N_14660);
nand U15276 (N_15276,N_14774,N_14712);
nor U15277 (N_15277,N_14679,N_14559);
and U15278 (N_15278,N_14576,N_14580);
or U15279 (N_15279,N_14524,N_14753);
nor U15280 (N_15280,N_14669,N_14878);
nand U15281 (N_15281,N_14731,N_14720);
xor U15282 (N_15282,N_14988,N_14870);
or U15283 (N_15283,N_14810,N_14631);
or U15284 (N_15284,N_14834,N_14920);
and U15285 (N_15285,N_14763,N_14540);
and U15286 (N_15286,N_14600,N_14980);
nor U15287 (N_15287,N_14881,N_14706);
or U15288 (N_15288,N_14918,N_14732);
nand U15289 (N_15289,N_14829,N_14722);
or U15290 (N_15290,N_14720,N_14756);
or U15291 (N_15291,N_14697,N_14551);
xnor U15292 (N_15292,N_14890,N_14643);
or U15293 (N_15293,N_14937,N_14995);
xnor U15294 (N_15294,N_14569,N_14646);
xor U15295 (N_15295,N_14835,N_14751);
nand U15296 (N_15296,N_14694,N_14971);
or U15297 (N_15297,N_14655,N_14967);
nor U15298 (N_15298,N_14788,N_14681);
nand U15299 (N_15299,N_14624,N_14852);
nand U15300 (N_15300,N_14868,N_14935);
or U15301 (N_15301,N_14948,N_14999);
and U15302 (N_15302,N_14691,N_14900);
xnor U15303 (N_15303,N_14811,N_14907);
nand U15304 (N_15304,N_14528,N_14987);
nor U15305 (N_15305,N_14831,N_14524);
nor U15306 (N_15306,N_14854,N_14798);
and U15307 (N_15307,N_14792,N_14735);
or U15308 (N_15308,N_14731,N_14953);
or U15309 (N_15309,N_14510,N_14525);
or U15310 (N_15310,N_14840,N_14524);
or U15311 (N_15311,N_14912,N_14947);
and U15312 (N_15312,N_14818,N_14986);
xor U15313 (N_15313,N_14920,N_14702);
xnor U15314 (N_15314,N_14977,N_14767);
or U15315 (N_15315,N_14520,N_14970);
nor U15316 (N_15316,N_14689,N_14778);
and U15317 (N_15317,N_14955,N_14980);
and U15318 (N_15318,N_14973,N_14856);
and U15319 (N_15319,N_14633,N_14824);
nand U15320 (N_15320,N_14817,N_14857);
and U15321 (N_15321,N_14907,N_14626);
nand U15322 (N_15322,N_14674,N_14851);
or U15323 (N_15323,N_14812,N_14879);
xnor U15324 (N_15324,N_14620,N_14521);
and U15325 (N_15325,N_14592,N_14879);
nand U15326 (N_15326,N_14564,N_14993);
and U15327 (N_15327,N_14584,N_14630);
nand U15328 (N_15328,N_14788,N_14927);
xor U15329 (N_15329,N_14520,N_14985);
nand U15330 (N_15330,N_14543,N_14787);
nor U15331 (N_15331,N_14598,N_14766);
xnor U15332 (N_15332,N_14517,N_14575);
and U15333 (N_15333,N_14934,N_14857);
nand U15334 (N_15334,N_14501,N_14517);
xnor U15335 (N_15335,N_14703,N_14846);
nor U15336 (N_15336,N_14785,N_14989);
nand U15337 (N_15337,N_14881,N_14920);
nand U15338 (N_15338,N_14541,N_14576);
and U15339 (N_15339,N_14803,N_14937);
xor U15340 (N_15340,N_14941,N_14668);
nor U15341 (N_15341,N_14831,N_14557);
xor U15342 (N_15342,N_14524,N_14771);
nor U15343 (N_15343,N_14508,N_14703);
xor U15344 (N_15344,N_14745,N_14812);
nor U15345 (N_15345,N_14606,N_14559);
nand U15346 (N_15346,N_14998,N_14811);
and U15347 (N_15347,N_14803,N_14611);
nand U15348 (N_15348,N_14767,N_14868);
or U15349 (N_15349,N_14794,N_14969);
and U15350 (N_15350,N_14592,N_14917);
xor U15351 (N_15351,N_14594,N_14645);
xnor U15352 (N_15352,N_14741,N_14591);
or U15353 (N_15353,N_14957,N_14766);
nor U15354 (N_15354,N_14611,N_14573);
or U15355 (N_15355,N_14512,N_14929);
and U15356 (N_15356,N_14695,N_14857);
and U15357 (N_15357,N_14608,N_14711);
xor U15358 (N_15358,N_14804,N_14672);
xor U15359 (N_15359,N_14539,N_14778);
nor U15360 (N_15360,N_14789,N_14668);
nand U15361 (N_15361,N_14853,N_14929);
nand U15362 (N_15362,N_14875,N_14684);
and U15363 (N_15363,N_14636,N_14748);
xnor U15364 (N_15364,N_14830,N_14559);
xnor U15365 (N_15365,N_14713,N_14543);
xor U15366 (N_15366,N_14564,N_14715);
nor U15367 (N_15367,N_14709,N_14537);
nand U15368 (N_15368,N_14908,N_14750);
and U15369 (N_15369,N_14917,N_14565);
and U15370 (N_15370,N_14697,N_14624);
xnor U15371 (N_15371,N_14816,N_14945);
nor U15372 (N_15372,N_14576,N_14958);
xnor U15373 (N_15373,N_14588,N_14808);
or U15374 (N_15374,N_14854,N_14818);
and U15375 (N_15375,N_14893,N_14624);
and U15376 (N_15376,N_14511,N_14896);
or U15377 (N_15377,N_14941,N_14528);
nor U15378 (N_15378,N_14831,N_14961);
and U15379 (N_15379,N_14745,N_14596);
and U15380 (N_15380,N_14960,N_14736);
and U15381 (N_15381,N_14777,N_14690);
nand U15382 (N_15382,N_14958,N_14517);
nand U15383 (N_15383,N_14681,N_14781);
nor U15384 (N_15384,N_14535,N_14805);
nand U15385 (N_15385,N_14952,N_14594);
nor U15386 (N_15386,N_14631,N_14740);
xnor U15387 (N_15387,N_14501,N_14673);
xor U15388 (N_15388,N_14676,N_14554);
nand U15389 (N_15389,N_14794,N_14607);
nor U15390 (N_15390,N_14642,N_14686);
or U15391 (N_15391,N_14796,N_14628);
nand U15392 (N_15392,N_14639,N_14887);
nor U15393 (N_15393,N_14741,N_14537);
or U15394 (N_15394,N_14771,N_14575);
nor U15395 (N_15395,N_14787,N_14843);
nor U15396 (N_15396,N_14917,N_14550);
and U15397 (N_15397,N_14639,N_14975);
and U15398 (N_15398,N_14569,N_14598);
nor U15399 (N_15399,N_14740,N_14675);
nor U15400 (N_15400,N_14875,N_14970);
or U15401 (N_15401,N_14861,N_14712);
or U15402 (N_15402,N_14876,N_14920);
nor U15403 (N_15403,N_14750,N_14672);
nor U15404 (N_15404,N_14766,N_14889);
nand U15405 (N_15405,N_14725,N_14520);
nor U15406 (N_15406,N_14893,N_14917);
and U15407 (N_15407,N_14697,N_14692);
and U15408 (N_15408,N_14659,N_14802);
or U15409 (N_15409,N_14969,N_14607);
and U15410 (N_15410,N_14889,N_14768);
or U15411 (N_15411,N_14842,N_14634);
and U15412 (N_15412,N_14664,N_14973);
xor U15413 (N_15413,N_14585,N_14824);
xnor U15414 (N_15414,N_14992,N_14931);
nor U15415 (N_15415,N_14546,N_14531);
or U15416 (N_15416,N_14972,N_14807);
nor U15417 (N_15417,N_14500,N_14700);
nand U15418 (N_15418,N_14835,N_14865);
nand U15419 (N_15419,N_14900,N_14977);
nor U15420 (N_15420,N_14895,N_14841);
nand U15421 (N_15421,N_14761,N_14565);
xor U15422 (N_15422,N_14564,N_14729);
or U15423 (N_15423,N_14619,N_14730);
xor U15424 (N_15424,N_14718,N_14765);
nor U15425 (N_15425,N_14622,N_14769);
nor U15426 (N_15426,N_14806,N_14785);
or U15427 (N_15427,N_14783,N_14513);
xor U15428 (N_15428,N_14996,N_14914);
xor U15429 (N_15429,N_14545,N_14711);
nand U15430 (N_15430,N_14633,N_14720);
nand U15431 (N_15431,N_14707,N_14573);
nor U15432 (N_15432,N_14722,N_14698);
nor U15433 (N_15433,N_14906,N_14605);
nor U15434 (N_15434,N_14936,N_14789);
and U15435 (N_15435,N_14521,N_14909);
or U15436 (N_15436,N_14647,N_14855);
and U15437 (N_15437,N_14643,N_14967);
nor U15438 (N_15438,N_14911,N_14667);
and U15439 (N_15439,N_14893,N_14740);
and U15440 (N_15440,N_14580,N_14666);
nor U15441 (N_15441,N_14738,N_14974);
nor U15442 (N_15442,N_14600,N_14761);
and U15443 (N_15443,N_14640,N_14634);
xor U15444 (N_15444,N_14828,N_14929);
or U15445 (N_15445,N_14547,N_14698);
or U15446 (N_15446,N_14660,N_14921);
and U15447 (N_15447,N_14837,N_14878);
or U15448 (N_15448,N_14758,N_14872);
and U15449 (N_15449,N_14700,N_14646);
nand U15450 (N_15450,N_14505,N_14675);
xor U15451 (N_15451,N_14537,N_14885);
xnor U15452 (N_15452,N_14789,N_14579);
and U15453 (N_15453,N_14611,N_14632);
and U15454 (N_15454,N_14947,N_14951);
nor U15455 (N_15455,N_14600,N_14936);
nand U15456 (N_15456,N_14848,N_14979);
or U15457 (N_15457,N_14946,N_14506);
nand U15458 (N_15458,N_14896,N_14504);
and U15459 (N_15459,N_14522,N_14524);
and U15460 (N_15460,N_14564,N_14822);
nand U15461 (N_15461,N_14966,N_14555);
or U15462 (N_15462,N_14845,N_14959);
and U15463 (N_15463,N_14844,N_14656);
or U15464 (N_15464,N_14610,N_14756);
or U15465 (N_15465,N_14854,N_14847);
nand U15466 (N_15466,N_14752,N_14558);
xnor U15467 (N_15467,N_14761,N_14811);
or U15468 (N_15468,N_14954,N_14709);
xor U15469 (N_15469,N_14557,N_14684);
and U15470 (N_15470,N_14728,N_14894);
or U15471 (N_15471,N_14976,N_14956);
nand U15472 (N_15472,N_14843,N_14973);
nand U15473 (N_15473,N_14930,N_14993);
nor U15474 (N_15474,N_14778,N_14739);
and U15475 (N_15475,N_14686,N_14913);
or U15476 (N_15476,N_14520,N_14714);
nand U15477 (N_15477,N_14784,N_14712);
nand U15478 (N_15478,N_14584,N_14602);
and U15479 (N_15479,N_14781,N_14524);
xnor U15480 (N_15480,N_14822,N_14536);
xor U15481 (N_15481,N_14661,N_14644);
xnor U15482 (N_15482,N_14742,N_14682);
nand U15483 (N_15483,N_14811,N_14904);
nand U15484 (N_15484,N_14621,N_14769);
nor U15485 (N_15485,N_14907,N_14523);
nor U15486 (N_15486,N_14583,N_14641);
nor U15487 (N_15487,N_14695,N_14729);
xnor U15488 (N_15488,N_14900,N_14642);
xnor U15489 (N_15489,N_14742,N_14944);
or U15490 (N_15490,N_14587,N_14920);
or U15491 (N_15491,N_14541,N_14970);
nor U15492 (N_15492,N_14708,N_14923);
xor U15493 (N_15493,N_14803,N_14879);
nand U15494 (N_15494,N_14741,N_14897);
nand U15495 (N_15495,N_14510,N_14996);
nand U15496 (N_15496,N_14827,N_14969);
xnor U15497 (N_15497,N_14706,N_14806);
and U15498 (N_15498,N_14788,N_14558);
and U15499 (N_15499,N_14812,N_14602);
xnor U15500 (N_15500,N_15061,N_15014);
nand U15501 (N_15501,N_15112,N_15193);
xor U15502 (N_15502,N_15370,N_15135);
nor U15503 (N_15503,N_15401,N_15448);
xor U15504 (N_15504,N_15047,N_15085);
or U15505 (N_15505,N_15341,N_15044);
or U15506 (N_15506,N_15372,N_15146);
xor U15507 (N_15507,N_15223,N_15130);
and U15508 (N_15508,N_15490,N_15423);
xor U15509 (N_15509,N_15159,N_15081);
and U15510 (N_15510,N_15455,N_15416);
xnor U15511 (N_15511,N_15183,N_15017);
nor U15512 (N_15512,N_15400,N_15331);
and U15513 (N_15513,N_15247,N_15351);
nor U15514 (N_15514,N_15322,N_15239);
nand U15515 (N_15515,N_15116,N_15140);
nor U15516 (N_15516,N_15025,N_15069);
and U15517 (N_15517,N_15035,N_15408);
nand U15518 (N_15518,N_15115,N_15127);
nand U15519 (N_15519,N_15361,N_15210);
nand U15520 (N_15520,N_15198,N_15218);
nor U15521 (N_15521,N_15093,N_15141);
and U15522 (N_15522,N_15214,N_15373);
and U15523 (N_15523,N_15386,N_15224);
xor U15524 (N_15524,N_15182,N_15487);
nand U15525 (N_15525,N_15005,N_15368);
and U15526 (N_15526,N_15407,N_15104);
nor U15527 (N_15527,N_15212,N_15273);
nand U15528 (N_15528,N_15421,N_15467);
nand U15529 (N_15529,N_15452,N_15462);
and U15530 (N_15530,N_15028,N_15250);
and U15531 (N_15531,N_15275,N_15158);
and U15532 (N_15532,N_15260,N_15283);
nand U15533 (N_15533,N_15216,N_15168);
nor U15534 (N_15534,N_15279,N_15219);
xor U15535 (N_15535,N_15200,N_15019);
nor U15536 (N_15536,N_15466,N_15165);
nand U15537 (N_15537,N_15229,N_15397);
and U15538 (N_15538,N_15052,N_15011);
nor U15539 (N_15539,N_15123,N_15021);
xor U15540 (N_15540,N_15330,N_15381);
xor U15541 (N_15541,N_15451,N_15306);
nand U15542 (N_15542,N_15184,N_15226);
nand U15543 (N_15543,N_15084,N_15196);
or U15544 (N_15544,N_15228,N_15109);
or U15545 (N_15545,N_15234,N_15142);
and U15546 (N_15546,N_15113,N_15072);
nor U15547 (N_15547,N_15179,N_15491);
xnor U15548 (N_15548,N_15237,N_15268);
nor U15549 (N_15549,N_15043,N_15495);
nand U15550 (N_15550,N_15269,N_15354);
nor U15551 (N_15551,N_15288,N_15075);
and U15552 (N_15552,N_15329,N_15101);
nor U15553 (N_15553,N_15076,N_15441);
nand U15554 (N_15554,N_15055,N_15255);
or U15555 (N_15555,N_15050,N_15257);
nor U15556 (N_15556,N_15111,N_15024);
nor U15557 (N_15557,N_15305,N_15468);
or U15558 (N_15558,N_15125,N_15298);
or U15559 (N_15559,N_15153,N_15436);
or U15560 (N_15560,N_15427,N_15340);
xnor U15561 (N_15561,N_15256,N_15089);
and U15562 (N_15562,N_15435,N_15432);
xnor U15563 (N_15563,N_15302,N_15151);
nand U15564 (N_15564,N_15190,N_15059);
nand U15565 (N_15565,N_15001,N_15133);
nand U15566 (N_15566,N_15039,N_15171);
xnor U15567 (N_15567,N_15128,N_15197);
and U15568 (N_15568,N_15456,N_15316);
nand U15569 (N_15569,N_15206,N_15164);
nand U15570 (N_15570,N_15387,N_15012);
nand U15571 (N_15571,N_15318,N_15308);
nor U15572 (N_15572,N_15339,N_15355);
xor U15573 (N_15573,N_15481,N_15174);
nor U15574 (N_15574,N_15424,N_15057);
nand U15575 (N_15575,N_15328,N_15178);
nand U15576 (N_15576,N_15319,N_15307);
xnor U15577 (N_15577,N_15254,N_15045);
or U15578 (N_15578,N_15494,N_15327);
nor U15579 (N_15579,N_15120,N_15415);
or U15580 (N_15580,N_15169,N_15071);
and U15581 (N_15581,N_15332,N_15137);
nand U15582 (N_15582,N_15033,N_15476);
xor U15583 (N_15583,N_15412,N_15244);
nand U15584 (N_15584,N_15110,N_15439);
and U15585 (N_15585,N_15315,N_15245);
nand U15586 (N_15586,N_15067,N_15027);
nor U15587 (N_15587,N_15073,N_15472);
nand U15588 (N_15588,N_15366,N_15095);
nand U15589 (N_15589,N_15484,N_15003);
and U15590 (N_15590,N_15249,N_15395);
and U15591 (N_15591,N_15099,N_15020);
nor U15592 (N_15592,N_15409,N_15492);
xnor U15593 (N_15593,N_15177,N_15459);
or U15594 (N_15594,N_15480,N_15195);
and U15595 (N_15595,N_15263,N_15356);
xor U15596 (N_15596,N_15393,N_15161);
and U15597 (N_15597,N_15488,N_15342);
or U15598 (N_15598,N_15499,N_15231);
nand U15599 (N_15599,N_15261,N_15392);
nand U15600 (N_15600,N_15438,N_15497);
nand U15601 (N_15601,N_15086,N_15363);
nand U15602 (N_15602,N_15360,N_15049);
xnor U15603 (N_15603,N_15469,N_15388);
nor U15604 (N_15604,N_15292,N_15227);
xor U15605 (N_15605,N_15060,N_15425);
nor U15606 (N_15606,N_15270,N_15037);
nor U15607 (N_15607,N_15294,N_15242);
or U15608 (N_15608,N_15262,N_15038);
nor U15609 (N_15609,N_15285,N_15258);
xor U15610 (N_15610,N_15384,N_15296);
or U15611 (N_15611,N_15148,N_15192);
nand U15612 (N_15612,N_15465,N_15325);
xor U15613 (N_15613,N_15383,N_15326);
nand U15614 (N_15614,N_15471,N_15320);
nor U15615 (N_15615,N_15016,N_15083);
nand U15616 (N_15616,N_15442,N_15188);
or U15617 (N_15617,N_15313,N_15413);
nand U15618 (N_15618,N_15473,N_15460);
or U15619 (N_15619,N_15353,N_15345);
nand U15620 (N_15620,N_15160,N_15176);
nand U15621 (N_15621,N_15008,N_15002);
or U15622 (N_15622,N_15241,N_15291);
xor U15623 (N_15623,N_15121,N_15139);
nand U15624 (N_15624,N_15034,N_15079);
nor U15625 (N_15625,N_15259,N_15031);
nor U15626 (N_15626,N_15352,N_15478);
or U15627 (N_15627,N_15369,N_15201);
xnor U15628 (N_15628,N_15129,N_15006);
nor U15629 (N_15629,N_15007,N_15194);
xnor U15630 (N_15630,N_15280,N_15185);
nand U15631 (N_15631,N_15350,N_15243);
nand U15632 (N_15632,N_15082,N_15236);
or U15633 (N_15633,N_15094,N_15170);
and U15634 (N_15634,N_15264,N_15321);
and U15635 (N_15635,N_15347,N_15180);
or U15636 (N_15636,N_15163,N_15064);
nor U15637 (N_15637,N_15453,N_15138);
xor U15638 (N_15638,N_15364,N_15222);
and U15639 (N_15639,N_15394,N_15359);
or U15640 (N_15640,N_15404,N_15205);
nor U15641 (N_15641,N_15235,N_15346);
and U15642 (N_15642,N_15398,N_15091);
nor U15643 (N_15643,N_15217,N_15040);
nand U15644 (N_15644,N_15150,N_15365);
xor U15645 (N_15645,N_15446,N_15252);
nor U15646 (N_15646,N_15225,N_15117);
nor U15647 (N_15647,N_15207,N_15181);
nand U15648 (N_15648,N_15131,N_15303);
and U15649 (N_15649,N_15406,N_15100);
and U15650 (N_15650,N_15434,N_15209);
nor U15651 (N_15651,N_15385,N_15248);
nand U15652 (N_15652,N_15013,N_15486);
nor U15653 (N_15653,N_15087,N_15444);
and U15654 (N_15654,N_15417,N_15042);
xnor U15655 (N_15655,N_15167,N_15375);
nor U15656 (N_15656,N_15000,N_15485);
nand U15657 (N_15657,N_15274,N_15030);
nor U15658 (N_15658,N_15475,N_15483);
or U15659 (N_15659,N_15310,N_15051);
xnor U15660 (N_15660,N_15286,N_15058);
or U15661 (N_15661,N_15232,N_15080);
or U15662 (N_15662,N_15114,N_15389);
nand U15663 (N_15663,N_15449,N_15119);
or U15664 (N_15664,N_15103,N_15284);
and U15665 (N_15665,N_15046,N_15102);
xor U15666 (N_15666,N_15238,N_15134);
nand U15667 (N_15667,N_15418,N_15070);
nor U15668 (N_15668,N_15063,N_15479);
or U15669 (N_15669,N_15374,N_15297);
and U15670 (N_15670,N_15144,N_15272);
and U15671 (N_15671,N_15199,N_15376);
or U15672 (N_15672,N_15186,N_15032);
xor U15673 (N_15673,N_15379,N_15036);
or U15674 (N_15674,N_15145,N_15162);
xnor U15675 (N_15675,N_15090,N_15010);
and U15676 (N_15676,N_15204,N_15166);
and U15677 (N_15677,N_15132,N_15411);
nand U15678 (N_15678,N_15240,N_15362);
nand U15679 (N_15679,N_15477,N_15429);
xor U15680 (N_15680,N_15251,N_15314);
nor U15681 (N_15681,N_15018,N_15276);
xnor U15682 (N_15682,N_15191,N_15382);
and U15683 (N_15683,N_15147,N_15155);
or U15684 (N_15684,N_15221,N_15498);
or U15685 (N_15685,N_15312,N_15414);
and U15686 (N_15686,N_15367,N_15311);
or U15687 (N_15687,N_15143,N_15334);
or U15688 (N_15688,N_15287,N_15349);
or U15689 (N_15689,N_15066,N_15092);
and U15690 (N_15690,N_15156,N_15097);
nor U15691 (N_15691,N_15358,N_15157);
nand U15692 (N_15692,N_15396,N_15175);
xor U15693 (N_15693,N_15278,N_15056);
xor U15694 (N_15694,N_15420,N_15445);
or U15695 (N_15695,N_15317,N_15450);
or U15696 (N_15696,N_15323,N_15405);
xor U15697 (N_15697,N_15062,N_15118);
nand U15698 (N_15698,N_15422,N_15246);
or U15699 (N_15699,N_15344,N_15428);
nand U15700 (N_15700,N_15403,N_15433);
nand U15701 (N_15701,N_15022,N_15324);
or U15702 (N_15702,N_15202,N_15293);
and U15703 (N_15703,N_15458,N_15220);
xor U15704 (N_15704,N_15464,N_15333);
or U15705 (N_15705,N_15074,N_15009);
and U15706 (N_15706,N_15440,N_15096);
nor U15707 (N_15707,N_15004,N_15402);
and U15708 (N_15708,N_15053,N_15489);
nor U15709 (N_15709,N_15437,N_15187);
and U15710 (N_15710,N_15189,N_15309);
nand U15711 (N_15711,N_15271,N_15172);
and U15712 (N_15712,N_15474,N_15122);
nand U15713 (N_15713,N_15290,N_15300);
nor U15714 (N_15714,N_15496,N_15267);
nand U15715 (N_15715,N_15108,N_15088);
xor U15716 (N_15716,N_15265,N_15447);
or U15717 (N_15717,N_15041,N_15335);
nand U15718 (N_15718,N_15431,N_15152);
or U15719 (N_15719,N_15301,N_15105);
or U15720 (N_15720,N_15211,N_15023);
xor U15721 (N_15721,N_15338,N_15233);
nor U15722 (N_15722,N_15281,N_15493);
nand U15723 (N_15723,N_15289,N_15430);
or U15724 (N_15724,N_15173,N_15295);
nand U15725 (N_15725,N_15098,N_15282);
xnor U15726 (N_15726,N_15378,N_15337);
nor U15727 (N_15727,N_15077,N_15371);
and U15728 (N_15728,N_15348,N_15463);
xnor U15729 (N_15729,N_15215,N_15299);
and U15730 (N_15730,N_15107,N_15029);
nand U15731 (N_15731,N_15277,N_15336);
and U15732 (N_15732,N_15343,N_15136);
nand U15733 (N_15733,N_15410,N_15304);
nand U15734 (N_15734,N_15419,N_15357);
xor U15735 (N_15735,N_15454,N_15203);
or U15736 (N_15736,N_15253,N_15154);
and U15737 (N_15737,N_15482,N_15208);
and U15738 (N_15738,N_15078,N_15054);
nand U15739 (N_15739,N_15149,N_15426);
or U15740 (N_15740,N_15380,N_15461);
nor U15741 (N_15741,N_15457,N_15213);
and U15742 (N_15742,N_15026,N_15065);
nor U15743 (N_15743,N_15399,N_15391);
nor U15744 (N_15744,N_15048,N_15068);
nor U15745 (N_15745,N_15106,N_15377);
nand U15746 (N_15746,N_15266,N_15015);
nor U15747 (N_15747,N_15230,N_15470);
xnor U15748 (N_15748,N_15443,N_15390);
or U15749 (N_15749,N_15124,N_15126);
nor U15750 (N_15750,N_15496,N_15401);
xor U15751 (N_15751,N_15020,N_15495);
and U15752 (N_15752,N_15045,N_15197);
nor U15753 (N_15753,N_15248,N_15480);
xor U15754 (N_15754,N_15048,N_15093);
xor U15755 (N_15755,N_15109,N_15191);
nand U15756 (N_15756,N_15359,N_15122);
and U15757 (N_15757,N_15343,N_15472);
nor U15758 (N_15758,N_15008,N_15459);
xnor U15759 (N_15759,N_15298,N_15404);
or U15760 (N_15760,N_15257,N_15013);
xor U15761 (N_15761,N_15368,N_15344);
nor U15762 (N_15762,N_15283,N_15228);
xor U15763 (N_15763,N_15084,N_15303);
xor U15764 (N_15764,N_15266,N_15279);
and U15765 (N_15765,N_15362,N_15170);
or U15766 (N_15766,N_15021,N_15371);
and U15767 (N_15767,N_15317,N_15154);
nand U15768 (N_15768,N_15156,N_15288);
or U15769 (N_15769,N_15067,N_15399);
nor U15770 (N_15770,N_15490,N_15122);
and U15771 (N_15771,N_15166,N_15317);
xor U15772 (N_15772,N_15285,N_15441);
or U15773 (N_15773,N_15178,N_15393);
nand U15774 (N_15774,N_15205,N_15428);
nand U15775 (N_15775,N_15439,N_15423);
xor U15776 (N_15776,N_15156,N_15039);
xnor U15777 (N_15777,N_15392,N_15218);
xnor U15778 (N_15778,N_15180,N_15087);
nand U15779 (N_15779,N_15067,N_15003);
and U15780 (N_15780,N_15335,N_15157);
nand U15781 (N_15781,N_15100,N_15314);
nor U15782 (N_15782,N_15099,N_15208);
and U15783 (N_15783,N_15101,N_15398);
nor U15784 (N_15784,N_15490,N_15081);
or U15785 (N_15785,N_15357,N_15463);
xor U15786 (N_15786,N_15334,N_15361);
or U15787 (N_15787,N_15358,N_15219);
or U15788 (N_15788,N_15339,N_15273);
and U15789 (N_15789,N_15053,N_15008);
nand U15790 (N_15790,N_15265,N_15362);
nor U15791 (N_15791,N_15063,N_15104);
and U15792 (N_15792,N_15020,N_15467);
and U15793 (N_15793,N_15476,N_15471);
nor U15794 (N_15794,N_15195,N_15345);
or U15795 (N_15795,N_15243,N_15044);
xnor U15796 (N_15796,N_15206,N_15293);
or U15797 (N_15797,N_15237,N_15259);
nor U15798 (N_15798,N_15268,N_15058);
or U15799 (N_15799,N_15264,N_15233);
xor U15800 (N_15800,N_15134,N_15467);
and U15801 (N_15801,N_15228,N_15344);
nand U15802 (N_15802,N_15477,N_15090);
nand U15803 (N_15803,N_15223,N_15119);
xor U15804 (N_15804,N_15471,N_15285);
nand U15805 (N_15805,N_15039,N_15168);
or U15806 (N_15806,N_15416,N_15305);
or U15807 (N_15807,N_15316,N_15337);
nand U15808 (N_15808,N_15280,N_15089);
xor U15809 (N_15809,N_15407,N_15304);
or U15810 (N_15810,N_15384,N_15369);
nand U15811 (N_15811,N_15416,N_15189);
and U15812 (N_15812,N_15458,N_15415);
nor U15813 (N_15813,N_15250,N_15258);
xor U15814 (N_15814,N_15292,N_15340);
nand U15815 (N_15815,N_15225,N_15476);
xnor U15816 (N_15816,N_15388,N_15177);
xor U15817 (N_15817,N_15282,N_15421);
xnor U15818 (N_15818,N_15326,N_15082);
or U15819 (N_15819,N_15170,N_15229);
nor U15820 (N_15820,N_15411,N_15412);
nand U15821 (N_15821,N_15483,N_15305);
and U15822 (N_15822,N_15257,N_15464);
xnor U15823 (N_15823,N_15437,N_15118);
and U15824 (N_15824,N_15228,N_15150);
xor U15825 (N_15825,N_15126,N_15075);
and U15826 (N_15826,N_15187,N_15129);
xnor U15827 (N_15827,N_15467,N_15439);
xor U15828 (N_15828,N_15489,N_15163);
xnor U15829 (N_15829,N_15495,N_15247);
xnor U15830 (N_15830,N_15175,N_15119);
xnor U15831 (N_15831,N_15392,N_15120);
nand U15832 (N_15832,N_15452,N_15232);
nor U15833 (N_15833,N_15141,N_15209);
nand U15834 (N_15834,N_15184,N_15166);
xor U15835 (N_15835,N_15081,N_15043);
nor U15836 (N_15836,N_15428,N_15272);
nand U15837 (N_15837,N_15144,N_15425);
nor U15838 (N_15838,N_15430,N_15284);
and U15839 (N_15839,N_15445,N_15348);
xnor U15840 (N_15840,N_15116,N_15185);
nand U15841 (N_15841,N_15197,N_15212);
xnor U15842 (N_15842,N_15298,N_15266);
and U15843 (N_15843,N_15030,N_15314);
or U15844 (N_15844,N_15176,N_15125);
xnor U15845 (N_15845,N_15336,N_15106);
and U15846 (N_15846,N_15246,N_15261);
or U15847 (N_15847,N_15273,N_15168);
and U15848 (N_15848,N_15016,N_15076);
nor U15849 (N_15849,N_15147,N_15217);
xor U15850 (N_15850,N_15029,N_15317);
nor U15851 (N_15851,N_15253,N_15242);
nor U15852 (N_15852,N_15269,N_15288);
xnor U15853 (N_15853,N_15164,N_15221);
nor U15854 (N_15854,N_15245,N_15314);
and U15855 (N_15855,N_15496,N_15114);
or U15856 (N_15856,N_15339,N_15054);
nand U15857 (N_15857,N_15299,N_15122);
or U15858 (N_15858,N_15133,N_15209);
nor U15859 (N_15859,N_15120,N_15090);
and U15860 (N_15860,N_15270,N_15265);
xnor U15861 (N_15861,N_15426,N_15268);
nor U15862 (N_15862,N_15139,N_15097);
xnor U15863 (N_15863,N_15074,N_15086);
nand U15864 (N_15864,N_15162,N_15449);
nor U15865 (N_15865,N_15410,N_15359);
and U15866 (N_15866,N_15497,N_15371);
xnor U15867 (N_15867,N_15348,N_15014);
and U15868 (N_15868,N_15261,N_15322);
nor U15869 (N_15869,N_15240,N_15117);
and U15870 (N_15870,N_15397,N_15075);
xnor U15871 (N_15871,N_15101,N_15126);
nand U15872 (N_15872,N_15096,N_15227);
or U15873 (N_15873,N_15276,N_15190);
nand U15874 (N_15874,N_15317,N_15111);
nand U15875 (N_15875,N_15016,N_15430);
and U15876 (N_15876,N_15356,N_15331);
nor U15877 (N_15877,N_15087,N_15381);
nand U15878 (N_15878,N_15369,N_15158);
nor U15879 (N_15879,N_15267,N_15084);
nor U15880 (N_15880,N_15374,N_15474);
or U15881 (N_15881,N_15268,N_15096);
nand U15882 (N_15882,N_15489,N_15439);
and U15883 (N_15883,N_15394,N_15442);
xor U15884 (N_15884,N_15443,N_15340);
nor U15885 (N_15885,N_15274,N_15298);
nand U15886 (N_15886,N_15255,N_15160);
nor U15887 (N_15887,N_15020,N_15308);
nor U15888 (N_15888,N_15061,N_15033);
nor U15889 (N_15889,N_15443,N_15290);
or U15890 (N_15890,N_15247,N_15340);
nor U15891 (N_15891,N_15007,N_15051);
nand U15892 (N_15892,N_15004,N_15016);
nor U15893 (N_15893,N_15042,N_15298);
xnor U15894 (N_15894,N_15138,N_15125);
nand U15895 (N_15895,N_15192,N_15305);
and U15896 (N_15896,N_15076,N_15461);
and U15897 (N_15897,N_15132,N_15307);
nand U15898 (N_15898,N_15053,N_15323);
nand U15899 (N_15899,N_15156,N_15133);
nand U15900 (N_15900,N_15216,N_15353);
nand U15901 (N_15901,N_15444,N_15411);
nor U15902 (N_15902,N_15306,N_15153);
or U15903 (N_15903,N_15131,N_15355);
or U15904 (N_15904,N_15056,N_15250);
and U15905 (N_15905,N_15395,N_15175);
nor U15906 (N_15906,N_15021,N_15129);
nand U15907 (N_15907,N_15195,N_15442);
nand U15908 (N_15908,N_15205,N_15011);
and U15909 (N_15909,N_15242,N_15292);
and U15910 (N_15910,N_15298,N_15062);
nand U15911 (N_15911,N_15238,N_15214);
and U15912 (N_15912,N_15185,N_15142);
and U15913 (N_15913,N_15233,N_15153);
xor U15914 (N_15914,N_15346,N_15091);
nor U15915 (N_15915,N_15004,N_15167);
and U15916 (N_15916,N_15423,N_15044);
nand U15917 (N_15917,N_15105,N_15219);
or U15918 (N_15918,N_15277,N_15453);
xnor U15919 (N_15919,N_15331,N_15054);
nand U15920 (N_15920,N_15475,N_15025);
xor U15921 (N_15921,N_15134,N_15315);
nor U15922 (N_15922,N_15070,N_15018);
and U15923 (N_15923,N_15480,N_15471);
nor U15924 (N_15924,N_15055,N_15023);
xnor U15925 (N_15925,N_15003,N_15434);
or U15926 (N_15926,N_15020,N_15336);
nand U15927 (N_15927,N_15321,N_15187);
xnor U15928 (N_15928,N_15450,N_15313);
and U15929 (N_15929,N_15443,N_15291);
nor U15930 (N_15930,N_15232,N_15329);
xor U15931 (N_15931,N_15422,N_15498);
or U15932 (N_15932,N_15120,N_15017);
nor U15933 (N_15933,N_15447,N_15404);
or U15934 (N_15934,N_15105,N_15277);
xnor U15935 (N_15935,N_15383,N_15299);
xor U15936 (N_15936,N_15348,N_15107);
or U15937 (N_15937,N_15160,N_15439);
nor U15938 (N_15938,N_15391,N_15488);
nor U15939 (N_15939,N_15011,N_15216);
xor U15940 (N_15940,N_15490,N_15184);
or U15941 (N_15941,N_15356,N_15336);
nor U15942 (N_15942,N_15316,N_15036);
nor U15943 (N_15943,N_15268,N_15166);
or U15944 (N_15944,N_15157,N_15384);
or U15945 (N_15945,N_15150,N_15246);
or U15946 (N_15946,N_15099,N_15082);
xnor U15947 (N_15947,N_15431,N_15054);
xnor U15948 (N_15948,N_15232,N_15030);
or U15949 (N_15949,N_15386,N_15353);
and U15950 (N_15950,N_15056,N_15328);
xnor U15951 (N_15951,N_15376,N_15227);
nor U15952 (N_15952,N_15328,N_15263);
xor U15953 (N_15953,N_15056,N_15492);
or U15954 (N_15954,N_15420,N_15211);
nand U15955 (N_15955,N_15011,N_15308);
nand U15956 (N_15956,N_15293,N_15163);
nand U15957 (N_15957,N_15185,N_15050);
nand U15958 (N_15958,N_15281,N_15003);
nor U15959 (N_15959,N_15137,N_15439);
nor U15960 (N_15960,N_15155,N_15350);
nand U15961 (N_15961,N_15136,N_15174);
nand U15962 (N_15962,N_15393,N_15257);
or U15963 (N_15963,N_15059,N_15317);
xor U15964 (N_15964,N_15006,N_15020);
and U15965 (N_15965,N_15097,N_15140);
and U15966 (N_15966,N_15013,N_15156);
nor U15967 (N_15967,N_15407,N_15165);
xnor U15968 (N_15968,N_15410,N_15288);
or U15969 (N_15969,N_15162,N_15070);
xnor U15970 (N_15970,N_15262,N_15372);
xnor U15971 (N_15971,N_15234,N_15432);
xnor U15972 (N_15972,N_15073,N_15196);
and U15973 (N_15973,N_15317,N_15005);
xnor U15974 (N_15974,N_15362,N_15320);
and U15975 (N_15975,N_15300,N_15351);
xnor U15976 (N_15976,N_15140,N_15127);
xor U15977 (N_15977,N_15355,N_15293);
nor U15978 (N_15978,N_15103,N_15490);
nand U15979 (N_15979,N_15113,N_15099);
nor U15980 (N_15980,N_15390,N_15202);
or U15981 (N_15981,N_15032,N_15446);
nand U15982 (N_15982,N_15296,N_15097);
xnor U15983 (N_15983,N_15008,N_15156);
nand U15984 (N_15984,N_15395,N_15345);
nor U15985 (N_15985,N_15332,N_15446);
or U15986 (N_15986,N_15135,N_15262);
xor U15987 (N_15987,N_15361,N_15371);
and U15988 (N_15988,N_15228,N_15469);
nor U15989 (N_15989,N_15421,N_15208);
or U15990 (N_15990,N_15271,N_15017);
nor U15991 (N_15991,N_15477,N_15292);
and U15992 (N_15992,N_15237,N_15276);
nor U15993 (N_15993,N_15484,N_15329);
nor U15994 (N_15994,N_15346,N_15119);
nor U15995 (N_15995,N_15183,N_15390);
xnor U15996 (N_15996,N_15474,N_15091);
and U15997 (N_15997,N_15174,N_15231);
and U15998 (N_15998,N_15182,N_15222);
nand U15999 (N_15999,N_15491,N_15174);
or U16000 (N_16000,N_15502,N_15968);
and U16001 (N_16001,N_15879,N_15826);
xnor U16002 (N_16002,N_15679,N_15907);
or U16003 (N_16003,N_15756,N_15747);
nand U16004 (N_16004,N_15840,N_15998);
nand U16005 (N_16005,N_15515,N_15769);
nand U16006 (N_16006,N_15867,N_15650);
or U16007 (N_16007,N_15711,N_15587);
and U16008 (N_16008,N_15675,N_15648);
and U16009 (N_16009,N_15746,N_15910);
nand U16010 (N_16010,N_15553,N_15970);
or U16011 (N_16011,N_15504,N_15703);
and U16012 (N_16012,N_15795,N_15512);
nor U16013 (N_16013,N_15584,N_15570);
xnor U16014 (N_16014,N_15734,N_15542);
or U16015 (N_16015,N_15993,N_15865);
xor U16016 (N_16016,N_15611,N_15996);
xnor U16017 (N_16017,N_15992,N_15561);
nor U16018 (N_16018,N_15702,N_15706);
nand U16019 (N_16019,N_15904,N_15645);
or U16020 (N_16020,N_15720,N_15919);
xnor U16021 (N_16021,N_15820,N_15972);
nor U16022 (N_16022,N_15667,N_15573);
nand U16023 (N_16023,N_15540,N_15912);
xor U16024 (N_16024,N_15770,N_15827);
and U16025 (N_16025,N_15959,N_15562);
nor U16026 (N_16026,N_15606,N_15958);
or U16027 (N_16027,N_15618,N_15614);
and U16028 (N_16028,N_15822,N_15724);
xnor U16029 (N_16029,N_15949,N_15790);
nand U16030 (N_16030,N_15523,N_15609);
or U16031 (N_16031,N_15565,N_15982);
nor U16032 (N_16032,N_15773,N_15913);
or U16033 (N_16033,N_15691,N_15537);
and U16034 (N_16034,N_15843,N_15709);
or U16035 (N_16035,N_15610,N_15903);
nor U16036 (N_16036,N_15593,N_15923);
nand U16037 (N_16037,N_15829,N_15776);
nor U16038 (N_16038,N_15988,N_15683);
or U16039 (N_16039,N_15571,N_15841);
nand U16040 (N_16040,N_15625,N_15851);
nor U16041 (N_16041,N_15941,N_15616);
nand U16042 (N_16042,N_15933,N_15596);
nand U16043 (N_16043,N_15588,N_15883);
nand U16044 (N_16044,N_15874,N_15716);
nand U16045 (N_16045,N_15527,N_15931);
or U16046 (N_16046,N_15856,N_15940);
and U16047 (N_16047,N_15877,N_15926);
or U16048 (N_16048,N_15695,N_15999);
nor U16049 (N_16049,N_15801,N_15550);
nor U16050 (N_16050,N_15644,N_15951);
nor U16051 (N_16051,N_15758,N_15661);
and U16052 (N_16052,N_15814,N_15783);
nor U16053 (N_16053,N_15973,N_15861);
or U16054 (N_16054,N_15705,N_15898);
xor U16055 (N_16055,N_15511,N_15902);
nor U16056 (N_16056,N_15965,N_15722);
nor U16057 (N_16057,N_15529,N_15536);
nand U16058 (N_16058,N_15738,N_15510);
xnor U16059 (N_16059,N_15894,N_15971);
nand U16060 (N_16060,N_15849,N_15725);
or U16061 (N_16061,N_15655,N_15567);
and U16062 (N_16062,N_15714,N_15892);
or U16063 (N_16063,N_15659,N_15761);
and U16064 (N_16064,N_15696,N_15805);
and U16065 (N_16065,N_15948,N_15925);
nand U16066 (N_16066,N_15522,N_15885);
or U16067 (N_16067,N_15600,N_15654);
nand U16068 (N_16068,N_15873,N_15799);
and U16069 (N_16069,N_15669,N_15953);
and U16070 (N_16070,N_15707,N_15938);
and U16071 (N_16071,N_15581,N_15665);
nand U16072 (N_16072,N_15742,N_15750);
and U16073 (N_16073,N_15560,N_15890);
or U16074 (N_16074,N_15721,N_15607);
nand U16075 (N_16075,N_15821,N_15528);
xor U16076 (N_16076,N_15979,N_15930);
or U16077 (N_16077,N_15863,N_15545);
nor U16078 (N_16078,N_15848,N_15842);
nor U16079 (N_16079,N_15525,N_15524);
xor U16080 (N_16080,N_15918,N_15859);
nor U16081 (N_16081,N_15623,N_15835);
nand U16082 (N_16082,N_15757,N_15880);
nor U16083 (N_16083,N_15539,N_15875);
nand U16084 (N_16084,N_15778,N_15768);
xnor U16085 (N_16085,N_15915,N_15909);
xnor U16086 (N_16086,N_15546,N_15765);
nor U16087 (N_16087,N_15637,N_15806);
nor U16088 (N_16088,N_15690,N_15628);
nor U16089 (N_16089,N_15647,N_15895);
or U16090 (N_16090,N_15983,N_15990);
xor U16091 (N_16091,N_15664,N_15824);
nand U16092 (N_16092,N_15929,N_15960);
nor U16093 (N_16093,N_15558,N_15576);
and U16094 (N_16094,N_15854,N_15678);
nand U16095 (N_16095,N_15878,N_15900);
nand U16096 (N_16096,N_15782,N_15615);
nand U16097 (N_16097,N_15891,N_15514);
nand U16098 (N_16098,N_15955,N_15518);
xnor U16099 (N_16099,N_15549,N_15597);
or U16100 (N_16100,N_15500,N_15694);
or U16101 (N_16101,N_15828,N_15501);
or U16102 (N_16102,N_15946,N_15741);
nor U16103 (N_16103,N_15533,N_15530);
and U16104 (N_16104,N_15568,N_15869);
nor U16105 (N_16105,N_15939,N_15882);
nor U16106 (N_16106,N_15643,N_15509);
and U16107 (N_16107,N_15737,N_15519);
xor U16108 (N_16108,N_15825,N_15864);
or U16109 (N_16109,N_15505,N_15781);
xnor U16110 (N_16110,N_15980,N_15839);
nand U16111 (N_16111,N_15927,N_15978);
or U16112 (N_16112,N_15922,N_15710);
and U16113 (N_16113,N_15956,N_15796);
nand U16114 (N_16114,N_15764,N_15870);
nand U16115 (N_16115,N_15771,N_15589);
nand U16116 (N_16116,N_15914,N_15893);
and U16117 (N_16117,N_15717,N_15866);
nand U16118 (N_16118,N_15962,N_15630);
and U16119 (N_16119,N_15816,N_15671);
nand U16120 (N_16120,N_15548,N_15754);
and U16121 (N_16121,N_15831,N_15957);
xor U16122 (N_16122,N_15640,N_15753);
or U16123 (N_16123,N_15833,N_15744);
nand U16124 (N_16124,N_15670,N_15845);
nor U16125 (N_16125,N_15622,N_15785);
and U16126 (N_16126,N_15850,N_15520);
nand U16127 (N_16127,N_15794,N_15743);
nor U16128 (N_16128,N_15563,N_15846);
or U16129 (N_16129,N_15674,N_15937);
nand U16130 (N_16130,N_15619,N_15692);
and U16131 (N_16131,N_15728,N_15547);
nor U16132 (N_16132,N_15852,N_15974);
and U16133 (N_16133,N_15911,N_15963);
nand U16134 (N_16134,N_15862,N_15652);
nand U16135 (N_16135,N_15975,N_15704);
xor U16136 (N_16136,N_15767,N_15759);
or U16137 (N_16137,N_15837,N_15700);
nor U16138 (N_16138,N_15748,N_15662);
nand U16139 (N_16139,N_15897,N_15855);
nand U16140 (N_16140,N_15689,N_15534);
and U16141 (N_16141,N_15802,N_15920);
or U16142 (N_16142,N_15556,N_15792);
nor U16143 (N_16143,N_15803,N_15888);
or U16144 (N_16144,N_15595,N_15574);
nor U16145 (N_16145,N_15755,N_15507);
xor U16146 (N_16146,N_15649,N_15967);
nand U16147 (N_16147,N_15774,N_15751);
or U16148 (N_16148,N_15809,N_15886);
or U16149 (N_16149,N_15513,N_15638);
or U16150 (N_16150,N_15994,N_15964);
or U16151 (N_16151,N_15777,N_15532);
nand U16152 (N_16152,N_15740,N_15881);
nor U16153 (N_16153,N_15995,N_15921);
xnor U16154 (N_16154,N_15876,N_15715);
xor U16155 (N_16155,N_15699,N_15541);
nor U16156 (N_16156,N_15604,N_15559);
nand U16157 (N_16157,N_15682,N_15749);
nand U16158 (N_16158,N_15543,N_15779);
xor U16159 (N_16159,N_15697,N_15853);
nor U16160 (N_16160,N_15732,N_15932);
nor U16161 (N_16161,N_15884,N_15653);
nand U16162 (N_16162,N_15812,N_15591);
and U16163 (N_16163,N_15733,N_15836);
or U16164 (N_16164,N_15585,N_15943);
or U16165 (N_16165,N_15631,N_15680);
xor U16166 (N_16166,N_15646,N_15656);
xor U16167 (N_16167,N_15658,N_15668);
or U16168 (N_16168,N_15813,N_15552);
nor U16169 (N_16169,N_15731,N_15544);
nand U16170 (N_16170,N_15791,N_15693);
nor U16171 (N_16171,N_15657,N_15997);
nor U16172 (N_16172,N_15569,N_15735);
and U16173 (N_16173,N_15760,N_15739);
nor U16174 (N_16174,N_15521,N_15917);
and U16175 (N_16175,N_15780,N_15896);
or U16176 (N_16176,N_15688,N_15599);
nor U16177 (N_16177,N_15935,N_15555);
or U16178 (N_16178,N_15551,N_15804);
and U16179 (N_16179,N_15617,N_15723);
nor U16180 (N_16180,N_15684,N_15517);
and U16181 (N_16181,N_15977,N_15626);
and U16182 (N_16182,N_15719,N_15908);
nand U16183 (N_16183,N_15676,N_15621);
nand U16184 (N_16184,N_15947,N_15984);
and U16185 (N_16185,N_15916,N_15590);
nand U16186 (N_16186,N_15905,N_15726);
xor U16187 (N_16187,N_15830,N_15819);
xnor U16188 (N_16188,N_15583,N_15698);
and U16189 (N_16189,N_15557,N_15800);
or U16190 (N_16190,N_15944,N_15627);
and U16191 (N_16191,N_15901,N_15887);
nand U16192 (N_16192,N_15868,N_15966);
nand U16193 (N_16193,N_15936,N_15538);
nand U16194 (N_16194,N_15899,N_15834);
xor U16195 (N_16195,N_15580,N_15817);
nor U16196 (N_16196,N_15808,N_15950);
nand U16197 (N_16197,N_15666,N_15579);
xor U16198 (N_16198,N_15981,N_15844);
nor U16199 (N_16199,N_15789,N_15681);
and U16200 (N_16200,N_15620,N_15807);
xnor U16201 (N_16201,N_15928,N_15531);
or U16202 (N_16202,N_15811,N_15976);
nor U16203 (N_16203,N_15858,N_15554);
xor U16204 (N_16204,N_15612,N_15663);
nand U16205 (N_16205,N_15763,N_15687);
nor U16206 (N_16206,N_15608,N_15634);
and U16207 (N_16207,N_15857,N_15651);
xor U16208 (N_16208,N_15686,N_15677);
xor U16209 (N_16209,N_15730,N_15642);
xnor U16210 (N_16210,N_15586,N_15577);
or U16211 (N_16211,N_15823,N_15578);
or U16212 (N_16212,N_15798,N_15632);
xor U16213 (N_16213,N_15815,N_15772);
or U16214 (N_16214,N_15685,N_15788);
and U16215 (N_16215,N_15673,N_15952);
nand U16216 (N_16216,N_15572,N_15605);
and U16217 (N_16217,N_15736,N_15745);
xor U16218 (N_16218,N_15989,N_15818);
xnor U16219 (N_16219,N_15832,N_15969);
xnor U16220 (N_16220,N_15526,N_15797);
or U16221 (N_16221,N_15872,N_15793);
nand U16222 (N_16222,N_15986,N_15592);
or U16223 (N_16223,N_15713,N_15871);
and U16224 (N_16224,N_15613,N_15889);
and U16225 (N_16225,N_15508,N_15639);
xnor U16226 (N_16226,N_15775,N_15945);
nand U16227 (N_16227,N_15660,N_15906);
xor U16228 (N_16228,N_15598,N_15810);
and U16229 (N_16229,N_15624,N_15942);
and U16230 (N_16230,N_15838,N_15603);
and U16231 (N_16231,N_15708,N_15641);
and U16232 (N_16232,N_15786,N_15934);
or U16233 (N_16233,N_15727,N_15712);
and U16234 (N_16234,N_15784,N_15762);
and U16235 (N_16235,N_15535,N_15961);
or U16236 (N_16236,N_15575,N_15729);
or U16237 (N_16237,N_15503,N_15718);
xor U16238 (N_16238,N_15701,N_15954);
and U16239 (N_16239,N_15860,N_15602);
xor U16240 (N_16240,N_15506,N_15601);
nor U16241 (N_16241,N_15629,N_15636);
nand U16242 (N_16242,N_15985,N_15516);
or U16243 (N_16243,N_15594,N_15991);
or U16244 (N_16244,N_15787,N_15672);
or U16245 (N_16245,N_15635,N_15847);
or U16246 (N_16246,N_15566,N_15564);
nor U16247 (N_16247,N_15582,N_15633);
nor U16248 (N_16248,N_15924,N_15752);
xnor U16249 (N_16249,N_15766,N_15987);
nand U16250 (N_16250,N_15885,N_15653);
or U16251 (N_16251,N_15970,N_15532);
xnor U16252 (N_16252,N_15761,N_15631);
nor U16253 (N_16253,N_15946,N_15931);
and U16254 (N_16254,N_15539,N_15966);
and U16255 (N_16255,N_15515,N_15862);
nand U16256 (N_16256,N_15514,N_15691);
nor U16257 (N_16257,N_15924,N_15543);
nor U16258 (N_16258,N_15555,N_15541);
nor U16259 (N_16259,N_15596,N_15763);
and U16260 (N_16260,N_15770,N_15911);
nor U16261 (N_16261,N_15803,N_15557);
and U16262 (N_16262,N_15766,N_15857);
nand U16263 (N_16263,N_15705,N_15697);
nor U16264 (N_16264,N_15762,N_15816);
and U16265 (N_16265,N_15858,N_15956);
or U16266 (N_16266,N_15964,N_15883);
or U16267 (N_16267,N_15558,N_15552);
xnor U16268 (N_16268,N_15859,N_15619);
xor U16269 (N_16269,N_15702,N_15933);
nand U16270 (N_16270,N_15747,N_15789);
and U16271 (N_16271,N_15653,N_15749);
or U16272 (N_16272,N_15615,N_15506);
xor U16273 (N_16273,N_15721,N_15549);
xor U16274 (N_16274,N_15785,N_15722);
nand U16275 (N_16275,N_15647,N_15870);
xnor U16276 (N_16276,N_15867,N_15597);
xor U16277 (N_16277,N_15843,N_15978);
and U16278 (N_16278,N_15894,N_15983);
and U16279 (N_16279,N_15869,N_15624);
and U16280 (N_16280,N_15592,N_15642);
or U16281 (N_16281,N_15895,N_15505);
nor U16282 (N_16282,N_15598,N_15672);
or U16283 (N_16283,N_15631,N_15774);
nor U16284 (N_16284,N_15724,N_15782);
or U16285 (N_16285,N_15563,N_15747);
nand U16286 (N_16286,N_15843,N_15866);
or U16287 (N_16287,N_15811,N_15925);
nor U16288 (N_16288,N_15760,N_15573);
and U16289 (N_16289,N_15697,N_15606);
xor U16290 (N_16290,N_15671,N_15921);
xnor U16291 (N_16291,N_15700,N_15876);
nand U16292 (N_16292,N_15670,N_15749);
xor U16293 (N_16293,N_15776,N_15779);
or U16294 (N_16294,N_15834,N_15626);
or U16295 (N_16295,N_15840,N_15669);
nand U16296 (N_16296,N_15720,N_15864);
xor U16297 (N_16297,N_15763,N_15830);
or U16298 (N_16298,N_15546,N_15735);
and U16299 (N_16299,N_15838,N_15745);
and U16300 (N_16300,N_15774,N_15544);
nor U16301 (N_16301,N_15584,N_15503);
nor U16302 (N_16302,N_15568,N_15622);
nand U16303 (N_16303,N_15779,N_15919);
xnor U16304 (N_16304,N_15904,N_15660);
nor U16305 (N_16305,N_15652,N_15960);
nand U16306 (N_16306,N_15715,N_15905);
xnor U16307 (N_16307,N_15708,N_15638);
nor U16308 (N_16308,N_15987,N_15563);
and U16309 (N_16309,N_15654,N_15987);
xor U16310 (N_16310,N_15749,N_15641);
or U16311 (N_16311,N_15508,N_15922);
xor U16312 (N_16312,N_15978,N_15646);
or U16313 (N_16313,N_15668,N_15751);
nand U16314 (N_16314,N_15634,N_15580);
xor U16315 (N_16315,N_15871,N_15533);
and U16316 (N_16316,N_15755,N_15870);
xnor U16317 (N_16317,N_15814,N_15660);
nand U16318 (N_16318,N_15582,N_15955);
or U16319 (N_16319,N_15601,N_15594);
nor U16320 (N_16320,N_15958,N_15836);
nor U16321 (N_16321,N_15795,N_15766);
and U16322 (N_16322,N_15765,N_15682);
and U16323 (N_16323,N_15594,N_15635);
xor U16324 (N_16324,N_15629,N_15714);
xnor U16325 (N_16325,N_15503,N_15873);
and U16326 (N_16326,N_15577,N_15842);
or U16327 (N_16327,N_15992,N_15664);
xnor U16328 (N_16328,N_15741,N_15824);
xor U16329 (N_16329,N_15980,N_15985);
xor U16330 (N_16330,N_15932,N_15753);
nand U16331 (N_16331,N_15562,N_15685);
nor U16332 (N_16332,N_15683,N_15635);
and U16333 (N_16333,N_15626,N_15702);
nor U16334 (N_16334,N_15693,N_15643);
and U16335 (N_16335,N_15763,N_15633);
xnor U16336 (N_16336,N_15654,N_15876);
and U16337 (N_16337,N_15545,N_15813);
nand U16338 (N_16338,N_15627,N_15821);
nor U16339 (N_16339,N_15997,N_15944);
or U16340 (N_16340,N_15652,N_15518);
nor U16341 (N_16341,N_15696,N_15841);
nor U16342 (N_16342,N_15646,N_15574);
nand U16343 (N_16343,N_15973,N_15953);
or U16344 (N_16344,N_15546,N_15956);
or U16345 (N_16345,N_15630,N_15509);
or U16346 (N_16346,N_15612,N_15644);
xor U16347 (N_16347,N_15898,N_15673);
or U16348 (N_16348,N_15683,N_15856);
xor U16349 (N_16349,N_15620,N_15756);
and U16350 (N_16350,N_15985,N_15768);
xor U16351 (N_16351,N_15785,N_15899);
nand U16352 (N_16352,N_15510,N_15777);
or U16353 (N_16353,N_15979,N_15921);
nand U16354 (N_16354,N_15895,N_15739);
xnor U16355 (N_16355,N_15650,N_15972);
and U16356 (N_16356,N_15877,N_15698);
and U16357 (N_16357,N_15705,N_15919);
and U16358 (N_16358,N_15558,N_15954);
and U16359 (N_16359,N_15969,N_15866);
xnor U16360 (N_16360,N_15556,N_15610);
xor U16361 (N_16361,N_15502,N_15918);
xor U16362 (N_16362,N_15750,N_15891);
nor U16363 (N_16363,N_15709,N_15686);
xor U16364 (N_16364,N_15683,N_15633);
nor U16365 (N_16365,N_15812,N_15959);
nor U16366 (N_16366,N_15831,N_15891);
xor U16367 (N_16367,N_15793,N_15685);
nand U16368 (N_16368,N_15948,N_15583);
nor U16369 (N_16369,N_15921,N_15545);
xor U16370 (N_16370,N_15967,N_15736);
xnor U16371 (N_16371,N_15848,N_15626);
xnor U16372 (N_16372,N_15768,N_15611);
or U16373 (N_16373,N_15688,N_15837);
nor U16374 (N_16374,N_15541,N_15520);
xor U16375 (N_16375,N_15830,N_15991);
nand U16376 (N_16376,N_15611,N_15573);
xnor U16377 (N_16377,N_15815,N_15867);
or U16378 (N_16378,N_15912,N_15545);
nor U16379 (N_16379,N_15902,N_15507);
nand U16380 (N_16380,N_15915,N_15535);
nand U16381 (N_16381,N_15817,N_15508);
or U16382 (N_16382,N_15911,N_15738);
nor U16383 (N_16383,N_15673,N_15909);
nand U16384 (N_16384,N_15889,N_15600);
or U16385 (N_16385,N_15562,N_15775);
and U16386 (N_16386,N_15843,N_15742);
nand U16387 (N_16387,N_15631,N_15836);
and U16388 (N_16388,N_15776,N_15798);
nor U16389 (N_16389,N_15658,N_15586);
and U16390 (N_16390,N_15672,N_15724);
nand U16391 (N_16391,N_15611,N_15960);
or U16392 (N_16392,N_15590,N_15799);
or U16393 (N_16393,N_15800,N_15661);
and U16394 (N_16394,N_15904,N_15651);
or U16395 (N_16395,N_15634,N_15985);
nand U16396 (N_16396,N_15839,N_15551);
nand U16397 (N_16397,N_15591,N_15880);
nor U16398 (N_16398,N_15585,N_15637);
nand U16399 (N_16399,N_15772,N_15508);
or U16400 (N_16400,N_15608,N_15785);
and U16401 (N_16401,N_15966,N_15928);
or U16402 (N_16402,N_15691,N_15884);
nor U16403 (N_16403,N_15639,N_15925);
and U16404 (N_16404,N_15816,N_15927);
nand U16405 (N_16405,N_15793,N_15570);
and U16406 (N_16406,N_15644,N_15786);
or U16407 (N_16407,N_15536,N_15859);
xnor U16408 (N_16408,N_15553,N_15599);
nor U16409 (N_16409,N_15895,N_15707);
xnor U16410 (N_16410,N_15988,N_15853);
xnor U16411 (N_16411,N_15857,N_15800);
and U16412 (N_16412,N_15883,N_15774);
or U16413 (N_16413,N_15945,N_15919);
nor U16414 (N_16414,N_15603,N_15817);
nor U16415 (N_16415,N_15794,N_15502);
and U16416 (N_16416,N_15501,N_15619);
nand U16417 (N_16417,N_15574,N_15506);
and U16418 (N_16418,N_15929,N_15958);
xnor U16419 (N_16419,N_15924,N_15844);
xnor U16420 (N_16420,N_15758,N_15764);
nand U16421 (N_16421,N_15521,N_15993);
and U16422 (N_16422,N_15671,N_15786);
nand U16423 (N_16423,N_15590,N_15971);
nor U16424 (N_16424,N_15518,N_15849);
xor U16425 (N_16425,N_15564,N_15506);
xnor U16426 (N_16426,N_15681,N_15868);
nand U16427 (N_16427,N_15962,N_15586);
nand U16428 (N_16428,N_15521,N_15999);
xor U16429 (N_16429,N_15531,N_15896);
nor U16430 (N_16430,N_15523,N_15692);
nand U16431 (N_16431,N_15976,N_15721);
and U16432 (N_16432,N_15932,N_15678);
and U16433 (N_16433,N_15512,N_15917);
nand U16434 (N_16434,N_15655,N_15879);
nor U16435 (N_16435,N_15565,N_15735);
nor U16436 (N_16436,N_15932,N_15685);
and U16437 (N_16437,N_15755,N_15915);
nor U16438 (N_16438,N_15780,N_15907);
nor U16439 (N_16439,N_15913,N_15882);
or U16440 (N_16440,N_15901,N_15601);
nor U16441 (N_16441,N_15857,N_15736);
nor U16442 (N_16442,N_15646,N_15897);
nand U16443 (N_16443,N_15784,N_15505);
and U16444 (N_16444,N_15668,N_15923);
xnor U16445 (N_16445,N_15624,N_15824);
nand U16446 (N_16446,N_15629,N_15892);
and U16447 (N_16447,N_15528,N_15889);
or U16448 (N_16448,N_15864,N_15608);
nand U16449 (N_16449,N_15690,N_15837);
nor U16450 (N_16450,N_15763,N_15866);
or U16451 (N_16451,N_15553,N_15974);
nand U16452 (N_16452,N_15782,N_15779);
xor U16453 (N_16453,N_15904,N_15662);
xnor U16454 (N_16454,N_15708,N_15524);
nor U16455 (N_16455,N_15955,N_15794);
nand U16456 (N_16456,N_15869,N_15857);
and U16457 (N_16457,N_15978,N_15508);
or U16458 (N_16458,N_15509,N_15594);
and U16459 (N_16459,N_15512,N_15854);
nand U16460 (N_16460,N_15508,N_15841);
and U16461 (N_16461,N_15585,N_15650);
and U16462 (N_16462,N_15770,N_15978);
nand U16463 (N_16463,N_15783,N_15749);
and U16464 (N_16464,N_15744,N_15737);
or U16465 (N_16465,N_15677,N_15966);
nor U16466 (N_16466,N_15799,N_15727);
nand U16467 (N_16467,N_15643,N_15792);
nand U16468 (N_16468,N_15721,N_15813);
nor U16469 (N_16469,N_15553,N_15570);
or U16470 (N_16470,N_15812,N_15687);
or U16471 (N_16471,N_15518,N_15555);
nor U16472 (N_16472,N_15813,N_15635);
or U16473 (N_16473,N_15930,N_15536);
nor U16474 (N_16474,N_15775,N_15538);
xor U16475 (N_16475,N_15704,N_15868);
xor U16476 (N_16476,N_15760,N_15552);
xnor U16477 (N_16477,N_15940,N_15632);
nor U16478 (N_16478,N_15570,N_15855);
and U16479 (N_16479,N_15573,N_15855);
or U16480 (N_16480,N_15501,N_15840);
nor U16481 (N_16481,N_15801,N_15807);
xor U16482 (N_16482,N_15742,N_15726);
nand U16483 (N_16483,N_15843,N_15829);
and U16484 (N_16484,N_15929,N_15846);
or U16485 (N_16485,N_15962,N_15923);
nand U16486 (N_16486,N_15679,N_15544);
and U16487 (N_16487,N_15757,N_15688);
xor U16488 (N_16488,N_15697,N_15592);
nand U16489 (N_16489,N_15802,N_15925);
nor U16490 (N_16490,N_15861,N_15769);
xor U16491 (N_16491,N_15940,N_15953);
nand U16492 (N_16492,N_15777,N_15840);
nor U16493 (N_16493,N_15839,N_15815);
or U16494 (N_16494,N_15728,N_15595);
xnor U16495 (N_16495,N_15632,N_15846);
nand U16496 (N_16496,N_15958,N_15685);
nor U16497 (N_16497,N_15941,N_15822);
nor U16498 (N_16498,N_15594,N_15840);
xnor U16499 (N_16499,N_15836,N_15788);
nor U16500 (N_16500,N_16264,N_16321);
nand U16501 (N_16501,N_16282,N_16211);
nand U16502 (N_16502,N_16440,N_16146);
nand U16503 (N_16503,N_16431,N_16187);
nand U16504 (N_16504,N_16009,N_16061);
or U16505 (N_16505,N_16023,N_16201);
nand U16506 (N_16506,N_16136,N_16276);
and U16507 (N_16507,N_16481,N_16249);
and U16508 (N_16508,N_16286,N_16089);
nand U16509 (N_16509,N_16169,N_16407);
xor U16510 (N_16510,N_16058,N_16491);
and U16511 (N_16511,N_16190,N_16356);
nand U16512 (N_16512,N_16304,N_16138);
nor U16513 (N_16513,N_16322,N_16067);
or U16514 (N_16514,N_16480,N_16175);
nor U16515 (N_16515,N_16127,N_16162);
nor U16516 (N_16516,N_16002,N_16066);
or U16517 (N_16517,N_16100,N_16053);
and U16518 (N_16518,N_16297,N_16438);
nor U16519 (N_16519,N_16306,N_16004);
or U16520 (N_16520,N_16395,N_16316);
xor U16521 (N_16521,N_16313,N_16192);
xnor U16522 (N_16522,N_16318,N_16019);
nand U16523 (N_16523,N_16013,N_16011);
nand U16524 (N_16524,N_16236,N_16258);
nand U16525 (N_16525,N_16433,N_16291);
nand U16526 (N_16526,N_16307,N_16254);
or U16527 (N_16527,N_16308,N_16470);
or U16528 (N_16528,N_16271,N_16101);
and U16529 (N_16529,N_16107,N_16241);
nand U16530 (N_16530,N_16404,N_16498);
xor U16531 (N_16531,N_16422,N_16419);
nand U16532 (N_16532,N_16208,N_16221);
nor U16533 (N_16533,N_16060,N_16281);
nand U16534 (N_16534,N_16256,N_16283);
and U16535 (N_16535,N_16430,N_16094);
and U16536 (N_16536,N_16025,N_16046);
or U16537 (N_16537,N_16115,N_16080);
xnor U16538 (N_16538,N_16263,N_16425);
and U16539 (N_16539,N_16257,N_16156);
xor U16540 (N_16540,N_16397,N_16451);
nor U16541 (N_16541,N_16062,N_16212);
or U16542 (N_16542,N_16015,N_16197);
and U16543 (N_16543,N_16075,N_16409);
or U16544 (N_16544,N_16096,N_16170);
and U16545 (N_16545,N_16145,N_16469);
and U16546 (N_16546,N_16355,N_16396);
and U16547 (N_16547,N_16006,N_16091);
nor U16548 (N_16548,N_16045,N_16383);
or U16549 (N_16549,N_16434,N_16064);
xnor U16550 (N_16550,N_16132,N_16171);
nor U16551 (N_16551,N_16366,N_16044);
nand U16552 (N_16552,N_16479,N_16387);
xor U16553 (N_16553,N_16389,N_16376);
and U16554 (N_16554,N_16377,N_16134);
or U16555 (N_16555,N_16348,N_16268);
xnor U16556 (N_16556,N_16110,N_16184);
nor U16557 (N_16557,N_16166,N_16074);
or U16558 (N_16558,N_16453,N_16230);
nand U16559 (N_16559,N_16022,N_16029);
nand U16560 (N_16560,N_16168,N_16000);
and U16561 (N_16561,N_16144,N_16153);
xor U16562 (N_16562,N_16375,N_16259);
nor U16563 (N_16563,N_16421,N_16070);
or U16564 (N_16564,N_16027,N_16465);
or U16565 (N_16565,N_16418,N_16370);
nand U16566 (N_16566,N_16051,N_16243);
nor U16567 (N_16567,N_16069,N_16391);
nor U16568 (N_16568,N_16054,N_16467);
and U16569 (N_16569,N_16328,N_16447);
xor U16570 (N_16570,N_16113,N_16333);
xnor U16571 (N_16571,N_16084,N_16079);
nand U16572 (N_16572,N_16476,N_16103);
or U16573 (N_16573,N_16309,N_16394);
xnor U16574 (N_16574,N_16408,N_16129);
nand U16575 (N_16575,N_16194,N_16008);
and U16576 (N_16576,N_16233,N_16179);
nand U16577 (N_16577,N_16336,N_16018);
xor U16578 (N_16578,N_16373,N_16047);
nand U16579 (N_16579,N_16454,N_16260);
nand U16580 (N_16580,N_16350,N_16059);
xnor U16581 (N_16581,N_16287,N_16120);
nor U16582 (N_16582,N_16381,N_16317);
nor U16583 (N_16583,N_16458,N_16003);
nand U16584 (N_16584,N_16403,N_16483);
nor U16585 (N_16585,N_16083,N_16463);
xor U16586 (N_16586,N_16439,N_16424);
nand U16587 (N_16587,N_16489,N_16126);
or U16588 (N_16588,N_16442,N_16130);
or U16589 (N_16589,N_16477,N_16152);
nor U16590 (N_16590,N_16493,N_16455);
and U16591 (N_16591,N_16246,N_16315);
and U16592 (N_16592,N_16423,N_16154);
and U16593 (N_16593,N_16217,N_16332);
and U16594 (N_16594,N_16147,N_16114);
nor U16595 (N_16595,N_16160,N_16310);
xor U16596 (N_16596,N_16071,N_16385);
nand U16597 (N_16597,N_16035,N_16123);
and U16598 (N_16598,N_16106,N_16104);
xor U16599 (N_16599,N_16231,N_16343);
nand U16600 (N_16600,N_16405,N_16415);
nor U16601 (N_16601,N_16349,N_16224);
xnor U16602 (N_16602,N_16068,N_16228);
xnor U16603 (N_16603,N_16295,N_16048);
and U16604 (N_16604,N_16119,N_16368);
nor U16605 (N_16605,N_16226,N_16326);
nand U16606 (N_16606,N_16420,N_16176);
nor U16607 (N_16607,N_16195,N_16347);
or U16608 (N_16608,N_16116,N_16300);
and U16609 (N_16609,N_16040,N_16063);
nor U16610 (N_16610,N_16320,N_16112);
or U16611 (N_16611,N_16081,N_16225);
nand U16612 (N_16612,N_16010,N_16327);
nand U16613 (N_16613,N_16234,N_16237);
nor U16614 (N_16614,N_16255,N_16329);
and U16615 (N_16615,N_16494,N_16473);
or U16616 (N_16616,N_16398,N_16095);
nand U16617 (N_16617,N_16238,N_16242);
xor U16618 (N_16618,N_16272,N_16191);
and U16619 (N_16619,N_16173,N_16001);
nor U16620 (N_16620,N_16369,N_16325);
nand U16621 (N_16621,N_16247,N_16189);
and U16622 (N_16622,N_16352,N_16390);
and U16623 (N_16623,N_16038,N_16078);
or U16624 (N_16624,N_16105,N_16335);
or U16625 (N_16625,N_16155,N_16359);
nand U16626 (N_16626,N_16097,N_16188);
xnor U16627 (N_16627,N_16092,N_16266);
nand U16628 (N_16628,N_16109,N_16161);
xnor U16629 (N_16629,N_16198,N_16043);
xor U16630 (N_16630,N_16401,N_16026);
and U16631 (N_16631,N_16185,N_16486);
and U16632 (N_16632,N_16371,N_16049);
and U16633 (N_16633,N_16496,N_16305);
or U16634 (N_16634,N_16361,N_16073);
nand U16635 (N_16635,N_16471,N_16034);
nand U16636 (N_16636,N_16250,N_16285);
nor U16637 (N_16637,N_16388,N_16290);
nand U16638 (N_16638,N_16111,N_16065);
nand U16639 (N_16639,N_16088,N_16055);
and U16640 (N_16640,N_16086,N_16319);
nand U16641 (N_16641,N_16151,N_16267);
and U16642 (N_16642,N_16178,N_16449);
nand U16643 (N_16643,N_16344,N_16174);
nor U16644 (N_16644,N_16219,N_16461);
or U16645 (N_16645,N_16362,N_16206);
xnor U16646 (N_16646,N_16202,N_16222);
or U16647 (N_16647,N_16444,N_16417);
nand U16648 (N_16648,N_16386,N_16143);
xnor U16649 (N_16649,N_16482,N_16142);
nand U16650 (N_16650,N_16057,N_16165);
nor U16651 (N_16651,N_16252,N_16363);
or U16652 (N_16652,N_16342,N_16122);
or U16653 (N_16653,N_16411,N_16484);
and U16654 (N_16654,N_16452,N_16090);
and U16655 (N_16655,N_16076,N_16137);
nor U16656 (N_16656,N_16157,N_16167);
xnor U16657 (N_16657,N_16159,N_16302);
nor U16658 (N_16658,N_16245,N_16032);
and U16659 (N_16659,N_16207,N_16232);
nor U16660 (N_16660,N_16312,N_16036);
xnor U16661 (N_16661,N_16412,N_16478);
nand U16662 (N_16662,N_16098,N_16284);
xnor U16663 (N_16663,N_16495,N_16042);
nand U16664 (N_16664,N_16253,N_16414);
nand U16665 (N_16665,N_16031,N_16181);
and U16666 (N_16666,N_16445,N_16041);
nor U16667 (N_16667,N_16164,N_16331);
nand U16668 (N_16668,N_16339,N_16492);
nor U16669 (N_16669,N_16399,N_16210);
xor U16670 (N_16670,N_16186,N_16223);
nor U16671 (N_16671,N_16436,N_16292);
and U16672 (N_16672,N_16301,N_16082);
and U16673 (N_16673,N_16273,N_16270);
nor U16674 (N_16674,N_16262,N_16372);
and U16675 (N_16675,N_16072,N_16204);
nor U16676 (N_16676,N_16200,N_16121);
and U16677 (N_16677,N_16400,N_16466);
or U16678 (N_16678,N_16416,N_16012);
nand U16679 (N_16679,N_16056,N_16450);
or U16680 (N_16680,N_16149,N_16472);
xor U16681 (N_16681,N_16085,N_16269);
xnor U16682 (N_16682,N_16220,N_16296);
or U16683 (N_16683,N_16117,N_16261);
and U16684 (N_16684,N_16443,N_16357);
and U16685 (N_16685,N_16158,N_16150);
nand U16686 (N_16686,N_16488,N_16028);
nand U16687 (N_16687,N_16183,N_16037);
or U16688 (N_16688,N_16214,N_16340);
xnor U16689 (N_16689,N_16360,N_16213);
xor U16690 (N_16690,N_16163,N_16406);
xnor U16691 (N_16691,N_16141,N_16227);
nand U16692 (N_16692,N_16099,N_16148);
or U16693 (N_16693,N_16402,N_16393);
nor U16694 (N_16694,N_16133,N_16351);
or U16695 (N_16695,N_16490,N_16474);
xor U16696 (N_16696,N_16384,N_16378);
xor U16697 (N_16697,N_16077,N_16193);
or U16698 (N_16698,N_16118,N_16215);
or U16699 (N_16699,N_16140,N_16240);
nand U16700 (N_16700,N_16275,N_16135);
or U16701 (N_16701,N_16209,N_16341);
nand U16702 (N_16702,N_16364,N_16182);
xnor U16703 (N_16703,N_16475,N_16280);
xor U16704 (N_16704,N_16125,N_16303);
xor U16705 (N_16705,N_16050,N_16435);
or U16706 (N_16706,N_16274,N_16456);
or U16707 (N_16707,N_16311,N_16139);
nand U16708 (N_16708,N_16446,N_16017);
nor U16709 (N_16709,N_16354,N_16177);
and U16710 (N_16710,N_16108,N_16180);
nor U16711 (N_16711,N_16033,N_16014);
and U16712 (N_16712,N_16235,N_16102);
xor U16713 (N_16713,N_16410,N_16239);
xnor U16714 (N_16714,N_16374,N_16468);
or U16715 (N_16715,N_16172,N_16459);
nand U16716 (N_16716,N_16279,N_16131);
nor U16717 (N_16717,N_16203,N_16196);
xnor U16718 (N_16718,N_16426,N_16338);
and U16719 (N_16719,N_16248,N_16294);
and U16720 (N_16720,N_16487,N_16379);
and U16721 (N_16721,N_16427,N_16030);
or U16722 (N_16722,N_16289,N_16464);
and U16723 (N_16723,N_16216,N_16288);
nor U16724 (N_16724,N_16298,N_16392);
nor U16725 (N_16725,N_16460,N_16278);
nor U16726 (N_16726,N_16293,N_16330);
and U16727 (N_16727,N_16277,N_16346);
and U16728 (N_16728,N_16345,N_16432);
nor U16729 (N_16729,N_16358,N_16353);
nor U16730 (N_16730,N_16429,N_16428);
xnor U16731 (N_16731,N_16039,N_16441);
or U16732 (N_16732,N_16005,N_16007);
or U16733 (N_16733,N_16365,N_16457);
or U16734 (N_16734,N_16380,N_16021);
nand U16735 (N_16735,N_16323,N_16093);
nor U16736 (N_16736,N_16020,N_16205);
nor U16737 (N_16737,N_16314,N_16324);
and U16738 (N_16738,N_16087,N_16016);
xnor U16739 (N_16739,N_16448,N_16334);
nand U16740 (N_16740,N_16462,N_16024);
nand U16741 (N_16741,N_16497,N_16382);
or U16742 (N_16742,N_16299,N_16265);
or U16743 (N_16743,N_16499,N_16229);
xor U16744 (N_16744,N_16052,N_16413);
or U16745 (N_16745,N_16485,N_16437);
and U16746 (N_16746,N_16367,N_16244);
or U16747 (N_16747,N_16199,N_16337);
nor U16748 (N_16748,N_16124,N_16128);
and U16749 (N_16749,N_16218,N_16251);
nand U16750 (N_16750,N_16169,N_16164);
and U16751 (N_16751,N_16462,N_16393);
nor U16752 (N_16752,N_16380,N_16113);
or U16753 (N_16753,N_16436,N_16273);
xor U16754 (N_16754,N_16351,N_16409);
nand U16755 (N_16755,N_16068,N_16205);
or U16756 (N_16756,N_16380,N_16024);
nand U16757 (N_16757,N_16267,N_16028);
xnor U16758 (N_16758,N_16425,N_16475);
xnor U16759 (N_16759,N_16415,N_16157);
and U16760 (N_16760,N_16082,N_16361);
xor U16761 (N_16761,N_16494,N_16463);
or U16762 (N_16762,N_16042,N_16251);
nand U16763 (N_16763,N_16487,N_16408);
nor U16764 (N_16764,N_16204,N_16054);
nor U16765 (N_16765,N_16194,N_16245);
and U16766 (N_16766,N_16404,N_16422);
and U16767 (N_16767,N_16319,N_16287);
or U16768 (N_16768,N_16117,N_16078);
xnor U16769 (N_16769,N_16220,N_16354);
and U16770 (N_16770,N_16344,N_16411);
nand U16771 (N_16771,N_16249,N_16318);
nor U16772 (N_16772,N_16102,N_16163);
or U16773 (N_16773,N_16033,N_16438);
nand U16774 (N_16774,N_16034,N_16138);
nor U16775 (N_16775,N_16477,N_16225);
and U16776 (N_16776,N_16157,N_16344);
nor U16777 (N_16777,N_16063,N_16007);
xor U16778 (N_16778,N_16304,N_16074);
xnor U16779 (N_16779,N_16052,N_16299);
or U16780 (N_16780,N_16408,N_16314);
and U16781 (N_16781,N_16134,N_16331);
nor U16782 (N_16782,N_16241,N_16410);
or U16783 (N_16783,N_16341,N_16348);
xor U16784 (N_16784,N_16332,N_16131);
nand U16785 (N_16785,N_16052,N_16378);
nand U16786 (N_16786,N_16482,N_16404);
nand U16787 (N_16787,N_16053,N_16393);
and U16788 (N_16788,N_16126,N_16187);
nand U16789 (N_16789,N_16276,N_16182);
nand U16790 (N_16790,N_16267,N_16449);
and U16791 (N_16791,N_16151,N_16413);
nor U16792 (N_16792,N_16115,N_16093);
xor U16793 (N_16793,N_16057,N_16051);
nor U16794 (N_16794,N_16297,N_16177);
or U16795 (N_16795,N_16347,N_16337);
or U16796 (N_16796,N_16442,N_16453);
or U16797 (N_16797,N_16354,N_16249);
nand U16798 (N_16798,N_16045,N_16288);
or U16799 (N_16799,N_16093,N_16306);
nand U16800 (N_16800,N_16421,N_16387);
xnor U16801 (N_16801,N_16062,N_16057);
or U16802 (N_16802,N_16127,N_16301);
or U16803 (N_16803,N_16041,N_16199);
and U16804 (N_16804,N_16269,N_16126);
nor U16805 (N_16805,N_16040,N_16039);
nor U16806 (N_16806,N_16133,N_16331);
nand U16807 (N_16807,N_16284,N_16385);
nor U16808 (N_16808,N_16179,N_16454);
or U16809 (N_16809,N_16182,N_16154);
nand U16810 (N_16810,N_16172,N_16133);
and U16811 (N_16811,N_16438,N_16153);
xnor U16812 (N_16812,N_16420,N_16386);
nor U16813 (N_16813,N_16320,N_16181);
nor U16814 (N_16814,N_16457,N_16262);
nor U16815 (N_16815,N_16132,N_16257);
nand U16816 (N_16816,N_16055,N_16425);
nor U16817 (N_16817,N_16283,N_16263);
nor U16818 (N_16818,N_16255,N_16394);
xnor U16819 (N_16819,N_16053,N_16210);
nor U16820 (N_16820,N_16142,N_16126);
and U16821 (N_16821,N_16326,N_16014);
xnor U16822 (N_16822,N_16356,N_16222);
xnor U16823 (N_16823,N_16234,N_16326);
xnor U16824 (N_16824,N_16423,N_16020);
nand U16825 (N_16825,N_16043,N_16057);
nand U16826 (N_16826,N_16160,N_16442);
xor U16827 (N_16827,N_16105,N_16108);
xor U16828 (N_16828,N_16228,N_16273);
xnor U16829 (N_16829,N_16482,N_16416);
or U16830 (N_16830,N_16194,N_16449);
and U16831 (N_16831,N_16339,N_16239);
nand U16832 (N_16832,N_16124,N_16029);
nand U16833 (N_16833,N_16194,N_16161);
nor U16834 (N_16834,N_16004,N_16426);
xnor U16835 (N_16835,N_16457,N_16232);
or U16836 (N_16836,N_16125,N_16326);
and U16837 (N_16837,N_16408,N_16086);
nor U16838 (N_16838,N_16405,N_16332);
xor U16839 (N_16839,N_16316,N_16421);
nand U16840 (N_16840,N_16106,N_16082);
nand U16841 (N_16841,N_16371,N_16269);
nand U16842 (N_16842,N_16070,N_16198);
nor U16843 (N_16843,N_16366,N_16252);
or U16844 (N_16844,N_16042,N_16436);
nand U16845 (N_16845,N_16205,N_16025);
or U16846 (N_16846,N_16426,N_16137);
xnor U16847 (N_16847,N_16358,N_16097);
and U16848 (N_16848,N_16159,N_16404);
nand U16849 (N_16849,N_16153,N_16313);
and U16850 (N_16850,N_16489,N_16066);
nor U16851 (N_16851,N_16354,N_16306);
nor U16852 (N_16852,N_16364,N_16268);
or U16853 (N_16853,N_16215,N_16389);
nand U16854 (N_16854,N_16075,N_16192);
nand U16855 (N_16855,N_16347,N_16067);
or U16856 (N_16856,N_16207,N_16410);
and U16857 (N_16857,N_16285,N_16188);
nand U16858 (N_16858,N_16437,N_16231);
and U16859 (N_16859,N_16479,N_16271);
or U16860 (N_16860,N_16354,N_16395);
nand U16861 (N_16861,N_16021,N_16154);
nand U16862 (N_16862,N_16114,N_16227);
nor U16863 (N_16863,N_16380,N_16193);
xnor U16864 (N_16864,N_16466,N_16358);
and U16865 (N_16865,N_16130,N_16180);
nor U16866 (N_16866,N_16290,N_16227);
and U16867 (N_16867,N_16135,N_16255);
nand U16868 (N_16868,N_16079,N_16117);
or U16869 (N_16869,N_16030,N_16098);
nand U16870 (N_16870,N_16233,N_16318);
or U16871 (N_16871,N_16085,N_16218);
and U16872 (N_16872,N_16372,N_16397);
nor U16873 (N_16873,N_16352,N_16443);
nor U16874 (N_16874,N_16214,N_16291);
or U16875 (N_16875,N_16444,N_16003);
xnor U16876 (N_16876,N_16064,N_16159);
and U16877 (N_16877,N_16001,N_16452);
or U16878 (N_16878,N_16234,N_16253);
nor U16879 (N_16879,N_16089,N_16494);
nand U16880 (N_16880,N_16211,N_16168);
nand U16881 (N_16881,N_16155,N_16318);
nor U16882 (N_16882,N_16070,N_16045);
and U16883 (N_16883,N_16453,N_16061);
or U16884 (N_16884,N_16126,N_16178);
nor U16885 (N_16885,N_16237,N_16318);
nor U16886 (N_16886,N_16398,N_16350);
nand U16887 (N_16887,N_16140,N_16165);
nand U16888 (N_16888,N_16100,N_16378);
nand U16889 (N_16889,N_16233,N_16312);
xor U16890 (N_16890,N_16188,N_16417);
xnor U16891 (N_16891,N_16346,N_16311);
xor U16892 (N_16892,N_16465,N_16302);
nor U16893 (N_16893,N_16259,N_16362);
nor U16894 (N_16894,N_16155,N_16219);
xor U16895 (N_16895,N_16141,N_16096);
xnor U16896 (N_16896,N_16292,N_16111);
or U16897 (N_16897,N_16463,N_16133);
xnor U16898 (N_16898,N_16405,N_16380);
xor U16899 (N_16899,N_16322,N_16207);
nand U16900 (N_16900,N_16254,N_16342);
and U16901 (N_16901,N_16035,N_16497);
nor U16902 (N_16902,N_16428,N_16166);
and U16903 (N_16903,N_16142,N_16268);
nor U16904 (N_16904,N_16194,N_16089);
or U16905 (N_16905,N_16001,N_16157);
or U16906 (N_16906,N_16090,N_16008);
or U16907 (N_16907,N_16158,N_16196);
and U16908 (N_16908,N_16152,N_16475);
or U16909 (N_16909,N_16114,N_16219);
and U16910 (N_16910,N_16374,N_16194);
and U16911 (N_16911,N_16119,N_16236);
nand U16912 (N_16912,N_16011,N_16367);
nor U16913 (N_16913,N_16041,N_16081);
xor U16914 (N_16914,N_16178,N_16483);
or U16915 (N_16915,N_16224,N_16298);
xnor U16916 (N_16916,N_16060,N_16236);
nand U16917 (N_16917,N_16206,N_16222);
nand U16918 (N_16918,N_16277,N_16419);
and U16919 (N_16919,N_16481,N_16312);
nor U16920 (N_16920,N_16487,N_16321);
nand U16921 (N_16921,N_16284,N_16253);
xor U16922 (N_16922,N_16126,N_16333);
nor U16923 (N_16923,N_16480,N_16395);
nand U16924 (N_16924,N_16269,N_16022);
xnor U16925 (N_16925,N_16176,N_16102);
nand U16926 (N_16926,N_16026,N_16021);
nand U16927 (N_16927,N_16281,N_16353);
nand U16928 (N_16928,N_16462,N_16423);
nor U16929 (N_16929,N_16355,N_16362);
nor U16930 (N_16930,N_16080,N_16097);
and U16931 (N_16931,N_16350,N_16447);
or U16932 (N_16932,N_16165,N_16315);
xor U16933 (N_16933,N_16259,N_16236);
nor U16934 (N_16934,N_16328,N_16299);
nor U16935 (N_16935,N_16216,N_16204);
nand U16936 (N_16936,N_16256,N_16447);
nor U16937 (N_16937,N_16124,N_16221);
and U16938 (N_16938,N_16239,N_16342);
and U16939 (N_16939,N_16231,N_16236);
xor U16940 (N_16940,N_16356,N_16226);
or U16941 (N_16941,N_16214,N_16176);
or U16942 (N_16942,N_16358,N_16170);
or U16943 (N_16943,N_16007,N_16014);
or U16944 (N_16944,N_16138,N_16132);
xor U16945 (N_16945,N_16189,N_16345);
nor U16946 (N_16946,N_16328,N_16303);
and U16947 (N_16947,N_16253,N_16141);
nand U16948 (N_16948,N_16080,N_16170);
nor U16949 (N_16949,N_16095,N_16122);
or U16950 (N_16950,N_16353,N_16240);
xnor U16951 (N_16951,N_16168,N_16017);
or U16952 (N_16952,N_16413,N_16274);
xor U16953 (N_16953,N_16196,N_16026);
xnor U16954 (N_16954,N_16301,N_16493);
nor U16955 (N_16955,N_16315,N_16175);
and U16956 (N_16956,N_16482,N_16454);
nor U16957 (N_16957,N_16202,N_16072);
or U16958 (N_16958,N_16052,N_16482);
or U16959 (N_16959,N_16090,N_16336);
and U16960 (N_16960,N_16037,N_16281);
or U16961 (N_16961,N_16064,N_16418);
and U16962 (N_16962,N_16014,N_16061);
xor U16963 (N_16963,N_16046,N_16244);
or U16964 (N_16964,N_16183,N_16196);
nand U16965 (N_16965,N_16448,N_16083);
nor U16966 (N_16966,N_16089,N_16353);
nor U16967 (N_16967,N_16070,N_16442);
and U16968 (N_16968,N_16453,N_16497);
xor U16969 (N_16969,N_16279,N_16370);
or U16970 (N_16970,N_16480,N_16125);
or U16971 (N_16971,N_16374,N_16120);
nor U16972 (N_16972,N_16320,N_16073);
and U16973 (N_16973,N_16492,N_16063);
or U16974 (N_16974,N_16161,N_16237);
and U16975 (N_16975,N_16277,N_16431);
nand U16976 (N_16976,N_16150,N_16292);
nor U16977 (N_16977,N_16227,N_16345);
or U16978 (N_16978,N_16119,N_16380);
or U16979 (N_16979,N_16418,N_16192);
nor U16980 (N_16980,N_16194,N_16323);
nor U16981 (N_16981,N_16132,N_16121);
xor U16982 (N_16982,N_16413,N_16142);
nor U16983 (N_16983,N_16300,N_16190);
nor U16984 (N_16984,N_16200,N_16317);
xnor U16985 (N_16985,N_16307,N_16347);
and U16986 (N_16986,N_16300,N_16348);
nand U16987 (N_16987,N_16267,N_16442);
nor U16988 (N_16988,N_16046,N_16275);
and U16989 (N_16989,N_16187,N_16136);
nor U16990 (N_16990,N_16083,N_16361);
nand U16991 (N_16991,N_16140,N_16125);
xnor U16992 (N_16992,N_16476,N_16411);
and U16993 (N_16993,N_16163,N_16219);
nor U16994 (N_16994,N_16406,N_16035);
nand U16995 (N_16995,N_16218,N_16069);
xnor U16996 (N_16996,N_16407,N_16460);
nand U16997 (N_16997,N_16474,N_16001);
xnor U16998 (N_16998,N_16175,N_16216);
nor U16999 (N_16999,N_16323,N_16177);
nand U17000 (N_17000,N_16514,N_16679);
nand U17001 (N_17001,N_16928,N_16548);
nor U17002 (N_17002,N_16525,N_16870);
and U17003 (N_17003,N_16619,N_16644);
nor U17004 (N_17004,N_16827,N_16549);
or U17005 (N_17005,N_16746,N_16797);
xnor U17006 (N_17006,N_16999,N_16680);
or U17007 (N_17007,N_16925,N_16979);
or U17008 (N_17008,N_16556,N_16992);
nand U17009 (N_17009,N_16778,N_16875);
nand U17010 (N_17010,N_16840,N_16788);
nor U17011 (N_17011,N_16735,N_16758);
or U17012 (N_17012,N_16555,N_16537);
or U17013 (N_17013,N_16609,N_16569);
nand U17014 (N_17014,N_16906,N_16536);
xnor U17015 (N_17015,N_16707,N_16576);
or U17016 (N_17016,N_16708,N_16553);
xor U17017 (N_17017,N_16658,N_16752);
nor U17018 (N_17018,N_16688,N_16581);
and U17019 (N_17019,N_16937,N_16511);
nor U17020 (N_17020,N_16828,N_16844);
nor U17021 (N_17021,N_16886,N_16820);
and U17022 (N_17022,N_16868,N_16583);
or U17023 (N_17023,N_16584,N_16878);
nor U17024 (N_17024,N_16572,N_16745);
and U17025 (N_17025,N_16803,N_16712);
nand U17026 (N_17026,N_16736,N_16591);
xor U17027 (N_17027,N_16653,N_16987);
and U17028 (N_17028,N_16869,N_16633);
nor U17029 (N_17029,N_16782,N_16718);
and U17030 (N_17030,N_16675,N_16663);
nand U17031 (N_17031,N_16903,N_16952);
and U17032 (N_17032,N_16704,N_16655);
or U17033 (N_17033,N_16622,N_16734);
nor U17034 (N_17034,N_16770,N_16682);
nand U17035 (N_17035,N_16776,N_16777);
nand U17036 (N_17036,N_16931,N_16709);
nor U17037 (N_17037,N_16919,N_16687);
nor U17038 (N_17038,N_16713,N_16754);
xnor U17039 (N_17039,N_16836,N_16551);
and U17040 (N_17040,N_16528,N_16898);
and U17041 (N_17041,N_16970,N_16599);
nor U17042 (N_17042,N_16539,N_16524);
nand U17043 (N_17043,N_16699,N_16690);
or U17044 (N_17044,N_16966,N_16516);
and U17045 (N_17045,N_16637,N_16862);
and U17046 (N_17046,N_16825,N_16748);
nand U17047 (N_17047,N_16535,N_16888);
and U17048 (N_17048,N_16686,N_16676);
xnor U17049 (N_17049,N_16985,N_16720);
or U17050 (N_17050,N_16550,N_16650);
and U17051 (N_17051,N_16726,N_16911);
xor U17052 (N_17052,N_16649,N_16916);
and U17053 (N_17053,N_16750,N_16672);
xor U17054 (N_17054,N_16849,N_16697);
and U17055 (N_17055,N_16765,N_16645);
nor U17056 (N_17056,N_16821,N_16538);
nand U17057 (N_17057,N_16560,N_16808);
nand U17058 (N_17058,N_16507,N_16625);
nand U17059 (N_17059,N_16744,N_16900);
or U17060 (N_17060,N_16986,N_16833);
and U17061 (N_17061,N_16968,N_16879);
nand U17062 (N_17062,N_16795,N_16781);
or U17063 (N_17063,N_16897,N_16700);
nand U17064 (N_17064,N_16544,N_16978);
and U17065 (N_17065,N_16580,N_16755);
nor U17066 (N_17066,N_16729,N_16960);
nand U17067 (N_17067,N_16895,N_16670);
nor U17068 (N_17068,N_16956,N_16927);
or U17069 (N_17069,N_16858,N_16905);
nand U17070 (N_17070,N_16856,N_16739);
nand U17071 (N_17071,N_16588,N_16640);
and U17072 (N_17072,N_16958,N_16684);
and U17073 (N_17073,N_16520,N_16772);
xnor U17074 (N_17074,N_16989,N_16616);
or U17075 (N_17075,N_16972,N_16817);
and U17076 (N_17076,N_16936,N_16711);
and U17077 (N_17077,N_16839,N_16554);
nand U17078 (N_17078,N_16872,N_16501);
or U17079 (N_17079,N_16615,N_16894);
and U17080 (N_17080,N_16998,N_16961);
or U17081 (N_17081,N_16683,N_16922);
and U17082 (N_17082,N_16887,N_16692);
xor U17083 (N_17083,N_16941,N_16620);
nor U17084 (N_17084,N_16882,N_16678);
and U17085 (N_17085,N_16890,N_16757);
and U17086 (N_17086,N_16863,N_16626);
xnor U17087 (N_17087,N_16629,N_16673);
and U17088 (N_17088,N_16769,N_16592);
nor U17089 (N_17089,N_16610,N_16988);
nor U17090 (N_17090,N_16871,N_16908);
or U17091 (N_17091,N_16743,N_16723);
xor U17092 (N_17092,N_16587,N_16603);
and U17093 (N_17093,N_16873,N_16502);
or U17094 (N_17094,N_16984,N_16607);
nor U17095 (N_17095,N_16510,N_16977);
nor U17096 (N_17096,N_16593,N_16740);
nor U17097 (N_17097,N_16864,N_16799);
xnor U17098 (N_17098,N_16768,N_16913);
or U17099 (N_17099,N_16693,N_16598);
nor U17100 (N_17100,N_16596,N_16793);
and U17101 (N_17101,N_16563,N_16889);
nor U17102 (N_17102,N_16847,N_16689);
and U17103 (N_17103,N_16706,N_16855);
or U17104 (N_17104,N_16866,N_16814);
or U17105 (N_17105,N_16842,N_16737);
and U17106 (N_17106,N_16834,N_16955);
xnor U17107 (N_17107,N_16945,N_16741);
xor U17108 (N_17108,N_16585,N_16660);
nand U17109 (N_17109,N_16606,N_16786);
and U17110 (N_17110,N_16779,N_16874);
or U17111 (N_17111,N_16509,N_16976);
and U17112 (N_17112,N_16921,N_16618);
nor U17113 (N_17113,N_16896,N_16621);
xnor U17114 (N_17114,N_16794,N_16969);
nor U17115 (N_17115,N_16807,N_16639);
xor U17116 (N_17116,N_16933,N_16954);
or U17117 (N_17117,N_16943,N_16613);
and U17118 (N_17118,N_16738,N_16843);
and U17119 (N_17119,N_16796,N_16590);
and U17120 (N_17120,N_16751,N_16506);
or U17121 (N_17121,N_16865,N_16608);
nand U17122 (N_17122,N_16651,N_16627);
nor U17123 (N_17123,N_16950,N_16915);
or U17124 (N_17124,N_16791,N_16631);
and U17125 (N_17125,N_16767,N_16891);
nand U17126 (N_17126,N_16717,N_16567);
and U17127 (N_17127,N_16540,N_16636);
nor U17128 (N_17128,N_16574,N_16910);
nor U17129 (N_17129,N_16851,N_16532);
and U17130 (N_17130,N_16826,N_16545);
nand U17131 (N_17131,N_16932,N_16527);
or U17132 (N_17132,N_16638,N_16760);
and U17133 (N_17133,N_16668,N_16573);
or U17134 (N_17134,N_16824,N_16561);
and U17135 (N_17135,N_16694,N_16727);
xor U17136 (N_17136,N_16732,N_16703);
nor U17137 (N_17137,N_16991,N_16518);
nor U17138 (N_17138,N_16918,N_16806);
nand U17139 (N_17139,N_16946,N_16594);
or U17140 (N_17140,N_16996,N_16800);
or U17141 (N_17141,N_16571,N_16657);
and U17142 (N_17142,N_16881,N_16531);
or U17143 (N_17143,N_16812,N_16541);
or U17144 (N_17144,N_16964,N_16790);
xnor U17145 (N_17145,N_16747,N_16696);
xnor U17146 (N_17146,N_16837,N_16530);
nand U17147 (N_17147,N_16677,N_16938);
xor U17148 (N_17148,N_16764,N_16801);
xnor U17149 (N_17149,N_16517,N_16995);
xor U17150 (N_17150,N_16940,N_16893);
and U17151 (N_17151,N_16939,N_16892);
and U17152 (N_17152,N_16522,N_16601);
nand U17153 (N_17153,N_16733,N_16557);
or U17154 (N_17154,N_16597,N_16646);
or U17155 (N_17155,N_16611,N_16722);
nand U17156 (N_17156,N_16953,N_16762);
nor U17157 (N_17157,N_16578,N_16665);
or U17158 (N_17158,N_16831,N_16546);
or U17159 (N_17159,N_16914,N_16787);
xnor U17160 (N_17160,N_16512,N_16813);
and U17161 (N_17161,N_16965,N_16508);
or U17162 (N_17162,N_16789,N_16642);
or U17163 (N_17163,N_16835,N_16997);
nand U17164 (N_17164,N_16829,N_16771);
or U17165 (N_17165,N_16920,N_16529);
and U17166 (N_17166,N_16761,N_16785);
xnor U17167 (N_17167,N_16500,N_16861);
nand U17168 (N_17168,N_16853,N_16804);
nor U17169 (N_17169,N_16564,N_16917);
nand U17170 (N_17170,N_16542,N_16568);
and U17171 (N_17171,N_16774,N_16515);
or U17172 (N_17172,N_16852,N_16521);
xor U17173 (N_17173,N_16652,N_16883);
nand U17174 (N_17174,N_16749,N_16805);
nor U17175 (N_17175,N_16662,N_16559);
and U17176 (N_17176,N_16582,N_16702);
nand U17177 (N_17177,N_16534,N_16533);
and U17178 (N_17178,N_16565,N_16698);
or U17179 (N_17179,N_16595,N_16973);
and U17180 (N_17180,N_16763,N_16980);
or U17181 (N_17181,N_16884,N_16605);
and U17182 (N_17182,N_16944,N_16635);
nand U17183 (N_17183,N_16957,N_16775);
and U17184 (N_17184,N_16959,N_16859);
nand U17185 (N_17185,N_16586,N_16513);
and U17186 (N_17186,N_16730,N_16523);
nor U17187 (N_17187,N_16857,N_16691);
or U17188 (N_17188,N_16876,N_16798);
nand U17189 (N_17189,N_16543,N_16634);
nand U17190 (N_17190,N_16845,N_16783);
xnor U17191 (N_17191,N_16671,N_16681);
nand U17192 (N_17192,N_16742,N_16600);
and U17193 (N_17193,N_16810,N_16784);
xnor U17194 (N_17194,N_16942,N_16867);
xor U17195 (N_17195,N_16721,N_16624);
xor U17196 (N_17196,N_16664,N_16714);
nand U17197 (N_17197,N_16983,N_16562);
and U17198 (N_17198,N_16674,N_16641);
xor U17199 (N_17199,N_16811,N_16993);
or U17200 (N_17200,N_16885,N_16981);
nor U17201 (N_17201,N_16930,N_16899);
nor U17202 (N_17202,N_16630,N_16850);
nor U17203 (N_17203,N_16552,N_16654);
nor U17204 (N_17204,N_16659,N_16759);
or U17205 (N_17205,N_16710,N_16728);
nand U17206 (N_17206,N_16623,N_16695);
and U17207 (N_17207,N_16628,N_16909);
or U17208 (N_17208,N_16602,N_16974);
nand U17209 (N_17209,N_16948,N_16614);
and U17210 (N_17210,N_16612,N_16715);
nand U17211 (N_17211,N_16832,N_16926);
xnor U17212 (N_17212,N_16830,N_16815);
xnor U17213 (N_17213,N_16773,N_16971);
xnor U17214 (N_17214,N_16951,N_16724);
or U17215 (N_17215,N_16579,N_16802);
and U17216 (N_17216,N_16823,N_16575);
or U17217 (N_17217,N_16648,N_16901);
and U17218 (N_17218,N_16780,N_16547);
or U17219 (N_17219,N_16846,N_16725);
nor U17220 (N_17220,N_16577,N_16990);
or U17221 (N_17221,N_16617,N_16935);
and U17222 (N_17222,N_16841,N_16570);
or U17223 (N_17223,N_16589,N_16904);
and U17224 (N_17224,N_16902,N_16912);
and U17225 (N_17225,N_16719,N_16854);
and U17226 (N_17226,N_16505,N_16822);
nor U17227 (N_17227,N_16924,N_16818);
nor U17228 (N_17228,N_16923,N_16604);
nor U17229 (N_17229,N_16967,N_16656);
nand U17230 (N_17230,N_16929,N_16982);
or U17231 (N_17231,N_16877,N_16643);
nand U17232 (N_17232,N_16766,N_16949);
and U17233 (N_17233,N_16809,N_16962);
or U17234 (N_17234,N_16566,N_16819);
nand U17235 (N_17235,N_16963,N_16503);
and U17236 (N_17236,N_16792,N_16848);
and U17237 (N_17237,N_16753,N_16731);
and U17238 (N_17238,N_16716,N_16816);
xnor U17239 (N_17239,N_16504,N_16685);
and U17240 (N_17240,N_16669,N_16934);
nor U17241 (N_17241,N_16975,N_16666);
xor U17242 (N_17242,N_16705,N_16667);
nor U17243 (N_17243,N_16661,N_16860);
xnor U17244 (N_17244,N_16838,N_16880);
xor U17245 (N_17245,N_16526,N_16701);
nand U17246 (N_17246,N_16519,N_16994);
and U17247 (N_17247,N_16632,N_16907);
or U17248 (N_17248,N_16558,N_16647);
nand U17249 (N_17249,N_16756,N_16947);
nor U17250 (N_17250,N_16710,N_16810);
nor U17251 (N_17251,N_16703,N_16669);
nand U17252 (N_17252,N_16772,N_16662);
nor U17253 (N_17253,N_16968,N_16712);
and U17254 (N_17254,N_16670,N_16746);
xnor U17255 (N_17255,N_16522,N_16941);
xnor U17256 (N_17256,N_16627,N_16706);
xnor U17257 (N_17257,N_16805,N_16523);
nand U17258 (N_17258,N_16593,N_16953);
nand U17259 (N_17259,N_16848,N_16548);
or U17260 (N_17260,N_16978,N_16547);
and U17261 (N_17261,N_16648,N_16885);
xnor U17262 (N_17262,N_16653,N_16526);
nor U17263 (N_17263,N_16814,N_16549);
xor U17264 (N_17264,N_16907,N_16669);
nand U17265 (N_17265,N_16518,N_16724);
xnor U17266 (N_17266,N_16808,N_16781);
nor U17267 (N_17267,N_16781,N_16585);
and U17268 (N_17268,N_16587,N_16869);
nand U17269 (N_17269,N_16792,N_16881);
and U17270 (N_17270,N_16927,N_16901);
nand U17271 (N_17271,N_16811,N_16676);
xnor U17272 (N_17272,N_16925,N_16816);
or U17273 (N_17273,N_16694,N_16622);
nor U17274 (N_17274,N_16578,N_16851);
nand U17275 (N_17275,N_16890,N_16689);
and U17276 (N_17276,N_16644,N_16786);
nor U17277 (N_17277,N_16544,N_16888);
nor U17278 (N_17278,N_16898,N_16505);
xnor U17279 (N_17279,N_16903,N_16853);
xnor U17280 (N_17280,N_16681,N_16632);
or U17281 (N_17281,N_16543,N_16677);
nor U17282 (N_17282,N_16925,N_16524);
xor U17283 (N_17283,N_16574,N_16997);
or U17284 (N_17284,N_16894,N_16624);
nand U17285 (N_17285,N_16930,N_16738);
and U17286 (N_17286,N_16924,N_16962);
or U17287 (N_17287,N_16937,N_16860);
or U17288 (N_17288,N_16934,N_16742);
and U17289 (N_17289,N_16537,N_16533);
nor U17290 (N_17290,N_16516,N_16510);
xor U17291 (N_17291,N_16853,N_16717);
and U17292 (N_17292,N_16634,N_16771);
xor U17293 (N_17293,N_16909,N_16820);
xor U17294 (N_17294,N_16562,N_16515);
nor U17295 (N_17295,N_16924,N_16632);
xnor U17296 (N_17296,N_16516,N_16588);
nand U17297 (N_17297,N_16559,N_16586);
or U17298 (N_17298,N_16880,N_16819);
xnor U17299 (N_17299,N_16984,N_16516);
or U17300 (N_17300,N_16863,N_16577);
or U17301 (N_17301,N_16631,N_16570);
xor U17302 (N_17302,N_16869,N_16912);
nand U17303 (N_17303,N_16757,N_16623);
and U17304 (N_17304,N_16944,N_16649);
and U17305 (N_17305,N_16512,N_16888);
or U17306 (N_17306,N_16689,N_16738);
xnor U17307 (N_17307,N_16597,N_16561);
xnor U17308 (N_17308,N_16901,N_16643);
nor U17309 (N_17309,N_16850,N_16949);
or U17310 (N_17310,N_16986,N_16602);
xor U17311 (N_17311,N_16572,N_16962);
nand U17312 (N_17312,N_16695,N_16982);
nand U17313 (N_17313,N_16500,N_16548);
and U17314 (N_17314,N_16875,N_16666);
nor U17315 (N_17315,N_16992,N_16598);
or U17316 (N_17316,N_16611,N_16687);
and U17317 (N_17317,N_16668,N_16927);
nand U17318 (N_17318,N_16779,N_16650);
nand U17319 (N_17319,N_16817,N_16871);
or U17320 (N_17320,N_16823,N_16983);
xor U17321 (N_17321,N_16562,N_16533);
or U17322 (N_17322,N_16648,N_16934);
or U17323 (N_17323,N_16957,N_16823);
xnor U17324 (N_17324,N_16569,N_16671);
nand U17325 (N_17325,N_16673,N_16780);
or U17326 (N_17326,N_16716,N_16774);
xnor U17327 (N_17327,N_16786,N_16594);
nor U17328 (N_17328,N_16835,N_16634);
and U17329 (N_17329,N_16806,N_16614);
nor U17330 (N_17330,N_16515,N_16518);
or U17331 (N_17331,N_16975,N_16848);
or U17332 (N_17332,N_16686,N_16632);
xnor U17333 (N_17333,N_16914,N_16819);
nand U17334 (N_17334,N_16596,N_16531);
or U17335 (N_17335,N_16758,N_16700);
xor U17336 (N_17336,N_16989,N_16819);
nor U17337 (N_17337,N_16990,N_16890);
or U17338 (N_17338,N_16995,N_16548);
or U17339 (N_17339,N_16960,N_16864);
nand U17340 (N_17340,N_16656,N_16773);
xnor U17341 (N_17341,N_16622,N_16838);
and U17342 (N_17342,N_16962,N_16708);
and U17343 (N_17343,N_16600,N_16530);
nand U17344 (N_17344,N_16735,N_16772);
and U17345 (N_17345,N_16914,N_16540);
xor U17346 (N_17346,N_16734,N_16737);
xnor U17347 (N_17347,N_16879,N_16999);
nor U17348 (N_17348,N_16811,N_16891);
or U17349 (N_17349,N_16604,N_16581);
nor U17350 (N_17350,N_16736,N_16800);
nor U17351 (N_17351,N_16939,N_16582);
and U17352 (N_17352,N_16626,N_16514);
and U17353 (N_17353,N_16539,N_16919);
xor U17354 (N_17354,N_16885,N_16770);
nand U17355 (N_17355,N_16924,N_16862);
xnor U17356 (N_17356,N_16696,N_16644);
and U17357 (N_17357,N_16955,N_16600);
nand U17358 (N_17358,N_16593,N_16952);
or U17359 (N_17359,N_16706,N_16715);
or U17360 (N_17360,N_16906,N_16966);
nand U17361 (N_17361,N_16681,N_16850);
nand U17362 (N_17362,N_16885,N_16891);
nand U17363 (N_17363,N_16599,N_16808);
nand U17364 (N_17364,N_16972,N_16769);
xor U17365 (N_17365,N_16550,N_16644);
nand U17366 (N_17366,N_16820,N_16731);
and U17367 (N_17367,N_16579,N_16790);
or U17368 (N_17368,N_16693,N_16663);
nor U17369 (N_17369,N_16995,N_16920);
or U17370 (N_17370,N_16721,N_16789);
and U17371 (N_17371,N_16815,N_16841);
nand U17372 (N_17372,N_16661,N_16520);
nand U17373 (N_17373,N_16746,N_16936);
or U17374 (N_17374,N_16769,N_16747);
nor U17375 (N_17375,N_16666,N_16932);
nand U17376 (N_17376,N_16715,N_16831);
or U17377 (N_17377,N_16643,N_16891);
or U17378 (N_17378,N_16832,N_16923);
xnor U17379 (N_17379,N_16566,N_16542);
nand U17380 (N_17380,N_16838,N_16912);
and U17381 (N_17381,N_16828,N_16684);
xor U17382 (N_17382,N_16671,N_16888);
or U17383 (N_17383,N_16868,N_16532);
nand U17384 (N_17384,N_16906,N_16988);
nor U17385 (N_17385,N_16502,N_16843);
and U17386 (N_17386,N_16833,N_16670);
or U17387 (N_17387,N_16959,N_16609);
xnor U17388 (N_17388,N_16646,N_16755);
and U17389 (N_17389,N_16609,N_16655);
xnor U17390 (N_17390,N_16739,N_16661);
and U17391 (N_17391,N_16958,N_16651);
or U17392 (N_17392,N_16968,N_16999);
nor U17393 (N_17393,N_16851,N_16850);
nand U17394 (N_17394,N_16949,N_16505);
or U17395 (N_17395,N_16573,N_16716);
xor U17396 (N_17396,N_16514,N_16983);
nor U17397 (N_17397,N_16873,N_16874);
nor U17398 (N_17398,N_16933,N_16699);
nor U17399 (N_17399,N_16686,N_16866);
xor U17400 (N_17400,N_16856,N_16776);
nor U17401 (N_17401,N_16842,N_16962);
xor U17402 (N_17402,N_16885,N_16760);
xor U17403 (N_17403,N_16682,N_16543);
nand U17404 (N_17404,N_16797,N_16901);
nor U17405 (N_17405,N_16708,N_16641);
and U17406 (N_17406,N_16501,N_16570);
nand U17407 (N_17407,N_16773,N_16597);
nor U17408 (N_17408,N_16813,N_16917);
or U17409 (N_17409,N_16617,N_16994);
nand U17410 (N_17410,N_16931,N_16873);
nand U17411 (N_17411,N_16540,N_16527);
nand U17412 (N_17412,N_16795,N_16578);
or U17413 (N_17413,N_16816,N_16536);
xor U17414 (N_17414,N_16576,N_16834);
nor U17415 (N_17415,N_16722,N_16714);
and U17416 (N_17416,N_16920,N_16619);
or U17417 (N_17417,N_16921,N_16508);
xnor U17418 (N_17418,N_16855,N_16808);
xor U17419 (N_17419,N_16702,N_16686);
or U17420 (N_17420,N_16531,N_16640);
nor U17421 (N_17421,N_16672,N_16500);
xor U17422 (N_17422,N_16873,N_16946);
nand U17423 (N_17423,N_16604,N_16516);
xor U17424 (N_17424,N_16567,N_16582);
nor U17425 (N_17425,N_16667,N_16826);
and U17426 (N_17426,N_16778,N_16761);
or U17427 (N_17427,N_16816,N_16791);
and U17428 (N_17428,N_16508,N_16745);
or U17429 (N_17429,N_16648,N_16672);
and U17430 (N_17430,N_16672,N_16983);
nor U17431 (N_17431,N_16694,N_16784);
or U17432 (N_17432,N_16511,N_16833);
xor U17433 (N_17433,N_16725,N_16553);
or U17434 (N_17434,N_16994,N_16704);
or U17435 (N_17435,N_16864,N_16844);
or U17436 (N_17436,N_16598,N_16999);
and U17437 (N_17437,N_16635,N_16670);
nor U17438 (N_17438,N_16986,N_16615);
nor U17439 (N_17439,N_16573,N_16871);
and U17440 (N_17440,N_16877,N_16893);
or U17441 (N_17441,N_16834,N_16803);
xnor U17442 (N_17442,N_16783,N_16549);
and U17443 (N_17443,N_16780,N_16786);
nor U17444 (N_17444,N_16975,N_16586);
or U17445 (N_17445,N_16842,N_16548);
and U17446 (N_17446,N_16555,N_16660);
xnor U17447 (N_17447,N_16633,N_16934);
or U17448 (N_17448,N_16897,N_16871);
xor U17449 (N_17449,N_16600,N_16860);
nor U17450 (N_17450,N_16664,N_16606);
nand U17451 (N_17451,N_16708,N_16647);
and U17452 (N_17452,N_16651,N_16695);
nor U17453 (N_17453,N_16969,N_16921);
or U17454 (N_17454,N_16771,N_16804);
and U17455 (N_17455,N_16960,N_16795);
or U17456 (N_17456,N_16800,N_16603);
and U17457 (N_17457,N_16893,N_16658);
and U17458 (N_17458,N_16663,N_16743);
nand U17459 (N_17459,N_16825,N_16936);
xor U17460 (N_17460,N_16545,N_16960);
nand U17461 (N_17461,N_16589,N_16809);
or U17462 (N_17462,N_16776,N_16871);
nor U17463 (N_17463,N_16993,N_16518);
and U17464 (N_17464,N_16841,N_16616);
nand U17465 (N_17465,N_16839,N_16858);
and U17466 (N_17466,N_16773,N_16945);
xor U17467 (N_17467,N_16961,N_16816);
or U17468 (N_17468,N_16682,N_16518);
nand U17469 (N_17469,N_16638,N_16689);
xnor U17470 (N_17470,N_16758,N_16592);
nor U17471 (N_17471,N_16835,N_16661);
or U17472 (N_17472,N_16650,N_16704);
nand U17473 (N_17473,N_16618,N_16598);
and U17474 (N_17474,N_16674,N_16900);
nand U17475 (N_17475,N_16801,N_16633);
and U17476 (N_17476,N_16910,N_16601);
or U17477 (N_17477,N_16537,N_16991);
or U17478 (N_17478,N_16919,N_16950);
and U17479 (N_17479,N_16885,N_16641);
nor U17480 (N_17480,N_16817,N_16558);
nor U17481 (N_17481,N_16737,N_16954);
or U17482 (N_17482,N_16550,N_16593);
xor U17483 (N_17483,N_16939,N_16710);
nand U17484 (N_17484,N_16807,N_16664);
nor U17485 (N_17485,N_16680,N_16916);
or U17486 (N_17486,N_16862,N_16645);
nand U17487 (N_17487,N_16789,N_16621);
xnor U17488 (N_17488,N_16544,N_16559);
xnor U17489 (N_17489,N_16846,N_16762);
and U17490 (N_17490,N_16832,N_16804);
and U17491 (N_17491,N_16957,N_16809);
or U17492 (N_17492,N_16999,N_16739);
or U17493 (N_17493,N_16681,N_16669);
nor U17494 (N_17494,N_16558,N_16573);
nor U17495 (N_17495,N_16622,N_16998);
xnor U17496 (N_17496,N_16956,N_16851);
and U17497 (N_17497,N_16720,N_16983);
nand U17498 (N_17498,N_16940,N_16793);
xnor U17499 (N_17499,N_16911,N_16559);
and U17500 (N_17500,N_17305,N_17052);
or U17501 (N_17501,N_17449,N_17046);
xnor U17502 (N_17502,N_17341,N_17183);
nor U17503 (N_17503,N_17056,N_17169);
nor U17504 (N_17504,N_17379,N_17243);
and U17505 (N_17505,N_17357,N_17035);
and U17506 (N_17506,N_17293,N_17426);
or U17507 (N_17507,N_17415,N_17176);
nand U17508 (N_17508,N_17041,N_17421);
or U17509 (N_17509,N_17155,N_17478);
xor U17510 (N_17510,N_17318,N_17100);
or U17511 (N_17511,N_17441,N_17322);
or U17512 (N_17512,N_17022,N_17213);
nor U17513 (N_17513,N_17099,N_17185);
or U17514 (N_17514,N_17334,N_17209);
and U17515 (N_17515,N_17181,N_17374);
or U17516 (N_17516,N_17292,N_17034);
nand U17517 (N_17517,N_17417,N_17274);
or U17518 (N_17518,N_17385,N_17028);
nor U17519 (N_17519,N_17167,N_17211);
nand U17520 (N_17520,N_17164,N_17290);
xnor U17521 (N_17521,N_17073,N_17189);
nand U17522 (N_17522,N_17496,N_17342);
nor U17523 (N_17523,N_17231,N_17260);
nor U17524 (N_17524,N_17472,N_17002);
xnor U17525 (N_17525,N_17451,N_17029);
xor U17526 (N_17526,N_17372,N_17266);
nor U17527 (N_17527,N_17406,N_17326);
and U17528 (N_17528,N_17188,N_17126);
nor U17529 (N_17529,N_17066,N_17287);
nor U17530 (N_17530,N_17259,N_17152);
nand U17531 (N_17531,N_17497,N_17068);
and U17532 (N_17532,N_17456,N_17197);
nand U17533 (N_17533,N_17229,N_17377);
nor U17534 (N_17534,N_17013,N_17368);
xnor U17535 (N_17535,N_17378,N_17074);
nand U17536 (N_17536,N_17195,N_17224);
xnor U17537 (N_17537,N_17355,N_17257);
nand U17538 (N_17538,N_17036,N_17284);
and U17539 (N_17539,N_17043,N_17180);
xnor U17540 (N_17540,N_17413,N_17148);
nor U17541 (N_17541,N_17006,N_17475);
and U17542 (N_17542,N_17236,N_17050);
nand U17543 (N_17543,N_17241,N_17348);
or U17544 (N_17544,N_17248,N_17075);
nand U17545 (N_17545,N_17222,N_17303);
nor U17546 (N_17546,N_17463,N_17389);
nand U17547 (N_17547,N_17190,N_17016);
or U17548 (N_17548,N_17218,N_17157);
nand U17549 (N_17549,N_17246,N_17080);
and U17550 (N_17550,N_17216,N_17346);
nand U17551 (N_17551,N_17301,N_17384);
xor U17552 (N_17552,N_17249,N_17156);
nand U17553 (N_17553,N_17051,N_17324);
xnor U17554 (N_17554,N_17380,N_17004);
xnor U17555 (N_17555,N_17261,N_17135);
xnor U17556 (N_17556,N_17174,N_17172);
and U17557 (N_17557,N_17267,N_17273);
nand U17558 (N_17558,N_17098,N_17399);
and U17559 (N_17559,N_17170,N_17161);
and U17560 (N_17560,N_17032,N_17306);
nand U17561 (N_17561,N_17001,N_17452);
nand U17562 (N_17562,N_17239,N_17309);
nand U17563 (N_17563,N_17465,N_17200);
or U17564 (N_17564,N_17280,N_17467);
nand U17565 (N_17565,N_17408,N_17125);
xnor U17566 (N_17566,N_17017,N_17455);
xor U17567 (N_17567,N_17281,N_17479);
xor U17568 (N_17568,N_17210,N_17140);
xor U17569 (N_17569,N_17354,N_17272);
nand U17570 (N_17570,N_17150,N_17228);
nand U17571 (N_17571,N_17336,N_17205);
nand U17572 (N_17572,N_17076,N_17403);
and U17573 (N_17573,N_17038,N_17483);
or U17574 (N_17574,N_17347,N_17042);
nor U17575 (N_17575,N_17420,N_17476);
xor U17576 (N_17576,N_17323,N_17160);
nor U17577 (N_17577,N_17079,N_17250);
xor U17578 (N_17578,N_17162,N_17247);
nand U17579 (N_17579,N_17393,N_17445);
or U17580 (N_17580,N_17095,N_17296);
nand U17581 (N_17581,N_17102,N_17428);
or U17582 (N_17582,N_17337,N_17443);
xor U17583 (N_17583,N_17439,N_17493);
nand U17584 (N_17584,N_17270,N_17430);
nor U17585 (N_17585,N_17492,N_17448);
or U17586 (N_17586,N_17414,N_17008);
nand U17587 (N_17587,N_17119,N_17025);
nor U17588 (N_17588,N_17044,N_17178);
nor U17589 (N_17589,N_17388,N_17071);
xor U17590 (N_17590,N_17136,N_17314);
nand U17591 (N_17591,N_17225,N_17457);
and U17592 (N_17592,N_17431,N_17360);
and U17593 (N_17593,N_17235,N_17412);
or U17594 (N_17594,N_17113,N_17254);
nor U17595 (N_17595,N_17444,N_17325);
nor U17596 (N_17596,N_17376,N_17327);
and U17597 (N_17597,N_17468,N_17143);
nor U17598 (N_17598,N_17486,N_17215);
nor U17599 (N_17599,N_17137,N_17395);
nand U17600 (N_17600,N_17437,N_17319);
and U17601 (N_17601,N_17397,N_17130);
or U17602 (N_17602,N_17107,N_17300);
nor U17603 (N_17603,N_17061,N_17147);
nor U17604 (N_17604,N_17091,N_17485);
xnor U17605 (N_17605,N_17312,N_17089);
nand U17606 (N_17606,N_17227,N_17361);
nand U17607 (N_17607,N_17154,N_17409);
or U17608 (N_17608,N_17067,N_17165);
or U17609 (N_17609,N_17366,N_17432);
xnor U17610 (N_17610,N_17462,N_17026);
or U17611 (N_17611,N_17132,N_17477);
or U17612 (N_17612,N_17277,N_17434);
nand U17613 (N_17613,N_17391,N_17124);
and U17614 (N_17614,N_17392,N_17410);
nor U17615 (N_17615,N_17332,N_17304);
nor U17616 (N_17616,N_17440,N_17382);
or U17617 (N_17617,N_17386,N_17233);
xnor U17618 (N_17618,N_17010,N_17144);
and U17619 (N_17619,N_17003,N_17453);
or U17620 (N_17620,N_17356,N_17111);
xor U17621 (N_17621,N_17122,N_17490);
or U17622 (N_17622,N_17442,N_17031);
nor U17623 (N_17623,N_17398,N_17315);
nor U17624 (N_17624,N_17268,N_17244);
or U17625 (N_17625,N_17184,N_17134);
nand U17626 (N_17626,N_17471,N_17383);
nand U17627 (N_17627,N_17158,N_17092);
nand U17628 (N_17628,N_17110,N_17353);
xnor U17629 (N_17629,N_17207,N_17234);
nor U17630 (N_17630,N_17049,N_17230);
nand U17631 (N_17631,N_17037,N_17271);
nand U17632 (N_17632,N_17129,N_17297);
or U17633 (N_17633,N_17352,N_17242);
or U17634 (N_17634,N_17473,N_17459);
or U17635 (N_17635,N_17310,N_17163);
xnor U17636 (N_17636,N_17394,N_17015);
nor U17637 (N_17637,N_17454,N_17018);
and U17638 (N_17638,N_17105,N_17466);
and U17639 (N_17639,N_17123,N_17367);
nand U17640 (N_17640,N_17220,N_17240);
or U17641 (N_17641,N_17117,N_17116);
nand U17642 (N_17642,N_17065,N_17020);
nor U17643 (N_17643,N_17369,N_17206);
nor U17644 (N_17644,N_17182,N_17402);
or U17645 (N_17645,N_17208,N_17438);
or U17646 (N_17646,N_17151,N_17407);
or U17647 (N_17647,N_17316,N_17464);
or U17648 (N_17648,N_17429,N_17194);
or U17649 (N_17649,N_17064,N_17159);
nand U17650 (N_17650,N_17411,N_17153);
or U17651 (N_17651,N_17494,N_17401);
xor U17652 (N_17652,N_17404,N_17350);
nor U17653 (N_17653,N_17109,N_17217);
or U17654 (N_17654,N_17237,N_17351);
nor U17655 (N_17655,N_17335,N_17416);
or U17656 (N_17656,N_17264,N_17145);
nor U17657 (N_17657,N_17302,N_17498);
and U17658 (N_17658,N_17187,N_17371);
and U17659 (N_17659,N_17470,N_17375);
nand U17660 (N_17660,N_17390,N_17138);
xnor U17661 (N_17661,N_17062,N_17487);
and U17662 (N_17662,N_17364,N_17345);
nor U17663 (N_17663,N_17196,N_17339);
or U17664 (N_17664,N_17232,N_17255);
nand U17665 (N_17665,N_17427,N_17285);
or U17666 (N_17666,N_17000,N_17057);
nor U17667 (N_17667,N_17317,N_17058);
nor U17668 (N_17668,N_17276,N_17328);
and U17669 (N_17669,N_17104,N_17387);
xor U17670 (N_17670,N_17094,N_17023);
and U17671 (N_17671,N_17084,N_17146);
nor U17672 (N_17672,N_17083,N_17482);
nor U17673 (N_17673,N_17495,N_17149);
xnor U17674 (N_17674,N_17005,N_17054);
or U17675 (N_17675,N_17030,N_17373);
and U17676 (N_17676,N_17458,N_17175);
nor U17677 (N_17677,N_17214,N_17333);
nor U17678 (N_17678,N_17115,N_17400);
nor U17679 (N_17679,N_17060,N_17294);
or U17680 (N_17680,N_17489,N_17085);
nand U17681 (N_17681,N_17072,N_17168);
nor U17682 (N_17682,N_17338,N_17418);
and U17683 (N_17683,N_17329,N_17363);
and U17684 (N_17684,N_17423,N_17330);
nand U17685 (N_17685,N_17033,N_17106);
and U17686 (N_17686,N_17245,N_17112);
nand U17687 (N_17687,N_17460,N_17021);
nand U17688 (N_17688,N_17223,N_17045);
xnor U17689 (N_17689,N_17081,N_17212);
xnor U17690 (N_17690,N_17131,N_17425);
and U17691 (N_17691,N_17491,N_17088);
nor U17692 (N_17692,N_17007,N_17253);
nor U17693 (N_17693,N_17278,N_17093);
nor U17694 (N_17694,N_17202,N_17474);
and U17695 (N_17695,N_17047,N_17405);
or U17696 (N_17696,N_17024,N_17450);
xnor U17697 (N_17697,N_17219,N_17291);
xor U17698 (N_17698,N_17127,N_17078);
xor U17699 (N_17699,N_17480,N_17461);
and U17700 (N_17700,N_17433,N_17370);
nor U17701 (N_17701,N_17048,N_17435);
or U17702 (N_17702,N_17108,N_17469);
or U17703 (N_17703,N_17070,N_17258);
nor U17704 (N_17704,N_17142,N_17313);
nand U17705 (N_17705,N_17331,N_17396);
or U17706 (N_17706,N_17308,N_17082);
nand U17707 (N_17707,N_17256,N_17193);
or U17708 (N_17708,N_17289,N_17286);
or U17709 (N_17709,N_17365,N_17359);
or U17710 (N_17710,N_17238,N_17090);
or U17711 (N_17711,N_17499,N_17262);
xnor U17712 (N_17712,N_17320,N_17128);
nand U17713 (N_17713,N_17344,N_17179);
or U17714 (N_17714,N_17436,N_17488);
xnor U17715 (N_17715,N_17204,N_17192);
or U17716 (N_17716,N_17019,N_17481);
or U17717 (N_17717,N_17321,N_17201);
nor U17718 (N_17718,N_17299,N_17171);
nand U17719 (N_17719,N_17251,N_17059);
and U17720 (N_17720,N_17120,N_17141);
xor U17721 (N_17721,N_17226,N_17282);
or U17722 (N_17722,N_17358,N_17027);
xor U17723 (N_17723,N_17419,N_17191);
nand U17724 (N_17724,N_17166,N_17199);
nand U17725 (N_17725,N_17139,N_17307);
and U17726 (N_17726,N_17343,N_17288);
nand U17727 (N_17727,N_17087,N_17096);
and U17728 (N_17728,N_17053,N_17446);
xnor U17729 (N_17729,N_17009,N_17298);
nor U17730 (N_17730,N_17362,N_17040);
and U17731 (N_17731,N_17295,N_17447);
nand U17732 (N_17732,N_17381,N_17311);
nor U17733 (N_17733,N_17263,N_17484);
and U17734 (N_17734,N_17077,N_17340);
or U17735 (N_17735,N_17349,N_17011);
nand U17736 (N_17736,N_17012,N_17069);
or U17737 (N_17737,N_17252,N_17279);
and U17738 (N_17738,N_17177,N_17424);
nand U17739 (N_17739,N_17422,N_17103);
xor U17740 (N_17740,N_17121,N_17221);
xnor U17741 (N_17741,N_17133,N_17198);
and U17742 (N_17742,N_17055,N_17097);
nor U17743 (N_17743,N_17039,N_17063);
or U17744 (N_17744,N_17283,N_17114);
and U17745 (N_17745,N_17203,N_17173);
xor U17746 (N_17746,N_17086,N_17275);
nor U17747 (N_17747,N_17269,N_17101);
xor U17748 (N_17748,N_17118,N_17265);
and U17749 (N_17749,N_17186,N_17014);
xor U17750 (N_17750,N_17039,N_17237);
and U17751 (N_17751,N_17174,N_17063);
nor U17752 (N_17752,N_17307,N_17038);
xor U17753 (N_17753,N_17160,N_17441);
or U17754 (N_17754,N_17291,N_17343);
nand U17755 (N_17755,N_17423,N_17057);
nand U17756 (N_17756,N_17146,N_17007);
xor U17757 (N_17757,N_17066,N_17035);
and U17758 (N_17758,N_17068,N_17308);
nand U17759 (N_17759,N_17301,N_17309);
and U17760 (N_17760,N_17118,N_17340);
nor U17761 (N_17761,N_17109,N_17049);
nand U17762 (N_17762,N_17123,N_17048);
xnor U17763 (N_17763,N_17157,N_17196);
xor U17764 (N_17764,N_17059,N_17230);
xnor U17765 (N_17765,N_17264,N_17469);
nand U17766 (N_17766,N_17228,N_17463);
xor U17767 (N_17767,N_17010,N_17233);
or U17768 (N_17768,N_17314,N_17409);
or U17769 (N_17769,N_17029,N_17408);
or U17770 (N_17770,N_17474,N_17147);
or U17771 (N_17771,N_17204,N_17496);
nand U17772 (N_17772,N_17312,N_17443);
xnor U17773 (N_17773,N_17027,N_17103);
nand U17774 (N_17774,N_17026,N_17388);
and U17775 (N_17775,N_17134,N_17160);
and U17776 (N_17776,N_17315,N_17170);
xnor U17777 (N_17777,N_17207,N_17353);
and U17778 (N_17778,N_17134,N_17431);
or U17779 (N_17779,N_17044,N_17302);
xnor U17780 (N_17780,N_17491,N_17135);
and U17781 (N_17781,N_17069,N_17345);
xnor U17782 (N_17782,N_17441,N_17102);
nand U17783 (N_17783,N_17115,N_17453);
nand U17784 (N_17784,N_17435,N_17050);
and U17785 (N_17785,N_17147,N_17121);
or U17786 (N_17786,N_17102,N_17442);
or U17787 (N_17787,N_17404,N_17434);
xnor U17788 (N_17788,N_17298,N_17284);
or U17789 (N_17789,N_17020,N_17194);
or U17790 (N_17790,N_17153,N_17323);
xor U17791 (N_17791,N_17174,N_17208);
nand U17792 (N_17792,N_17453,N_17093);
xnor U17793 (N_17793,N_17136,N_17446);
or U17794 (N_17794,N_17062,N_17099);
xor U17795 (N_17795,N_17037,N_17177);
nor U17796 (N_17796,N_17245,N_17424);
xor U17797 (N_17797,N_17094,N_17441);
or U17798 (N_17798,N_17409,N_17157);
nand U17799 (N_17799,N_17060,N_17379);
nand U17800 (N_17800,N_17170,N_17347);
and U17801 (N_17801,N_17112,N_17222);
nor U17802 (N_17802,N_17411,N_17072);
or U17803 (N_17803,N_17211,N_17158);
and U17804 (N_17804,N_17162,N_17340);
xor U17805 (N_17805,N_17314,N_17004);
or U17806 (N_17806,N_17266,N_17111);
xor U17807 (N_17807,N_17334,N_17202);
and U17808 (N_17808,N_17093,N_17038);
xor U17809 (N_17809,N_17481,N_17448);
nor U17810 (N_17810,N_17008,N_17424);
xor U17811 (N_17811,N_17491,N_17207);
nand U17812 (N_17812,N_17151,N_17142);
xnor U17813 (N_17813,N_17218,N_17073);
xnor U17814 (N_17814,N_17169,N_17034);
nor U17815 (N_17815,N_17471,N_17361);
nand U17816 (N_17816,N_17357,N_17471);
and U17817 (N_17817,N_17380,N_17120);
xor U17818 (N_17818,N_17315,N_17052);
and U17819 (N_17819,N_17401,N_17481);
xor U17820 (N_17820,N_17234,N_17001);
or U17821 (N_17821,N_17186,N_17071);
and U17822 (N_17822,N_17252,N_17370);
xor U17823 (N_17823,N_17175,N_17133);
nor U17824 (N_17824,N_17069,N_17329);
nor U17825 (N_17825,N_17301,N_17252);
nor U17826 (N_17826,N_17321,N_17074);
xor U17827 (N_17827,N_17275,N_17468);
and U17828 (N_17828,N_17368,N_17089);
or U17829 (N_17829,N_17139,N_17356);
and U17830 (N_17830,N_17335,N_17270);
nor U17831 (N_17831,N_17308,N_17321);
or U17832 (N_17832,N_17062,N_17164);
nand U17833 (N_17833,N_17470,N_17003);
nand U17834 (N_17834,N_17477,N_17362);
nand U17835 (N_17835,N_17050,N_17471);
and U17836 (N_17836,N_17162,N_17478);
or U17837 (N_17837,N_17351,N_17435);
nand U17838 (N_17838,N_17422,N_17202);
and U17839 (N_17839,N_17442,N_17187);
or U17840 (N_17840,N_17209,N_17359);
nor U17841 (N_17841,N_17295,N_17441);
xnor U17842 (N_17842,N_17283,N_17187);
xor U17843 (N_17843,N_17411,N_17467);
or U17844 (N_17844,N_17080,N_17074);
nor U17845 (N_17845,N_17378,N_17109);
xnor U17846 (N_17846,N_17121,N_17352);
and U17847 (N_17847,N_17302,N_17434);
or U17848 (N_17848,N_17333,N_17477);
xor U17849 (N_17849,N_17110,N_17465);
nor U17850 (N_17850,N_17252,N_17183);
and U17851 (N_17851,N_17103,N_17359);
or U17852 (N_17852,N_17431,N_17086);
nor U17853 (N_17853,N_17186,N_17141);
nand U17854 (N_17854,N_17353,N_17127);
nor U17855 (N_17855,N_17443,N_17054);
nand U17856 (N_17856,N_17346,N_17422);
nor U17857 (N_17857,N_17443,N_17128);
or U17858 (N_17858,N_17226,N_17212);
and U17859 (N_17859,N_17434,N_17082);
nor U17860 (N_17860,N_17042,N_17174);
and U17861 (N_17861,N_17131,N_17225);
and U17862 (N_17862,N_17278,N_17273);
and U17863 (N_17863,N_17369,N_17111);
nor U17864 (N_17864,N_17227,N_17450);
nor U17865 (N_17865,N_17125,N_17314);
and U17866 (N_17866,N_17201,N_17027);
nor U17867 (N_17867,N_17182,N_17235);
nand U17868 (N_17868,N_17105,N_17464);
or U17869 (N_17869,N_17247,N_17064);
nor U17870 (N_17870,N_17466,N_17108);
and U17871 (N_17871,N_17459,N_17128);
or U17872 (N_17872,N_17075,N_17388);
and U17873 (N_17873,N_17004,N_17360);
nor U17874 (N_17874,N_17329,N_17499);
and U17875 (N_17875,N_17200,N_17105);
xor U17876 (N_17876,N_17290,N_17027);
or U17877 (N_17877,N_17272,N_17494);
or U17878 (N_17878,N_17398,N_17023);
or U17879 (N_17879,N_17120,N_17156);
nor U17880 (N_17880,N_17153,N_17455);
nor U17881 (N_17881,N_17463,N_17420);
nand U17882 (N_17882,N_17115,N_17452);
xor U17883 (N_17883,N_17162,N_17013);
or U17884 (N_17884,N_17171,N_17413);
nor U17885 (N_17885,N_17471,N_17491);
and U17886 (N_17886,N_17112,N_17020);
or U17887 (N_17887,N_17154,N_17243);
and U17888 (N_17888,N_17373,N_17045);
nand U17889 (N_17889,N_17156,N_17247);
or U17890 (N_17890,N_17247,N_17315);
nand U17891 (N_17891,N_17270,N_17138);
or U17892 (N_17892,N_17167,N_17322);
and U17893 (N_17893,N_17424,N_17175);
xnor U17894 (N_17894,N_17070,N_17404);
nand U17895 (N_17895,N_17428,N_17138);
and U17896 (N_17896,N_17147,N_17002);
nand U17897 (N_17897,N_17330,N_17466);
nand U17898 (N_17898,N_17173,N_17109);
and U17899 (N_17899,N_17154,N_17084);
nand U17900 (N_17900,N_17019,N_17264);
and U17901 (N_17901,N_17435,N_17216);
nand U17902 (N_17902,N_17145,N_17011);
or U17903 (N_17903,N_17064,N_17177);
nor U17904 (N_17904,N_17135,N_17000);
and U17905 (N_17905,N_17494,N_17186);
nor U17906 (N_17906,N_17315,N_17211);
nand U17907 (N_17907,N_17036,N_17471);
xor U17908 (N_17908,N_17163,N_17052);
nor U17909 (N_17909,N_17478,N_17135);
xnor U17910 (N_17910,N_17362,N_17484);
and U17911 (N_17911,N_17077,N_17150);
and U17912 (N_17912,N_17066,N_17099);
nor U17913 (N_17913,N_17052,N_17238);
nor U17914 (N_17914,N_17048,N_17452);
and U17915 (N_17915,N_17233,N_17209);
xnor U17916 (N_17916,N_17499,N_17180);
and U17917 (N_17917,N_17393,N_17187);
xor U17918 (N_17918,N_17246,N_17429);
or U17919 (N_17919,N_17013,N_17063);
nor U17920 (N_17920,N_17228,N_17416);
and U17921 (N_17921,N_17330,N_17251);
nand U17922 (N_17922,N_17092,N_17028);
nor U17923 (N_17923,N_17369,N_17379);
xor U17924 (N_17924,N_17028,N_17474);
or U17925 (N_17925,N_17320,N_17274);
or U17926 (N_17926,N_17305,N_17274);
nand U17927 (N_17927,N_17436,N_17240);
nand U17928 (N_17928,N_17267,N_17459);
nor U17929 (N_17929,N_17415,N_17158);
and U17930 (N_17930,N_17180,N_17387);
xor U17931 (N_17931,N_17090,N_17048);
nand U17932 (N_17932,N_17134,N_17033);
nor U17933 (N_17933,N_17427,N_17486);
nand U17934 (N_17934,N_17057,N_17213);
or U17935 (N_17935,N_17064,N_17153);
and U17936 (N_17936,N_17170,N_17081);
and U17937 (N_17937,N_17016,N_17449);
xnor U17938 (N_17938,N_17463,N_17167);
nand U17939 (N_17939,N_17065,N_17003);
nor U17940 (N_17940,N_17384,N_17027);
or U17941 (N_17941,N_17379,N_17086);
xnor U17942 (N_17942,N_17009,N_17130);
xnor U17943 (N_17943,N_17275,N_17423);
xor U17944 (N_17944,N_17496,N_17304);
nand U17945 (N_17945,N_17307,N_17312);
xor U17946 (N_17946,N_17101,N_17282);
or U17947 (N_17947,N_17236,N_17258);
and U17948 (N_17948,N_17207,N_17005);
nand U17949 (N_17949,N_17437,N_17192);
or U17950 (N_17950,N_17052,N_17416);
xnor U17951 (N_17951,N_17290,N_17237);
and U17952 (N_17952,N_17335,N_17180);
nor U17953 (N_17953,N_17366,N_17270);
xor U17954 (N_17954,N_17476,N_17292);
nand U17955 (N_17955,N_17279,N_17344);
nand U17956 (N_17956,N_17400,N_17210);
nand U17957 (N_17957,N_17076,N_17377);
xnor U17958 (N_17958,N_17204,N_17462);
or U17959 (N_17959,N_17408,N_17139);
nor U17960 (N_17960,N_17380,N_17420);
and U17961 (N_17961,N_17152,N_17065);
or U17962 (N_17962,N_17090,N_17071);
or U17963 (N_17963,N_17412,N_17288);
nand U17964 (N_17964,N_17201,N_17388);
and U17965 (N_17965,N_17077,N_17193);
and U17966 (N_17966,N_17280,N_17099);
and U17967 (N_17967,N_17233,N_17440);
or U17968 (N_17968,N_17275,N_17330);
xnor U17969 (N_17969,N_17158,N_17153);
and U17970 (N_17970,N_17091,N_17435);
or U17971 (N_17971,N_17093,N_17354);
nor U17972 (N_17972,N_17493,N_17056);
xor U17973 (N_17973,N_17146,N_17079);
nor U17974 (N_17974,N_17464,N_17159);
nand U17975 (N_17975,N_17089,N_17233);
nor U17976 (N_17976,N_17261,N_17490);
nor U17977 (N_17977,N_17392,N_17121);
nand U17978 (N_17978,N_17490,N_17367);
nand U17979 (N_17979,N_17341,N_17379);
xnor U17980 (N_17980,N_17307,N_17446);
nand U17981 (N_17981,N_17069,N_17175);
or U17982 (N_17982,N_17275,N_17281);
or U17983 (N_17983,N_17004,N_17199);
and U17984 (N_17984,N_17284,N_17228);
or U17985 (N_17985,N_17092,N_17452);
nand U17986 (N_17986,N_17286,N_17256);
nor U17987 (N_17987,N_17016,N_17436);
nor U17988 (N_17988,N_17024,N_17216);
and U17989 (N_17989,N_17285,N_17224);
nand U17990 (N_17990,N_17250,N_17492);
nor U17991 (N_17991,N_17108,N_17206);
nand U17992 (N_17992,N_17033,N_17320);
or U17993 (N_17993,N_17040,N_17434);
or U17994 (N_17994,N_17134,N_17385);
nor U17995 (N_17995,N_17397,N_17479);
and U17996 (N_17996,N_17139,N_17344);
xnor U17997 (N_17997,N_17235,N_17110);
nor U17998 (N_17998,N_17312,N_17327);
xnor U17999 (N_17999,N_17389,N_17415);
nor U18000 (N_18000,N_17778,N_17540);
and U18001 (N_18001,N_17872,N_17943);
nor U18002 (N_18002,N_17728,N_17622);
xor U18003 (N_18003,N_17779,N_17867);
and U18004 (N_18004,N_17678,N_17987);
nand U18005 (N_18005,N_17534,N_17653);
nor U18006 (N_18006,N_17595,N_17966);
nor U18007 (N_18007,N_17766,N_17915);
xnor U18008 (N_18008,N_17860,N_17865);
or U18009 (N_18009,N_17507,N_17814);
nand U18010 (N_18010,N_17866,N_17536);
nand U18011 (N_18011,N_17942,N_17813);
or U18012 (N_18012,N_17679,N_17510);
xor U18013 (N_18013,N_17952,N_17807);
and U18014 (N_18014,N_17928,N_17722);
or U18015 (N_18015,N_17840,N_17771);
or U18016 (N_18016,N_17881,N_17919);
nand U18017 (N_18017,N_17996,N_17922);
xor U18018 (N_18018,N_17597,N_17879);
nor U18019 (N_18019,N_17926,N_17542);
xor U18020 (N_18020,N_17941,N_17627);
xnor U18021 (N_18021,N_17822,N_17982);
xor U18022 (N_18022,N_17832,N_17786);
xor U18023 (N_18023,N_17702,N_17620);
or U18024 (N_18024,N_17868,N_17890);
xnor U18025 (N_18025,N_17748,N_17632);
nor U18026 (N_18026,N_17703,N_17818);
nand U18027 (N_18027,N_17961,N_17921);
xor U18028 (N_18028,N_17774,N_17810);
and U18029 (N_18029,N_17658,N_17972);
nor U18030 (N_18030,N_17637,N_17916);
xnor U18031 (N_18031,N_17660,N_17856);
nand U18032 (N_18032,N_17859,N_17671);
and U18033 (N_18033,N_17694,N_17553);
or U18034 (N_18034,N_17842,N_17739);
xor U18035 (N_18035,N_17635,N_17517);
and U18036 (N_18036,N_17955,N_17712);
or U18037 (N_18037,N_17654,N_17543);
and U18038 (N_18038,N_17600,N_17614);
and U18039 (N_18039,N_17924,N_17985);
nor U18040 (N_18040,N_17834,N_17648);
xor U18041 (N_18041,N_17572,N_17850);
nand U18042 (N_18042,N_17613,N_17874);
xor U18043 (N_18043,N_17537,N_17788);
nand U18044 (N_18044,N_17724,N_17900);
nand U18045 (N_18045,N_17812,N_17997);
and U18046 (N_18046,N_17773,N_17646);
nand U18047 (N_18047,N_17563,N_17599);
or U18048 (N_18048,N_17845,N_17524);
or U18049 (N_18049,N_17701,N_17768);
nand U18050 (N_18050,N_17615,N_17677);
nor U18051 (N_18051,N_17887,N_17501);
or U18052 (N_18052,N_17947,N_17820);
nor U18053 (N_18053,N_17761,N_17640);
or U18054 (N_18054,N_17516,N_17905);
xnor U18055 (N_18055,N_17970,N_17617);
xnor U18056 (N_18056,N_17690,N_17932);
and U18057 (N_18057,N_17885,N_17755);
xnor U18058 (N_18058,N_17623,N_17806);
or U18059 (N_18059,N_17571,N_17706);
and U18060 (N_18060,N_17621,N_17716);
xor U18061 (N_18061,N_17583,N_17601);
nand U18062 (N_18062,N_17664,N_17847);
nor U18063 (N_18063,N_17741,N_17667);
and U18064 (N_18064,N_17532,N_17995);
and U18065 (N_18065,N_17696,N_17817);
xor U18066 (N_18066,N_17781,N_17695);
nand U18067 (N_18067,N_17562,N_17959);
and U18068 (N_18068,N_17514,N_17732);
nor U18069 (N_18069,N_17522,N_17809);
nor U18070 (N_18070,N_17629,N_17914);
xnor U18071 (N_18071,N_17992,N_17541);
xnor U18072 (N_18072,N_17760,N_17849);
xnor U18073 (N_18073,N_17854,N_17544);
or U18074 (N_18074,N_17642,N_17857);
nor U18075 (N_18075,N_17911,N_17593);
nor U18076 (N_18076,N_17986,N_17631);
or U18077 (N_18077,N_17675,N_17580);
nand U18078 (N_18078,N_17795,N_17962);
nor U18079 (N_18079,N_17945,N_17826);
nor U18080 (N_18080,N_17588,N_17616);
nor U18081 (N_18081,N_17519,N_17670);
nor U18082 (N_18082,N_17692,N_17843);
xor U18083 (N_18083,N_17949,N_17568);
xnor U18084 (N_18084,N_17883,N_17909);
nor U18085 (N_18085,N_17512,N_17937);
xnor U18086 (N_18086,N_17711,N_17977);
and U18087 (N_18087,N_17935,N_17521);
nor U18088 (N_18088,N_17686,N_17533);
nand U18089 (N_18089,N_17668,N_17901);
nand U18090 (N_18090,N_17983,N_17683);
or U18091 (N_18091,N_17659,N_17780);
and U18092 (N_18092,N_17802,N_17956);
or U18093 (N_18093,N_17567,N_17720);
xor U18094 (N_18094,N_17772,N_17697);
nor U18095 (N_18095,N_17518,N_17609);
nor U18096 (N_18096,N_17757,N_17882);
or U18097 (N_18097,N_17550,N_17875);
nor U18098 (N_18098,N_17902,N_17746);
xnor U18099 (N_18099,N_17950,N_17792);
xnor U18100 (N_18100,N_17828,N_17651);
xnor U18101 (N_18101,N_17994,N_17946);
or U18102 (N_18102,N_17893,N_17699);
or U18103 (N_18103,N_17889,N_17661);
and U18104 (N_18104,N_17500,N_17693);
nor U18105 (N_18105,N_17734,N_17633);
xnor U18106 (N_18106,N_17839,N_17819);
and U18107 (N_18107,N_17573,N_17698);
nor U18108 (N_18108,N_17687,N_17569);
nor U18109 (N_18109,N_17624,N_17570);
nand U18110 (N_18110,N_17823,N_17731);
and U18111 (N_18111,N_17899,N_17884);
or U18112 (N_18112,N_17581,N_17608);
and U18113 (N_18113,N_17863,N_17681);
xnor U18114 (N_18114,N_17709,N_17841);
and U18115 (N_18115,N_17531,N_17846);
nand U18116 (N_18116,N_17509,N_17689);
and U18117 (N_18117,N_17894,N_17829);
xnor U18118 (N_18118,N_17577,N_17645);
xnor U18119 (N_18119,N_17896,N_17762);
nor U18120 (N_18120,N_17564,N_17933);
or U18121 (N_18121,N_17920,N_17628);
or U18122 (N_18122,N_17643,N_17736);
xor U18123 (N_18123,N_17805,N_17951);
and U18124 (N_18124,N_17862,N_17619);
or U18125 (N_18125,N_17576,N_17979);
xor U18126 (N_18126,N_17864,N_17725);
and U18127 (N_18127,N_17506,N_17684);
or U18128 (N_18128,N_17747,N_17527);
or U18129 (N_18129,N_17816,N_17906);
or U18130 (N_18130,N_17682,N_17944);
nand U18131 (N_18131,N_17723,N_17844);
nor U18132 (N_18132,N_17777,N_17871);
and U18133 (N_18133,N_17783,N_17662);
nor U18134 (N_18134,N_17708,N_17851);
nand U18135 (N_18135,N_17606,N_17821);
xnor U18136 (N_18136,N_17878,N_17790);
nand U18137 (N_18137,N_17713,N_17930);
or U18138 (N_18138,N_17877,N_17674);
nor U18139 (N_18139,N_17796,N_17744);
or U18140 (N_18140,N_17538,N_17803);
and U18141 (N_18141,N_17529,N_17759);
and U18142 (N_18142,N_17511,N_17891);
nand U18143 (N_18143,N_17910,N_17742);
or U18144 (N_18144,N_17785,N_17825);
or U18145 (N_18145,N_17912,N_17974);
xnor U18146 (N_18146,N_17547,N_17650);
xnor U18147 (N_18147,N_17753,N_17958);
or U18148 (N_18148,N_17784,N_17688);
xor U18149 (N_18149,N_17663,N_17641);
nand U18150 (N_18150,N_17673,N_17980);
xnor U18151 (N_18151,N_17908,N_17749);
nand U18152 (N_18152,N_17726,N_17833);
and U18153 (N_18153,N_17556,N_17848);
nor U18154 (N_18154,N_17978,N_17528);
nand U18155 (N_18155,N_17793,N_17764);
and U18156 (N_18156,N_17903,N_17858);
xnor U18157 (N_18157,N_17590,N_17665);
nand U18158 (N_18158,N_17680,N_17605);
and U18159 (N_18159,N_17552,N_17936);
and U18160 (N_18160,N_17656,N_17676);
nand U18161 (N_18161,N_17582,N_17776);
or U18162 (N_18162,N_17791,N_17503);
xnor U18163 (N_18163,N_17603,N_17561);
nor U18164 (N_18164,N_17895,N_17575);
and U18165 (N_18165,N_17523,N_17602);
and U18166 (N_18166,N_17775,N_17797);
nand U18167 (N_18167,N_17535,N_17504);
xnor U18168 (N_18168,N_17756,N_17586);
and U18169 (N_18169,N_17923,N_17960);
nor U18170 (N_18170,N_17855,N_17707);
nand U18171 (N_18171,N_17546,N_17515);
nor U18172 (N_18172,N_17824,N_17957);
and U18173 (N_18173,N_17876,N_17918);
xor U18174 (N_18174,N_17559,N_17618);
nand U18175 (N_18175,N_17591,N_17968);
and U18176 (N_18176,N_17880,N_17636);
nor U18177 (N_18177,N_17525,N_17827);
and U18178 (N_18178,N_17520,N_17666);
xnor U18179 (N_18179,N_17811,N_17897);
nand U18180 (N_18180,N_17799,N_17963);
or U18181 (N_18181,N_17738,N_17969);
and U18182 (N_18182,N_17578,N_17815);
nand U18183 (N_18183,N_17989,N_17929);
and U18184 (N_18184,N_17873,N_17794);
and U18185 (N_18185,N_17769,N_17740);
xnor U18186 (N_18186,N_17967,N_17513);
nor U18187 (N_18187,N_17630,N_17938);
and U18188 (N_18188,N_17727,N_17730);
xor U18189 (N_18189,N_17735,N_17888);
xnor U18190 (N_18190,N_17870,N_17508);
nand U18191 (N_18191,N_17718,N_17612);
nand U18192 (N_18192,N_17971,N_17652);
and U18193 (N_18193,N_17789,N_17754);
or U18194 (N_18194,N_17587,N_17988);
and U18195 (N_18195,N_17558,N_17729);
xor U18196 (N_18196,N_17505,N_17752);
and U18197 (N_18197,N_17981,N_17604);
xor U18198 (N_18198,N_17639,N_17964);
nand U18199 (N_18199,N_17931,N_17917);
and U18200 (N_18200,N_17714,N_17808);
xor U18201 (N_18201,N_17904,N_17589);
nor U18202 (N_18202,N_17991,N_17763);
nand U18203 (N_18203,N_17626,N_17649);
and U18204 (N_18204,N_17999,N_17526);
and U18205 (N_18205,N_17973,N_17838);
and U18206 (N_18206,N_17548,N_17555);
nand U18207 (N_18207,N_17554,N_17551);
nor U18208 (N_18208,N_17976,N_17767);
and U18209 (N_18209,N_17717,N_17737);
nand U18210 (N_18210,N_17557,N_17565);
nand U18211 (N_18211,N_17831,N_17719);
xor U18212 (N_18212,N_17710,N_17998);
or U18213 (N_18213,N_17948,N_17672);
xor U18214 (N_18214,N_17657,N_17704);
and U18215 (N_18215,N_17954,N_17644);
xnor U18216 (N_18216,N_17907,N_17560);
nor U18217 (N_18217,N_17853,N_17852);
xnor U18218 (N_18218,N_17733,N_17939);
xor U18219 (N_18219,N_17610,N_17993);
nor U18220 (N_18220,N_17647,N_17940);
xnor U18221 (N_18221,N_17700,N_17715);
and U18222 (N_18222,N_17743,N_17549);
nor U18223 (N_18223,N_17685,N_17721);
nor U18224 (N_18224,N_17835,N_17965);
xor U18225 (N_18225,N_17782,N_17886);
or U18226 (N_18226,N_17990,N_17953);
nor U18227 (N_18227,N_17861,N_17545);
or U18228 (N_18228,N_17830,N_17638);
nor U18229 (N_18229,N_17745,N_17634);
xor U18230 (N_18230,N_17579,N_17607);
xnor U18231 (N_18231,N_17655,N_17758);
or U18232 (N_18232,N_17598,N_17898);
nand U18233 (N_18233,N_17800,N_17691);
or U18234 (N_18234,N_17502,N_17801);
nor U18235 (N_18235,N_17770,N_17574);
nor U18236 (N_18236,N_17596,N_17625);
nor U18237 (N_18237,N_17705,N_17611);
or U18238 (N_18238,N_17669,N_17585);
or U18239 (N_18239,N_17934,N_17892);
nor U18240 (N_18240,N_17927,N_17566);
nand U18241 (N_18241,N_17539,N_17787);
or U18242 (N_18242,N_17975,N_17584);
nand U18243 (N_18243,N_17869,N_17750);
nand U18244 (N_18244,N_17594,N_17925);
and U18245 (N_18245,N_17913,N_17530);
nor U18246 (N_18246,N_17837,N_17765);
nand U18247 (N_18247,N_17804,N_17836);
nand U18248 (N_18248,N_17798,N_17984);
nand U18249 (N_18249,N_17592,N_17751);
nor U18250 (N_18250,N_17679,N_17952);
and U18251 (N_18251,N_17919,N_17799);
nand U18252 (N_18252,N_17987,N_17897);
xor U18253 (N_18253,N_17653,N_17748);
nand U18254 (N_18254,N_17599,N_17742);
nor U18255 (N_18255,N_17612,N_17512);
nand U18256 (N_18256,N_17507,N_17981);
nor U18257 (N_18257,N_17992,N_17792);
nand U18258 (N_18258,N_17532,N_17692);
nor U18259 (N_18259,N_17601,N_17892);
and U18260 (N_18260,N_17978,N_17836);
nor U18261 (N_18261,N_17546,N_17766);
and U18262 (N_18262,N_17583,N_17799);
nor U18263 (N_18263,N_17575,N_17736);
nor U18264 (N_18264,N_17986,N_17998);
nand U18265 (N_18265,N_17726,N_17639);
and U18266 (N_18266,N_17940,N_17692);
and U18267 (N_18267,N_17571,N_17924);
nor U18268 (N_18268,N_17606,N_17970);
xnor U18269 (N_18269,N_17798,N_17509);
nand U18270 (N_18270,N_17971,N_17983);
xor U18271 (N_18271,N_17518,N_17658);
and U18272 (N_18272,N_17795,N_17932);
and U18273 (N_18273,N_17955,N_17951);
nor U18274 (N_18274,N_17903,N_17515);
and U18275 (N_18275,N_17683,N_17897);
and U18276 (N_18276,N_17784,N_17892);
or U18277 (N_18277,N_17576,N_17684);
nand U18278 (N_18278,N_17904,N_17905);
xnor U18279 (N_18279,N_17992,N_17899);
nor U18280 (N_18280,N_17788,N_17765);
xor U18281 (N_18281,N_17641,N_17785);
xor U18282 (N_18282,N_17914,N_17983);
nor U18283 (N_18283,N_17861,N_17843);
nand U18284 (N_18284,N_17942,N_17642);
nand U18285 (N_18285,N_17742,N_17779);
xor U18286 (N_18286,N_17983,N_17734);
xnor U18287 (N_18287,N_17826,N_17724);
or U18288 (N_18288,N_17806,N_17931);
or U18289 (N_18289,N_17734,N_17657);
nand U18290 (N_18290,N_17955,N_17730);
or U18291 (N_18291,N_17749,N_17594);
or U18292 (N_18292,N_17637,N_17893);
nor U18293 (N_18293,N_17722,N_17530);
or U18294 (N_18294,N_17913,N_17583);
xor U18295 (N_18295,N_17724,N_17756);
nor U18296 (N_18296,N_17753,N_17964);
xor U18297 (N_18297,N_17778,N_17564);
xor U18298 (N_18298,N_17971,N_17623);
xnor U18299 (N_18299,N_17503,N_17845);
xor U18300 (N_18300,N_17689,N_17965);
xnor U18301 (N_18301,N_17846,N_17864);
xnor U18302 (N_18302,N_17689,N_17989);
and U18303 (N_18303,N_17703,N_17982);
nand U18304 (N_18304,N_17864,N_17666);
nor U18305 (N_18305,N_17712,N_17817);
nand U18306 (N_18306,N_17973,N_17979);
nand U18307 (N_18307,N_17610,N_17758);
nand U18308 (N_18308,N_17526,N_17514);
xnor U18309 (N_18309,N_17904,N_17630);
xnor U18310 (N_18310,N_17965,N_17913);
nor U18311 (N_18311,N_17962,N_17642);
nand U18312 (N_18312,N_17887,N_17942);
and U18313 (N_18313,N_17546,N_17580);
xor U18314 (N_18314,N_17695,N_17804);
and U18315 (N_18315,N_17608,N_17504);
or U18316 (N_18316,N_17655,N_17533);
and U18317 (N_18317,N_17587,N_17828);
or U18318 (N_18318,N_17975,N_17544);
nor U18319 (N_18319,N_17929,N_17855);
xnor U18320 (N_18320,N_17997,N_17752);
or U18321 (N_18321,N_17553,N_17806);
or U18322 (N_18322,N_17916,N_17650);
nand U18323 (N_18323,N_17641,N_17528);
xor U18324 (N_18324,N_17646,N_17577);
xnor U18325 (N_18325,N_17669,N_17985);
nor U18326 (N_18326,N_17588,N_17678);
or U18327 (N_18327,N_17607,N_17726);
or U18328 (N_18328,N_17821,N_17890);
and U18329 (N_18329,N_17636,N_17945);
and U18330 (N_18330,N_17643,N_17894);
xor U18331 (N_18331,N_17689,N_17854);
xnor U18332 (N_18332,N_17774,N_17675);
nand U18333 (N_18333,N_17612,N_17586);
or U18334 (N_18334,N_17623,N_17603);
nand U18335 (N_18335,N_17581,N_17981);
nand U18336 (N_18336,N_17689,N_17645);
or U18337 (N_18337,N_17907,N_17795);
xor U18338 (N_18338,N_17846,N_17905);
and U18339 (N_18339,N_17740,N_17647);
xnor U18340 (N_18340,N_17636,N_17576);
nand U18341 (N_18341,N_17829,N_17972);
nor U18342 (N_18342,N_17551,N_17866);
or U18343 (N_18343,N_17827,N_17501);
and U18344 (N_18344,N_17964,N_17642);
xor U18345 (N_18345,N_17753,N_17901);
nor U18346 (N_18346,N_17800,N_17923);
xnor U18347 (N_18347,N_17579,N_17838);
or U18348 (N_18348,N_17628,N_17980);
nand U18349 (N_18349,N_17795,N_17596);
and U18350 (N_18350,N_17649,N_17803);
nor U18351 (N_18351,N_17698,N_17816);
nor U18352 (N_18352,N_17720,N_17633);
and U18353 (N_18353,N_17738,N_17728);
xnor U18354 (N_18354,N_17848,N_17855);
nand U18355 (N_18355,N_17705,N_17691);
and U18356 (N_18356,N_17801,N_17752);
xor U18357 (N_18357,N_17710,N_17723);
nand U18358 (N_18358,N_17752,N_17950);
and U18359 (N_18359,N_17775,N_17983);
xor U18360 (N_18360,N_17628,N_17543);
nor U18361 (N_18361,N_17902,N_17611);
or U18362 (N_18362,N_17516,N_17894);
xor U18363 (N_18363,N_17573,N_17891);
or U18364 (N_18364,N_17796,N_17973);
nor U18365 (N_18365,N_17782,N_17931);
and U18366 (N_18366,N_17676,N_17867);
or U18367 (N_18367,N_17764,N_17548);
xnor U18368 (N_18368,N_17916,N_17517);
or U18369 (N_18369,N_17812,N_17501);
or U18370 (N_18370,N_17954,N_17532);
or U18371 (N_18371,N_17816,N_17833);
or U18372 (N_18372,N_17533,N_17711);
or U18373 (N_18373,N_17960,N_17652);
nor U18374 (N_18374,N_17958,N_17550);
nor U18375 (N_18375,N_17521,N_17561);
or U18376 (N_18376,N_17779,N_17631);
or U18377 (N_18377,N_17638,N_17866);
or U18378 (N_18378,N_17646,N_17979);
and U18379 (N_18379,N_17660,N_17570);
xor U18380 (N_18380,N_17723,N_17801);
nor U18381 (N_18381,N_17923,N_17994);
nor U18382 (N_18382,N_17786,N_17948);
nor U18383 (N_18383,N_17585,N_17647);
or U18384 (N_18384,N_17997,N_17796);
nand U18385 (N_18385,N_17616,N_17644);
nor U18386 (N_18386,N_17666,N_17930);
xnor U18387 (N_18387,N_17771,N_17548);
nand U18388 (N_18388,N_17728,N_17548);
nand U18389 (N_18389,N_17678,N_17547);
and U18390 (N_18390,N_17621,N_17637);
nand U18391 (N_18391,N_17997,N_17776);
xnor U18392 (N_18392,N_17758,N_17741);
nand U18393 (N_18393,N_17934,N_17672);
and U18394 (N_18394,N_17873,N_17972);
and U18395 (N_18395,N_17736,N_17928);
or U18396 (N_18396,N_17813,N_17889);
nor U18397 (N_18397,N_17967,N_17510);
nand U18398 (N_18398,N_17538,N_17759);
or U18399 (N_18399,N_17735,N_17593);
and U18400 (N_18400,N_17823,N_17686);
nor U18401 (N_18401,N_17697,N_17928);
nor U18402 (N_18402,N_17683,N_17759);
xor U18403 (N_18403,N_17576,N_17873);
xor U18404 (N_18404,N_17821,N_17954);
nand U18405 (N_18405,N_17891,N_17897);
xor U18406 (N_18406,N_17677,N_17602);
nand U18407 (N_18407,N_17904,N_17620);
nand U18408 (N_18408,N_17715,N_17716);
xnor U18409 (N_18409,N_17746,N_17677);
nor U18410 (N_18410,N_17807,N_17765);
or U18411 (N_18411,N_17979,N_17565);
xnor U18412 (N_18412,N_17983,N_17876);
xnor U18413 (N_18413,N_17691,N_17572);
nand U18414 (N_18414,N_17552,N_17755);
and U18415 (N_18415,N_17566,N_17812);
or U18416 (N_18416,N_17704,N_17552);
and U18417 (N_18417,N_17733,N_17774);
xor U18418 (N_18418,N_17820,N_17725);
nand U18419 (N_18419,N_17906,N_17701);
xnor U18420 (N_18420,N_17558,N_17819);
nor U18421 (N_18421,N_17768,N_17950);
or U18422 (N_18422,N_17875,N_17603);
and U18423 (N_18423,N_17777,N_17970);
xnor U18424 (N_18424,N_17694,N_17504);
nand U18425 (N_18425,N_17725,N_17736);
nand U18426 (N_18426,N_17578,N_17924);
xor U18427 (N_18427,N_17642,N_17752);
nor U18428 (N_18428,N_17797,N_17976);
and U18429 (N_18429,N_17857,N_17803);
or U18430 (N_18430,N_17853,N_17930);
or U18431 (N_18431,N_17784,N_17717);
nand U18432 (N_18432,N_17945,N_17785);
nand U18433 (N_18433,N_17626,N_17742);
or U18434 (N_18434,N_17556,N_17797);
or U18435 (N_18435,N_17925,N_17775);
xnor U18436 (N_18436,N_17784,N_17634);
nor U18437 (N_18437,N_17826,N_17877);
nor U18438 (N_18438,N_17921,N_17927);
nor U18439 (N_18439,N_17643,N_17987);
xnor U18440 (N_18440,N_17660,N_17974);
nand U18441 (N_18441,N_17939,N_17958);
and U18442 (N_18442,N_17806,N_17747);
nand U18443 (N_18443,N_17905,N_17548);
or U18444 (N_18444,N_17628,N_17684);
nor U18445 (N_18445,N_17782,N_17951);
xor U18446 (N_18446,N_17870,N_17881);
and U18447 (N_18447,N_17788,N_17879);
and U18448 (N_18448,N_17575,N_17844);
xor U18449 (N_18449,N_17996,N_17693);
nand U18450 (N_18450,N_17645,N_17858);
nor U18451 (N_18451,N_17660,N_17757);
and U18452 (N_18452,N_17538,N_17598);
xor U18453 (N_18453,N_17848,N_17594);
xor U18454 (N_18454,N_17580,N_17844);
nand U18455 (N_18455,N_17550,N_17541);
nor U18456 (N_18456,N_17896,N_17617);
nor U18457 (N_18457,N_17945,N_17976);
nor U18458 (N_18458,N_17886,N_17928);
nor U18459 (N_18459,N_17890,N_17776);
xor U18460 (N_18460,N_17943,N_17751);
nand U18461 (N_18461,N_17803,N_17541);
and U18462 (N_18462,N_17572,N_17891);
xor U18463 (N_18463,N_17584,N_17516);
or U18464 (N_18464,N_17704,N_17990);
xnor U18465 (N_18465,N_17839,N_17674);
and U18466 (N_18466,N_17548,N_17511);
xor U18467 (N_18467,N_17591,N_17751);
xnor U18468 (N_18468,N_17917,N_17592);
nand U18469 (N_18469,N_17915,N_17898);
and U18470 (N_18470,N_17856,N_17553);
nor U18471 (N_18471,N_17607,N_17915);
or U18472 (N_18472,N_17858,N_17574);
or U18473 (N_18473,N_17891,N_17752);
or U18474 (N_18474,N_17543,N_17982);
and U18475 (N_18475,N_17990,N_17797);
and U18476 (N_18476,N_17625,N_17699);
or U18477 (N_18477,N_17692,N_17881);
or U18478 (N_18478,N_17819,N_17620);
xor U18479 (N_18479,N_17744,N_17758);
nand U18480 (N_18480,N_17516,N_17790);
nor U18481 (N_18481,N_17660,N_17518);
nor U18482 (N_18482,N_17792,N_17563);
xor U18483 (N_18483,N_17802,N_17795);
nand U18484 (N_18484,N_17834,N_17532);
or U18485 (N_18485,N_17618,N_17625);
or U18486 (N_18486,N_17608,N_17578);
xor U18487 (N_18487,N_17674,N_17944);
nor U18488 (N_18488,N_17968,N_17846);
nand U18489 (N_18489,N_17705,N_17844);
or U18490 (N_18490,N_17704,N_17738);
nor U18491 (N_18491,N_17708,N_17538);
xor U18492 (N_18492,N_17910,N_17736);
or U18493 (N_18493,N_17617,N_17612);
nor U18494 (N_18494,N_17705,N_17840);
and U18495 (N_18495,N_17532,N_17958);
nand U18496 (N_18496,N_17586,N_17632);
nor U18497 (N_18497,N_17962,N_17720);
xor U18498 (N_18498,N_17553,N_17911);
nand U18499 (N_18499,N_17650,N_17761);
xor U18500 (N_18500,N_18163,N_18369);
nand U18501 (N_18501,N_18094,N_18437);
xnor U18502 (N_18502,N_18071,N_18418);
nand U18503 (N_18503,N_18151,N_18357);
nand U18504 (N_18504,N_18431,N_18183);
or U18505 (N_18505,N_18073,N_18347);
nor U18506 (N_18506,N_18080,N_18399);
xor U18507 (N_18507,N_18489,N_18336);
nor U18508 (N_18508,N_18350,N_18309);
nor U18509 (N_18509,N_18424,N_18259);
nand U18510 (N_18510,N_18435,N_18119);
xor U18511 (N_18511,N_18129,N_18430);
and U18512 (N_18512,N_18219,N_18199);
nor U18513 (N_18513,N_18333,N_18480);
and U18514 (N_18514,N_18009,N_18019);
or U18515 (N_18515,N_18149,N_18014);
xnor U18516 (N_18516,N_18257,N_18345);
nor U18517 (N_18517,N_18474,N_18058);
and U18518 (N_18518,N_18290,N_18069);
nor U18519 (N_18519,N_18239,N_18203);
xnor U18520 (N_18520,N_18220,N_18132);
or U18521 (N_18521,N_18067,N_18024);
and U18522 (N_18522,N_18479,N_18329);
nand U18523 (N_18523,N_18439,N_18248);
xnor U18524 (N_18524,N_18256,N_18332);
nand U18525 (N_18525,N_18314,N_18361);
nand U18526 (N_18526,N_18134,N_18478);
nand U18527 (N_18527,N_18408,N_18005);
xnor U18528 (N_18528,N_18318,N_18485);
nor U18529 (N_18529,N_18139,N_18288);
xnor U18530 (N_18530,N_18008,N_18270);
and U18531 (N_18531,N_18242,N_18082);
and U18532 (N_18532,N_18040,N_18292);
nand U18533 (N_18533,N_18227,N_18059);
nor U18534 (N_18534,N_18229,N_18156);
nor U18535 (N_18535,N_18091,N_18170);
or U18536 (N_18536,N_18048,N_18160);
nor U18537 (N_18537,N_18216,N_18483);
xnor U18538 (N_18538,N_18407,N_18057);
xnor U18539 (N_18539,N_18497,N_18204);
and U18540 (N_18540,N_18244,N_18412);
or U18541 (N_18541,N_18240,N_18364);
nor U18542 (N_18542,N_18167,N_18371);
and U18543 (N_18543,N_18453,N_18362);
nor U18544 (N_18544,N_18377,N_18344);
and U18545 (N_18545,N_18238,N_18291);
and U18546 (N_18546,N_18271,N_18026);
or U18547 (N_18547,N_18277,N_18098);
nor U18548 (N_18548,N_18002,N_18223);
nor U18549 (N_18549,N_18015,N_18092);
or U18550 (N_18550,N_18150,N_18342);
nor U18551 (N_18551,N_18102,N_18245);
xnor U18552 (N_18552,N_18034,N_18116);
or U18553 (N_18553,N_18299,N_18231);
nor U18554 (N_18554,N_18384,N_18317);
nand U18555 (N_18555,N_18293,N_18012);
or U18556 (N_18556,N_18427,N_18442);
xnor U18557 (N_18557,N_18189,N_18035);
or U18558 (N_18558,N_18233,N_18348);
nand U18559 (N_18559,N_18236,N_18081);
xnor U18560 (N_18560,N_18454,N_18246);
nor U18561 (N_18561,N_18051,N_18083);
and U18562 (N_18562,N_18054,N_18247);
xnor U18563 (N_18563,N_18452,N_18396);
nor U18564 (N_18564,N_18389,N_18436);
nor U18565 (N_18565,N_18066,N_18494);
nor U18566 (N_18566,N_18086,N_18370);
and U18567 (N_18567,N_18016,N_18037);
xor U18568 (N_18568,N_18117,N_18459);
nor U18569 (N_18569,N_18473,N_18481);
xnor U18570 (N_18570,N_18420,N_18255);
or U18571 (N_18571,N_18367,N_18027);
nor U18572 (N_18572,N_18072,N_18105);
and U18573 (N_18573,N_18045,N_18328);
nor U18574 (N_18574,N_18295,N_18187);
nor U18575 (N_18575,N_18038,N_18079);
and U18576 (N_18576,N_18077,N_18155);
nor U18577 (N_18577,N_18202,N_18488);
and U18578 (N_18578,N_18148,N_18060);
nor U18579 (N_18579,N_18487,N_18410);
nor U18580 (N_18580,N_18153,N_18477);
or U18581 (N_18581,N_18089,N_18375);
xor U18582 (N_18582,N_18267,N_18433);
xnor U18583 (N_18583,N_18432,N_18177);
and U18584 (N_18584,N_18450,N_18282);
nor U18585 (N_18585,N_18266,N_18421);
and U18586 (N_18586,N_18275,N_18272);
nor U18587 (N_18587,N_18097,N_18251);
xnor U18588 (N_18588,N_18394,N_18111);
nor U18589 (N_18589,N_18249,N_18196);
nand U18590 (N_18590,N_18208,N_18122);
and U18591 (N_18591,N_18075,N_18010);
xnor U18592 (N_18592,N_18104,N_18032);
and U18593 (N_18593,N_18491,N_18327);
and U18594 (N_18594,N_18268,N_18180);
nor U18595 (N_18595,N_18360,N_18402);
xnor U18596 (N_18596,N_18315,N_18209);
xnor U18597 (N_18597,N_18434,N_18230);
nor U18598 (N_18598,N_18106,N_18182);
nor U18599 (N_18599,N_18064,N_18398);
xor U18600 (N_18600,N_18237,N_18354);
nor U18601 (N_18601,N_18062,N_18212);
and U18602 (N_18602,N_18368,N_18162);
nand U18603 (N_18603,N_18294,N_18004);
and U18604 (N_18604,N_18222,N_18286);
or U18605 (N_18605,N_18326,N_18274);
and U18606 (N_18606,N_18197,N_18118);
nor U18607 (N_18607,N_18235,N_18319);
and U18608 (N_18608,N_18047,N_18356);
nand U18609 (N_18609,N_18184,N_18385);
xor U18610 (N_18610,N_18260,N_18449);
and U18611 (N_18611,N_18093,N_18387);
xor U18612 (N_18612,N_18090,N_18164);
nand U18613 (N_18613,N_18337,N_18076);
and U18614 (N_18614,N_18046,N_18021);
xor U18615 (N_18615,N_18269,N_18099);
nand U18616 (N_18616,N_18313,N_18128);
xnor U18617 (N_18617,N_18417,N_18096);
xnor U18618 (N_18618,N_18391,N_18095);
xnor U18619 (N_18619,N_18401,N_18320);
and U18620 (N_18620,N_18440,N_18353);
xnor U18621 (N_18621,N_18300,N_18100);
or U18622 (N_18622,N_18341,N_18158);
and U18623 (N_18623,N_18154,N_18419);
and U18624 (N_18624,N_18425,N_18176);
xor U18625 (N_18625,N_18108,N_18492);
and U18626 (N_18626,N_18469,N_18053);
nand U18627 (N_18627,N_18415,N_18446);
nor U18628 (N_18628,N_18381,N_18355);
or U18629 (N_18629,N_18261,N_18224);
and U18630 (N_18630,N_18006,N_18388);
and U18631 (N_18631,N_18486,N_18476);
nand U18632 (N_18632,N_18438,N_18133);
xor U18633 (N_18633,N_18030,N_18284);
nand U18634 (N_18634,N_18358,N_18495);
xor U18635 (N_18635,N_18413,N_18068);
nor U18636 (N_18636,N_18173,N_18186);
nor U18637 (N_18637,N_18428,N_18470);
or U18638 (N_18638,N_18346,N_18039);
xor U18639 (N_18639,N_18339,N_18141);
or U18640 (N_18640,N_18215,N_18289);
or U18641 (N_18641,N_18144,N_18441);
nor U18642 (N_18642,N_18120,N_18498);
or U18643 (N_18643,N_18316,N_18340);
and U18644 (N_18644,N_18201,N_18429);
or U18645 (N_18645,N_18262,N_18475);
xor U18646 (N_18646,N_18192,N_18382);
or U18647 (N_18647,N_18351,N_18403);
nor U18648 (N_18648,N_18137,N_18018);
or U18649 (N_18649,N_18025,N_18043);
or U18650 (N_18650,N_18458,N_18028);
nor U18651 (N_18651,N_18135,N_18422);
xnor U18652 (N_18652,N_18308,N_18188);
nand U18653 (N_18653,N_18022,N_18264);
nor U18654 (N_18654,N_18460,N_18378);
xor U18655 (N_18655,N_18392,N_18365);
or U18656 (N_18656,N_18221,N_18185);
or U18657 (N_18657,N_18101,N_18124);
and U18658 (N_18658,N_18088,N_18338);
nand U18659 (N_18659,N_18457,N_18456);
nand U18660 (N_18660,N_18296,N_18250);
and U18661 (N_18661,N_18307,N_18065);
nand U18662 (N_18662,N_18056,N_18029);
xnor U18663 (N_18663,N_18049,N_18213);
and U18664 (N_18664,N_18297,N_18363);
xor U18665 (N_18665,N_18322,N_18330);
nand U18666 (N_18666,N_18178,N_18145);
nor U18667 (N_18667,N_18131,N_18190);
nor U18668 (N_18668,N_18279,N_18390);
and U18669 (N_18669,N_18252,N_18405);
xnor U18670 (N_18670,N_18114,N_18397);
or U18671 (N_18671,N_18455,N_18234);
nand U18672 (N_18672,N_18138,N_18359);
nand U18673 (N_18673,N_18301,N_18445);
xnor U18674 (N_18674,N_18146,N_18409);
nor U18675 (N_18675,N_18020,N_18303);
nor U18676 (N_18676,N_18383,N_18334);
nor U18677 (N_18677,N_18263,N_18042);
or U18678 (N_18678,N_18311,N_18136);
nor U18679 (N_18679,N_18325,N_18463);
or U18680 (N_18680,N_18205,N_18011);
or U18681 (N_18681,N_18130,N_18200);
or U18682 (N_18682,N_18107,N_18447);
nand U18683 (N_18683,N_18499,N_18052);
and U18684 (N_18684,N_18254,N_18193);
nor U18685 (N_18685,N_18312,N_18305);
or U18686 (N_18686,N_18044,N_18142);
nand U18687 (N_18687,N_18411,N_18207);
and U18688 (N_18688,N_18226,N_18243);
and U18689 (N_18689,N_18461,N_18493);
xnor U18690 (N_18690,N_18147,N_18000);
xor U18691 (N_18691,N_18007,N_18464);
or U18692 (N_18692,N_18276,N_18017);
and U18693 (N_18693,N_18416,N_18281);
nand U18694 (N_18694,N_18084,N_18121);
or U18695 (N_18695,N_18165,N_18406);
xnor U18696 (N_18696,N_18050,N_18331);
and U18697 (N_18697,N_18143,N_18087);
nand U18698 (N_18698,N_18125,N_18241);
or U18699 (N_18699,N_18055,N_18191);
and U18700 (N_18700,N_18126,N_18112);
and U18701 (N_18701,N_18298,N_18306);
nor U18702 (N_18702,N_18172,N_18159);
xnor U18703 (N_18703,N_18157,N_18304);
nor U18704 (N_18704,N_18490,N_18161);
and U18705 (N_18705,N_18414,N_18324);
and U18706 (N_18706,N_18217,N_18280);
xnor U18707 (N_18707,N_18287,N_18444);
xnor U18708 (N_18708,N_18343,N_18013);
or U18709 (N_18709,N_18194,N_18206);
nor U18710 (N_18710,N_18074,N_18426);
nor U18711 (N_18711,N_18210,N_18225);
and U18712 (N_18712,N_18462,N_18152);
and U18713 (N_18713,N_18109,N_18078);
nand U18714 (N_18714,N_18310,N_18181);
xnor U18715 (N_18715,N_18465,N_18036);
or U18716 (N_18716,N_18171,N_18395);
and U18717 (N_18717,N_18352,N_18366);
xor U18718 (N_18718,N_18386,N_18085);
or U18719 (N_18719,N_18166,N_18467);
nor U18720 (N_18720,N_18253,N_18265);
or U18721 (N_18721,N_18423,N_18041);
nand U18722 (N_18722,N_18321,N_18110);
or U18723 (N_18723,N_18404,N_18103);
and U18724 (N_18724,N_18063,N_18179);
xor U18725 (N_18725,N_18031,N_18400);
or U18726 (N_18726,N_18379,N_18061);
and U18727 (N_18727,N_18228,N_18349);
and U18728 (N_18728,N_18169,N_18484);
nor U18729 (N_18729,N_18175,N_18123);
nor U18730 (N_18730,N_18482,N_18258);
and U18731 (N_18731,N_18140,N_18372);
or U18732 (N_18732,N_18232,N_18393);
nand U18733 (N_18733,N_18285,N_18335);
or U18734 (N_18734,N_18218,N_18380);
or U18735 (N_18735,N_18323,N_18451);
nor U18736 (N_18736,N_18302,N_18273);
or U18737 (N_18737,N_18373,N_18448);
nor U18738 (N_18738,N_18001,N_18496);
xor U18739 (N_18739,N_18115,N_18471);
nand U18740 (N_18740,N_18376,N_18466);
or U18741 (N_18741,N_18214,N_18127);
or U18742 (N_18742,N_18113,N_18195);
nor U18743 (N_18743,N_18211,N_18174);
and U18744 (N_18744,N_18198,N_18023);
xor U18745 (N_18745,N_18168,N_18070);
and U18746 (N_18746,N_18468,N_18374);
xnor U18747 (N_18747,N_18003,N_18443);
xnor U18748 (N_18748,N_18033,N_18283);
nand U18749 (N_18749,N_18472,N_18278);
nor U18750 (N_18750,N_18023,N_18083);
nand U18751 (N_18751,N_18197,N_18059);
nor U18752 (N_18752,N_18227,N_18320);
xor U18753 (N_18753,N_18384,N_18248);
xor U18754 (N_18754,N_18110,N_18146);
nor U18755 (N_18755,N_18289,N_18259);
nor U18756 (N_18756,N_18208,N_18041);
or U18757 (N_18757,N_18058,N_18186);
and U18758 (N_18758,N_18436,N_18227);
nand U18759 (N_18759,N_18484,N_18028);
nor U18760 (N_18760,N_18214,N_18360);
and U18761 (N_18761,N_18012,N_18443);
or U18762 (N_18762,N_18268,N_18347);
nand U18763 (N_18763,N_18482,N_18056);
or U18764 (N_18764,N_18382,N_18221);
nor U18765 (N_18765,N_18267,N_18020);
xor U18766 (N_18766,N_18360,N_18019);
nor U18767 (N_18767,N_18495,N_18024);
nor U18768 (N_18768,N_18344,N_18013);
xnor U18769 (N_18769,N_18043,N_18120);
and U18770 (N_18770,N_18154,N_18183);
nor U18771 (N_18771,N_18381,N_18210);
nand U18772 (N_18772,N_18317,N_18086);
nor U18773 (N_18773,N_18230,N_18400);
and U18774 (N_18774,N_18286,N_18349);
nor U18775 (N_18775,N_18261,N_18292);
xnor U18776 (N_18776,N_18259,N_18371);
nand U18777 (N_18777,N_18193,N_18382);
nand U18778 (N_18778,N_18036,N_18375);
xor U18779 (N_18779,N_18142,N_18199);
or U18780 (N_18780,N_18310,N_18194);
or U18781 (N_18781,N_18398,N_18499);
or U18782 (N_18782,N_18340,N_18169);
or U18783 (N_18783,N_18036,N_18145);
xor U18784 (N_18784,N_18128,N_18412);
or U18785 (N_18785,N_18101,N_18048);
nand U18786 (N_18786,N_18067,N_18193);
and U18787 (N_18787,N_18340,N_18315);
nand U18788 (N_18788,N_18185,N_18286);
nand U18789 (N_18789,N_18243,N_18142);
xnor U18790 (N_18790,N_18301,N_18417);
or U18791 (N_18791,N_18295,N_18411);
or U18792 (N_18792,N_18100,N_18210);
and U18793 (N_18793,N_18223,N_18265);
or U18794 (N_18794,N_18098,N_18166);
nor U18795 (N_18795,N_18300,N_18015);
nor U18796 (N_18796,N_18482,N_18217);
nor U18797 (N_18797,N_18250,N_18303);
and U18798 (N_18798,N_18401,N_18357);
and U18799 (N_18799,N_18167,N_18385);
or U18800 (N_18800,N_18356,N_18072);
nand U18801 (N_18801,N_18016,N_18175);
nand U18802 (N_18802,N_18451,N_18316);
and U18803 (N_18803,N_18202,N_18382);
nor U18804 (N_18804,N_18456,N_18093);
xnor U18805 (N_18805,N_18055,N_18384);
nor U18806 (N_18806,N_18407,N_18170);
xnor U18807 (N_18807,N_18059,N_18338);
and U18808 (N_18808,N_18005,N_18214);
and U18809 (N_18809,N_18383,N_18479);
nand U18810 (N_18810,N_18375,N_18488);
or U18811 (N_18811,N_18121,N_18218);
nand U18812 (N_18812,N_18423,N_18360);
or U18813 (N_18813,N_18009,N_18448);
nor U18814 (N_18814,N_18394,N_18138);
or U18815 (N_18815,N_18226,N_18409);
nor U18816 (N_18816,N_18299,N_18125);
nand U18817 (N_18817,N_18480,N_18012);
nor U18818 (N_18818,N_18105,N_18383);
or U18819 (N_18819,N_18273,N_18143);
nand U18820 (N_18820,N_18417,N_18161);
or U18821 (N_18821,N_18229,N_18178);
or U18822 (N_18822,N_18442,N_18075);
nor U18823 (N_18823,N_18228,N_18099);
xor U18824 (N_18824,N_18416,N_18078);
and U18825 (N_18825,N_18299,N_18000);
xnor U18826 (N_18826,N_18279,N_18374);
nor U18827 (N_18827,N_18230,N_18175);
and U18828 (N_18828,N_18414,N_18044);
and U18829 (N_18829,N_18405,N_18473);
or U18830 (N_18830,N_18080,N_18242);
nor U18831 (N_18831,N_18479,N_18386);
xor U18832 (N_18832,N_18178,N_18318);
and U18833 (N_18833,N_18370,N_18209);
xnor U18834 (N_18834,N_18461,N_18354);
and U18835 (N_18835,N_18466,N_18001);
nor U18836 (N_18836,N_18451,N_18414);
nand U18837 (N_18837,N_18129,N_18420);
or U18838 (N_18838,N_18073,N_18262);
nand U18839 (N_18839,N_18216,N_18480);
xnor U18840 (N_18840,N_18061,N_18412);
nand U18841 (N_18841,N_18084,N_18386);
nor U18842 (N_18842,N_18349,N_18439);
and U18843 (N_18843,N_18288,N_18241);
nor U18844 (N_18844,N_18216,N_18006);
nor U18845 (N_18845,N_18190,N_18126);
or U18846 (N_18846,N_18013,N_18414);
and U18847 (N_18847,N_18359,N_18122);
nor U18848 (N_18848,N_18271,N_18291);
nand U18849 (N_18849,N_18282,N_18006);
or U18850 (N_18850,N_18379,N_18467);
and U18851 (N_18851,N_18354,N_18161);
or U18852 (N_18852,N_18153,N_18133);
or U18853 (N_18853,N_18210,N_18034);
nor U18854 (N_18854,N_18313,N_18011);
xor U18855 (N_18855,N_18162,N_18223);
or U18856 (N_18856,N_18368,N_18308);
xnor U18857 (N_18857,N_18371,N_18340);
nor U18858 (N_18858,N_18200,N_18239);
nand U18859 (N_18859,N_18401,N_18476);
and U18860 (N_18860,N_18225,N_18144);
or U18861 (N_18861,N_18109,N_18418);
nand U18862 (N_18862,N_18011,N_18132);
and U18863 (N_18863,N_18370,N_18222);
nand U18864 (N_18864,N_18374,N_18491);
nor U18865 (N_18865,N_18292,N_18470);
xor U18866 (N_18866,N_18081,N_18215);
or U18867 (N_18867,N_18204,N_18342);
and U18868 (N_18868,N_18382,N_18346);
and U18869 (N_18869,N_18033,N_18055);
or U18870 (N_18870,N_18275,N_18137);
xnor U18871 (N_18871,N_18330,N_18238);
and U18872 (N_18872,N_18306,N_18223);
or U18873 (N_18873,N_18129,N_18279);
or U18874 (N_18874,N_18181,N_18002);
nand U18875 (N_18875,N_18230,N_18200);
nor U18876 (N_18876,N_18008,N_18227);
and U18877 (N_18877,N_18458,N_18478);
nand U18878 (N_18878,N_18112,N_18217);
xor U18879 (N_18879,N_18072,N_18424);
xnor U18880 (N_18880,N_18002,N_18304);
or U18881 (N_18881,N_18366,N_18445);
nand U18882 (N_18882,N_18252,N_18258);
nand U18883 (N_18883,N_18429,N_18358);
nand U18884 (N_18884,N_18412,N_18095);
nor U18885 (N_18885,N_18206,N_18002);
nand U18886 (N_18886,N_18415,N_18285);
nand U18887 (N_18887,N_18423,N_18354);
nor U18888 (N_18888,N_18352,N_18317);
nor U18889 (N_18889,N_18368,N_18460);
xnor U18890 (N_18890,N_18193,N_18021);
and U18891 (N_18891,N_18136,N_18155);
and U18892 (N_18892,N_18203,N_18207);
nand U18893 (N_18893,N_18248,N_18204);
nor U18894 (N_18894,N_18360,N_18227);
or U18895 (N_18895,N_18234,N_18185);
or U18896 (N_18896,N_18367,N_18309);
or U18897 (N_18897,N_18431,N_18094);
xnor U18898 (N_18898,N_18357,N_18194);
nand U18899 (N_18899,N_18290,N_18064);
nor U18900 (N_18900,N_18233,N_18086);
nand U18901 (N_18901,N_18396,N_18381);
xnor U18902 (N_18902,N_18304,N_18452);
nor U18903 (N_18903,N_18297,N_18166);
nor U18904 (N_18904,N_18414,N_18151);
nor U18905 (N_18905,N_18317,N_18206);
xnor U18906 (N_18906,N_18051,N_18104);
or U18907 (N_18907,N_18288,N_18400);
xnor U18908 (N_18908,N_18209,N_18415);
and U18909 (N_18909,N_18217,N_18191);
and U18910 (N_18910,N_18431,N_18088);
nand U18911 (N_18911,N_18144,N_18248);
or U18912 (N_18912,N_18203,N_18197);
xor U18913 (N_18913,N_18283,N_18187);
and U18914 (N_18914,N_18289,N_18357);
xnor U18915 (N_18915,N_18193,N_18374);
and U18916 (N_18916,N_18146,N_18411);
or U18917 (N_18917,N_18276,N_18364);
xor U18918 (N_18918,N_18390,N_18347);
xor U18919 (N_18919,N_18332,N_18097);
and U18920 (N_18920,N_18351,N_18469);
nand U18921 (N_18921,N_18016,N_18339);
xnor U18922 (N_18922,N_18409,N_18496);
xor U18923 (N_18923,N_18375,N_18429);
xor U18924 (N_18924,N_18260,N_18421);
nand U18925 (N_18925,N_18271,N_18243);
nand U18926 (N_18926,N_18494,N_18159);
or U18927 (N_18927,N_18481,N_18301);
and U18928 (N_18928,N_18156,N_18207);
or U18929 (N_18929,N_18309,N_18300);
and U18930 (N_18930,N_18402,N_18168);
and U18931 (N_18931,N_18446,N_18095);
nand U18932 (N_18932,N_18150,N_18208);
or U18933 (N_18933,N_18253,N_18199);
nor U18934 (N_18934,N_18427,N_18050);
or U18935 (N_18935,N_18395,N_18339);
nand U18936 (N_18936,N_18001,N_18028);
and U18937 (N_18937,N_18480,N_18415);
nor U18938 (N_18938,N_18332,N_18394);
nor U18939 (N_18939,N_18055,N_18031);
nor U18940 (N_18940,N_18254,N_18135);
and U18941 (N_18941,N_18496,N_18295);
and U18942 (N_18942,N_18464,N_18282);
and U18943 (N_18943,N_18067,N_18299);
or U18944 (N_18944,N_18459,N_18172);
nand U18945 (N_18945,N_18337,N_18216);
nor U18946 (N_18946,N_18358,N_18485);
nand U18947 (N_18947,N_18139,N_18335);
nor U18948 (N_18948,N_18277,N_18481);
xnor U18949 (N_18949,N_18313,N_18271);
or U18950 (N_18950,N_18499,N_18131);
or U18951 (N_18951,N_18461,N_18095);
and U18952 (N_18952,N_18104,N_18268);
nand U18953 (N_18953,N_18057,N_18424);
and U18954 (N_18954,N_18279,N_18379);
nor U18955 (N_18955,N_18446,N_18325);
nor U18956 (N_18956,N_18209,N_18369);
nand U18957 (N_18957,N_18070,N_18109);
nand U18958 (N_18958,N_18482,N_18200);
xor U18959 (N_18959,N_18348,N_18291);
xnor U18960 (N_18960,N_18297,N_18142);
nand U18961 (N_18961,N_18003,N_18107);
nand U18962 (N_18962,N_18270,N_18163);
xnor U18963 (N_18963,N_18457,N_18079);
xnor U18964 (N_18964,N_18401,N_18015);
and U18965 (N_18965,N_18496,N_18478);
and U18966 (N_18966,N_18431,N_18471);
nor U18967 (N_18967,N_18351,N_18409);
nor U18968 (N_18968,N_18252,N_18428);
or U18969 (N_18969,N_18216,N_18415);
and U18970 (N_18970,N_18006,N_18191);
nor U18971 (N_18971,N_18084,N_18047);
xnor U18972 (N_18972,N_18056,N_18499);
nor U18973 (N_18973,N_18401,N_18452);
or U18974 (N_18974,N_18112,N_18116);
nor U18975 (N_18975,N_18420,N_18421);
and U18976 (N_18976,N_18410,N_18190);
or U18977 (N_18977,N_18487,N_18248);
and U18978 (N_18978,N_18388,N_18485);
nand U18979 (N_18979,N_18186,N_18205);
xnor U18980 (N_18980,N_18104,N_18178);
nor U18981 (N_18981,N_18224,N_18472);
xor U18982 (N_18982,N_18424,N_18069);
or U18983 (N_18983,N_18188,N_18085);
or U18984 (N_18984,N_18313,N_18365);
or U18985 (N_18985,N_18108,N_18296);
nor U18986 (N_18986,N_18415,N_18418);
nand U18987 (N_18987,N_18319,N_18337);
nand U18988 (N_18988,N_18318,N_18150);
and U18989 (N_18989,N_18046,N_18437);
and U18990 (N_18990,N_18389,N_18051);
or U18991 (N_18991,N_18091,N_18491);
xor U18992 (N_18992,N_18290,N_18482);
nor U18993 (N_18993,N_18029,N_18349);
or U18994 (N_18994,N_18148,N_18381);
and U18995 (N_18995,N_18339,N_18204);
and U18996 (N_18996,N_18058,N_18177);
nand U18997 (N_18997,N_18309,N_18204);
xor U18998 (N_18998,N_18204,N_18344);
and U18999 (N_18999,N_18417,N_18284);
or U19000 (N_19000,N_18965,N_18775);
or U19001 (N_19001,N_18570,N_18741);
or U19002 (N_19002,N_18746,N_18514);
or U19003 (N_19003,N_18503,N_18760);
nor U19004 (N_19004,N_18858,N_18949);
nor U19005 (N_19005,N_18914,N_18950);
and U19006 (N_19006,N_18656,N_18872);
nand U19007 (N_19007,N_18921,N_18876);
or U19008 (N_19008,N_18716,N_18789);
and U19009 (N_19009,N_18601,N_18887);
nand U19010 (N_19010,N_18569,N_18770);
or U19011 (N_19011,N_18518,N_18962);
and U19012 (N_19012,N_18780,N_18946);
xor U19013 (N_19013,N_18587,N_18952);
nor U19014 (N_19014,N_18596,N_18781);
xor U19015 (N_19015,N_18571,N_18862);
and U19016 (N_19016,N_18642,N_18592);
or U19017 (N_19017,N_18523,N_18891);
nand U19018 (N_19018,N_18820,N_18925);
xnor U19019 (N_19019,N_18702,N_18577);
or U19020 (N_19020,N_18609,N_18634);
and U19021 (N_19021,N_18703,N_18699);
and U19022 (N_19022,N_18648,N_18755);
and U19023 (N_19023,N_18815,N_18590);
and U19024 (N_19024,N_18606,N_18524);
nor U19025 (N_19025,N_18611,N_18813);
xor U19026 (N_19026,N_18961,N_18973);
nor U19027 (N_19027,N_18974,N_18776);
nor U19028 (N_19028,N_18883,N_18995);
or U19029 (N_19029,N_18810,N_18796);
nor U19030 (N_19030,N_18807,N_18607);
nor U19031 (N_19031,N_18839,N_18672);
or U19032 (N_19032,N_18764,N_18725);
xnor U19033 (N_19033,N_18993,N_18855);
and U19034 (N_19034,N_18882,N_18941);
and U19035 (N_19035,N_18561,N_18701);
nand U19036 (N_19036,N_18976,N_18557);
nor U19037 (N_19037,N_18693,N_18720);
nor U19038 (N_19038,N_18553,N_18654);
nand U19039 (N_19039,N_18541,N_18788);
xnor U19040 (N_19040,N_18738,N_18920);
nand U19041 (N_19041,N_18660,N_18830);
nor U19042 (N_19042,N_18522,N_18826);
nand U19043 (N_19043,N_18762,N_18836);
nand U19044 (N_19044,N_18657,N_18893);
and U19045 (N_19045,N_18564,N_18583);
xnor U19046 (N_19046,N_18581,N_18774);
or U19047 (N_19047,N_18797,N_18875);
nand U19048 (N_19048,N_18623,N_18852);
xor U19049 (N_19049,N_18512,N_18558);
xor U19050 (N_19050,N_18707,N_18566);
nand U19051 (N_19051,N_18972,N_18730);
xor U19052 (N_19052,N_18911,N_18689);
and U19053 (N_19053,N_18799,N_18683);
and U19054 (N_19054,N_18595,N_18958);
or U19055 (N_19055,N_18842,N_18975);
xnor U19056 (N_19056,N_18812,N_18988);
or U19057 (N_19057,N_18837,N_18533);
nor U19058 (N_19058,N_18579,N_18981);
xor U19059 (N_19059,N_18968,N_18767);
and U19060 (N_19060,N_18506,N_18772);
or U19061 (N_19061,N_18804,N_18632);
nand U19062 (N_19062,N_18681,N_18625);
xnor U19063 (N_19063,N_18884,N_18873);
nand U19064 (N_19064,N_18684,N_18811);
nor U19065 (N_19065,N_18889,N_18602);
and U19066 (N_19066,N_18863,N_18795);
and U19067 (N_19067,N_18585,N_18906);
and U19068 (N_19068,N_18990,N_18828);
nor U19069 (N_19069,N_18645,N_18881);
nand U19070 (N_19070,N_18675,N_18713);
nor U19071 (N_19071,N_18752,N_18859);
xor U19072 (N_19072,N_18792,N_18868);
or U19073 (N_19073,N_18616,N_18535);
nand U19074 (N_19074,N_18886,N_18817);
and U19075 (N_19075,N_18531,N_18897);
nand U19076 (N_19076,N_18998,N_18662);
xor U19077 (N_19077,N_18655,N_18549);
or U19078 (N_19078,N_18945,N_18546);
nand U19079 (N_19079,N_18930,N_18710);
nor U19080 (N_19080,N_18668,N_18633);
nand U19081 (N_19081,N_18980,N_18850);
or U19082 (N_19082,N_18833,N_18615);
nor U19083 (N_19083,N_18635,N_18900);
nand U19084 (N_19084,N_18849,N_18790);
nor U19085 (N_19085,N_18773,N_18860);
and U19086 (N_19086,N_18761,N_18907);
nand U19087 (N_19087,N_18905,N_18644);
nand U19088 (N_19088,N_18674,N_18992);
or U19089 (N_19089,N_18769,N_18794);
nand U19090 (N_19090,N_18621,N_18745);
nand U19091 (N_19091,N_18622,N_18798);
nor U19092 (N_19092,N_18573,N_18680);
and U19093 (N_19093,N_18824,N_18779);
nand U19094 (N_19094,N_18664,N_18909);
xor U19095 (N_19095,N_18538,N_18584);
nand U19096 (N_19096,N_18869,N_18574);
or U19097 (N_19097,N_18526,N_18898);
xnor U19098 (N_19098,N_18866,N_18731);
nor U19099 (N_19099,N_18617,N_18955);
nor U19100 (N_19100,N_18540,N_18959);
xor U19101 (N_19101,N_18562,N_18696);
xnor U19102 (N_19102,N_18953,N_18782);
nand U19103 (N_19103,N_18971,N_18578);
nor U19104 (N_19104,N_18851,N_18588);
nor U19105 (N_19105,N_18537,N_18610);
nand U19106 (N_19106,N_18509,N_18697);
or U19107 (N_19107,N_18986,N_18880);
or U19108 (N_19108,N_18960,N_18966);
and U19109 (N_19109,N_18737,N_18519);
and U19110 (N_19110,N_18723,N_18676);
nor U19111 (N_19111,N_18791,N_18597);
xnor U19112 (N_19112,N_18977,N_18806);
nand U19113 (N_19113,N_18923,N_18848);
and U19114 (N_19114,N_18671,N_18756);
nor U19115 (N_19115,N_18888,N_18834);
nor U19116 (N_19116,N_18910,N_18832);
or U19117 (N_19117,N_18734,N_18547);
or U19118 (N_19118,N_18554,N_18690);
xor U19119 (N_19119,N_18517,N_18515);
nand U19120 (N_19120,N_18525,N_18908);
and U19121 (N_19121,N_18957,N_18678);
nand U19122 (N_19122,N_18765,N_18661);
nand U19123 (N_19123,N_18956,N_18922);
xor U19124 (N_19124,N_18864,N_18530);
nand U19125 (N_19125,N_18800,N_18840);
nor U19126 (N_19126,N_18695,N_18637);
xor U19127 (N_19127,N_18704,N_18529);
and U19128 (N_19128,N_18709,N_18626);
nor U19129 (N_19129,N_18721,N_18739);
nand U19130 (N_19130,N_18801,N_18895);
xnor U19131 (N_19131,N_18854,N_18935);
nand U19132 (N_19132,N_18827,N_18989);
and U19133 (N_19133,N_18636,N_18614);
or U19134 (N_19134,N_18659,N_18736);
nor U19135 (N_19135,N_18630,N_18818);
nor U19136 (N_19136,N_18777,N_18631);
nand U19137 (N_19137,N_18857,N_18802);
or U19138 (N_19138,N_18618,N_18933);
and U19139 (N_19139,N_18712,N_18890);
nor U19140 (N_19140,N_18539,N_18983);
or U19141 (N_19141,N_18843,N_18751);
and U19142 (N_19142,N_18663,N_18867);
or U19143 (N_19143,N_18567,N_18521);
or U19144 (N_19144,N_18809,N_18901);
nand U19145 (N_19145,N_18786,N_18542);
xnor U19146 (N_19146,N_18768,N_18722);
nor U19147 (N_19147,N_18604,N_18728);
xnor U19148 (N_19148,N_18706,N_18576);
xnor U19149 (N_19149,N_18670,N_18856);
and U19150 (N_19150,N_18766,N_18744);
and U19151 (N_19151,N_18698,N_18679);
xnor U19152 (N_19152,N_18673,N_18692);
nor U19153 (N_19153,N_18532,N_18651);
xnor U19154 (N_19154,N_18669,N_18686);
or U19155 (N_19155,N_18598,N_18917);
nand U19156 (N_19156,N_18892,N_18783);
xor U19157 (N_19157,N_18613,N_18719);
and U19158 (N_19158,N_18999,N_18551);
and U19159 (N_19159,N_18740,N_18653);
or U19160 (N_19160,N_18778,N_18688);
and U19161 (N_19161,N_18919,N_18628);
or U19162 (N_19162,N_18500,N_18527);
nor U19163 (N_19163,N_18967,N_18808);
nor U19164 (N_19164,N_18505,N_18639);
nand U19165 (N_19165,N_18853,N_18511);
or U19166 (N_19166,N_18787,N_18589);
nand U19167 (N_19167,N_18847,N_18507);
and U19168 (N_19168,N_18726,N_18685);
or U19169 (N_19169,N_18915,N_18708);
nand U19170 (N_19170,N_18575,N_18705);
xnor U19171 (N_19171,N_18711,N_18927);
nor U19172 (N_19172,N_18580,N_18603);
nand U19173 (N_19173,N_18885,N_18552);
nand U19174 (N_19174,N_18819,N_18504);
and U19175 (N_19175,N_18757,N_18643);
and U19176 (N_19176,N_18743,N_18687);
xor U19177 (N_19177,N_18665,N_18940);
or U19178 (N_19178,N_18534,N_18560);
xor U19179 (N_19179,N_18793,N_18870);
or U19180 (N_19180,N_18929,N_18555);
xnor U19181 (N_19181,N_18572,N_18608);
nand U19182 (N_19182,N_18510,N_18994);
and U19183 (N_19183,N_18831,N_18638);
xor U19184 (N_19184,N_18987,N_18747);
and U19185 (N_19185,N_18829,N_18931);
and U19186 (N_19186,N_18948,N_18846);
or U19187 (N_19187,N_18700,N_18677);
nand U19188 (N_19188,N_18822,N_18785);
or U19189 (N_19189,N_18733,N_18821);
and U19190 (N_19190,N_18896,N_18691);
and U19191 (N_19191,N_18928,N_18620);
xor U19192 (N_19192,N_18913,N_18749);
and U19193 (N_19193,N_18682,N_18624);
and U19194 (N_19194,N_18874,N_18825);
xnor U19195 (N_19195,N_18528,N_18649);
nor U19196 (N_19196,N_18586,N_18784);
or U19197 (N_19197,N_18964,N_18750);
nand U19198 (N_19198,N_18865,N_18543);
or U19199 (N_19199,N_18666,N_18904);
nor U19200 (N_19200,N_18600,N_18916);
nor U19201 (N_19201,N_18970,N_18985);
and U19202 (N_19202,N_18902,N_18984);
or U19203 (N_19203,N_18715,N_18939);
nor U19204 (N_19204,N_18894,N_18727);
nand U19205 (N_19205,N_18835,N_18877);
xor U19206 (N_19206,N_18568,N_18758);
or U19207 (N_19207,N_18627,N_18763);
xnor U19208 (N_19208,N_18501,N_18878);
and U19209 (N_19209,N_18997,N_18803);
nand U19210 (N_19210,N_18871,N_18978);
xor U19211 (N_19211,N_18742,N_18718);
and U19212 (N_19212,N_18924,N_18646);
nand U19213 (N_19213,N_18748,N_18550);
or U19214 (N_19214,N_18918,N_18816);
nor U19215 (N_19215,N_18934,N_18947);
or U19216 (N_19216,N_18544,N_18963);
nor U19217 (N_19217,N_18735,N_18667);
and U19218 (N_19218,N_18841,N_18814);
xor U19219 (N_19219,N_18838,N_18593);
or U19220 (N_19220,N_18516,N_18753);
nand U19221 (N_19221,N_18520,N_18938);
or U19222 (N_19222,N_18942,N_18943);
or U19223 (N_19223,N_18605,N_18556);
or U19224 (N_19224,N_18652,N_18844);
nor U19225 (N_19225,N_18951,N_18619);
and U19226 (N_19226,N_18612,N_18658);
and U19227 (N_19227,N_18640,N_18944);
nand U19228 (N_19228,N_18879,N_18805);
nand U19229 (N_19229,N_18650,N_18508);
and U19230 (N_19230,N_18926,N_18641);
nor U19231 (N_19231,N_18724,N_18823);
nor U19232 (N_19232,N_18502,N_18717);
nand U19233 (N_19233,N_18565,N_18759);
nand U19234 (N_19234,N_18754,N_18647);
and U19235 (N_19235,N_18932,N_18845);
and U19236 (N_19236,N_18969,N_18937);
and U19237 (N_19237,N_18861,N_18714);
nand U19238 (N_19238,N_18979,N_18594);
nor U19239 (N_19239,N_18513,N_18563);
and U19240 (N_19240,N_18936,N_18771);
xnor U19241 (N_19241,N_18954,N_18629);
or U19242 (N_19242,N_18545,N_18991);
nor U19243 (N_19243,N_18599,N_18548);
and U19244 (N_19244,N_18996,N_18732);
and U19245 (N_19245,N_18694,N_18729);
nor U19246 (N_19246,N_18982,N_18559);
nor U19247 (N_19247,N_18899,N_18912);
nor U19248 (N_19248,N_18582,N_18591);
nand U19249 (N_19249,N_18903,N_18536);
nand U19250 (N_19250,N_18533,N_18555);
and U19251 (N_19251,N_18904,N_18550);
and U19252 (N_19252,N_18545,N_18624);
xnor U19253 (N_19253,N_18596,N_18759);
or U19254 (N_19254,N_18787,N_18797);
nor U19255 (N_19255,N_18836,N_18802);
xor U19256 (N_19256,N_18588,N_18716);
nand U19257 (N_19257,N_18989,N_18794);
and U19258 (N_19258,N_18936,N_18548);
and U19259 (N_19259,N_18717,N_18929);
and U19260 (N_19260,N_18908,N_18858);
or U19261 (N_19261,N_18891,N_18636);
and U19262 (N_19262,N_18847,N_18849);
or U19263 (N_19263,N_18635,N_18777);
or U19264 (N_19264,N_18821,N_18855);
or U19265 (N_19265,N_18648,N_18761);
xnor U19266 (N_19266,N_18826,N_18552);
xnor U19267 (N_19267,N_18784,N_18688);
xor U19268 (N_19268,N_18835,N_18843);
or U19269 (N_19269,N_18669,N_18561);
xnor U19270 (N_19270,N_18828,N_18862);
xor U19271 (N_19271,N_18652,N_18740);
or U19272 (N_19272,N_18636,N_18867);
nor U19273 (N_19273,N_18801,N_18755);
and U19274 (N_19274,N_18749,N_18801);
nand U19275 (N_19275,N_18996,N_18894);
and U19276 (N_19276,N_18514,N_18901);
nand U19277 (N_19277,N_18837,N_18547);
nand U19278 (N_19278,N_18996,N_18544);
nor U19279 (N_19279,N_18846,N_18635);
xor U19280 (N_19280,N_18996,N_18648);
or U19281 (N_19281,N_18541,N_18744);
nor U19282 (N_19282,N_18611,N_18994);
or U19283 (N_19283,N_18727,N_18653);
nand U19284 (N_19284,N_18908,N_18506);
and U19285 (N_19285,N_18618,N_18954);
nor U19286 (N_19286,N_18900,N_18861);
or U19287 (N_19287,N_18573,N_18540);
nand U19288 (N_19288,N_18772,N_18935);
nand U19289 (N_19289,N_18808,N_18565);
xor U19290 (N_19290,N_18615,N_18855);
nor U19291 (N_19291,N_18727,N_18872);
or U19292 (N_19292,N_18982,N_18892);
or U19293 (N_19293,N_18927,N_18856);
nor U19294 (N_19294,N_18674,N_18618);
or U19295 (N_19295,N_18753,N_18969);
xor U19296 (N_19296,N_18684,N_18820);
nor U19297 (N_19297,N_18707,N_18746);
xnor U19298 (N_19298,N_18580,N_18944);
xor U19299 (N_19299,N_18967,N_18664);
or U19300 (N_19300,N_18637,N_18948);
nor U19301 (N_19301,N_18758,N_18908);
nor U19302 (N_19302,N_18878,N_18989);
nor U19303 (N_19303,N_18928,N_18824);
or U19304 (N_19304,N_18519,N_18787);
or U19305 (N_19305,N_18555,N_18677);
xor U19306 (N_19306,N_18772,N_18944);
xnor U19307 (N_19307,N_18797,N_18538);
nor U19308 (N_19308,N_18912,N_18525);
and U19309 (N_19309,N_18628,N_18528);
xnor U19310 (N_19310,N_18621,N_18846);
nand U19311 (N_19311,N_18598,N_18784);
nor U19312 (N_19312,N_18868,N_18534);
and U19313 (N_19313,N_18842,N_18844);
nand U19314 (N_19314,N_18553,N_18617);
xnor U19315 (N_19315,N_18875,N_18835);
or U19316 (N_19316,N_18812,N_18678);
or U19317 (N_19317,N_18679,N_18660);
nand U19318 (N_19318,N_18588,N_18994);
nand U19319 (N_19319,N_18569,N_18926);
xnor U19320 (N_19320,N_18842,N_18947);
xor U19321 (N_19321,N_18732,N_18573);
nor U19322 (N_19322,N_18958,N_18849);
xor U19323 (N_19323,N_18769,N_18721);
xnor U19324 (N_19324,N_18926,N_18839);
or U19325 (N_19325,N_18954,N_18675);
nor U19326 (N_19326,N_18696,N_18504);
xnor U19327 (N_19327,N_18565,N_18677);
and U19328 (N_19328,N_18688,N_18924);
nor U19329 (N_19329,N_18757,N_18525);
nand U19330 (N_19330,N_18646,N_18770);
and U19331 (N_19331,N_18700,N_18716);
nor U19332 (N_19332,N_18958,N_18861);
and U19333 (N_19333,N_18555,N_18820);
and U19334 (N_19334,N_18730,N_18848);
xor U19335 (N_19335,N_18691,N_18743);
or U19336 (N_19336,N_18508,N_18930);
nand U19337 (N_19337,N_18843,N_18867);
or U19338 (N_19338,N_18896,N_18664);
nand U19339 (N_19339,N_18631,N_18514);
nor U19340 (N_19340,N_18849,N_18583);
nor U19341 (N_19341,N_18879,N_18815);
nor U19342 (N_19342,N_18565,N_18912);
xnor U19343 (N_19343,N_18756,N_18805);
xor U19344 (N_19344,N_18767,N_18679);
xor U19345 (N_19345,N_18608,N_18871);
and U19346 (N_19346,N_18522,N_18899);
xor U19347 (N_19347,N_18881,N_18836);
nand U19348 (N_19348,N_18727,N_18816);
xnor U19349 (N_19349,N_18649,N_18667);
or U19350 (N_19350,N_18610,N_18814);
nor U19351 (N_19351,N_18908,N_18594);
or U19352 (N_19352,N_18793,N_18726);
nand U19353 (N_19353,N_18712,N_18738);
or U19354 (N_19354,N_18806,N_18810);
nand U19355 (N_19355,N_18545,N_18756);
xnor U19356 (N_19356,N_18786,N_18818);
and U19357 (N_19357,N_18655,N_18925);
xor U19358 (N_19358,N_18925,N_18957);
nand U19359 (N_19359,N_18830,N_18965);
nor U19360 (N_19360,N_18618,N_18714);
nand U19361 (N_19361,N_18888,N_18531);
or U19362 (N_19362,N_18930,N_18671);
nand U19363 (N_19363,N_18721,N_18875);
or U19364 (N_19364,N_18928,N_18720);
or U19365 (N_19365,N_18810,N_18938);
or U19366 (N_19366,N_18623,N_18986);
nor U19367 (N_19367,N_18919,N_18570);
xnor U19368 (N_19368,N_18632,N_18612);
and U19369 (N_19369,N_18687,N_18948);
nor U19370 (N_19370,N_18640,N_18976);
or U19371 (N_19371,N_18784,N_18535);
and U19372 (N_19372,N_18961,N_18629);
or U19373 (N_19373,N_18669,N_18521);
nor U19374 (N_19374,N_18938,N_18963);
nor U19375 (N_19375,N_18709,N_18777);
and U19376 (N_19376,N_18664,N_18575);
and U19377 (N_19377,N_18790,N_18573);
and U19378 (N_19378,N_18940,N_18637);
nor U19379 (N_19379,N_18866,N_18605);
and U19380 (N_19380,N_18849,N_18730);
nand U19381 (N_19381,N_18524,N_18659);
nand U19382 (N_19382,N_18650,N_18952);
nor U19383 (N_19383,N_18825,N_18575);
nand U19384 (N_19384,N_18969,N_18725);
nand U19385 (N_19385,N_18787,N_18615);
and U19386 (N_19386,N_18540,N_18517);
nor U19387 (N_19387,N_18641,N_18514);
nand U19388 (N_19388,N_18871,N_18758);
xor U19389 (N_19389,N_18841,N_18502);
and U19390 (N_19390,N_18791,N_18965);
xnor U19391 (N_19391,N_18521,N_18846);
and U19392 (N_19392,N_18517,N_18502);
xor U19393 (N_19393,N_18561,N_18789);
nor U19394 (N_19394,N_18609,N_18773);
nand U19395 (N_19395,N_18876,N_18924);
xnor U19396 (N_19396,N_18567,N_18695);
xor U19397 (N_19397,N_18542,N_18521);
nor U19398 (N_19398,N_18855,N_18755);
nor U19399 (N_19399,N_18584,N_18592);
or U19400 (N_19400,N_18963,N_18513);
or U19401 (N_19401,N_18579,N_18532);
nand U19402 (N_19402,N_18837,N_18551);
xnor U19403 (N_19403,N_18833,N_18896);
nand U19404 (N_19404,N_18793,N_18953);
and U19405 (N_19405,N_18626,N_18797);
nand U19406 (N_19406,N_18640,N_18557);
nand U19407 (N_19407,N_18815,N_18857);
nor U19408 (N_19408,N_18634,N_18776);
and U19409 (N_19409,N_18759,N_18775);
or U19410 (N_19410,N_18726,N_18523);
or U19411 (N_19411,N_18633,N_18858);
or U19412 (N_19412,N_18695,N_18513);
or U19413 (N_19413,N_18512,N_18601);
and U19414 (N_19414,N_18705,N_18526);
or U19415 (N_19415,N_18833,N_18911);
nand U19416 (N_19416,N_18542,N_18718);
or U19417 (N_19417,N_18563,N_18535);
xnor U19418 (N_19418,N_18967,N_18506);
and U19419 (N_19419,N_18804,N_18703);
nand U19420 (N_19420,N_18509,N_18958);
or U19421 (N_19421,N_18800,N_18716);
nand U19422 (N_19422,N_18991,N_18578);
xor U19423 (N_19423,N_18665,N_18529);
nor U19424 (N_19424,N_18970,N_18822);
nand U19425 (N_19425,N_18821,N_18546);
nor U19426 (N_19426,N_18881,N_18695);
nor U19427 (N_19427,N_18821,N_18903);
nand U19428 (N_19428,N_18946,N_18653);
nand U19429 (N_19429,N_18695,N_18940);
and U19430 (N_19430,N_18725,N_18684);
nor U19431 (N_19431,N_18966,N_18729);
xor U19432 (N_19432,N_18677,N_18725);
or U19433 (N_19433,N_18834,N_18578);
nor U19434 (N_19434,N_18946,N_18792);
nor U19435 (N_19435,N_18554,N_18511);
xor U19436 (N_19436,N_18697,N_18586);
nor U19437 (N_19437,N_18652,N_18939);
nor U19438 (N_19438,N_18667,N_18746);
xor U19439 (N_19439,N_18998,N_18983);
or U19440 (N_19440,N_18892,N_18724);
xor U19441 (N_19441,N_18666,N_18782);
xor U19442 (N_19442,N_18771,N_18923);
xnor U19443 (N_19443,N_18507,N_18989);
xnor U19444 (N_19444,N_18567,N_18838);
xnor U19445 (N_19445,N_18500,N_18868);
nor U19446 (N_19446,N_18887,N_18732);
and U19447 (N_19447,N_18956,N_18706);
nand U19448 (N_19448,N_18547,N_18996);
xnor U19449 (N_19449,N_18549,N_18821);
nand U19450 (N_19450,N_18866,N_18660);
and U19451 (N_19451,N_18821,N_18697);
nand U19452 (N_19452,N_18737,N_18949);
nor U19453 (N_19453,N_18926,N_18993);
xnor U19454 (N_19454,N_18994,N_18993);
nand U19455 (N_19455,N_18571,N_18570);
nor U19456 (N_19456,N_18706,N_18783);
xnor U19457 (N_19457,N_18979,N_18618);
nor U19458 (N_19458,N_18925,N_18559);
xor U19459 (N_19459,N_18880,N_18742);
and U19460 (N_19460,N_18864,N_18519);
and U19461 (N_19461,N_18543,N_18957);
xor U19462 (N_19462,N_18562,N_18751);
nor U19463 (N_19463,N_18624,N_18953);
nand U19464 (N_19464,N_18588,N_18714);
nor U19465 (N_19465,N_18559,N_18823);
nand U19466 (N_19466,N_18868,N_18842);
xnor U19467 (N_19467,N_18995,N_18673);
nand U19468 (N_19468,N_18719,N_18820);
nand U19469 (N_19469,N_18679,N_18858);
nor U19470 (N_19470,N_18635,N_18932);
and U19471 (N_19471,N_18725,N_18540);
or U19472 (N_19472,N_18700,N_18995);
nand U19473 (N_19473,N_18901,N_18936);
and U19474 (N_19474,N_18688,N_18841);
xor U19475 (N_19475,N_18650,N_18825);
nor U19476 (N_19476,N_18665,N_18736);
nor U19477 (N_19477,N_18794,N_18538);
and U19478 (N_19478,N_18525,N_18603);
or U19479 (N_19479,N_18903,N_18874);
nor U19480 (N_19480,N_18913,N_18757);
or U19481 (N_19481,N_18545,N_18828);
and U19482 (N_19482,N_18957,N_18975);
nand U19483 (N_19483,N_18755,N_18820);
nor U19484 (N_19484,N_18716,N_18875);
or U19485 (N_19485,N_18923,N_18745);
and U19486 (N_19486,N_18955,N_18770);
xor U19487 (N_19487,N_18784,N_18945);
xnor U19488 (N_19488,N_18778,N_18842);
or U19489 (N_19489,N_18602,N_18654);
xnor U19490 (N_19490,N_18567,N_18950);
nor U19491 (N_19491,N_18805,N_18624);
xor U19492 (N_19492,N_18917,N_18766);
and U19493 (N_19493,N_18936,N_18963);
nand U19494 (N_19494,N_18816,N_18782);
nor U19495 (N_19495,N_18922,N_18609);
xor U19496 (N_19496,N_18555,N_18694);
and U19497 (N_19497,N_18669,N_18864);
nand U19498 (N_19498,N_18820,N_18544);
xnor U19499 (N_19499,N_18545,N_18787);
nor U19500 (N_19500,N_19475,N_19195);
nor U19501 (N_19501,N_19393,N_19367);
nand U19502 (N_19502,N_19117,N_19217);
and U19503 (N_19503,N_19280,N_19123);
and U19504 (N_19504,N_19069,N_19019);
nor U19505 (N_19505,N_19040,N_19423);
nand U19506 (N_19506,N_19115,N_19318);
nand U19507 (N_19507,N_19490,N_19452);
nand U19508 (N_19508,N_19128,N_19396);
nand U19509 (N_19509,N_19402,N_19350);
nand U19510 (N_19510,N_19205,N_19065);
and U19511 (N_19511,N_19159,N_19200);
or U19512 (N_19512,N_19301,N_19213);
or U19513 (N_19513,N_19204,N_19493);
or U19514 (N_19514,N_19339,N_19078);
xor U19515 (N_19515,N_19351,N_19068);
nor U19516 (N_19516,N_19429,N_19267);
nor U19517 (N_19517,N_19037,N_19137);
xor U19518 (N_19518,N_19212,N_19265);
and U19519 (N_19519,N_19394,N_19100);
nand U19520 (N_19520,N_19033,N_19438);
xnor U19521 (N_19521,N_19409,N_19197);
nor U19522 (N_19522,N_19106,N_19361);
and U19523 (N_19523,N_19164,N_19118);
nor U19524 (N_19524,N_19007,N_19229);
nand U19525 (N_19525,N_19447,N_19162);
xor U19526 (N_19526,N_19016,N_19463);
and U19527 (N_19527,N_19306,N_19485);
nor U19528 (N_19528,N_19253,N_19290);
xnor U19529 (N_19529,N_19289,N_19122);
or U19530 (N_19530,N_19376,N_19093);
or U19531 (N_19531,N_19021,N_19334);
nand U19532 (N_19532,N_19488,N_19067);
xnor U19533 (N_19533,N_19154,N_19134);
and U19534 (N_19534,N_19096,N_19145);
and U19535 (N_19535,N_19222,N_19446);
and U19536 (N_19536,N_19331,N_19214);
nor U19537 (N_19537,N_19435,N_19398);
nor U19538 (N_19538,N_19010,N_19104);
and U19539 (N_19539,N_19101,N_19340);
xnor U19540 (N_19540,N_19170,N_19043);
or U19541 (N_19541,N_19032,N_19410);
or U19542 (N_19542,N_19129,N_19413);
and U19543 (N_19543,N_19184,N_19120);
and U19544 (N_19544,N_19173,N_19035);
nor U19545 (N_19545,N_19194,N_19210);
and U19546 (N_19546,N_19342,N_19270);
nand U19547 (N_19547,N_19277,N_19023);
nand U19548 (N_19548,N_19076,N_19260);
and U19549 (N_19549,N_19244,N_19360);
xor U19550 (N_19550,N_19044,N_19415);
nor U19551 (N_19551,N_19223,N_19450);
xnor U19552 (N_19552,N_19169,N_19070);
nor U19553 (N_19553,N_19264,N_19378);
and U19554 (N_19554,N_19356,N_19155);
nand U19555 (N_19555,N_19457,N_19333);
and U19556 (N_19556,N_19309,N_19209);
and U19557 (N_19557,N_19303,N_19110);
nor U19558 (N_19558,N_19077,N_19433);
nand U19559 (N_19559,N_19114,N_19291);
and U19560 (N_19560,N_19001,N_19241);
xor U19561 (N_19561,N_19025,N_19317);
and U19562 (N_19562,N_19481,N_19235);
or U19563 (N_19563,N_19284,N_19363);
xor U19564 (N_19564,N_19458,N_19300);
nand U19565 (N_19565,N_19431,N_19066);
or U19566 (N_19566,N_19151,N_19332);
nand U19567 (N_19567,N_19233,N_19304);
nand U19568 (N_19568,N_19459,N_19052);
or U19569 (N_19569,N_19246,N_19368);
xor U19570 (N_19570,N_19183,N_19256);
nor U19571 (N_19571,N_19091,N_19479);
xor U19572 (N_19572,N_19116,N_19236);
nor U19573 (N_19573,N_19072,N_19189);
nor U19574 (N_19574,N_19422,N_19056);
xor U19575 (N_19575,N_19299,N_19421);
and U19576 (N_19576,N_19330,N_19337);
and U19577 (N_19577,N_19392,N_19175);
nand U19578 (N_19578,N_19105,N_19387);
and U19579 (N_19579,N_19397,N_19419);
nor U19580 (N_19580,N_19036,N_19403);
and U19581 (N_19581,N_19441,N_19090);
or U19582 (N_19582,N_19168,N_19268);
nor U19583 (N_19583,N_19219,N_19092);
and U19584 (N_19584,N_19171,N_19028);
nor U19585 (N_19585,N_19266,N_19257);
or U19586 (N_19586,N_19487,N_19058);
or U19587 (N_19587,N_19095,N_19180);
nand U19588 (N_19588,N_19187,N_19167);
and U19589 (N_19589,N_19443,N_19478);
nand U19590 (N_19590,N_19285,N_19074);
xor U19591 (N_19591,N_19430,N_19460);
nor U19592 (N_19592,N_19152,N_19148);
nand U19593 (N_19593,N_19375,N_19005);
or U19594 (N_19594,N_19373,N_19472);
xor U19595 (N_19595,N_19379,N_19407);
nand U19596 (N_19596,N_19225,N_19081);
and U19597 (N_19597,N_19172,N_19130);
or U19598 (N_19598,N_19160,N_19377);
nor U19599 (N_19599,N_19055,N_19121);
xor U19600 (N_19600,N_19020,N_19372);
or U19601 (N_19601,N_19254,N_19243);
nand U19602 (N_19602,N_19495,N_19370);
and U19603 (N_19603,N_19408,N_19251);
or U19604 (N_19604,N_19271,N_19305);
and U19605 (N_19605,N_19030,N_19302);
and U19606 (N_19606,N_19085,N_19287);
nor U19607 (N_19607,N_19136,N_19412);
nor U19608 (N_19608,N_19494,N_19111);
or U19609 (N_19609,N_19215,N_19467);
nor U19610 (N_19610,N_19158,N_19341);
and U19611 (N_19611,N_19426,N_19273);
or U19612 (N_19612,N_19144,N_19073);
nand U19613 (N_19613,N_19462,N_19324);
xor U19614 (N_19614,N_19099,N_19456);
or U19615 (N_19615,N_19046,N_19424);
xor U19616 (N_19616,N_19064,N_19322);
xnor U19617 (N_19617,N_19464,N_19161);
nand U19618 (N_19618,N_19261,N_19147);
nor U19619 (N_19619,N_19027,N_19166);
nand U19620 (N_19620,N_19211,N_19482);
or U19621 (N_19621,N_19432,N_19060);
nor U19622 (N_19622,N_19124,N_19202);
xor U19623 (N_19623,N_19362,N_19442);
nand U19624 (N_19624,N_19477,N_19142);
or U19625 (N_19625,N_19262,N_19000);
or U19626 (N_19626,N_19017,N_19191);
xnor U19627 (N_19627,N_19269,N_19371);
or U19628 (N_19628,N_19050,N_19240);
xnor U19629 (N_19629,N_19496,N_19181);
nor U19630 (N_19630,N_19230,N_19112);
nand U19631 (N_19631,N_19084,N_19366);
and U19632 (N_19632,N_19102,N_19454);
xnor U19633 (N_19633,N_19048,N_19150);
nand U19634 (N_19634,N_19216,N_19185);
xnor U19635 (N_19635,N_19358,N_19059);
xor U19636 (N_19636,N_19042,N_19400);
nor U19637 (N_19637,N_19208,N_19497);
or U19638 (N_19638,N_19338,N_19193);
xnor U19639 (N_19639,N_19390,N_19250);
xor U19640 (N_19640,N_19468,N_19153);
nor U19641 (N_19641,N_19247,N_19119);
and U19642 (N_19642,N_19307,N_19355);
xor U19643 (N_19643,N_19486,N_19440);
or U19644 (N_19644,N_19080,N_19312);
nand U19645 (N_19645,N_19483,N_19013);
nand U19646 (N_19646,N_19245,N_19038);
or U19647 (N_19647,N_19022,N_19049);
and U19648 (N_19648,N_19418,N_19420);
xnor U19649 (N_19649,N_19428,N_19316);
nor U19650 (N_19650,N_19138,N_19224);
or U19651 (N_19651,N_19239,N_19006);
and U19652 (N_19652,N_19258,N_19218);
nand U19653 (N_19653,N_19346,N_19344);
nand U19654 (N_19654,N_19113,N_19369);
nand U19655 (N_19655,N_19404,N_19276);
xnor U19656 (N_19656,N_19480,N_19384);
xnor U19657 (N_19657,N_19131,N_19201);
xnor U19658 (N_19658,N_19034,N_19009);
or U19659 (N_19659,N_19436,N_19226);
or U19660 (N_19660,N_19414,N_19071);
nor U19661 (N_19661,N_19045,N_19125);
nor U19662 (N_19662,N_19374,N_19295);
nor U19663 (N_19663,N_19274,N_19278);
and U19664 (N_19664,N_19026,N_19308);
nand U19665 (N_19665,N_19087,N_19177);
xor U19666 (N_19666,N_19190,N_19263);
nand U19667 (N_19667,N_19015,N_19383);
xor U19668 (N_19668,N_19051,N_19196);
and U19669 (N_19669,N_19326,N_19186);
nand U19670 (N_19670,N_19364,N_19089);
nor U19671 (N_19671,N_19465,N_19395);
nor U19672 (N_19672,N_19365,N_19109);
and U19673 (N_19673,N_19381,N_19206);
or U19674 (N_19674,N_19416,N_19434);
or U19675 (N_19675,N_19149,N_19437);
or U19676 (N_19676,N_19199,N_19139);
nor U19677 (N_19677,N_19335,N_19461);
or U19678 (N_19678,N_19179,N_19126);
nor U19679 (N_19679,N_19391,N_19327);
and U19680 (N_19680,N_19328,N_19231);
and U19681 (N_19681,N_19228,N_19348);
nand U19682 (N_19682,N_19029,N_19024);
and U19683 (N_19683,N_19275,N_19135);
xor U19684 (N_19684,N_19491,N_19476);
nor U19685 (N_19685,N_19140,N_19207);
nor U19686 (N_19686,N_19133,N_19062);
or U19687 (N_19687,N_19313,N_19174);
xnor U19688 (N_19688,N_19314,N_19469);
nor U19689 (N_19689,N_19405,N_19054);
xnor U19690 (N_19690,N_19382,N_19473);
nand U19691 (N_19691,N_19227,N_19088);
nand U19692 (N_19692,N_19466,N_19484);
nor U19693 (N_19693,N_19315,N_19498);
and U19694 (N_19694,N_19012,N_19310);
nor U19695 (N_19695,N_19386,N_19141);
nor U19696 (N_19696,N_19293,N_19083);
or U19697 (N_19697,N_19347,N_19425);
nor U19698 (N_19698,N_19079,N_19325);
nor U19699 (N_19699,N_19272,N_19041);
or U19700 (N_19700,N_19323,N_19232);
and U19701 (N_19701,N_19321,N_19132);
nor U19702 (N_19702,N_19470,N_19234);
nor U19703 (N_19703,N_19444,N_19345);
or U19704 (N_19704,N_19255,N_19453);
nor U19705 (N_19705,N_19127,N_19259);
and U19706 (N_19706,N_19489,N_19288);
and U19707 (N_19707,N_19082,N_19357);
and U19708 (N_19708,N_19075,N_19439);
and U19709 (N_19709,N_19283,N_19039);
nor U19710 (N_19710,N_19455,N_19242);
and U19711 (N_19711,N_19349,N_19448);
or U19712 (N_19712,N_19192,N_19279);
and U19713 (N_19713,N_19417,N_19352);
nor U19714 (N_19714,N_19427,N_19451);
xnor U19715 (N_19715,N_19198,N_19004);
and U19716 (N_19716,N_19203,N_19146);
nor U19717 (N_19717,N_19343,N_19380);
or U19718 (N_19718,N_19108,N_19406);
or U19719 (N_19719,N_19249,N_19003);
xor U19720 (N_19720,N_19094,N_19389);
nor U19721 (N_19721,N_19086,N_19336);
xnor U19722 (N_19722,N_19103,N_19499);
xnor U19723 (N_19723,N_19047,N_19311);
or U19724 (N_19724,N_19238,N_19297);
and U19725 (N_19725,N_19031,N_19292);
nand U19726 (N_19726,N_19008,N_19097);
and U19727 (N_19727,N_19165,N_19296);
or U19728 (N_19728,N_19359,N_19237);
nand U19729 (N_19729,N_19063,N_19220);
nand U19730 (N_19730,N_19298,N_19182);
nor U19731 (N_19731,N_19018,N_19353);
xor U19732 (N_19732,N_19320,N_19445);
xnor U19733 (N_19733,N_19011,N_19002);
and U19734 (N_19734,N_19107,N_19057);
and U19735 (N_19735,N_19282,N_19176);
nor U19736 (N_19736,N_19156,N_19143);
and U19737 (N_19737,N_19471,N_19474);
and U19738 (N_19738,N_19401,N_19157);
nor U19739 (N_19739,N_19053,N_19492);
or U19740 (N_19740,N_19286,N_19221);
and U19741 (N_19741,N_19329,N_19385);
or U19742 (N_19742,N_19248,N_19399);
nand U19743 (N_19743,N_19061,N_19281);
or U19744 (N_19744,N_19188,N_19098);
xor U19745 (N_19745,N_19178,N_19411);
and U19746 (N_19746,N_19014,N_19294);
and U19747 (N_19747,N_19449,N_19163);
xor U19748 (N_19748,N_19252,N_19388);
or U19749 (N_19749,N_19319,N_19354);
or U19750 (N_19750,N_19384,N_19272);
nand U19751 (N_19751,N_19328,N_19445);
or U19752 (N_19752,N_19426,N_19435);
nand U19753 (N_19753,N_19260,N_19024);
nor U19754 (N_19754,N_19491,N_19047);
and U19755 (N_19755,N_19251,N_19382);
and U19756 (N_19756,N_19307,N_19054);
xor U19757 (N_19757,N_19436,N_19170);
nand U19758 (N_19758,N_19473,N_19460);
nand U19759 (N_19759,N_19311,N_19076);
xnor U19760 (N_19760,N_19023,N_19092);
nor U19761 (N_19761,N_19002,N_19463);
or U19762 (N_19762,N_19089,N_19155);
nor U19763 (N_19763,N_19452,N_19181);
nor U19764 (N_19764,N_19314,N_19173);
nor U19765 (N_19765,N_19068,N_19386);
nand U19766 (N_19766,N_19203,N_19490);
nor U19767 (N_19767,N_19029,N_19113);
and U19768 (N_19768,N_19298,N_19215);
nor U19769 (N_19769,N_19346,N_19364);
and U19770 (N_19770,N_19417,N_19445);
nor U19771 (N_19771,N_19169,N_19290);
xnor U19772 (N_19772,N_19160,N_19375);
and U19773 (N_19773,N_19333,N_19114);
or U19774 (N_19774,N_19280,N_19362);
nor U19775 (N_19775,N_19341,N_19260);
and U19776 (N_19776,N_19090,N_19377);
nand U19777 (N_19777,N_19158,N_19018);
or U19778 (N_19778,N_19360,N_19319);
and U19779 (N_19779,N_19211,N_19022);
nor U19780 (N_19780,N_19419,N_19170);
xor U19781 (N_19781,N_19356,N_19016);
or U19782 (N_19782,N_19126,N_19262);
xor U19783 (N_19783,N_19306,N_19182);
nor U19784 (N_19784,N_19307,N_19019);
nor U19785 (N_19785,N_19406,N_19301);
xor U19786 (N_19786,N_19409,N_19230);
nor U19787 (N_19787,N_19011,N_19393);
and U19788 (N_19788,N_19404,N_19259);
xor U19789 (N_19789,N_19462,N_19480);
nand U19790 (N_19790,N_19148,N_19007);
nor U19791 (N_19791,N_19183,N_19260);
or U19792 (N_19792,N_19499,N_19488);
and U19793 (N_19793,N_19262,N_19001);
nor U19794 (N_19794,N_19487,N_19347);
xnor U19795 (N_19795,N_19086,N_19176);
or U19796 (N_19796,N_19329,N_19194);
or U19797 (N_19797,N_19095,N_19434);
or U19798 (N_19798,N_19177,N_19404);
xor U19799 (N_19799,N_19351,N_19434);
nor U19800 (N_19800,N_19277,N_19009);
or U19801 (N_19801,N_19068,N_19141);
or U19802 (N_19802,N_19313,N_19365);
or U19803 (N_19803,N_19394,N_19283);
xnor U19804 (N_19804,N_19132,N_19242);
or U19805 (N_19805,N_19125,N_19216);
nor U19806 (N_19806,N_19165,N_19131);
and U19807 (N_19807,N_19209,N_19059);
nor U19808 (N_19808,N_19117,N_19350);
or U19809 (N_19809,N_19271,N_19236);
xor U19810 (N_19810,N_19350,N_19220);
nand U19811 (N_19811,N_19334,N_19112);
and U19812 (N_19812,N_19215,N_19197);
xnor U19813 (N_19813,N_19312,N_19088);
nor U19814 (N_19814,N_19179,N_19338);
or U19815 (N_19815,N_19100,N_19004);
nand U19816 (N_19816,N_19069,N_19315);
nor U19817 (N_19817,N_19275,N_19129);
nand U19818 (N_19818,N_19010,N_19110);
nor U19819 (N_19819,N_19458,N_19367);
nor U19820 (N_19820,N_19179,N_19334);
or U19821 (N_19821,N_19429,N_19153);
and U19822 (N_19822,N_19381,N_19155);
and U19823 (N_19823,N_19320,N_19144);
and U19824 (N_19824,N_19390,N_19375);
or U19825 (N_19825,N_19210,N_19151);
xnor U19826 (N_19826,N_19426,N_19246);
or U19827 (N_19827,N_19054,N_19417);
nand U19828 (N_19828,N_19133,N_19057);
nand U19829 (N_19829,N_19482,N_19496);
or U19830 (N_19830,N_19269,N_19099);
nand U19831 (N_19831,N_19254,N_19164);
nor U19832 (N_19832,N_19469,N_19321);
or U19833 (N_19833,N_19011,N_19126);
or U19834 (N_19834,N_19029,N_19073);
or U19835 (N_19835,N_19416,N_19072);
and U19836 (N_19836,N_19305,N_19100);
or U19837 (N_19837,N_19387,N_19096);
nor U19838 (N_19838,N_19170,N_19213);
nand U19839 (N_19839,N_19043,N_19016);
or U19840 (N_19840,N_19224,N_19245);
xor U19841 (N_19841,N_19376,N_19454);
or U19842 (N_19842,N_19378,N_19450);
or U19843 (N_19843,N_19376,N_19442);
xnor U19844 (N_19844,N_19094,N_19452);
nand U19845 (N_19845,N_19390,N_19165);
or U19846 (N_19846,N_19210,N_19424);
nand U19847 (N_19847,N_19282,N_19077);
xnor U19848 (N_19848,N_19372,N_19157);
or U19849 (N_19849,N_19194,N_19086);
xor U19850 (N_19850,N_19453,N_19461);
xor U19851 (N_19851,N_19339,N_19315);
or U19852 (N_19852,N_19262,N_19278);
nor U19853 (N_19853,N_19337,N_19438);
nand U19854 (N_19854,N_19440,N_19028);
and U19855 (N_19855,N_19258,N_19493);
or U19856 (N_19856,N_19285,N_19011);
and U19857 (N_19857,N_19297,N_19472);
and U19858 (N_19858,N_19331,N_19028);
or U19859 (N_19859,N_19307,N_19241);
xor U19860 (N_19860,N_19072,N_19107);
nor U19861 (N_19861,N_19251,N_19469);
or U19862 (N_19862,N_19309,N_19379);
and U19863 (N_19863,N_19300,N_19364);
or U19864 (N_19864,N_19243,N_19441);
xor U19865 (N_19865,N_19382,N_19274);
nand U19866 (N_19866,N_19092,N_19255);
nor U19867 (N_19867,N_19137,N_19128);
nor U19868 (N_19868,N_19098,N_19002);
or U19869 (N_19869,N_19486,N_19341);
and U19870 (N_19870,N_19379,N_19429);
and U19871 (N_19871,N_19378,N_19350);
or U19872 (N_19872,N_19284,N_19421);
nor U19873 (N_19873,N_19471,N_19089);
xor U19874 (N_19874,N_19210,N_19308);
nor U19875 (N_19875,N_19355,N_19268);
and U19876 (N_19876,N_19329,N_19407);
or U19877 (N_19877,N_19252,N_19000);
and U19878 (N_19878,N_19208,N_19094);
and U19879 (N_19879,N_19285,N_19054);
xnor U19880 (N_19880,N_19140,N_19425);
nor U19881 (N_19881,N_19321,N_19113);
nor U19882 (N_19882,N_19397,N_19207);
and U19883 (N_19883,N_19110,N_19036);
and U19884 (N_19884,N_19448,N_19333);
nor U19885 (N_19885,N_19375,N_19399);
xnor U19886 (N_19886,N_19408,N_19126);
nor U19887 (N_19887,N_19017,N_19096);
and U19888 (N_19888,N_19061,N_19403);
nor U19889 (N_19889,N_19023,N_19132);
or U19890 (N_19890,N_19421,N_19038);
and U19891 (N_19891,N_19020,N_19111);
xor U19892 (N_19892,N_19433,N_19325);
and U19893 (N_19893,N_19338,N_19160);
xor U19894 (N_19894,N_19219,N_19018);
and U19895 (N_19895,N_19177,N_19389);
xnor U19896 (N_19896,N_19114,N_19167);
and U19897 (N_19897,N_19262,N_19037);
nand U19898 (N_19898,N_19328,N_19018);
xor U19899 (N_19899,N_19341,N_19342);
or U19900 (N_19900,N_19498,N_19018);
nand U19901 (N_19901,N_19397,N_19132);
nand U19902 (N_19902,N_19360,N_19446);
xor U19903 (N_19903,N_19472,N_19349);
xnor U19904 (N_19904,N_19164,N_19374);
xnor U19905 (N_19905,N_19244,N_19286);
xnor U19906 (N_19906,N_19063,N_19132);
nand U19907 (N_19907,N_19019,N_19024);
xor U19908 (N_19908,N_19401,N_19321);
xor U19909 (N_19909,N_19492,N_19207);
nand U19910 (N_19910,N_19423,N_19435);
xor U19911 (N_19911,N_19044,N_19150);
xor U19912 (N_19912,N_19498,N_19389);
nand U19913 (N_19913,N_19082,N_19148);
xnor U19914 (N_19914,N_19495,N_19325);
and U19915 (N_19915,N_19498,N_19479);
xor U19916 (N_19916,N_19138,N_19195);
and U19917 (N_19917,N_19023,N_19123);
nor U19918 (N_19918,N_19045,N_19274);
and U19919 (N_19919,N_19140,N_19041);
nand U19920 (N_19920,N_19013,N_19373);
nand U19921 (N_19921,N_19055,N_19220);
nand U19922 (N_19922,N_19050,N_19489);
and U19923 (N_19923,N_19278,N_19234);
or U19924 (N_19924,N_19101,N_19344);
xnor U19925 (N_19925,N_19070,N_19025);
nor U19926 (N_19926,N_19074,N_19262);
nor U19927 (N_19927,N_19193,N_19499);
nand U19928 (N_19928,N_19288,N_19024);
and U19929 (N_19929,N_19151,N_19059);
xor U19930 (N_19930,N_19350,N_19261);
or U19931 (N_19931,N_19137,N_19272);
or U19932 (N_19932,N_19348,N_19034);
nand U19933 (N_19933,N_19203,N_19237);
or U19934 (N_19934,N_19063,N_19247);
nand U19935 (N_19935,N_19320,N_19237);
nand U19936 (N_19936,N_19114,N_19499);
or U19937 (N_19937,N_19393,N_19458);
and U19938 (N_19938,N_19432,N_19274);
or U19939 (N_19939,N_19222,N_19267);
and U19940 (N_19940,N_19421,N_19301);
nand U19941 (N_19941,N_19435,N_19027);
nor U19942 (N_19942,N_19369,N_19013);
xnor U19943 (N_19943,N_19259,N_19482);
nand U19944 (N_19944,N_19305,N_19343);
and U19945 (N_19945,N_19366,N_19385);
and U19946 (N_19946,N_19291,N_19353);
nand U19947 (N_19947,N_19159,N_19128);
xnor U19948 (N_19948,N_19439,N_19424);
and U19949 (N_19949,N_19293,N_19244);
or U19950 (N_19950,N_19379,N_19408);
nor U19951 (N_19951,N_19083,N_19457);
xor U19952 (N_19952,N_19463,N_19050);
nand U19953 (N_19953,N_19373,N_19414);
or U19954 (N_19954,N_19015,N_19111);
xnor U19955 (N_19955,N_19319,N_19085);
nand U19956 (N_19956,N_19173,N_19115);
xnor U19957 (N_19957,N_19345,N_19199);
xor U19958 (N_19958,N_19065,N_19372);
nor U19959 (N_19959,N_19189,N_19180);
nor U19960 (N_19960,N_19007,N_19163);
nor U19961 (N_19961,N_19164,N_19210);
and U19962 (N_19962,N_19465,N_19265);
nand U19963 (N_19963,N_19295,N_19104);
xor U19964 (N_19964,N_19344,N_19391);
nand U19965 (N_19965,N_19131,N_19241);
or U19966 (N_19966,N_19145,N_19454);
nand U19967 (N_19967,N_19034,N_19210);
and U19968 (N_19968,N_19226,N_19371);
nand U19969 (N_19969,N_19292,N_19475);
xor U19970 (N_19970,N_19146,N_19422);
nand U19971 (N_19971,N_19375,N_19175);
nand U19972 (N_19972,N_19488,N_19482);
nor U19973 (N_19973,N_19194,N_19324);
or U19974 (N_19974,N_19457,N_19335);
nor U19975 (N_19975,N_19088,N_19021);
or U19976 (N_19976,N_19094,N_19035);
nor U19977 (N_19977,N_19219,N_19295);
or U19978 (N_19978,N_19399,N_19213);
or U19979 (N_19979,N_19028,N_19252);
or U19980 (N_19980,N_19012,N_19295);
or U19981 (N_19981,N_19108,N_19243);
or U19982 (N_19982,N_19217,N_19397);
nand U19983 (N_19983,N_19026,N_19466);
and U19984 (N_19984,N_19215,N_19067);
and U19985 (N_19985,N_19463,N_19172);
or U19986 (N_19986,N_19280,N_19176);
and U19987 (N_19987,N_19362,N_19139);
nor U19988 (N_19988,N_19082,N_19334);
or U19989 (N_19989,N_19484,N_19415);
nand U19990 (N_19990,N_19228,N_19136);
nor U19991 (N_19991,N_19063,N_19315);
xnor U19992 (N_19992,N_19107,N_19296);
or U19993 (N_19993,N_19130,N_19357);
xor U19994 (N_19994,N_19441,N_19309);
or U19995 (N_19995,N_19374,N_19467);
nand U19996 (N_19996,N_19472,N_19193);
nor U19997 (N_19997,N_19498,N_19115);
nand U19998 (N_19998,N_19029,N_19483);
and U19999 (N_19999,N_19237,N_19370);
xnor U20000 (N_20000,N_19902,N_19958);
and U20001 (N_20001,N_19562,N_19676);
nor U20002 (N_20002,N_19677,N_19758);
or U20003 (N_20003,N_19834,N_19573);
and U20004 (N_20004,N_19514,N_19895);
or U20005 (N_20005,N_19539,N_19766);
and U20006 (N_20006,N_19957,N_19976);
and U20007 (N_20007,N_19732,N_19774);
xnor U20008 (N_20008,N_19639,N_19692);
xnor U20009 (N_20009,N_19517,N_19810);
nand U20010 (N_20010,N_19821,N_19854);
xnor U20011 (N_20011,N_19859,N_19634);
xnor U20012 (N_20012,N_19883,N_19581);
and U20013 (N_20013,N_19734,N_19983);
and U20014 (N_20014,N_19722,N_19901);
xnor U20015 (N_20015,N_19953,N_19659);
nor U20016 (N_20016,N_19724,N_19877);
or U20017 (N_20017,N_19952,N_19597);
and U20018 (N_20018,N_19754,N_19599);
or U20019 (N_20019,N_19835,N_19625);
and U20020 (N_20020,N_19836,N_19658);
xor U20021 (N_20021,N_19663,N_19791);
or U20022 (N_20022,N_19665,N_19532);
nand U20023 (N_20023,N_19997,N_19762);
nand U20024 (N_20024,N_19930,N_19541);
nand U20025 (N_20025,N_19784,N_19623);
xnor U20026 (N_20026,N_19905,N_19660);
xnor U20027 (N_20027,N_19914,N_19556);
nor U20028 (N_20028,N_19986,N_19887);
xnor U20029 (N_20029,N_19501,N_19678);
nor U20030 (N_20030,N_19866,N_19988);
and U20031 (N_20031,N_19884,N_19654);
nor U20032 (N_20032,N_19857,N_19811);
xnor U20033 (N_20033,N_19743,N_19959);
nand U20034 (N_20034,N_19742,N_19805);
nor U20035 (N_20035,N_19981,N_19596);
nor U20036 (N_20036,N_19993,N_19941);
or U20037 (N_20037,N_19519,N_19750);
or U20038 (N_20038,N_19846,N_19703);
or U20039 (N_20039,N_19558,N_19649);
or U20040 (N_20040,N_19557,N_19951);
xor U20041 (N_20041,N_19644,N_19571);
xnor U20042 (N_20042,N_19603,N_19511);
or U20043 (N_20043,N_19925,N_19605);
xnor U20044 (N_20044,N_19527,N_19820);
xor U20045 (N_20045,N_19554,N_19777);
or U20046 (N_20046,N_19770,N_19506);
nor U20047 (N_20047,N_19622,N_19847);
xor U20048 (N_20048,N_19830,N_19994);
and U20049 (N_20049,N_19707,N_19672);
xor U20050 (N_20050,N_19587,N_19995);
and U20051 (N_20051,N_19827,N_19667);
xnor U20052 (N_20052,N_19538,N_19711);
nor U20053 (N_20053,N_19746,N_19792);
or U20054 (N_20054,N_19646,N_19787);
xor U20055 (N_20055,N_19651,N_19813);
xnor U20056 (N_20056,N_19693,N_19867);
and U20057 (N_20057,N_19619,N_19701);
or U20058 (N_20058,N_19864,N_19923);
or U20059 (N_20059,N_19900,N_19535);
nor U20060 (N_20060,N_19794,N_19829);
and U20061 (N_20061,N_19688,N_19697);
nor U20062 (N_20062,N_19522,N_19781);
xnor U20063 (N_20063,N_19868,N_19909);
nor U20064 (N_20064,N_19767,N_19826);
and U20065 (N_20065,N_19823,N_19698);
or U20066 (N_20066,N_19771,N_19968);
nor U20067 (N_20067,N_19938,N_19899);
xnor U20068 (N_20068,N_19718,N_19662);
xor U20069 (N_20069,N_19635,N_19642);
or U20070 (N_20070,N_19931,N_19531);
or U20071 (N_20071,N_19949,N_19509);
or U20072 (N_20072,N_19727,N_19956);
nor U20073 (N_20073,N_19790,N_19542);
and U20074 (N_20074,N_19566,N_19606);
nor U20075 (N_20075,N_19897,N_19533);
or U20076 (N_20076,N_19741,N_19926);
nor U20077 (N_20077,N_19521,N_19626);
and U20078 (N_20078,N_19604,N_19761);
xor U20079 (N_20079,N_19840,N_19789);
nand U20080 (N_20080,N_19575,N_19929);
nand U20081 (N_20081,N_19973,N_19728);
nand U20082 (N_20082,N_19713,N_19648);
or U20083 (N_20083,N_19806,N_19747);
xor U20084 (N_20084,N_19888,N_19875);
nand U20085 (N_20085,N_19675,N_19971);
nor U20086 (N_20086,N_19779,N_19674);
nor U20087 (N_20087,N_19681,N_19808);
nor U20088 (N_20088,N_19853,N_19963);
xnor U20089 (N_20089,N_19894,N_19611);
nor U20090 (N_20090,N_19920,N_19704);
nand U20091 (N_20091,N_19512,N_19600);
nand U20092 (N_20092,N_19881,N_19955);
or U20093 (N_20093,N_19749,N_19756);
nand U20094 (N_20094,N_19621,N_19543);
nand U20095 (N_20095,N_19560,N_19924);
or U20096 (N_20096,N_19755,N_19773);
xnor U20097 (N_20097,N_19680,N_19892);
nor U20098 (N_20098,N_19882,N_19970);
xnor U20099 (N_20099,N_19526,N_19588);
or U20100 (N_20100,N_19992,N_19975);
xor U20101 (N_20101,N_19637,N_19669);
xnor U20102 (N_20102,N_19712,N_19801);
nor U20103 (N_20103,N_19855,N_19860);
nor U20104 (N_20104,N_19870,N_19641);
or U20105 (N_20105,N_19736,N_19708);
and U20106 (N_20106,N_19977,N_19764);
and U20107 (N_20107,N_19843,N_19928);
nor U20108 (N_20108,N_19601,N_19943);
or U20109 (N_20109,N_19536,N_19776);
xor U20110 (N_20110,N_19880,N_19653);
nand U20111 (N_20111,N_19735,N_19919);
nand U20112 (N_20112,N_19763,N_19630);
nor U20113 (N_20113,N_19567,N_19620);
nand U20114 (N_20114,N_19798,N_19967);
xor U20115 (N_20115,N_19879,N_19765);
or U20116 (N_20116,N_19748,N_19624);
nor U20117 (N_20117,N_19803,N_19578);
nor U20118 (N_20118,N_19655,N_19799);
or U20119 (N_20119,N_19964,N_19709);
or U20120 (N_20120,N_19769,N_19702);
nor U20121 (N_20121,N_19515,N_19710);
nand U20122 (N_20122,N_19996,N_19516);
or U20123 (N_20123,N_19679,N_19500);
nor U20124 (N_20124,N_19807,N_19856);
nand U20125 (N_20125,N_19814,N_19796);
nand U20126 (N_20126,N_19972,N_19832);
xnor U20127 (N_20127,N_19922,N_19927);
or U20128 (N_20128,N_19590,N_19686);
nor U20129 (N_20129,N_19844,N_19910);
nand U20130 (N_20130,N_19589,N_19872);
nor U20131 (N_20131,N_19613,N_19917);
and U20132 (N_20132,N_19574,N_19906);
nand U20133 (N_20133,N_19569,N_19858);
or U20134 (N_20134,N_19645,N_19564);
nor U20135 (N_20135,N_19565,N_19802);
and U20136 (N_20136,N_19640,N_19775);
nor U20137 (N_20137,N_19759,N_19552);
xnor U20138 (N_20138,N_19961,N_19528);
and U20139 (N_20139,N_19607,N_19595);
and U20140 (N_20140,N_19948,N_19740);
nand U20141 (N_20141,N_19714,N_19682);
or U20142 (N_20142,N_19785,N_19842);
xor U20143 (N_20143,N_19852,N_19800);
or U20144 (N_20144,N_19598,N_19631);
nor U20145 (N_20145,N_19730,N_19824);
and U20146 (N_20146,N_19966,N_19699);
nand U20147 (N_20147,N_19544,N_19939);
nand U20148 (N_20148,N_19982,N_19591);
nand U20149 (N_20149,N_19638,N_19664);
xor U20150 (N_20150,N_19984,N_19614);
and U20151 (N_20151,N_19999,N_19523);
or U20152 (N_20152,N_19585,N_19944);
xnor U20153 (N_20153,N_19918,N_19726);
nand U20154 (N_20154,N_19768,N_19705);
nand U20155 (N_20155,N_19694,N_19804);
and U20156 (N_20156,N_19998,N_19954);
nor U20157 (N_20157,N_19783,N_19819);
xor U20158 (N_20158,N_19795,N_19723);
and U20159 (N_20159,N_19561,N_19793);
or U20160 (N_20160,N_19617,N_19991);
xor U20161 (N_20161,N_19507,N_19584);
and U20162 (N_20162,N_19563,N_19960);
and U20163 (N_20163,N_19862,N_19530);
nor U20164 (N_20164,N_19540,N_19890);
or U20165 (N_20165,N_19656,N_19729);
nor U20166 (N_20166,N_19513,N_19576);
and U20167 (N_20167,N_19594,N_19898);
nand U20168 (N_20168,N_19572,N_19738);
and U20169 (N_20169,N_19700,N_19885);
or U20170 (N_20170,N_19666,N_19979);
or U20171 (N_20171,N_19815,N_19609);
and U20172 (N_20172,N_19845,N_19912);
nand U20173 (N_20173,N_19618,N_19851);
nand U20174 (N_20174,N_19989,N_19889);
xor U20175 (N_20175,N_19610,N_19833);
and U20176 (N_20176,N_19850,N_19546);
and U20177 (N_20177,N_19745,N_19932);
nor U20178 (N_20178,N_19848,N_19627);
or U20179 (N_20179,N_19668,N_19706);
xnor U20180 (N_20180,N_19893,N_19782);
or U20181 (N_20181,N_19551,N_19524);
xor U20182 (N_20182,N_19871,N_19828);
nor U20183 (N_20183,N_19838,N_19822);
and U20184 (N_20184,N_19592,N_19933);
xor U20185 (N_20185,N_19636,N_19744);
and U20186 (N_20186,N_19553,N_19547);
or U20187 (N_20187,N_19583,N_19650);
nand U20188 (N_20188,N_19849,N_19643);
xnor U20189 (N_20189,N_19934,N_19896);
and U20190 (N_20190,N_19760,N_19962);
and U20191 (N_20191,N_19751,N_19737);
nor U20192 (N_20192,N_19690,N_19947);
and U20193 (N_20193,N_19670,N_19683);
and U20194 (N_20194,N_19725,N_19548);
nor U20195 (N_20195,N_19633,N_19689);
xnor U20196 (N_20196,N_19869,N_19969);
nand U20197 (N_20197,N_19831,N_19647);
nand U20198 (N_20198,N_19915,N_19980);
nor U20199 (N_20199,N_19570,N_19945);
xor U20200 (N_20200,N_19525,N_19720);
nand U20201 (N_20201,N_19753,N_19673);
xor U20202 (N_20202,N_19937,N_19502);
xor U20203 (N_20203,N_19579,N_19817);
nand U20204 (N_20204,N_19593,N_19687);
xnor U20205 (N_20205,N_19695,N_19685);
nor U20206 (N_20206,N_19778,N_19950);
xnor U20207 (N_20207,N_19752,N_19629);
or U20208 (N_20208,N_19978,N_19861);
nand U20209 (N_20209,N_19510,N_19555);
nand U20210 (N_20210,N_19508,N_19863);
and U20211 (N_20211,N_19550,N_19816);
nand U20212 (N_20212,N_19913,N_19797);
nand U20213 (N_20213,N_19615,N_19661);
nor U20214 (N_20214,N_19965,N_19757);
or U20215 (N_20215,N_19602,N_19908);
and U20216 (N_20216,N_19987,N_19586);
and U20217 (N_20217,N_19990,N_19721);
nor U20218 (N_20218,N_19549,N_19911);
xor U20219 (N_20219,N_19812,N_19534);
or U20220 (N_20220,N_19545,N_19628);
and U20221 (N_20221,N_19568,N_19520);
or U20222 (N_20222,N_19825,N_19772);
and U20223 (N_20223,N_19691,N_19935);
xnor U20224 (N_20224,N_19874,N_19657);
xor U20225 (N_20225,N_19907,N_19974);
nand U20226 (N_20226,N_19529,N_19878);
or U20227 (N_20227,N_19616,N_19839);
xor U20228 (N_20228,N_19886,N_19865);
nand U20229 (N_20229,N_19788,N_19559);
xnor U20230 (N_20230,N_19612,N_19891);
or U20231 (N_20231,N_19518,N_19731);
xnor U20232 (N_20232,N_19684,N_19916);
nor U20233 (N_20233,N_19580,N_19904);
nor U20234 (N_20234,N_19717,N_19537);
nor U20235 (N_20235,N_19505,N_19719);
xor U20236 (N_20236,N_19818,N_19837);
nor U20237 (N_20237,N_19841,N_19936);
or U20238 (N_20238,N_19632,N_19608);
nand U20239 (N_20239,N_19946,N_19809);
nor U20240 (N_20240,N_19921,N_19903);
and U20241 (N_20241,N_19577,N_19671);
xnor U20242 (N_20242,N_19503,N_19582);
nor U20243 (N_20243,N_19652,N_19504);
and U20244 (N_20244,N_19716,N_19873);
and U20245 (N_20245,N_19780,N_19985);
nand U20246 (N_20246,N_19696,N_19786);
xor U20247 (N_20247,N_19715,N_19876);
or U20248 (N_20248,N_19940,N_19733);
nor U20249 (N_20249,N_19942,N_19739);
or U20250 (N_20250,N_19629,N_19678);
xor U20251 (N_20251,N_19929,N_19918);
xnor U20252 (N_20252,N_19733,N_19509);
xnor U20253 (N_20253,N_19979,N_19521);
or U20254 (N_20254,N_19885,N_19610);
nand U20255 (N_20255,N_19651,N_19930);
and U20256 (N_20256,N_19642,N_19759);
xor U20257 (N_20257,N_19697,N_19642);
xnor U20258 (N_20258,N_19510,N_19892);
nor U20259 (N_20259,N_19549,N_19976);
and U20260 (N_20260,N_19725,N_19611);
xor U20261 (N_20261,N_19796,N_19606);
xnor U20262 (N_20262,N_19500,N_19636);
nand U20263 (N_20263,N_19847,N_19995);
and U20264 (N_20264,N_19802,N_19950);
and U20265 (N_20265,N_19614,N_19521);
nor U20266 (N_20266,N_19519,N_19585);
nor U20267 (N_20267,N_19683,N_19827);
and U20268 (N_20268,N_19592,N_19656);
nand U20269 (N_20269,N_19810,N_19818);
nand U20270 (N_20270,N_19513,N_19626);
xnor U20271 (N_20271,N_19947,N_19886);
nand U20272 (N_20272,N_19510,N_19532);
or U20273 (N_20273,N_19850,N_19727);
xor U20274 (N_20274,N_19577,N_19845);
nand U20275 (N_20275,N_19907,N_19779);
nand U20276 (N_20276,N_19979,N_19936);
and U20277 (N_20277,N_19972,N_19708);
nor U20278 (N_20278,N_19804,N_19864);
nor U20279 (N_20279,N_19799,N_19681);
nand U20280 (N_20280,N_19810,N_19831);
or U20281 (N_20281,N_19784,N_19753);
or U20282 (N_20282,N_19729,N_19722);
and U20283 (N_20283,N_19704,N_19763);
xnor U20284 (N_20284,N_19707,N_19786);
or U20285 (N_20285,N_19517,N_19817);
nor U20286 (N_20286,N_19701,N_19686);
xor U20287 (N_20287,N_19794,N_19807);
nand U20288 (N_20288,N_19613,N_19655);
xnor U20289 (N_20289,N_19963,N_19966);
and U20290 (N_20290,N_19833,N_19865);
or U20291 (N_20291,N_19658,N_19673);
nand U20292 (N_20292,N_19566,N_19653);
and U20293 (N_20293,N_19809,N_19986);
and U20294 (N_20294,N_19969,N_19839);
xnor U20295 (N_20295,N_19963,N_19553);
or U20296 (N_20296,N_19849,N_19689);
and U20297 (N_20297,N_19521,N_19956);
nand U20298 (N_20298,N_19806,N_19963);
nor U20299 (N_20299,N_19553,N_19500);
and U20300 (N_20300,N_19918,N_19949);
and U20301 (N_20301,N_19712,N_19612);
xnor U20302 (N_20302,N_19529,N_19887);
nand U20303 (N_20303,N_19835,N_19511);
nor U20304 (N_20304,N_19722,N_19657);
nor U20305 (N_20305,N_19804,N_19821);
nor U20306 (N_20306,N_19560,N_19669);
or U20307 (N_20307,N_19851,N_19819);
nor U20308 (N_20308,N_19850,N_19912);
nor U20309 (N_20309,N_19773,N_19885);
nor U20310 (N_20310,N_19801,N_19539);
or U20311 (N_20311,N_19661,N_19596);
xor U20312 (N_20312,N_19672,N_19585);
and U20313 (N_20313,N_19955,N_19931);
and U20314 (N_20314,N_19633,N_19834);
or U20315 (N_20315,N_19614,N_19873);
nand U20316 (N_20316,N_19676,N_19568);
or U20317 (N_20317,N_19638,N_19789);
nand U20318 (N_20318,N_19638,N_19797);
nand U20319 (N_20319,N_19763,N_19913);
or U20320 (N_20320,N_19573,N_19538);
xor U20321 (N_20321,N_19676,N_19864);
nor U20322 (N_20322,N_19675,N_19549);
or U20323 (N_20323,N_19888,N_19987);
and U20324 (N_20324,N_19500,N_19745);
or U20325 (N_20325,N_19939,N_19512);
nor U20326 (N_20326,N_19677,N_19643);
nor U20327 (N_20327,N_19858,N_19601);
nor U20328 (N_20328,N_19776,N_19755);
nand U20329 (N_20329,N_19654,N_19927);
or U20330 (N_20330,N_19651,N_19583);
nand U20331 (N_20331,N_19802,N_19676);
nand U20332 (N_20332,N_19900,N_19996);
nand U20333 (N_20333,N_19617,N_19622);
and U20334 (N_20334,N_19898,N_19683);
xor U20335 (N_20335,N_19592,N_19906);
or U20336 (N_20336,N_19910,N_19615);
and U20337 (N_20337,N_19895,N_19957);
xnor U20338 (N_20338,N_19904,N_19618);
nor U20339 (N_20339,N_19924,N_19867);
nor U20340 (N_20340,N_19958,N_19777);
or U20341 (N_20341,N_19525,N_19876);
xnor U20342 (N_20342,N_19621,N_19823);
nor U20343 (N_20343,N_19887,N_19736);
nand U20344 (N_20344,N_19624,N_19825);
nand U20345 (N_20345,N_19743,N_19843);
nor U20346 (N_20346,N_19537,N_19626);
nand U20347 (N_20347,N_19658,N_19945);
nand U20348 (N_20348,N_19732,N_19890);
nand U20349 (N_20349,N_19685,N_19633);
nand U20350 (N_20350,N_19984,N_19923);
xor U20351 (N_20351,N_19595,N_19873);
nand U20352 (N_20352,N_19592,N_19665);
and U20353 (N_20353,N_19715,N_19844);
nor U20354 (N_20354,N_19894,N_19656);
nor U20355 (N_20355,N_19663,N_19994);
xor U20356 (N_20356,N_19895,N_19999);
nor U20357 (N_20357,N_19715,N_19918);
nor U20358 (N_20358,N_19576,N_19664);
xnor U20359 (N_20359,N_19930,N_19607);
nor U20360 (N_20360,N_19676,N_19792);
and U20361 (N_20361,N_19635,N_19688);
nor U20362 (N_20362,N_19532,N_19845);
nand U20363 (N_20363,N_19687,N_19666);
and U20364 (N_20364,N_19809,N_19854);
or U20365 (N_20365,N_19716,N_19897);
nor U20366 (N_20366,N_19961,N_19939);
and U20367 (N_20367,N_19986,N_19758);
nor U20368 (N_20368,N_19906,N_19864);
and U20369 (N_20369,N_19551,N_19813);
xor U20370 (N_20370,N_19761,N_19864);
and U20371 (N_20371,N_19763,N_19919);
xor U20372 (N_20372,N_19909,N_19996);
or U20373 (N_20373,N_19973,N_19552);
or U20374 (N_20374,N_19991,N_19649);
nor U20375 (N_20375,N_19577,N_19717);
nor U20376 (N_20376,N_19535,N_19855);
and U20377 (N_20377,N_19933,N_19886);
or U20378 (N_20378,N_19903,N_19969);
or U20379 (N_20379,N_19583,N_19728);
and U20380 (N_20380,N_19655,N_19693);
nor U20381 (N_20381,N_19505,N_19778);
xnor U20382 (N_20382,N_19511,N_19640);
and U20383 (N_20383,N_19919,N_19581);
nand U20384 (N_20384,N_19593,N_19618);
or U20385 (N_20385,N_19847,N_19853);
nand U20386 (N_20386,N_19971,N_19953);
nor U20387 (N_20387,N_19729,N_19736);
and U20388 (N_20388,N_19626,N_19807);
and U20389 (N_20389,N_19619,N_19770);
xor U20390 (N_20390,N_19682,N_19550);
or U20391 (N_20391,N_19901,N_19605);
nand U20392 (N_20392,N_19841,N_19740);
xor U20393 (N_20393,N_19767,N_19639);
and U20394 (N_20394,N_19805,N_19574);
nor U20395 (N_20395,N_19693,N_19509);
and U20396 (N_20396,N_19943,N_19810);
nand U20397 (N_20397,N_19880,N_19796);
or U20398 (N_20398,N_19812,N_19593);
and U20399 (N_20399,N_19529,N_19507);
xor U20400 (N_20400,N_19743,N_19597);
nor U20401 (N_20401,N_19733,N_19638);
xnor U20402 (N_20402,N_19994,N_19556);
nand U20403 (N_20403,N_19733,N_19997);
xnor U20404 (N_20404,N_19703,N_19771);
xnor U20405 (N_20405,N_19581,N_19750);
nand U20406 (N_20406,N_19797,N_19965);
xor U20407 (N_20407,N_19889,N_19891);
xor U20408 (N_20408,N_19802,N_19972);
or U20409 (N_20409,N_19666,N_19533);
and U20410 (N_20410,N_19932,N_19824);
xor U20411 (N_20411,N_19546,N_19733);
nand U20412 (N_20412,N_19512,N_19760);
nor U20413 (N_20413,N_19558,N_19900);
nand U20414 (N_20414,N_19535,N_19880);
or U20415 (N_20415,N_19661,N_19721);
nand U20416 (N_20416,N_19871,N_19882);
nor U20417 (N_20417,N_19836,N_19702);
or U20418 (N_20418,N_19619,N_19970);
nand U20419 (N_20419,N_19877,N_19810);
xnor U20420 (N_20420,N_19918,N_19866);
xor U20421 (N_20421,N_19870,N_19780);
nor U20422 (N_20422,N_19620,N_19858);
or U20423 (N_20423,N_19550,N_19637);
nand U20424 (N_20424,N_19602,N_19749);
or U20425 (N_20425,N_19997,N_19513);
or U20426 (N_20426,N_19767,N_19828);
nor U20427 (N_20427,N_19944,N_19738);
nand U20428 (N_20428,N_19574,N_19780);
and U20429 (N_20429,N_19714,N_19529);
xnor U20430 (N_20430,N_19838,N_19947);
nor U20431 (N_20431,N_19651,N_19831);
or U20432 (N_20432,N_19771,N_19922);
or U20433 (N_20433,N_19998,N_19734);
xor U20434 (N_20434,N_19942,N_19678);
nor U20435 (N_20435,N_19538,N_19832);
xor U20436 (N_20436,N_19874,N_19993);
and U20437 (N_20437,N_19623,N_19964);
and U20438 (N_20438,N_19547,N_19873);
xor U20439 (N_20439,N_19651,N_19869);
and U20440 (N_20440,N_19788,N_19856);
xnor U20441 (N_20441,N_19873,N_19804);
and U20442 (N_20442,N_19542,N_19535);
nand U20443 (N_20443,N_19960,N_19897);
and U20444 (N_20444,N_19756,N_19668);
and U20445 (N_20445,N_19978,N_19614);
and U20446 (N_20446,N_19509,N_19916);
and U20447 (N_20447,N_19943,N_19730);
and U20448 (N_20448,N_19695,N_19607);
nand U20449 (N_20449,N_19808,N_19887);
nand U20450 (N_20450,N_19745,N_19875);
xnor U20451 (N_20451,N_19761,N_19888);
nand U20452 (N_20452,N_19670,N_19850);
xor U20453 (N_20453,N_19959,N_19740);
xnor U20454 (N_20454,N_19858,N_19629);
and U20455 (N_20455,N_19749,N_19643);
or U20456 (N_20456,N_19658,N_19892);
nor U20457 (N_20457,N_19760,N_19630);
nor U20458 (N_20458,N_19653,N_19639);
or U20459 (N_20459,N_19832,N_19611);
and U20460 (N_20460,N_19980,N_19581);
xnor U20461 (N_20461,N_19873,N_19609);
xor U20462 (N_20462,N_19503,N_19989);
nand U20463 (N_20463,N_19538,N_19530);
nor U20464 (N_20464,N_19861,N_19649);
nor U20465 (N_20465,N_19831,N_19821);
nor U20466 (N_20466,N_19888,N_19606);
or U20467 (N_20467,N_19875,N_19774);
or U20468 (N_20468,N_19929,N_19619);
xnor U20469 (N_20469,N_19638,N_19811);
and U20470 (N_20470,N_19741,N_19959);
nand U20471 (N_20471,N_19626,N_19588);
nor U20472 (N_20472,N_19790,N_19610);
nor U20473 (N_20473,N_19864,N_19685);
and U20474 (N_20474,N_19890,N_19761);
xnor U20475 (N_20475,N_19709,N_19926);
or U20476 (N_20476,N_19981,N_19916);
nor U20477 (N_20477,N_19519,N_19803);
and U20478 (N_20478,N_19677,N_19985);
nand U20479 (N_20479,N_19564,N_19968);
nand U20480 (N_20480,N_19551,N_19839);
xor U20481 (N_20481,N_19508,N_19672);
and U20482 (N_20482,N_19787,N_19692);
nor U20483 (N_20483,N_19708,N_19902);
and U20484 (N_20484,N_19599,N_19562);
and U20485 (N_20485,N_19747,N_19768);
xor U20486 (N_20486,N_19846,N_19923);
and U20487 (N_20487,N_19780,N_19783);
xnor U20488 (N_20488,N_19543,N_19860);
nand U20489 (N_20489,N_19659,N_19580);
and U20490 (N_20490,N_19708,N_19567);
or U20491 (N_20491,N_19973,N_19763);
nor U20492 (N_20492,N_19986,N_19572);
xnor U20493 (N_20493,N_19583,N_19544);
xnor U20494 (N_20494,N_19505,N_19998);
xor U20495 (N_20495,N_19850,N_19612);
nand U20496 (N_20496,N_19550,N_19955);
nor U20497 (N_20497,N_19546,N_19539);
or U20498 (N_20498,N_19647,N_19902);
or U20499 (N_20499,N_19804,N_19716);
xor U20500 (N_20500,N_20244,N_20099);
xnor U20501 (N_20501,N_20154,N_20181);
nor U20502 (N_20502,N_20016,N_20261);
and U20503 (N_20503,N_20073,N_20416);
nand U20504 (N_20504,N_20380,N_20323);
or U20505 (N_20505,N_20036,N_20101);
xor U20506 (N_20506,N_20375,N_20346);
and U20507 (N_20507,N_20300,N_20234);
nand U20508 (N_20508,N_20427,N_20498);
or U20509 (N_20509,N_20053,N_20199);
and U20510 (N_20510,N_20390,N_20340);
nand U20511 (N_20511,N_20492,N_20172);
nand U20512 (N_20512,N_20135,N_20272);
xor U20513 (N_20513,N_20339,N_20382);
nand U20514 (N_20514,N_20214,N_20267);
xor U20515 (N_20515,N_20469,N_20421);
and U20516 (N_20516,N_20289,N_20413);
and U20517 (N_20517,N_20170,N_20160);
nor U20518 (N_20518,N_20259,N_20495);
xnor U20519 (N_20519,N_20316,N_20330);
nand U20520 (N_20520,N_20002,N_20363);
nor U20521 (N_20521,N_20046,N_20301);
nand U20522 (N_20522,N_20317,N_20168);
nor U20523 (N_20523,N_20219,N_20364);
xnor U20524 (N_20524,N_20249,N_20019);
and U20525 (N_20525,N_20367,N_20422);
nand U20526 (N_20526,N_20470,N_20408);
and U20527 (N_20527,N_20158,N_20447);
xor U20528 (N_20528,N_20049,N_20353);
or U20529 (N_20529,N_20263,N_20361);
and U20530 (N_20530,N_20403,N_20109);
and U20531 (N_20531,N_20349,N_20133);
nor U20532 (N_20532,N_20186,N_20277);
or U20533 (N_20533,N_20295,N_20080);
xnor U20534 (N_20534,N_20155,N_20430);
or U20535 (N_20535,N_20185,N_20088);
or U20536 (N_20536,N_20079,N_20078);
nor U20537 (N_20537,N_20038,N_20428);
nor U20538 (N_20538,N_20011,N_20311);
and U20539 (N_20539,N_20396,N_20494);
nor U20540 (N_20540,N_20001,N_20313);
and U20541 (N_20541,N_20114,N_20411);
or U20542 (N_20542,N_20304,N_20076);
or U20543 (N_20543,N_20452,N_20017);
xor U20544 (N_20544,N_20122,N_20281);
xor U20545 (N_20545,N_20128,N_20373);
xor U20546 (N_20546,N_20347,N_20478);
and U20547 (N_20547,N_20387,N_20131);
nand U20548 (N_20548,N_20153,N_20342);
nor U20549 (N_20549,N_20055,N_20488);
and U20550 (N_20550,N_20283,N_20298);
nor U20551 (N_20551,N_20231,N_20303);
nor U20552 (N_20552,N_20052,N_20041);
xnor U20553 (N_20553,N_20444,N_20265);
xor U20554 (N_20554,N_20013,N_20365);
xor U20555 (N_20555,N_20003,N_20157);
nor U20556 (N_20556,N_20381,N_20030);
xor U20557 (N_20557,N_20140,N_20275);
nor U20558 (N_20558,N_20391,N_20480);
and U20559 (N_20559,N_20207,N_20351);
or U20560 (N_20560,N_20412,N_20360);
nor U20561 (N_20561,N_20215,N_20376);
nor U20562 (N_20562,N_20178,N_20338);
nor U20563 (N_20563,N_20383,N_20393);
nand U20564 (N_20564,N_20320,N_20443);
xor U20565 (N_20565,N_20130,N_20042);
nor U20566 (N_20566,N_20167,N_20315);
nor U20567 (N_20567,N_20230,N_20125);
or U20568 (N_20568,N_20461,N_20032);
xor U20569 (N_20569,N_20145,N_20481);
and U20570 (N_20570,N_20379,N_20266);
nor U20571 (N_20571,N_20448,N_20308);
nand U20572 (N_20572,N_20009,N_20476);
or U20573 (N_20573,N_20108,N_20081);
nand U20574 (N_20574,N_20063,N_20325);
nand U20575 (N_20575,N_20483,N_20424);
nor U20576 (N_20576,N_20247,N_20243);
xnor U20577 (N_20577,N_20465,N_20450);
or U20578 (N_20578,N_20152,N_20429);
nand U20579 (N_20579,N_20439,N_20256);
xor U20580 (N_20580,N_20150,N_20056);
xor U20581 (N_20581,N_20296,N_20310);
or U20582 (N_20582,N_20290,N_20314);
nand U20583 (N_20583,N_20193,N_20358);
nor U20584 (N_20584,N_20064,N_20190);
nand U20585 (N_20585,N_20293,N_20202);
nor U20586 (N_20586,N_20400,N_20472);
xnor U20587 (N_20587,N_20370,N_20224);
nor U20588 (N_20588,N_20020,N_20348);
xor U20589 (N_20589,N_20218,N_20405);
nand U20590 (N_20590,N_20180,N_20018);
nor U20591 (N_20591,N_20384,N_20297);
or U20592 (N_20592,N_20216,N_20333);
xnor U20593 (N_20593,N_20033,N_20414);
nand U20594 (N_20594,N_20321,N_20060);
nand U20595 (N_20595,N_20149,N_20175);
nand U20596 (N_20596,N_20022,N_20473);
nand U20597 (N_20597,N_20436,N_20209);
xor U20598 (N_20598,N_20305,N_20139);
nor U20599 (N_20599,N_20229,N_20355);
nand U20600 (N_20600,N_20112,N_20394);
or U20601 (N_20601,N_20051,N_20402);
xnor U20602 (N_20602,N_20146,N_20235);
nor U20603 (N_20603,N_20457,N_20071);
xor U20604 (N_20604,N_20415,N_20183);
and U20605 (N_20605,N_20006,N_20499);
nor U20606 (N_20606,N_20327,N_20100);
xor U20607 (N_20607,N_20121,N_20095);
nor U20608 (N_20608,N_20169,N_20189);
and U20609 (N_20609,N_20442,N_20466);
or U20610 (N_20610,N_20262,N_20204);
and U20611 (N_20611,N_20120,N_20144);
nor U20612 (N_20612,N_20392,N_20226);
nor U20613 (N_20613,N_20270,N_20491);
and U20614 (N_20614,N_20048,N_20377);
nor U20615 (N_20615,N_20291,N_20035);
and U20616 (N_20616,N_20312,N_20433);
nand U20617 (N_20617,N_20386,N_20251);
xnor U20618 (N_20618,N_20434,N_20280);
and U20619 (N_20619,N_20047,N_20107);
and U20620 (N_20620,N_20082,N_20176);
nor U20621 (N_20621,N_20399,N_20104);
nor U20622 (N_20622,N_20138,N_20102);
and U20623 (N_20623,N_20287,N_20192);
and U20624 (N_20624,N_20173,N_20273);
nor U20625 (N_20625,N_20084,N_20083);
nor U20626 (N_20626,N_20407,N_20015);
nor U20627 (N_20627,N_20097,N_20123);
nand U20628 (N_20628,N_20012,N_20236);
nor U20629 (N_20629,N_20197,N_20057);
nor U20630 (N_20630,N_20490,N_20220);
xnor U20631 (N_20631,N_20369,N_20137);
and U20632 (N_20632,N_20184,N_20334);
xnor U20633 (N_20633,N_20441,N_20050);
xor U20634 (N_20634,N_20043,N_20420);
and U20635 (N_20635,N_20151,N_20241);
nand U20636 (N_20636,N_20067,N_20092);
xor U20637 (N_20637,N_20451,N_20200);
or U20638 (N_20638,N_20037,N_20459);
nor U20639 (N_20639,N_20171,N_20061);
nand U20640 (N_20640,N_20484,N_20028);
nand U20641 (N_20641,N_20460,N_20425);
and U20642 (N_20642,N_20350,N_20014);
and U20643 (N_20643,N_20212,N_20054);
xor U20644 (N_20644,N_20000,N_20217);
or U20645 (N_20645,N_20040,N_20468);
xnor U20646 (N_20646,N_20482,N_20010);
xor U20647 (N_20647,N_20438,N_20397);
xor U20648 (N_20648,N_20039,N_20326);
and U20649 (N_20649,N_20253,N_20329);
xnor U20650 (N_20650,N_20142,N_20113);
and U20651 (N_20651,N_20177,N_20237);
nor U20652 (N_20652,N_20248,N_20242);
or U20653 (N_20653,N_20264,N_20258);
nand U20654 (N_20654,N_20260,N_20410);
nor U20655 (N_20655,N_20257,N_20398);
or U20656 (N_20656,N_20233,N_20074);
nor U20657 (N_20657,N_20023,N_20285);
xnor U20658 (N_20658,N_20453,N_20194);
xor U20659 (N_20659,N_20423,N_20005);
xor U20660 (N_20660,N_20066,N_20129);
nand U20661 (N_20661,N_20045,N_20401);
xor U20662 (N_20662,N_20034,N_20222);
nand U20663 (N_20663,N_20201,N_20362);
or U20664 (N_20664,N_20206,N_20232);
nand U20665 (N_20665,N_20331,N_20458);
or U20666 (N_20666,N_20126,N_20250);
xnor U20667 (N_20667,N_20025,N_20007);
nand U20668 (N_20668,N_20366,N_20419);
and U20669 (N_20669,N_20276,N_20077);
nand U20670 (N_20670,N_20115,N_20445);
nand U20671 (N_20671,N_20162,N_20440);
and U20672 (N_20672,N_20096,N_20464);
or U20673 (N_20673,N_20294,N_20328);
or U20674 (N_20674,N_20134,N_20307);
nor U20675 (N_20675,N_20116,N_20198);
and U20676 (N_20676,N_20161,N_20119);
nor U20677 (N_20677,N_20409,N_20343);
and U20678 (N_20678,N_20069,N_20004);
and U20679 (N_20679,N_20371,N_20163);
and U20680 (N_20680,N_20378,N_20106);
nand U20681 (N_20681,N_20021,N_20467);
nor U20682 (N_20682,N_20487,N_20136);
nand U20683 (N_20683,N_20085,N_20024);
or U20684 (N_20684,N_20098,N_20255);
xnor U20685 (N_20685,N_20179,N_20345);
nand U20686 (N_20686,N_20324,N_20164);
or U20687 (N_20687,N_20431,N_20240);
xnor U20688 (N_20688,N_20059,N_20026);
xnor U20689 (N_20689,N_20065,N_20279);
nor U20690 (N_20690,N_20404,N_20463);
nor U20691 (N_20691,N_20159,N_20132);
xor U20692 (N_20692,N_20332,N_20174);
xnor U20693 (N_20693,N_20417,N_20309);
or U20694 (N_20694,N_20124,N_20356);
nor U20695 (N_20695,N_20027,N_20357);
and U20696 (N_20696,N_20489,N_20486);
nor U20697 (N_20697,N_20446,N_20406);
nor U20698 (N_20698,N_20493,N_20389);
xor U20699 (N_20699,N_20372,N_20288);
xor U20700 (N_20700,N_20426,N_20418);
or U20701 (N_20701,N_20091,N_20354);
or U20702 (N_20702,N_20008,N_20319);
xor U20703 (N_20703,N_20252,N_20395);
nor U20704 (N_20704,N_20117,N_20455);
or U20705 (N_20705,N_20166,N_20435);
xnor U20706 (N_20706,N_20147,N_20368);
and U20707 (N_20707,N_20485,N_20286);
or U20708 (N_20708,N_20211,N_20268);
nor U20709 (N_20709,N_20187,N_20182);
or U20710 (N_20710,N_20070,N_20062);
and U20711 (N_20711,N_20437,N_20497);
and U20712 (N_20712,N_20225,N_20118);
or U20713 (N_20713,N_20474,N_20031);
and U20714 (N_20714,N_20110,N_20087);
nor U20715 (N_20715,N_20322,N_20352);
nand U20716 (N_20716,N_20221,N_20210);
or U20717 (N_20717,N_20246,N_20385);
and U20718 (N_20718,N_20302,N_20086);
or U20719 (N_20719,N_20245,N_20284);
nand U20720 (N_20720,N_20359,N_20228);
nor U20721 (N_20721,N_20075,N_20292);
nand U20722 (N_20722,N_20271,N_20254);
nand U20723 (N_20723,N_20094,N_20223);
nand U20724 (N_20724,N_20089,N_20374);
nor U20725 (N_20725,N_20156,N_20227);
nand U20726 (N_20726,N_20205,N_20068);
xor U20727 (N_20727,N_20456,N_20341);
nand U20728 (N_20728,N_20195,N_20306);
and U20729 (N_20729,N_20238,N_20188);
xor U20730 (N_20730,N_20165,N_20475);
xnor U20731 (N_20731,N_20213,N_20274);
and U20732 (N_20732,N_20044,N_20479);
xor U20733 (N_20733,N_20335,N_20191);
and U20734 (N_20734,N_20449,N_20127);
nor U20735 (N_20735,N_20148,N_20462);
or U20736 (N_20736,N_20029,N_20203);
or U20737 (N_20737,N_20282,N_20471);
or U20738 (N_20738,N_20093,N_20477);
or U20739 (N_20739,N_20103,N_20090);
xnor U20740 (N_20740,N_20196,N_20299);
xor U20741 (N_20741,N_20432,N_20072);
or U20742 (N_20742,N_20388,N_20111);
and U20743 (N_20743,N_20454,N_20239);
nor U20744 (N_20744,N_20058,N_20105);
xnor U20745 (N_20745,N_20278,N_20337);
and U20746 (N_20746,N_20336,N_20143);
or U20747 (N_20747,N_20496,N_20344);
xnor U20748 (N_20748,N_20318,N_20208);
and U20749 (N_20749,N_20141,N_20269);
or U20750 (N_20750,N_20048,N_20282);
nand U20751 (N_20751,N_20285,N_20024);
nand U20752 (N_20752,N_20301,N_20314);
nor U20753 (N_20753,N_20385,N_20086);
or U20754 (N_20754,N_20285,N_20174);
or U20755 (N_20755,N_20224,N_20177);
or U20756 (N_20756,N_20322,N_20025);
nand U20757 (N_20757,N_20232,N_20335);
xnor U20758 (N_20758,N_20257,N_20406);
or U20759 (N_20759,N_20402,N_20319);
nor U20760 (N_20760,N_20289,N_20165);
and U20761 (N_20761,N_20449,N_20046);
xnor U20762 (N_20762,N_20445,N_20272);
xor U20763 (N_20763,N_20045,N_20380);
or U20764 (N_20764,N_20133,N_20421);
or U20765 (N_20765,N_20373,N_20466);
and U20766 (N_20766,N_20457,N_20173);
and U20767 (N_20767,N_20309,N_20256);
and U20768 (N_20768,N_20268,N_20431);
and U20769 (N_20769,N_20492,N_20075);
xnor U20770 (N_20770,N_20491,N_20292);
or U20771 (N_20771,N_20445,N_20192);
or U20772 (N_20772,N_20308,N_20276);
nor U20773 (N_20773,N_20323,N_20438);
nand U20774 (N_20774,N_20437,N_20142);
nor U20775 (N_20775,N_20186,N_20056);
and U20776 (N_20776,N_20065,N_20324);
or U20777 (N_20777,N_20183,N_20250);
and U20778 (N_20778,N_20359,N_20485);
or U20779 (N_20779,N_20206,N_20084);
nor U20780 (N_20780,N_20220,N_20447);
or U20781 (N_20781,N_20290,N_20010);
xnor U20782 (N_20782,N_20437,N_20457);
nand U20783 (N_20783,N_20136,N_20475);
nor U20784 (N_20784,N_20486,N_20346);
and U20785 (N_20785,N_20424,N_20380);
or U20786 (N_20786,N_20285,N_20094);
nor U20787 (N_20787,N_20156,N_20464);
xor U20788 (N_20788,N_20437,N_20116);
and U20789 (N_20789,N_20209,N_20044);
or U20790 (N_20790,N_20030,N_20457);
nor U20791 (N_20791,N_20149,N_20127);
xnor U20792 (N_20792,N_20075,N_20413);
and U20793 (N_20793,N_20383,N_20074);
nor U20794 (N_20794,N_20261,N_20381);
nor U20795 (N_20795,N_20211,N_20488);
nand U20796 (N_20796,N_20362,N_20136);
nand U20797 (N_20797,N_20490,N_20232);
or U20798 (N_20798,N_20317,N_20393);
nor U20799 (N_20799,N_20310,N_20157);
nor U20800 (N_20800,N_20039,N_20005);
xor U20801 (N_20801,N_20221,N_20282);
and U20802 (N_20802,N_20170,N_20331);
nor U20803 (N_20803,N_20337,N_20348);
xnor U20804 (N_20804,N_20148,N_20201);
or U20805 (N_20805,N_20048,N_20111);
or U20806 (N_20806,N_20197,N_20140);
or U20807 (N_20807,N_20334,N_20258);
and U20808 (N_20808,N_20344,N_20233);
or U20809 (N_20809,N_20054,N_20366);
and U20810 (N_20810,N_20034,N_20255);
or U20811 (N_20811,N_20273,N_20274);
nor U20812 (N_20812,N_20190,N_20357);
xor U20813 (N_20813,N_20160,N_20250);
or U20814 (N_20814,N_20464,N_20088);
nand U20815 (N_20815,N_20398,N_20197);
nand U20816 (N_20816,N_20050,N_20323);
xnor U20817 (N_20817,N_20298,N_20070);
nand U20818 (N_20818,N_20486,N_20482);
nand U20819 (N_20819,N_20287,N_20304);
and U20820 (N_20820,N_20296,N_20430);
xor U20821 (N_20821,N_20184,N_20287);
nor U20822 (N_20822,N_20267,N_20242);
and U20823 (N_20823,N_20446,N_20194);
xnor U20824 (N_20824,N_20078,N_20019);
or U20825 (N_20825,N_20013,N_20100);
xor U20826 (N_20826,N_20199,N_20449);
nor U20827 (N_20827,N_20330,N_20222);
or U20828 (N_20828,N_20169,N_20335);
or U20829 (N_20829,N_20376,N_20270);
nand U20830 (N_20830,N_20347,N_20442);
nor U20831 (N_20831,N_20313,N_20076);
nand U20832 (N_20832,N_20176,N_20043);
or U20833 (N_20833,N_20436,N_20340);
xnor U20834 (N_20834,N_20338,N_20329);
and U20835 (N_20835,N_20279,N_20312);
nor U20836 (N_20836,N_20195,N_20359);
nand U20837 (N_20837,N_20242,N_20466);
or U20838 (N_20838,N_20097,N_20422);
nand U20839 (N_20839,N_20146,N_20442);
and U20840 (N_20840,N_20106,N_20041);
nand U20841 (N_20841,N_20170,N_20105);
and U20842 (N_20842,N_20413,N_20381);
nor U20843 (N_20843,N_20433,N_20070);
nand U20844 (N_20844,N_20336,N_20008);
or U20845 (N_20845,N_20362,N_20038);
xnor U20846 (N_20846,N_20225,N_20206);
or U20847 (N_20847,N_20308,N_20477);
and U20848 (N_20848,N_20127,N_20308);
nor U20849 (N_20849,N_20292,N_20177);
and U20850 (N_20850,N_20263,N_20334);
nand U20851 (N_20851,N_20372,N_20012);
xor U20852 (N_20852,N_20494,N_20144);
nor U20853 (N_20853,N_20327,N_20283);
and U20854 (N_20854,N_20090,N_20427);
or U20855 (N_20855,N_20371,N_20161);
nor U20856 (N_20856,N_20157,N_20286);
nand U20857 (N_20857,N_20461,N_20046);
xor U20858 (N_20858,N_20033,N_20367);
xor U20859 (N_20859,N_20116,N_20067);
xnor U20860 (N_20860,N_20450,N_20274);
and U20861 (N_20861,N_20234,N_20268);
xor U20862 (N_20862,N_20339,N_20410);
nor U20863 (N_20863,N_20286,N_20359);
xnor U20864 (N_20864,N_20003,N_20333);
nand U20865 (N_20865,N_20370,N_20226);
xnor U20866 (N_20866,N_20456,N_20243);
xor U20867 (N_20867,N_20179,N_20461);
nor U20868 (N_20868,N_20039,N_20471);
xnor U20869 (N_20869,N_20222,N_20395);
xnor U20870 (N_20870,N_20049,N_20087);
xor U20871 (N_20871,N_20022,N_20456);
nor U20872 (N_20872,N_20499,N_20215);
nand U20873 (N_20873,N_20192,N_20067);
nand U20874 (N_20874,N_20338,N_20256);
or U20875 (N_20875,N_20478,N_20121);
nand U20876 (N_20876,N_20357,N_20054);
nand U20877 (N_20877,N_20278,N_20045);
or U20878 (N_20878,N_20452,N_20342);
and U20879 (N_20879,N_20447,N_20451);
nand U20880 (N_20880,N_20414,N_20208);
nand U20881 (N_20881,N_20198,N_20173);
and U20882 (N_20882,N_20075,N_20090);
or U20883 (N_20883,N_20130,N_20000);
or U20884 (N_20884,N_20258,N_20407);
nor U20885 (N_20885,N_20399,N_20419);
or U20886 (N_20886,N_20345,N_20356);
or U20887 (N_20887,N_20482,N_20025);
xor U20888 (N_20888,N_20118,N_20424);
and U20889 (N_20889,N_20067,N_20193);
nor U20890 (N_20890,N_20030,N_20467);
nand U20891 (N_20891,N_20138,N_20013);
or U20892 (N_20892,N_20223,N_20267);
or U20893 (N_20893,N_20137,N_20061);
and U20894 (N_20894,N_20067,N_20168);
xor U20895 (N_20895,N_20133,N_20366);
and U20896 (N_20896,N_20016,N_20308);
nor U20897 (N_20897,N_20224,N_20169);
xnor U20898 (N_20898,N_20293,N_20064);
nand U20899 (N_20899,N_20472,N_20345);
and U20900 (N_20900,N_20411,N_20133);
nand U20901 (N_20901,N_20172,N_20384);
or U20902 (N_20902,N_20030,N_20220);
xor U20903 (N_20903,N_20150,N_20070);
xor U20904 (N_20904,N_20454,N_20034);
xor U20905 (N_20905,N_20379,N_20276);
and U20906 (N_20906,N_20279,N_20154);
or U20907 (N_20907,N_20368,N_20465);
xnor U20908 (N_20908,N_20128,N_20389);
nor U20909 (N_20909,N_20387,N_20206);
and U20910 (N_20910,N_20318,N_20071);
xnor U20911 (N_20911,N_20189,N_20175);
or U20912 (N_20912,N_20393,N_20301);
and U20913 (N_20913,N_20253,N_20240);
or U20914 (N_20914,N_20288,N_20462);
or U20915 (N_20915,N_20174,N_20016);
or U20916 (N_20916,N_20236,N_20227);
nand U20917 (N_20917,N_20168,N_20489);
xnor U20918 (N_20918,N_20048,N_20356);
xnor U20919 (N_20919,N_20128,N_20105);
xnor U20920 (N_20920,N_20081,N_20383);
nor U20921 (N_20921,N_20200,N_20131);
and U20922 (N_20922,N_20463,N_20214);
or U20923 (N_20923,N_20225,N_20005);
and U20924 (N_20924,N_20372,N_20138);
and U20925 (N_20925,N_20138,N_20133);
nor U20926 (N_20926,N_20105,N_20323);
and U20927 (N_20927,N_20330,N_20125);
xor U20928 (N_20928,N_20220,N_20469);
nor U20929 (N_20929,N_20177,N_20405);
xnor U20930 (N_20930,N_20316,N_20096);
nand U20931 (N_20931,N_20243,N_20337);
xor U20932 (N_20932,N_20242,N_20027);
and U20933 (N_20933,N_20158,N_20220);
nand U20934 (N_20934,N_20423,N_20322);
xor U20935 (N_20935,N_20146,N_20485);
and U20936 (N_20936,N_20324,N_20493);
nand U20937 (N_20937,N_20463,N_20461);
or U20938 (N_20938,N_20066,N_20401);
and U20939 (N_20939,N_20222,N_20466);
nor U20940 (N_20940,N_20128,N_20375);
nand U20941 (N_20941,N_20480,N_20213);
and U20942 (N_20942,N_20400,N_20466);
nor U20943 (N_20943,N_20397,N_20127);
nor U20944 (N_20944,N_20169,N_20495);
nor U20945 (N_20945,N_20246,N_20343);
or U20946 (N_20946,N_20089,N_20261);
or U20947 (N_20947,N_20316,N_20468);
nand U20948 (N_20948,N_20407,N_20450);
and U20949 (N_20949,N_20111,N_20442);
and U20950 (N_20950,N_20418,N_20458);
xnor U20951 (N_20951,N_20254,N_20182);
nor U20952 (N_20952,N_20074,N_20227);
and U20953 (N_20953,N_20392,N_20234);
xnor U20954 (N_20954,N_20141,N_20461);
xor U20955 (N_20955,N_20380,N_20097);
and U20956 (N_20956,N_20231,N_20200);
nand U20957 (N_20957,N_20271,N_20395);
or U20958 (N_20958,N_20481,N_20415);
or U20959 (N_20959,N_20425,N_20251);
nor U20960 (N_20960,N_20133,N_20452);
or U20961 (N_20961,N_20136,N_20196);
or U20962 (N_20962,N_20159,N_20349);
xnor U20963 (N_20963,N_20004,N_20481);
or U20964 (N_20964,N_20181,N_20009);
nor U20965 (N_20965,N_20361,N_20275);
xor U20966 (N_20966,N_20280,N_20219);
or U20967 (N_20967,N_20079,N_20495);
xor U20968 (N_20968,N_20438,N_20147);
xnor U20969 (N_20969,N_20008,N_20441);
or U20970 (N_20970,N_20210,N_20134);
xor U20971 (N_20971,N_20052,N_20048);
and U20972 (N_20972,N_20013,N_20473);
xor U20973 (N_20973,N_20438,N_20050);
nand U20974 (N_20974,N_20276,N_20436);
or U20975 (N_20975,N_20451,N_20150);
or U20976 (N_20976,N_20184,N_20068);
and U20977 (N_20977,N_20469,N_20066);
and U20978 (N_20978,N_20461,N_20194);
or U20979 (N_20979,N_20102,N_20282);
xor U20980 (N_20980,N_20464,N_20082);
and U20981 (N_20981,N_20003,N_20249);
nor U20982 (N_20982,N_20139,N_20191);
nand U20983 (N_20983,N_20443,N_20111);
and U20984 (N_20984,N_20290,N_20286);
nand U20985 (N_20985,N_20034,N_20000);
nor U20986 (N_20986,N_20455,N_20259);
nand U20987 (N_20987,N_20115,N_20287);
nor U20988 (N_20988,N_20119,N_20110);
or U20989 (N_20989,N_20002,N_20223);
xor U20990 (N_20990,N_20332,N_20494);
nand U20991 (N_20991,N_20383,N_20474);
nor U20992 (N_20992,N_20230,N_20027);
nand U20993 (N_20993,N_20149,N_20441);
nor U20994 (N_20994,N_20038,N_20019);
nor U20995 (N_20995,N_20179,N_20358);
and U20996 (N_20996,N_20113,N_20257);
and U20997 (N_20997,N_20258,N_20462);
nor U20998 (N_20998,N_20147,N_20154);
nor U20999 (N_20999,N_20392,N_20379);
or U21000 (N_21000,N_20668,N_20678);
xor U21001 (N_21001,N_20955,N_20980);
or U21002 (N_21002,N_20610,N_20797);
nor U21003 (N_21003,N_20694,N_20585);
nor U21004 (N_21004,N_20855,N_20744);
xnor U21005 (N_21005,N_20530,N_20594);
and U21006 (N_21006,N_20776,N_20836);
or U21007 (N_21007,N_20539,N_20501);
nor U21008 (N_21008,N_20718,N_20684);
nor U21009 (N_21009,N_20764,N_20541);
xnor U21010 (N_21010,N_20620,N_20937);
and U21011 (N_21011,N_20535,N_20760);
nand U21012 (N_21012,N_20935,N_20833);
or U21013 (N_21013,N_20766,N_20685);
and U21014 (N_21014,N_20743,N_20555);
and U21015 (N_21015,N_20954,N_20985);
or U21016 (N_21016,N_20640,N_20564);
xnor U21017 (N_21017,N_20506,N_20545);
nand U21018 (N_21018,N_20952,N_20697);
nor U21019 (N_21019,N_20941,N_20614);
and U21020 (N_21020,N_20732,N_20831);
nor U21021 (N_21021,N_20580,N_20523);
nand U21022 (N_21022,N_20706,N_20522);
and U21023 (N_21023,N_20988,N_20548);
or U21024 (N_21024,N_20778,N_20606);
nand U21025 (N_21025,N_20999,N_20786);
xor U21026 (N_21026,N_20784,N_20666);
xnor U21027 (N_21027,N_20550,N_20802);
nor U21028 (N_21028,N_20559,N_20696);
nor U21029 (N_21029,N_20869,N_20946);
xor U21030 (N_21030,N_20630,N_20865);
nand U21031 (N_21031,N_20707,N_20572);
and U21032 (N_21032,N_20656,N_20790);
or U21033 (N_21033,N_20793,N_20789);
or U21034 (N_21034,N_20513,N_20839);
nor U21035 (N_21035,N_20834,N_20502);
nor U21036 (N_21036,N_20906,N_20704);
nor U21037 (N_21037,N_20714,N_20623);
or U21038 (N_21038,N_20611,N_20651);
xnor U21039 (N_21039,N_20960,N_20867);
nand U21040 (N_21040,N_20810,N_20991);
nor U21041 (N_21041,N_20526,N_20818);
and U21042 (N_21042,N_20726,N_20882);
nand U21043 (N_21043,N_20889,N_20801);
nand U21044 (N_21044,N_20687,N_20729);
or U21045 (N_21045,N_20929,N_20756);
nand U21046 (N_21046,N_20864,N_20986);
and U21047 (N_21047,N_20528,N_20939);
or U21048 (N_21048,N_20637,N_20984);
nand U21049 (N_21049,N_20874,N_20771);
or U21050 (N_21050,N_20933,N_20908);
or U21051 (N_21051,N_20748,N_20910);
and U21052 (N_21052,N_20827,N_20967);
or U21053 (N_21053,N_20773,N_20716);
xor U21054 (N_21054,N_20622,N_20664);
nor U21055 (N_21055,N_20949,N_20569);
nand U21056 (N_21056,N_20676,N_20537);
nor U21057 (N_21057,N_20521,N_20560);
xnor U21058 (N_21058,N_20953,N_20888);
nand U21059 (N_21059,N_20901,N_20853);
nand U21060 (N_21060,N_20915,N_20677);
nor U21061 (N_21061,N_20875,N_20657);
or U21062 (N_21062,N_20883,N_20824);
or U21063 (N_21063,N_20780,N_20503);
or U21064 (N_21064,N_20708,N_20540);
xnor U21065 (N_21065,N_20552,N_20649);
xor U21066 (N_21066,N_20663,N_20631);
xor U21067 (N_21067,N_20820,N_20507);
nand U21068 (N_21068,N_20994,N_20543);
xor U21069 (N_21069,N_20782,N_20893);
xor U21070 (N_21070,N_20654,N_20921);
nor U21071 (N_21071,N_20533,N_20500);
xnor U21072 (N_21072,N_20602,N_20742);
nand U21073 (N_21073,N_20795,N_20570);
and U21074 (N_21074,N_20926,N_20917);
nor U21075 (N_21075,N_20922,N_20591);
nor U21076 (N_21076,N_20613,N_20816);
nand U21077 (N_21077,N_20761,N_20616);
nand U21078 (N_21078,N_20813,N_20531);
or U21079 (N_21079,N_20730,N_20860);
and U21080 (N_21080,N_20607,N_20811);
nand U21081 (N_21081,N_20873,N_20675);
nor U21082 (N_21082,N_20823,N_20819);
and U21083 (N_21083,N_20632,N_20871);
nor U21084 (N_21084,N_20852,N_20951);
and U21085 (N_21085,N_20596,N_20931);
nor U21086 (N_21086,N_20592,N_20700);
nand U21087 (N_21087,N_20798,N_20775);
or U21088 (N_21088,N_20720,N_20682);
and U21089 (N_21089,N_20588,N_20963);
nand U21090 (N_21090,N_20642,N_20599);
nand U21091 (N_21091,N_20803,N_20619);
xnor U21092 (N_21092,N_20787,N_20680);
nand U21093 (N_21093,N_20876,N_20887);
and U21094 (N_21094,N_20753,N_20805);
nand U21095 (N_21095,N_20898,N_20574);
or U21096 (N_21096,N_20738,N_20538);
nor U21097 (N_21097,N_20907,N_20942);
and U21098 (N_21098,N_20512,N_20995);
xnor U21099 (N_21099,N_20544,N_20920);
nor U21100 (N_21100,N_20699,N_20733);
or U21101 (N_21101,N_20943,N_20737);
nand U21102 (N_21102,N_20542,N_20950);
or U21103 (N_21103,N_20968,N_20624);
and U21104 (N_21104,N_20520,N_20653);
and U21105 (N_21105,N_20551,N_20938);
or U21106 (N_21106,N_20846,N_20665);
xnor U21107 (N_21107,N_20768,N_20878);
nor U21108 (N_21108,N_20964,N_20711);
nor U21109 (N_21109,N_20600,N_20740);
nor U21110 (N_21110,N_20703,N_20830);
nand U21111 (N_21111,N_20840,N_20752);
and U21112 (N_21112,N_20576,N_20604);
nand U21113 (N_21113,N_20884,N_20828);
and U21114 (N_21114,N_20826,N_20965);
nand U21115 (N_21115,N_20791,N_20639);
nand U21116 (N_21116,N_20769,N_20959);
xor U21117 (N_21117,N_20681,N_20598);
nor U21118 (N_21118,N_20625,N_20977);
nand U21119 (N_21119,N_20851,N_20731);
nand U21120 (N_21120,N_20587,N_20843);
nor U21121 (N_21121,N_20809,N_20723);
and U21122 (N_21122,N_20563,N_20897);
nand U21123 (N_21123,N_20772,N_20998);
nand U21124 (N_21124,N_20796,N_20902);
and U21125 (N_21125,N_20962,N_20577);
nor U21126 (N_21126,N_20629,N_20751);
xnor U21127 (N_21127,N_20847,N_20862);
nand U21128 (N_21128,N_20721,N_20845);
or U21129 (N_21129,N_20932,N_20854);
or U21130 (N_21130,N_20568,N_20745);
xnor U21131 (N_21131,N_20841,N_20618);
or U21132 (N_21132,N_20844,N_20975);
nor U21133 (N_21133,N_20635,N_20701);
xnor U21134 (N_21134,N_20832,N_20573);
nand U21135 (N_21135,N_20688,N_20895);
nor U21136 (N_21136,N_20891,N_20582);
xor U21137 (N_21137,N_20662,N_20849);
or U21138 (N_21138,N_20728,N_20689);
and U21139 (N_21139,N_20800,N_20961);
or U21140 (N_21140,N_20597,N_20669);
xor U21141 (N_21141,N_20583,N_20736);
or U21142 (N_21142,N_20777,N_20658);
or U21143 (N_21143,N_20590,N_20673);
and U21144 (N_21144,N_20892,N_20627);
xnor U21145 (N_21145,N_20970,N_20822);
nand U21146 (N_21146,N_20628,N_20674);
nand U21147 (N_21147,N_20948,N_20866);
nor U21148 (N_21148,N_20947,N_20562);
nand U21149 (N_21149,N_20659,N_20525);
and U21150 (N_21150,N_20990,N_20636);
and U21151 (N_21151,N_20508,N_20527);
and U21152 (N_21152,N_20930,N_20925);
nor U21153 (N_21153,N_20992,N_20617);
and U21154 (N_21154,N_20971,N_20989);
nand U21155 (N_21155,N_20958,N_20671);
xor U21156 (N_21156,N_20670,N_20561);
or U21157 (N_21157,N_20595,N_20554);
xor U21158 (N_21158,N_20638,N_20812);
xnor U21159 (N_21159,N_20750,N_20565);
xor U21160 (N_21160,N_20660,N_20692);
or U21161 (N_21161,N_20605,N_20940);
and U21162 (N_21162,N_20927,N_20710);
nand U21163 (N_21163,N_20579,N_20698);
and U21164 (N_21164,N_20792,N_20667);
and U21165 (N_21165,N_20837,N_20806);
and U21166 (N_21166,N_20633,N_20709);
nor U21167 (N_21167,N_20783,N_20919);
nand U21168 (N_21168,N_20886,N_20974);
or U21169 (N_21169,N_20762,N_20848);
and U21170 (N_21170,N_20652,N_20510);
and U21171 (N_21171,N_20749,N_20880);
nand U21172 (N_21172,N_20646,N_20976);
or U21173 (N_21173,N_20566,N_20835);
xor U21174 (N_21174,N_20532,N_20996);
nor U21175 (N_21175,N_20615,N_20993);
xor U21176 (N_21176,N_20702,N_20896);
nand U21177 (N_21177,N_20767,N_20578);
nor U21178 (N_21178,N_20717,N_20524);
nand U21179 (N_21179,N_20912,N_20825);
nand U21180 (N_21180,N_20584,N_20982);
nor U21181 (N_21181,N_20807,N_20557);
or U21182 (N_21182,N_20739,N_20850);
or U21183 (N_21183,N_20799,N_20957);
and U21184 (N_21184,N_20546,N_20722);
or U21185 (N_21185,N_20788,N_20881);
nor U21186 (N_21186,N_20785,N_20981);
and U21187 (N_21187,N_20804,N_20567);
or U21188 (N_21188,N_20504,N_20944);
nor U21189 (N_21189,N_20724,N_20911);
xor U21190 (N_21190,N_20536,N_20894);
or U21191 (N_21191,N_20734,N_20549);
xor U21192 (N_21192,N_20603,N_20859);
and U21193 (N_21193,N_20586,N_20719);
xor U21194 (N_21194,N_20956,N_20774);
nor U21195 (N_21195,N_20519,N_20885);
xor U21196 (N_21196,N_20621,N_20899);
or U21197 (N_21197,N_20683,N_20715);
or U21198 (N_21198,N_20695,N_20593);
nand U21199 (N_21199,N_20969,N_20972);
and U21200 (N_21200,N_20529,N_20808);
and U21201 (N_21201,N_20817,N_20781);
and U21202 (N_21202,N_20755,N_20765);
and U21203 (N_21203,N_20547,N_20713);
nand U21204 (N_21204,N_20746,N_20966);
or U21205 (N_21205,N_20754,N_20691);
or U21206 (N_21206,N_20979,N_20918);
or U21207 (N_21207,N_20829,N_20641);
or U21208 (N_21208,N_20903,N_20648);
and U21209 (N_21209,N_20936,N_20747);
nand U21210 (N_21210,N_20644,N_20838);
or U21211 (N_21211,N_20857,N_20913);
or U21212 (N_21212,N_20877,N_20870);
and U21213 (N_21213,N_20924,N_20517);
nor U21214 (N_21214,N_20900,N_20815);
nor U21215 (N_21215,N_20909,N_20686);
nand U21216 (N_21216,N_20505,N_20916);
or U21217 (N_21217,N_20608,N_20589);
and U21218 (N_21218,N_20905,N_20770);
nor U21219 (N_21219,N_20856,N_20609);
or U21220 (N_21220,N_20712,N_20690);
or U21221 (N_21221,N_20553,N_20741);
nor U21222 (N_21222,N_20647,N_20779);
and U21223 (N_21223,N_20518,N_20534);
xor U21224 (N_21224,N_20987,N_20928);
nor U21225 (N_21225,N_20872,N_20556);
nand U21226 (N_21226,N_20879,N_20868);
and U21227 (N_21227,N_20842,N_20904);
or U21228 (N_21228,N_20558,N_20923);
nor U21229 (N_21229,N_20645,N_20516);
nor U21230 (N_21230,N_20758,N_20727);
or U21231 (N_21231,N_20705,N_20575);
nand U21232 (N_21232,N_20763,N_20601);
and U21233 (N_21233,N_20759,N_20997);
nor U21234 (N_21234,N_20634,N_20581);
xor U21235 (N_21235,N_20794,N_20983);
and U21236 (N_21236,N_20571,N_20511);
nand U21237 (N_21237,N_20626,N_20757);
xnor U21238 (N_21238,N_20973,N_20679);
nand U21239 (N_21239,N_20858,N_20509);
nand U21240 (N_21240,N_20693,N_20914);
nand U21241 (N_21241,N_20514,N_20735);
or U21242 (N_21242,N_20821,N_20725);
xor U21243 (N_21243,N_20890,N_20612);
xor U21244 (N_21244,N_20861,N_20672);
xor U21245 (N_21245,N_20661,N_20978);
xnor U21246 (N_21246,N_20814,N_20650);
and U21247 (N_21247,N_20863,N_20934);
nand U21248 (N_21248,N_20655,N_20945);
xor U21249 (N_21249,N_20515,N_20643);
nor U21250 (N_21250,N_20785,N_20730);
nor U21251 (N_21251,N_20763,N_20701);
xor U21252 (N_21252,N_20880,N_20814);
and U21253 (N_21253,N_20642,N_20540);
nand U21254 (N_21254,N_20543,N_20961);
nor U21255 (N_21255,N_20515,N_20772);
nand U21256 (N_21256,N_20997,N_20817);
nand U21257 (N_21257,N_20535,N_20753);
and U21258 (N_21258,N_20648,N_20885);
and U21259 (N_21259,N_20623,N_20907);
and U21260 (N_21260,N_20631,N_20861);
nor U21261 (N_21261,N_20886,N_20633);
nand U21262 (N_21262,N_20835,N_20562);
xnor U21263 (N_21263,N_20710,N_20918);
and U21264 (N_21264,N_20726,N_20694);
nor U21265 (N_21265,N_20590,N_20756);
nor U21266 (N_21266,N_20767,N_20635);
xnor U21267 (N_21267,N_20649,N_20838);
or U21268 (N_21268,N_20809,N_20885);
and U21269 (N_21269,N_20672,N_20961);
nand U21270 (N_21270,N_20902,N_20901);
nand U21271 (N_21271,N_20980,N_20887);
and U21272 (N_21272,N_20855,N_20525);
nand U21273 (N_21273,N_20636,N_20843);
and U21274 (N_21274,N_20688,N_20843);
or U21275 (N_21275,N_20607,N_20804);
nor U21276 (N_21276,N_20740,N_20811);
nor U21277 (N_21277,N_20873,N_20593);
xor U21278 (N_21278,N_20799,N_20728);
or U21279 (N_21279,N_20570,N_20755);
nor U21280 (N_21280,N_20776,N_20693);
nor U21281 (N_21281,N_20632,N_20997);
and U21282 (N_21282,N_20505,N_20722);
nand U21283 (N_21283,N_20784,N_20663);
or U21284 (N_21284,N_20686,N_20941);
or U21285 (N_21285,N_20593,N_20992);
or U21286 (N_21286,N_20636,N_20936);
or U21287 (N_21287,N_20715,N_20718);
nand U21288 (N_21288,N_20741,N_20727);
and U21289 (N_21289,N_20747,N_20781);
or U21290 (N_21290,N_20645,N_20949);
or U21291 (N_21291,N_20849,N_20760);
or U21292 (N_21292,N_20920,N_20750);
nor U21293 (N_21293,N_20853,N_20858);
nor U21294 (N_21294,N_20997,N_20565);
and U21295 (N_21295,N_20885,N_20902);
and U21296 (N_21296,N_20719,N_20931);
xnor U21297 (N_21297,N_20955,N_20584);
xor U21298 (N_21298,N_20842,N_20772);
nor U21299 (N_21299,N_20683,N_20553);
or U21300 (N_21300,N_20655,N_20723);
nand U21301 (N_21301,N_20815,N_20693);
xor U21302 (N_21302,N_20896,N_20634);
xor U21303 (N_21303,N_20821,N_20696);
nor U21304 (N_21304,N_20868,N_20522);
nor U21305 (N_21305,N_20695,N_20990);
xnor U21306 (N_21306,N_20801,N_20823);
xnor U21307 (N_21307,N_20931,N_20516);
and U21308 (N_21308,N_20528,N_20678);
or U21309 (N_21309,N_20976,N_20968);
and U21310 (N_21310,N_20952,N_20516);
nand U21311 (N_21311,N_20534,N_20958);
or U21312 (N_21312,N_20754,N_20893);
and U21313 (N_21313,N_20986,N_20723);
nor U21314 (N_21314,N_20711,N_20987);
xor U21315 (N_21315,N_20535,N_20748);
xnor U21316 (N_21316,N_20772,N_20605);
nand U21317 (N_21317,N_20573,N_20687);
xor U21318 (N_21318,N_20932,N_20961);
or U21319 (N_21319,N_20842,N_20869);
nand U21320 (N_21320,N_20848,N_20623);
nand U21321 (N_21321,N_20557,N_20722);
nor U21322 (N_21322,N_20748,N_20930);
nand U21323 (N_21323,N_20975,N_20776);
or U21324 (N_21324,N_20782,N_20967);
or U21325 (N_21325,N_20938,N_20806);
or U21326 (N_21326,N_20893,N_20664);
xnor U21327 (N_21327,N_20982,N_20693);
xor U21328 (N_21328,N_20744,N_20752);
nand U21329 (N_21329,N_20743,N_20516);
and U21330 (N_21330,N_20975,N_20976);
nand U21331 (N_21331,N_20578,N_20900);
xor U21332 (N_21332,N_20542,N_20729);
and U21333 (N_21333,N_20515,N_20770);
xnor U21334 (N_21334,N_20774,N_20621);
or U21335 (N_21335,N_20533,N_20978);
xnor U21336 (N_21336,N_20658,N_20557);
xor U21337 (N_21337,N_20593,N_20931);
xor U21338 (N_21338,N_20630,N_20526);
or U21339 (N_21339,N_20959,N_20636);
or U21340 (N_21340,N_20624,N_20588);
or U21341 (N_21341,N_20703,N_20998);
nor U21342 (N_21342,N_20713,N_20752);
or U21343 (N_21343,N_20841,N_20617);
and U21344 (N_21344,N_20673,N_20700);
xor U21345 (N_21345,N_20640,N_20577);
and U21346 (N_21346,N_20614,N_20718);
nor U21347 (N_21347,N_20535,N_20582);
and U21348 (N_21348,N_20692,N_20715);
nand U21349 (N_21349,N_20630,N_20584);
or U21350 (N_21350,N_20602,N_20992);
xor U21351 (N_21351,N_20710,N_20522);
nand U21352 (N_21352,N_20767,N_20756);
nand U21353 (N_21353,N_20650,N_20839);
or U21354 (N_21354,N_20539,N_20667);
or U21355 (N_21355,N_20927,N_20835);
nand U21356 (N_21356,N_20830,N_20587);
xor U21357 (N_21357,N_20645,N_20618);
or U21358 (N_21358,N_20932,N_20907);
nand U21359 (N_21359,N_20878,N_20606);
nor U21360 (N_21360,N_20854,N_20608);
and U21361 (N_21361,N_20728,N_20825);
and U21362 (N_21362,N_20994,N_20956);
nand U21363 (N_21363,N_20589,N_20667);
nor U21364 (N_21364,N_20901,N_20756);
or U21365 (N_21365,N_20512,N_20557);
nand U21366 (N_21366,N_20826,N_20767);
or U21367 (N_21367,N_20739,N_20682);
nand U21368 (N_21368,N_20878,N_20686);
and U21369 (N_21369,N_20984,N_20888);
nor U21370 (N_21370,N_20645,N_20584);
nand U21371 (N_21371,N_20563,N_20556);
and U21372 (N_21372,N_20549,N_20937);
or U21373 (N_21373,N_20540,N_20777);
nor U21374 (N_21374,N_20685,N_20932);
nand U21375 (N_21375,N_20750,N_20754);
nor U21376 (N_21376,N_20518,N_20769);
xnor U21377 (N_21377,N_20624,N_20931);
nand U21378 (N_21378,N_20500,N_20623);
or U21379 (N_21379,N_20651,N_20902);
and U21380 (N_21380,N_20534,N_20501);
nor U21381 (N_21381,N_20983,N_20776);
and U21382 (N_21382,N_20570,N_20597);
and U21383 (N_21383,N_20652,N_20623);
nor U21384 (N_21384,N_20585,N_20967);
and U21385 (N_21385,N_20680,N_20786);
xor U21386 (N_21386,N_20600,N_20717);
xor U21387 (N_21387,N_20526,N_20873);
xor U21388 (N_21388,N_20527,N_20885);
and U21389 (N_21389,N_20669,N_20877);
and U21390 (N_21390,N_20715,N_20950);
xor U21391 (N_21391,N_20854,N_20578);
nor U21392 (N_21392,N_20966,N_20964);
xnor U21393 (N_21393,N_20873,N_20869);
and U21394 (N_21394,N_20806,N_20654);
and U21395 (N_21395,N_20547,N_20748);
xor U21396 (N_21396,N_20732,N_20730);
or U21397 (N_21397,N_20850,N_20756);
and U21398 (N_21398,N_20594,N_20699);
nand U21399 (N_21399,N_20820,N_20515);
and U21400 (N_21400,N_20713,N_20962);
or U21401 (N_21401,N_20665,N_20521);
or U21402 (N_21402,N_20549,N_20755);
and U21403 (N_21403,N_20764,N_20720);
xor U21404 (N_21404,N_20946,N_20814);
nand U21405 (N_21405,N_20722,N_20789);
nor U21406 (N_21406,N_20619,N_20889);
and U21407 (N_21407,N_20905,N_20956);
or U21408 (N_21408,N_20675,N_20636);
xor U21409 (N_21409,N_20605,N_20692);
xor U21410 (N_21410,N_20671,N_20762);
nand U21411 (N_21411,N_20568,N_20755);
nor U21412 (N_21412,N_20766,N_20695);
xnor U21413 (N_21413,N_20779,N_20577);
nor U21414 (N_21414,N_20685,N_20563);
or U21415 (N_21415,N_20684,N_20637);
and U21416 (N_21416,N_20510,N_20632);
or U21417 (N_21417,N_20717,N_20988);
or U21418 (N_21418,N_20695,N_20636);
nand U21419 (N_21419,N_20737,N_20789);
and U21420 (N_21420,N_20975,N_20918);
xnor U21421 (N_21421,N_20874,N_20992);
or U21422 (N_21422,N_20839,N_20591);
or U21423 (N_21423,N_20806,N_20812);
and U21424 (N_21424,N_20602,N_20889);
and U21425 (N_21425,N_20868,N_20950);
or U21426 (N_21426,N_20783,N_20595);
nor U21427 (N_21427,N_20738,N_20639);
and U21428 (N_21428,N_20868,N_20997);
xnor U21429 (N_21429,N_20594,N_20723);
and U21430 (N_21430,N_20661,N_20502);
nand U21431 (N_21431,N_20924,N_20729);
nand U21432 (N_21432,N_20579,N_20860);
nor U21433 (N_21433,N_20725,N_20967);
or U21434 (N_21434,N_20595,N_20769);
nand U21435 (N_21435,N_20739,N_20700);
or U21436 (N_21436,N_20820,N_20852);
and U21437 (N_21437,N_20805,N_20748);
nand U21438 (N_21438,N_20695,N_20619);
nor U21439 (N_21439,N_20712,N_20689);
nor U21440 (N_21440,N_20601,N_20748);
or U21441 (N_21441,N_20717,N_20609);
and U21442 (N_21442,N_20765,N_20963);
xor U21443 (N_21443,N_20802,N_20662);
xnor U21444 (N_21444,N_20800,N_20830);
nor U21445 (N_21445,N_20696,N_20845);
and U21446 (N_21446,N_20564,N_20649);
xnor U21447 (N_21447,N_20911,N_20843);
nand U21448 (N_21448,N_20938,N_20845);
or U21449 (N_21449,N_20756,N_20963);
xnor U21450 (N_21450,N_20922,N_20910);
or U21451 (N_21451,N_20727,N_20792);
and U21452 (N_21452,N_20962,N_20629);
nand U21453 (N_21453,N_20846,N_20611);
and U21454 (N_21454,N_20704,N_20821);
nor U21455 (N_21455,N_20558,N_20752);
and U21456 (N_21456,N_20867,N_20733);
nand U21457 (N_21457,N_20983,N_20886);
and U21458 (N_21458,N_20773,N_20643);
xor U21459 (N_21459,N_20502,N_20588);
and U21460 (N_21460,N_20618,N_20960);
nor U21461 (N_21461,N_20740,N_20732);
nand U21462 (N_21462,N_20796,N_20724);
xor U21463 (N_21463,N_20797,N_20628);
nor U21464 (N_21464,N_20814,N_20542);
or U21465 (N_21465,N_20931,N_20580);
and U21466 (N_21466,N_20751,N_20602);
nor U21467 (N_21467,N_20800,N_20979);
nand U21468 (N_21468,N_20736,N_20694);
xor U21469 (N_21469,N_20719,N_20613);
nand U21470 (N_21470,N_20723,N_20650);
nand U21471 (N_21471,N_20840,N_20812);
and U21472 (N_21472,N_20700,N_20807);
nand U21473 (N_21473,N_20817,N_20696);
nor U21474 (N_21474,N_20977,N_20894);
xor U21475 (N_21475,N_20773,N_20554);
xnor U21476 (N_21476,N_20960,N_20663);
xnor U21477 (N_21477,N_20920,N_20991);
nor U21478 (N_21478,N_20659,N_20959);
nand U21479 (N_21479,N_20914,N_20837);
and U21480 (N_21480,N_20643,N_20686);
xor U21481 (N_21481,N_20707,N_20683);
nand U21482 (N_21482,N_20766,N_20609);
and U21483 (N_21483,N_20831,N_20579);
and U21484 (N_21484,N_20795,N_20979);
xnor U21485 (N_21485,N_20868,N_20687);
nor U21486 (N_21486,N_20900,N_20596);
nor U21487 (N_21487,N_20667,N_20986);
nand U21488 (N_21488,N_20521,N_20692);
and U21489 (N_21489,N_20947,N_20859);
nor U21490 (N_21490,N_20562,N_20744);
nor U21491 (N_21491,N_20722,N_20783);
xnor U21492 (N_21492,N_20513,N_20645);
or U21493 (N_21493,N_20955,N_20987);
or U21494 (N_21494,N_20742,N_20872);
nor U21495 (N_21495,N_20738,N_20905);
and U21496 (N_21496,N_20750,N_20809);
nand U21497 (N_21497,N_20735,N_20575);
nor U21498 (N_21498,N_20533,N_20998);
xor U21499 (N_21499,N_20643,N_20633);
nand U21500 (N_21500,N_21402,N_21307);
or U21501 (N_21501,N_21429,N_21432);
or U21502 (N_21502,N_21103,N_21342);
or U21503 (N_21503,N_21020,N_21072);
or U21504 (N_21504,N_21406,N_21431);
nand U21505 (N_21505,N_21233,N_21065);
or U21506 (N_21506,N_21074,N_21355);
and U21507 (N_21507,N_21029,N_21470);
xnor U21508 (N_21508,N_21267,N_21392);
and U21509 (N_21509,N_21326,N_21138);
nand U21510 (N_21510,N_21395,N_21259);
and U21511 (N_21511,N_21021,N_21136);
xnor U21512 (N_21512,N_21057,N_21046);
and U21513 (N_21513,N_21078,N_21086);
nand U21514 (N_21514,N_21033,N_21062);
nand U21515 (N_21515,N_21039,N_21323);
and U21516 (N_21516,N_21423,N_21195);
xor U21517 (N_21517,N_21480,N_21214);
nand U21518 (N_21518,N_21120,N_21230);
and U21519 (N_21519,N_21094,N_21393);
nor U21520 (N_21520,N_21114,N_21102);
nor U21521 (N_21521,N_21475,N_21206);
or U21522 (N_21522,N_21009,N_21171);
or U21523 (N_21523,N_21331,N_21116);
and U21524 (N_21524,N_21239,N_21347);
nor U21525 (N_21525,N_21128,N_21388);
nand U21526 (N_21526,N_21236,N_21436);
xnor U21527 (N_21527,N_21411,N_21237);
nand U21528 (N_21528,N_21364,N_21165);
or U21529 (N_21529,N_21224,N_21129);
nand U21530 (N_21530,N_21211,N_21053);
xnor U21531 (N_21531,N_21407,N_21182);
xnor U21532 (N_21532,N_21014,N_21369);
or U21533 (N_21533,N_21194,N_21338);
and U21534 (N_21534,N_21275,N_21111);
nand U21535 (N_21535,N_21435,N_21131);
nand U21536 (N_21536,N_21210,N_21274);
xor U21537 (N_21537,N_21006,N_21445);
and U21538 (N_21538,N_21169,N_21117);
nor U21539 (N_21539,N_21042,N_21066);
nand U21540 (N_21540,N_21321,N_21220);
or U21541 (N_21541,N_21306,N_21499);
or U21542 (N_21542,N_21430,N_21419);
and U21543 (N_21543,N_21213,N_21036);
or U21544 (N_21544,N_21121,N_21461);
and U21545 (N_21545,N_21426,N_21200);
nand U21546 (N_21546,N_21202,N_21399);
or U21547 (N_21547,N_21095,N_21277);
nor U21548 (N_21548,N_21408,N_21290);
or U21549 (N_21549,N_21007,N_21334);
xnor U21550 (N_21550,N_21428,N_21273);
nand U21551 (N_21551,N_21345,N_21447);
xnor U21552 (N_21552,N_21442,N_21023);
or U21553 (N_21553,N_21391,N_21264);
xor U21554 (N_21554,N_21293,N_21088);
or U21555 (N_21555,N_21105,N_21018);
xnor U21556 (N_21556,N_21135,N_21357);
nand U21557 (N_21557,N_21418,N_21374);
nor U21558 (N_21558,N_21226,N_21025);
or U21559 (N_21559,N_21350,N_21485);
nor U21560 (N_21560,N_21263,N_21150);
nor U21561 (N_21561,N_21246,N_21360);
or U21562 (N_21562,N_21482,N_21449);
or U21563 (N_21563,N_21467,N_21484);
nand U21564 (N_21564,N_21143,N_21058);
and U21565 (N_21565,N_21381,N_21166);
nor U21566 (N_21566,N_21162,N_21225);
and U21567 (N_21567,N_21261,N_21311);
and U21568 (N_21568,N_21157,N_21107);
nor U21569 (N_21569,N_21320,N_21075);
nor U21570 (N_21570,N_21285,N_21330);
nand U21571 (N_21571,N_21444,N_21379);
xnor U21572 (N_21572,N_21298,N_21177);
nor U21573 (N_21573,N_21440,N_21145);
or U21574 (N_21574,N_21147,N_21076);
xor U21575 (N_21575,N_21139,N_21005);
or U21576 (N_21576,N_21077,N_21151);
xor U21577 (N_21577,N_21141,N_21368);
xnor U21578 (N_21578,N_21375,N_21011);
or U21579 (N_21579,N_21133,N_21329);
and U21580 (N_21580,N_21056,N_21314);
xor U21581 (N_21581,N_21003,N_21333);
nor U21582 (N_21582,N_21457,N_21284);
xnor U21583 (N_21583,N_21271,N_21371);
or U21584 (N_21584,N_21491,N_21174);
nand U21585 (N_21585,N_21251,N_21473);
nor U21586 (N_21586,N_21041,N_21420);
xnor U21587 (N_21587,N_21010,N_21322);
nand U21588 (N_21588,N_21398,N_21051);
and U21589 (N_21589,N_21451,N_21175);
nand U21590 (N_21590,N_21389,N_21110);
nand U21591 (N_21591,N_21181,N_21292);
xor U21592 (N_21592,N_21097,N_21037);
or U21593 (N_21593,N_21409,N_21082);
nor U21594 (N_21594,N_21497,N_21244);
nor U21595 (N_21595,N_21280,N_21093);
nand U21596 (N_21596,N_21125,N_21235);
and U21597 (N_21597,N_21462,N_21034);
nand U21598 (N_21598,N_21043,N_21257);
nor U21599 (N_21599,N_21336,N_21365);
and U21600 (N_21600,N_21026,N_21463);
or U21601 (N_21601,N_21223,N_21348);
nand U21602 (N_21602,N_21495,N_21212);
and U21603 (N_21603,N_21363,N_21327);
xor U21604 (N_21604,N_21084,N_21173);
xor U21605 (N_21605,N_21413,N_21061);
nand U21606 (N_21606,N_21193,N_21013);
nor U21607 (N_21607,N_21112,N_21178);
or U21608 (N_21608,N_21332,N_21247);
nor U21609 (N_21609,N_21179,N_21291);
nor U21610 (N_21610,N_21064,N_21164);
and U21611 (N_21611,N_21149,N_21070);
and U21612 (N_21612,N_21113,N_21299);
nor U21613 (N_21613,N_21305,N_21241);
nor U21614 (N_21614,N_21486,N_21337);
and U21615 (N_21615,N_21468,N_21035);
nand U21616 (N_21616,N_21146,N_21481);
and U21617 (N_21617,N_21281,N_21203);
xnor U21618 (N_21618,N_21049,N_21303);
and U21619 (N_21619,N_21438,N_21301);
and U21620 (N_21620,N_21324,N_21390);
and U21621 (N_21621,N_21489,N_21498);
nand U21622 (N_21622,N_21243,N_21249);
nand U21623 (N_21623,N_21276,N_21268);
or U21624 (N_21624,N_21354,N_21073);
nand U21625 (N_21625,N_21218,N_21404);
nand U21626 (N_21626,N_21450,N_21279);
and U21627 (N_21627,N_21190,N_21297);
xor U21628 (N_21628,N_21192,N_21490);
nor U21629 (N_21629,N_21158,N_21401);
nand U21630 (N_21630,N_21340,N_21109);
nor U21631 (N_21631,N_21343,N_21159);
and U21632 (N_21632,N_21328,N_21400);
xor U21633 (N_21633,N_21130,N_21221);
and U21634 (N_21634,N_21469,N_21176);
xor U21635 (N_21635,N_21319,N_21378);
and U21636 (N_21636,N_21229,N_21022);
xor U21637 (N_21637,N_21416,N_21201);
and U21638 (N_21638,N_21119,N_21361);
xnor U21639 (N_21639,N_21253,N_21424);
and U21640 (N_21640,N_21232,N_21060);
nor U21641 (N_21641,N_21358,N_21197);
nor U21642 (N_21642,N_21155,N_21096);
and U21643 (N_21643,N_21494,N_21465);
or U21644 (N_21644,N_21087,N_21068);
and U21645 (N_21645,N_21312,N_21038);
xnor U21646 (N_21646,N_21403,N_21483);
and U21647 (N_21647,N_21100,N_21044);
xor U21648 (N_21648,N_21433,N_21474);
nor U21649 (N_21649,N_21460,N_21367);
or U21650 (N_21650,N_21069,N_21180);
nor U21651 (N_21651,N_21228,N_21089);
nor U21652 (N_21652,N_21118,N_21050);
nor U21653 (N_21653,N_21287,N_21387);
xor U21654 (N_21654,N_21380,N_21122);
nand U21655 (N_21655,N_21161,N_21017);
nor U21656 (N_21656,N_21153,N_21288);
nand U21657 (N_21657,N_21488,N_21079);
xor U21658 (N_21658,N_21040,N_21417);
xor U21659 (N_21659,N_21487,N_21466);
nor U21660 (N_21660,N_21170,N_21370);
xnor U21661 (N_21661,N_21304,N_21001);
xnor U21662 (N_21662,N_21030,N_21313);
nand U21663 (N_21663,N_21148,N_21152);
and U21664 (N_21664,N_21382,N_21356);
nand U21665 (N_21665,N_21351,N_21059);
and U21666 (N_21666,N_21300,N_21083);
xnor U21667 (N_21667,N_21296,N_21372);
xnor U21668 (N_21668,N_21405,N_21027);
or U21669 (N_21669,N_21415,N_21004);
xnor U21670 (N_21670,N_21455,N_21002);
nor U21671 (N_21671,N_21231,N_21278);
nand U21672 (N_21672,N_21384,N_21184);
or U21673 (N_21673,N_21071,N_21383);
nor U21674 (N_21674,N_21132,N_21217);
nor U21675 (N_21675,N_21309,N_21472);
or U21676 (N_21676,N_21453,N_21185);
and U21677 (N_21677,N_21396,N_21047);
xnor U21678 (N_21678,N_21349,N_21476);
nor U21679 (N_21679,N_21126,N_21208);
or U21680 (N_21680,N_21448,N_21352);
or U21681 (N_21681,N_21242,N_21421);
xnor U21682 (N_21682,N_21295,N_21191);
nor U21683 (N_21683,N_21492,N_21204);
nor U21684 (N_21684,N_21439,N_21199);
and U21685 (N_21685,N_21090,N_21187);
nor U21686 (N_21686,N_21254,N_21394);
or U21687 (N_21687,N_21386,N_21456);
or U21688 (N_21688,N_21373,N_21250);
xnor U21689 (N_21689,N_21067,N_21353);
xnor U21690 (N_21690,N_21265,N_21359);
xnor U21691 (N_21691,N_21063,N_21286);
and U21692 (N_21692,N_21142,N_21283);
nor U21693 (N_21693,N_21366,N_21479);
nand U21694 (N_21694,N_21317,N_21028);
and U21695 (N_21695,N_21144,N_21471);
or U21696 (N_21696,N_21092,N_21458);
and U21697 (N_21697,N_21346,N_21454);
or U21698 (N_21698,N_21140,N_21052);
nand U21699 (N_21699,N_21422,N_21252);
nand U21700 (N_21700,N_21315,N_21167);
xor U21701 (N_21701,N_21452,N_21183);
or U21702 (N_21702,N_21310,N_21446);
xnor U21703 (N_21703,N_21425,N_21362);
and U21704 (N_21704,N_21376,N_21186);
and U21705 (N_21705,N_21410,N_21024);
and U21706 (N_21706,N_21219,N_21012);
xnor U21707 (N_21707,N_21289,N_21108);
and U21708 (N_21708,N_21335,N_21019);
or U21709 (N_21709,N_21101,N_21085);
nor U21710 (N_21710,N_21016,N_21282);
and U21711 (N_21711,N_21216,N_21248);
nor U21712 (N_21712,N_21344,N_21015);
and U21713 (N_21713,N_21000,N_21339);
and U21714 (N_21714,N_21255,N_21104);
nor U21715 (N_21715,N_21256,N_21316);
nor U21716 (N_21716,N_21272,N_21269);
nand U21717 (N_21717,N_21106,N_21124);
or U21718 (N_21718,N_21154,N_21091);
or U21719 (N_21719,N_21385,N_21160);
nand U21720 (N_21720,N_21127,N_21080);
nor U21721 (N_21721,N_21464,N_21434);
nand U21722 (N_21722,N_21397,N_21054);
nor U21723 (N_21723,N_21168,N_21207);
or U21724 (N_21724,N_21443,N_21262);
xnor U21725 (N_21725,N_21266,N_21055);
xnor U21726 (N_21726,N_21008,N_21032);
nor U21727 (N_21727,N_21325,N_21115);
nand U21728 (N_21728,N_21031,N_21294);
xnor U21729 (N_21729,N_21198,N_21318);
or U21730 (N_21730,N_21437,N_21496);
nand U21731 (N_21731,N_21098,N_21123);
and U21732 (N_21732,N_21302,N_21478);
and U21733 (N_21733,N_21459,N_21441);
or U21734 (N_21734,N_21137,N_21215);
nand U21735 (N_21735,N_21341,N_21477);
nor U21736 (N_21736,N_21414,N_21209);
nand U21737 (N_21737,N_21045,N_21189);
and U21738 (N_21738,N_21156,N_21260);
or U21739 (N_21739,N_21240,N_21081);
or U21740 (N_21740,N_21196,N_21245);
xnor U21741 (N_21741,N_21427,N_21099);
xnor U21742 (N_21742,N_21377,N_21258);
xnor U21743 (N_21743,N_21205,N_21412);
or U21744 (N_21744,N_21227,N_21188);
nor U21745 (N_21745,N_21048,N_21172);
or U21746 (N_21746,N_21222,N_21270);
or U21747 (N_21747,N_21163,N_21308);
and U21748 (N_21748,N_21493,N_21238);
or U21749 (N_21749,N_21134,N_21234);
nor U21750 (N_21750,N_21057,N_21139);
or U21751 (N_21751,N_21062,N_21462);
xnor U21752 (N_21752,N_21468,N_21213);
nand U21753 (N_21753,N_21362,N_21407);
or U21754 (N_21754,N_21341,N_21372);
xor U21755 (N_21755,N_21108,N_21343);
nand U21756 (N_21756,N_21101,N_21199);
nand U21757 (N_21757,N_21488,N_21469);
and U21758 (N_21758,N_21010,N_21235);
xor U21759 (N_21759,N_21046,N_21210);
and U21760 (N_21760,N_21150,N_21187);
nor U21761 (N_21761,N_21189,N_21355);
nor U21762 (N_21762,N_21137,N_21136);
or U21763 (N_21763,N_21474,N_21337);
and U21764 (N_21764,N_21433,N_21212);
nand U21765 (N_21765,N_21296,N_21248);
and U21766 (N_21766,N_21142,N_21207);
nand U21767 (N_21767,N_21134,N_21381);
nor U21768 (N_21768,N_21384,N_21395);
nand U21769 (N_21769,N_21003,N_21048);
nand U21770 (N_21770,N_21015,N_21471);
xor U21771 (N_21771,N_21027,N_21166);
nor U21772 (N_21772,N_21124,N_21205);
or U21773 (N_21773,N_21205,N_21239);
and U21774 (N_21774,N_21344,N_21465);
nand U21775 (N_21775,N_21344,N_21162);
xnor U21776 (N_21776,N_21164,N_21388);
nor U21777 (N_21777,N_21094,N_21293);
nand U21778 (N_21778,N_21172,N_21474);
nor U21779 (N_21779,N_21059,N_21354);
and U21780 (N_21780,N_21186,N_21217);
nand U21781 (N_21781,N_21364,N_21464);
or U21782 (N_21782,N_21076,N_21027);
nand U21783 (N_21783,N_21120,N_21028);
xnor U21784 (N_21784,N_21253,N_21483);
nand U21785 (N_21785,N_21284,N_21156);
or U21786 (N_21786,N_21312,N_21423);
nor U21787 (N_21787,N_21100,N_21482);
xor U21788 (N_21788,N_21400,N_21407);
nand U21789 (N_21789,N_21450,N_21386);
and U21790 (N_21790,N_21172,N_21026);
or U21791 (N_21791,N_21129,N_21310);
nor U21792 (N_21792,N_21342,N_21391);
nor U21793 (N_21793,N_21285,N_21336);
or U21794 (N_21794,N_21114,N_21210);
xnor U21795 (N_21795,N_21239,N_21076);
nor U21796 (N_21796,N_21085,N_21034);
nand U21797 (N_21797,N_21054,N_21098);
xnor U21798 (N_21798,N_21011,N_21344);
nand U21799 (N_21799,N_21328,N_21138);
xnor U21800 (N_21800,N_21167,N_21454);
or U21801 (N_21801,N_21035,N_21452);
xor U21802 (N_21802,N_21251,N_21348);
and U21803 (N_21803,N_21126,N_21421);
nor U21804 (N_21804,N_21301,N_21312);
xnor U21805 (N_21805,N_21389,N_21164);
xor U21806 (N_21806,N_21418,N_21451);
nor U21807 (N_21807,N_21439,N_21429);
nand U21808 (N_21808,N_21110,N_21452);
nor U21809 (N_21809,N_21360,N_21075);
nand U21810 (N_21810,N_21268,N_21303);
and U21811 (N_21811,N_21436,N_21027);
or U21812 (N_21812,N_21402,N_21051);
nor U21813 (N_21813,N_21386,N_21245);
nor U21814 (N_21814,N_21094,N_21162);
and U21815 (N_21815,N_21394,N_21068);
or U21816 (N_21816,N_21220,N_21377);
nand U21817 (N_21817,N_21006,N_21335);
nor U21818 (N_21818,N_21493,N_21002);
and U21819 (N_21819,N_21414,N_21475);
or U21820 (N_21820,N_21463,N_21406);
xnor U21821 (N_21821,N_21258,N_21379);
and U21822 (N_21822,N_21454,N_21185);
nor U21823 (N_21823,N_21212,N_21180);
and U21824 (N_21824,N_21183,N_21189);
and U21825 (N_21825,N_21398,N_21387);
and U21826 (N_21826,N_21141,N_21394);
nor U21827 (N_21827,N_21399,N_21418);
nand U21828 (N_21828,N_21265,N_21399);
nand U21829 (N_21829,N_21491,N_21494);
nand U21830 (N_21830,N_21480,N_21258);
nand U21831 (N_21831,N_21463,N_21034);
or U21832 (N_21832,N_21490,N_21427);
nor U21833 (N_21833,N_21227,N_21397);
xnor U21834 (N_21834,N_21036,N_21250);
or U21835 (N_21835,N_21193,N_21469);
or U21836 (N_21836,N_21420,N_21020);
xor U21837 (N_21837,N_21263,N_21318);
or U21838 (N_21838,N_21366,N_21036);
and U21839 (N_21839,N_21106,N_21428);
and U21840 (N_21840,N_21007,N_21079);
or U21841 (N_21841,N_21305,N_21080);
xnor U21842 (N_21842,N_21187,N_21460);
xnor U21843 (N_21843,N_21200,N_21217);
and U21844 (N_21844,N_21296,N_21219);
or U21845 (N_21845,N_21339,N_21046);
or U21846 (N_21846,N_21268,N_21150);
and U21847 (N_21847,N_21070,N_21383);
nor U21848 (N_21848,N_21377,N_21047);
nor U21849 (N_21849,N_21168,N_21249);
and U21850 (N_21850,N_21052,N_21465);
or U21851 (N_21851,N_21269,N_21126);
nand U21852 (N_21852,N_21240,N_21417);
and U21853 (N_21853,N_21167,N_21246);
xnor U21854 (N_21854,N_21293,N_21499);
nor U21855 (N_21855,N_21276,N_21124);
or U21856 (N_21856,N_21347,N_21331);
nand U21857 (N_21857,N_21036,N_21314);
xor U21858 (N_21858,N_21215,N_21098);
nor U21859 (N_21859,N_21115,N_21314);
or U21860 (N_21860,N_21190,N_21470);
or U21861 (N_21861,N_21092,N_21401);
nor U21862 (N_21862,N_21351,N_21360);
or U21863 (N_21863,N_21354,N_21322);
xnor U21864 (N_21864,N_21176,N_21113);
and U21865 (N_21865,N_21346,N_21457);
and U21866 (N_21866,N_21313,N_21117);
nand U21867 (N_21867,N_21078,N_21353);
nand U21868 (N_21868,N_21249,N_21228);
and U21869 (N_21869,N_21116,N_21389);
and U21870 (N_21870,N_21031,N_21211);
nand U21871 (N_21871,N_21428,N_21174);
nor U21872 (N_21872,N_21175,N_21187);
or U21873 (N_21873,N_21224,N_21043);
or U21874 (N_21874,N_21007,N_21171);
and U21875 (N_21875,N_21490,N_21023);
nand U21876 (N_21876,N_21308,N_21463);
and U21877 (N_21877,N_21048,N_21022);
nor U21878 (N_21878,N_21220,N_21173);
and U21879 (N_21879,N_21337,N_21340);
nand U21880 (N_21880,N_21361,N_21286);
nor U21881 (N_21881,N_21445,N_21071);
nor U21882 (N_21882,N_21110,N_21314);
and U21883 (N_21883,N_21069,N_21303);
and U21884 (N_21884,N_21388,N_21110);
nand U21885 (N_21885,N_21093,N_21102);
nand U21886 (N_21886,N_21322,N_21145);
nor U21887 (N_21887,N_21433,N_21421);
or U21888 (N_21888,N_21295,N_21445);
nor U21889 (N_21889,N_21280,N_21326);
nor U21890 (N_21890,N_21448,N_21337);
or U21891 (N_21891,N_21300,N_21064);
xor U21892 (N_21892,N_21321,N_21291);
and U21893 (N_21893,N_21481,N_21044);
nand U21894 (N_21894,N_21339,N_21154);
nor U21895 (N_21895,N_21422,N_21297);
xor U21896 (N_21896,N_21393,N_21481);
nor U21897 (N_21897,N_21258,N_21221);
nor U21898 (N_21898,N_21429,N_21153);
nor U21899 (N_21899,N_21334,N_21092);
xor U21900 (N_21900,N_21098,N_21425);
and U21901 (N_21901,N_21155,N_21357);
or U21902 (N_21902,N_21303,N_21139);
and U21903 (N_21903,N_21160,N_21101);
xor U21904 (N_21904,N_21066,N_21465);
nor U21905 (N_21905,N_21205,N_21287);
nand U21906 (N_21906,N_21015,N_21118);
nor U21907 (N_21907,N_21114,N_21326);
nor U21908 (N_21908,N_21375,N_21027);
and U21909 (N_21909,N_21152,N_21331);
or U21910 (N_21910,N_21296,N_21344);
nor U21911 (N_21911,N_21190,N_21463);
nand U21912 (N_21912,N_21239,N_21228);
xnor U21913 (N_21913,N_21359,N_21012);
and U21914 (N_21914,N_21438,N_21332);
nor U21915 (N_21915,N_21398,N_21213);
or U21916 (N_21916,N_21461,N_21009);
nor U21917 (N_21917,N_21472,N_21213);
nor U21918 (N_21918,N_21075,N_21127);
xor U21919 (N_21919,N_21038,N_21085);
nor U21920 (N_21920,N_21035,N_21309);
nand U21921 (N_21921,N_21117,N_21183);
nor U21922 (N_21922,N_21014,N_21057);
or U21923 (N_21923,N_21304,N_21075);
and U21924 (N_21924,N_21300,N_21249);
and U21925 (N_21925,N_21340,N_21243);
xnor U21926 (N_21926,N_21456,N_21088);
xor U21927 (N_21927,N_21244,N_21408);
nor U21928 (N_21928,N_21105,N_21062);
nand U21929 (N_21929,N_21088,N_21148);
or U21930 (N_21930,N_21236,N_21255);
nand U21931 (N_21931,N_21492,N_21446);
or U21932 (N_21932,N_21138,N_21389);
nor U21933 (N_21933,N_21475,N_21000);
and U21934 (N_21934,N_21227,N_21411);
nor U21935 (N_21935,N_21102,N_21097);
nor U21936 (N_21936,N_21318,N_21001);
or U21937 (N_21937,N_21264,N_21447);
nor U21938 (N_21938,N_21266,N_21425);
nand U21939 (N_21939,N_21419,N_21318);
or U21940 (N_21940,N_21371,N_21107);
or U21941 (N_21941,N_21388,N_21209);
and U21942 (N_21942,N_21146,N_21308);
nor U21943 (N_21943,N_21305,N_21412);
or U21944 (N_21944,N_21476,N_21236);
nand U21945 (N_21945,N_21164,N_21041);
and U21946 (N_21946,N_21089,N_21078);
nor U21947 (N_21947,N_21322,N_21458);
nand U21948 (N_21948,N_21403,N_21375);
and U21949 (N_21949,N_21127,N_21021);
and U21950 (N_21950,N_21289,N_21453);
or U21951 (N_21951,N_21185,N_21129);
nor U21952 (N_21952,N_21205,N_21003);
nand U21953 (N_21953,N_21413,N_21249);
and U21954 (N_21954,N_21310,N_21134);
and U21955 (N_21955,N_21309,N_21257);
nor U21956 (N_21956,N_21248,N_21074);
or U21957 (N_21957,N_21191,N_21236);
or U21958 (N_21958,N_21374,N_21271);
nor U21959 (N_21959,N_21407,N_21096);
nand U21960 (N_21960,N_21268,N_21106);
or U21961 (N_21961,N_21339,N_21024);
xor U21962 (N_21962,N_21319,N_21075);
xnor U21963 (N_21963,N_21275,N_21306);
nor U21964 (N_21964,N_21228,N_21032);
xnor U21965 (N_21965,N_21178,N_21498);
nand U21966 (N_21966,N_21007,N_21145);
or U21967 (N_21967,N_21018,N_21174);
and U21968 (N_21968,N_21357,N_21193);
or U21969 (N_21969,N_21466,N_21397);
xnor U21970 (N_21970,N_21405,N_21111);
or U21971 (N_21971,N_21146,N_21307);
xnor U21972 (N_21972,N_21237,N_21153);
nand U21973 (N_21973,N_21415,N_21057);
xor U21974 (N_21974,N_21255,N_21009);
nand U21975 (N_21975,N_21485,N_21035);
nor U21976 (N_21976,N_21074,N_21479);
xor U21977 (N_21977,N_21248,N_21155);
and U21978 (N_21978,N_21037,N_21127);
or U21979 (N_21979,N_21032,N_21412);
nor U21980 (N_21980,N_21462,N_21496);
and U21981 (N_21981,N_21365,N_21174);
xnor U21982 (N_21982,N_21339,N_21438);
nand U21983 (N_21983,N_21026,N_21011);
or U21984 (N_21984,N_21141,N_21031);
nand U21985 (N_21985,N_21404,N_21210);
nand U21986 (N_21986,N_21370,N_21230);
nand U21987 (N_21987,N_21109,N_21302);
nand U21988 (N_21988,N_21154,N_21382);
nor U21989 (N_21989,N_21037,N_21007);
or U21990 (N_21990,N_21488,N_21374);
or U21991 (N_21991,N_21303,N_21218);
or U21992 (N_21992,N_21228,N_21361);
and U21993 (N_21993,N_21436,N_21172);
or U21994 (N_21994,N_21296,N_21493);
nor U21995 (N_21995,N_21497,N_21276);
xnor U21996 (N_21996,N_21090,N_21344);
xnor U21997 (N_21997,N_21447,N_21165);
or U21998 (N_21998,N_21078,N_21137);
or U21999 (N_21999,N_21205,N_21206);
nor U22000 (N_22000,N_21558,N_21873);
and U22001 (N_22001,N_21637,N_21806);
and U22002 (N_22002,N_21963,N_21703);
nand U22003 (N_22003,N_21933,N_21762);
xor U22004 (N_22004,N_21601,N_21970);
or U22005 (N_22005,N_21555,N_21512);
and U22006 (N_22006,N_21736,N_21774);
nor U22007 (N_22007,N_21866,N_21804);
nand U22008 (N_22008,N_21548,N_21683);
xor U22009 (N_22009,N_21900,N_21631);
or U22010 (N_22010,N_21645,N_21602);
nand U22011 (N_22011,N_21968,N_21655);
nand U22012 (N_22012,N_21597,N_21923);
and U22013 (N_22013,N_21792,N_21693);
nand U22014 (N_22014,N_21583,N_21921);
and U22015 (N_22015,N_21687,N_21901);
or U22016 (N_22016,N_21725,N_21985);
xnor U22017 (N_22017,N_21584,N_21864);
nor U22018 (N_22018,N_21625,N_21672);
or U22019 (N_22019,N_21952,N_21750);
nor U22020 (N_22020,N_21909,N_21653);
or U22021 (N_22021,N_21695,N_21786);
nor U22022 (N_22022,N_21814,N_21887);
nor U22023 (N_22023,N_21528,N_21825);
nor U22024 (N_22024,N_21839,N_21519);
xor U22025 (N_22025,N_21841,N_21675);
and U22026 (N_22026,N_21958,N_21521);
nand U22027 (N_22027,N_21808,N_21545);
or U22028 (N_22028,N_21605,N_21799);
nor U22029 (N_22029,N_21892,N_21656);
and U22030 (N_22030,N_21707,N_21940);
nand U22031 (N_22031,N_21938,N_21710);
and U22032 (N_22032,N_21904,N_21905);
nor U22033 (N_22033,N_21777,N_21794);
and U22034 (N_22034,N_21859,N_21827);
nor U22035 (N_22035,N_21701,N_21824);
and U22036 (N_22036,N_21998,N_21907);
nand U22037 (N_22037,N_21882,N_21870);
nand U22038 (N_22038,N_21834,N_21778);
or U22039 (N_22039,N_21747,N_21678);
nand U22040 (N_22040,N_21634,N_21805);
or U22041 (N_22041,N_21833,N_21871);
xor U22042 (N_22042,N_21630,N_21667);
nor U22043 (N_22043,N_21628,N_21680);
nor U22044 (N_22044,N_21809,N_21977);
nor U22045 (N_22045,N_21767,N_21636);
xnor U22046 (N_22046,N_21535,N_21781);
xnor U22047 (N_22047,N_21945,N_21649);
and U22048 (N_22048,N_21527,N_21543);
xor U22049 (N_22049,N_21925,N_21991);
and U22050 (N_22050,N_21658,N_21592);
xor U22051 (N_22051,N_21650,N_21522);
or U22052 (N_22052,N_21638,N_21537);
nand U22053 (N_22053,N_21622,N_21606);
xor U22054 (N_22054,N_21632,N_21503);
nor U22055 (N_22055,N_21876,N_21946);
nand U22056 (N_22056,N_21699,N_21937);
and U22057 (N_22057,N_21594,N_21782);
nor U22058 (N_22058,N_21593,N_21640);
nor U22059 (N_22059,N_21821,N_21560);
or U22060 (N_22060,N_21844,N_21980);
xor U22061 (N_22061,N_21990,N_21950);
nor U22062 (N_22062,N_21916,N_21822);
xor U22063 (N_22063,N_21588,N_21847);
xnor U22064 (N_22064,N_21738,N_21557);
nor U22065 (N_22065,N_21639,N_21926);
nor U22066 (N_22066,N_21677,N_21981);
nor U22067 (N_22067,N_21727,N_21733);
nand U22068 (N_22068,N_21501,N_21595);
nand U22069 (N_22069,N_21754,N_21918);
nand U22070 (N_22070,N_21800,N_21563);
and U22071 (N_22071,N_21642,N_21723);
nand U22072 (N_22072,N_21765,N_21883);
or U22073 (N_22073,N_21797,N_21550);
and U22074 (N_22074,N_21886,N_21694);
nand U22075 (N_22075,N_21944,N_21586);
and U22076 (N_22076,N_21720,N_21947);
or U22077 (N_22077,N_21609,N_21801);
or U22078 (N_22078,N_21831,N_21547);
and U22079 (N_22079,N_21552,N_21994);
nor U22080 (N_22080,N_21791,N_21965);
nand U22081 (N_22081,N_21744,N_21542);
xor U22082 (N_22082,N_21518,N_21881);
xor U22083 (N_22083,N_21955,N_21964);
nand U22084 (N_22084,N_21856,N_21995);
xnor U22085 (N_22085,N_21816,N_21686);
nand U22086 (N_22086,N_21961,N_21534);
or U22087 (N_22087,N_21743,N_21908);
nand U22088 (N_22088,N_21599,N_21889);
nand U22089 (N_22089,N_21697,N_21561);
and U22090 (N_22090,N_21681,N_21633);
and U22091 (N_22091,N_21842,N_21539);
nand U22092 (N_22092,N_21540,N_21529);
xnor U22093 (N_22093,N_21861,N_21502);
nor U22094 (N_22094,N_21993,N_21611);
xor U22095 (N_22095,N_21932,N_21807);
or U22096 (N_22096,N_21776,N_21910);
xor U22097 (N_22097,N_21721,N_21505);
nand U22098 (N_22098,N_21811,N_21868);
or U22099 (N_22099,N_21741,N_21784);
xor U22100 (N_22100,N_21812,N_21986);
nand U22101 (N_22101,N_21924,N_21732);
xor U22102 (N_22102,N_21511,N_21884);
or U22103 (N_22103,N_21549,N_21971);
nor U22104 (N_22104,N_21624,N_21897);
or U22105 (N_22105,N_21851,N_21795);
nand U22106 (N_22106,N_21587,N_21929);
nor U22107 (N_22107,N_21559,N_21838);
xnor U22108 (N_22108,N_21737,N_21880);
xnor U22109 (N_22109,N_21755,N_21676);
and U22110 (N_22110,N_21620,N_21914);
or U22111 (N_22111,N_21513,N_21953);
nand U22112 (N_22112,N_21793,N_21532);
or U22113 (N_22113,N_21858,N_21665);
and U22114 (N_22114,N_21819,N_21878);
xor U22115 (N_22115,N_21846,N_21618);
xnor U22116 (N_22116,N_21917,N_21617);
or U22117 (N_22117,N_21523,N_21506);
and U22118 (N_22118,N_21959,N_21850);
xor U22119 (N_22119,N_21810,N_21531);
or U22120 (N_22120,N_21826,N_21629);
or U22121 (N_22121,N_21504,N_21753);
and U22122 (N_22122,N_21714,N_21668);
and U22123 (N_22123,N_21891,N_21582);
or U22124 (N_22124,N_21930,N_21690);
nand U22125 (N_22125,N_21571,N_21516);
and U22126 (N_22126,N_21698,N_21644);
and U22127 (N_22127,N_21853,N_21722);
nand U22128 (N_22128,N_21840,N_21979);
xnor U22129 (N_22129,N_21724,N_21942);
and U22130 (N_22130,N_21612,N_21987);
xor U22131 (N_22131,N_21818,N_21578);
nor U22132 (N_22132,N_21713,N_21775);
nand U22133 (N_22133,N_21912,N_21514);
nor U22134 (N_22134,N_21948,N_21978);
or U22135 (N_22135,N_21689,N_21659);
xor U22136 (N_22136,N_21780,N_21598);
nor U22137 (N_22137,N_21553,N_21757);
nor U22138 (N_22138,N_21614,N_21888);
xor U22139 (N_22139,N_21957,N_21748);
nor U22140 (N_22140,N_21673,N_21515);
or U22141 (N_22141,N_21976,N_21734);
and U22142 (N_22142,N_21815,N_21789);
or U22143 (N_22143,N_21541,N_21773);
or U22144 (N_22144,N_21788,N_21684);
or U22145 (N_22145,N_21662,N_21719);
nand U22146 (N_22146,N_21544,N_21735);
and U22147 (N_22147,N_21829,N_21798);
nor U22148 (N_22148,N_21621,N_21607);
xnor U22149 (N_22149,N_21657,N_21603);
nand U22150 (N_22150,N_21641,N_21726);
nand U22151 (N_22151,N_21845,N_21749);
or U22152 (N_22152,N_21709,N_21761);
and U22153 (N_22153,N_21654,N_21813);
xor U22154 (N_22154,N_21565,N_21783);
nor U22155 (N_22155,N_21943,N_21573);
and U22156 (N_22156,N_21567,N_21854);
xor U22157 (N_22157,N_21664,N_21837);
nand U22158 (N_22158,N_21759,N_21685);
or U22159 (N_22159,N_21860,N_21520);
xnor U22160 (N_22160,N_21615,N_21890);
or U22161 (N_22161,N_21715,N_21712);
nor U22162 (N_22162,N_21731,N_21973);
xor U22163 (N_22163,N_21752,N_21613);
and U22164 (N_22164,N_21652,N_21817);
and U22165 (N_22165,N_21989,N_21779);
nand U22166 (N_22166,N_21982,N_21770);
nand U22167 (N_22167,N_21646,N_21857);
or U22168 (N_22168,N_21764,N_21936);
nor U22169 (N_22169,N_21716,N_21619);
nor U22170 (N_22170,N_21577,N_21832);
or U22171 (N_22171,N_21627,N_21526);
nand U22172 (N_22172,N_21863,N_21702);
and U22173 (N_22173,N_21556,N_21705);
nand U22174 (N_22174,N_21579,N_21533);
or U22175 (N_22175,N_21751,N_21706);
or U22176 (N_22176,N_21576,N_21530);
nand U22177 (N_22177,N_21729,N_21906);
or U22178 (N_22178,N_21865,N_21670);
xor U22179 (N_22179,N_21745,N_21769);
nor U22180 (N_22180,N_21972,N_21960);
or U22181 (N_22181,N_21728,N_21575);
nand U22182 (N_22182,N_21939,N_21700);
nor U22183 (N_22183,N_21796,N_21554);
nand U22184 (N_22184,N_21828,N_21691);
nand U22185 (N_22185,N_21830,N_21580);
nor U22186 (N_22186,N_21951,N_21651);
or U22187 (N_22187,N_21803,N_21843);
xor U22188 (N_22188,N_21999,N_21635);
or U22189 (N_22189,N_21682,N_21967);
and U22190 (N_22190,N_21975,N_21517);
xnor U22191 (N_22191,N_21927,N_21708);
xor U22192 (N_22192,N_21772,N_21836);
nor U22193 (N_22193,N_21756,N_21524);
nor U22194 (N_22194,N_21935,N_21974);
xor U22195 (N_22195,N_21768,N_21902);
or U22196 (N_22196,N_21536,N_21894);
or U22197 (N_22197,N_21903,N_21570);
and U22198 (N_22198,N_21546,N_21647);
nor U22199 (N_22199,N_21867,N_21616);
xnor U22200 (N_22200,N_21855,N_21604);
and U22201 (N_22201,N_21872,N_21941);
nand U22202 (N_22202,N_21671,N_21898);
nor U22203 (N_22203,N_21608,N_21823);
xor U22204 (N_22204,N_21988,N_21997);
xnor U22205 (N_22205,N_21643,N_21996);
nand U22206 (N_22206,N_21913,N_21954);
nand U22207 (N_22207,N_21669,N_21984);
nand U22208 (N_22208,N_21983,N_21802);
nand U22209 (N_22209,N_21717,N_21848);
nor U22210 (N_22210,N_21568,N_21696);
or U22211 (N_22211,N_21895,N_21875);
xnor U22212 (N_22212,N_21896,N_21581);
nand U22213 (N_22213,N_21648,N_21911);
nand U22214 (N_22214,N_21666,N_21688);
or U22215 (N_22215,N_21885,N_21739);
xnor U22216 (N_22216,N_21785,N_21852);
nor U22217 (N_22217,N_21787,N_21572);
and U22218 (N_22218,N_21869,N_21574);
xor U22219 (N_22219,N_21591,N_21835);
nor U22220 (N_22220,N_21934,N_21956);
xnor U22221 (N_22221,N_21730,N_21589);
nor U22222 (N_22222,N_21596,N_21711);
or U22223 (N_22223,N_21566,N_21899);
or U22224 (N_22224,N_21525,N_21509);
or U22225 (N_22225,N_21663,N_21766);
and U22226 (N_22226,N_21623,N_21915);
and U22227 (N_22227,N_21551,N_21874);
and U22228 (N_22228,N_21877,N_21674);
xor U22229 (N_22229,N_21679,N_21742);
nand U22230 (N_22230,N_21562,N_21564);
xnor U22231 (N_22231,N_21600,N_21500);
xnor U22232 (N_22232,N_21569,N_21771);
nand U22233 (N_22233,N_21969,N_21718);
nor U22234 (N_22234,N_21820,N_21538);
xnor U22235 (N_22235,N_21931,N_21758);
and U22236 (N_22236,N_21928,N_21660);
nor U22237 (N_22237,N_21966,N_21704);
and U22238 (N_22238,N_21763,N_21590);
nand U22239 (N_22239,N_21661,N_21862);
xor U22240 (N_22240,N_21740,N_21790);
nand U22241 (N_22241,N_21919,N_21508);
and U22242 (N_22242,N_21992,N_21585);
or U22243 (N_22243,N_21610,N_21849);
or U22244 (N_22244,N_21692,N_21922);
nor U22245 (N_22245,N_21760,N_21962);
or U22246 (N_22246,N_21510,N_21507);
nand U22247 (N_22247,N_21893,N_21879);
xor U22248 (N_22248,N_21949,N_21746);
or U22249 (N_22249,N_21626,N_21920);
and U22250 (N_22250,N_21597,N_21645);
nor U22251 (N_22251,N_21817,N_21866);
and U22252 (N_22252,N_21600,N_21976);
and U22253 (N_22253,N_21676,N_21748);
and U22254 (N_22254,N_21622,N_21911);
nor U22255 (N_22255,N_21772,N_21688);
and U22256 (N_22256,N_21722,N_21841);
nand U22257 (N_22257,N_21804,N_21538);
xor U22258 (N_22258,N_21949,N_21880);
or U22259 (N_22259,N_21885,N_21800);
nand U22260 (N_22260,N_21632,N_21669);
nor U22261 (N_22261,N_21689,N_21555);
or U22262 (N_22262,N_21628,N_21616);
xnor U22263 (N_22263,N_21757,N_21794);
or U22264 (N_22264,N_21685,N_21997);
nand U22265 (N_22265,N_21515,N_21710);
or U22266 (N_22266,N_21507,N_21985);
and U22267 (N_22267,N_21761,N_21692);
nand U22268 (N_22268,N_21626,N_21509);
nor U22269 (N_22269,N_21555,N_21739);
nor U22270 (N_22270,N_21818,N_21506);
or U22271 (N_22271,N_21782,N_21506);
and U22272 (N_22272,N_21592,N_21945);
or U22273 (N_22273,N_21662,N_21689);
xor U22274 (N_22274,N_21742,N_21737);
nand U22275 (N_22275,N_21784,N_21832);
nand U22276 (N_22276,N_21543,N_21948);
and U22277 (N_22277,N_21768,N_21840);
or U22278 (N_22278,N_21695,N_21937);
nand U22279 (N_22279,N_21723,N_21779);
or U22280 (N_22280,N_21887,N_21828);
or U22281 (N_22281,N_21612,N_21585);
nand U22282 (N_22282,N_21521,N_21730);
or U22283 (N_22283,N_21581,N_21729);
nand U22284 (N_22284,N_21994,N_21790);
or U22285 (N_22285,N_21622,N_21528);
nor U22286 (N_22286,N_21744,N_21724);
or U22287 (N_22287,N_21561,N_21705);
or U22288 (N_22288,N_21687,N_21550);
nand U22289 (N_22289,N_21920,N_21660);
xnor U22290 (N_22290,N_21993,N_21931);
nand U22291 (N_22291,N_21765,N_21658);
or U22292 (N_22292,N_21627,N_21937);
and U22293 (N_22293,N_21881,N_21999);
and U22294 (N_22294,N_21858,N_21650);
nor U22295 (N_22295,N_21603,N_21755);
nand U22296 (N_22296,N_21530,N_21685);
nand U22297 (N_22297,N_21670,N_21614);
nand U22298 (N_22298,N_21992,N_21741);
nand U22299 (N_22299,N_21518,N_21560);
nand U22300 (N_22300,N_21715,N_21515);
xor U22301 (N_22301,N_21516,N_21945);
xor U22302 (N_22302,N_21609,N_21728);
and U22303 (N_22303,N_21843,N_21564);
xnor U22304 (N_22304,N_21693,N_21680);
xor U22305 (N_22305,N_21550,N_21875);
or U22306 (N_22306,N_21969,N_21706);
xor U22307 (N_22307,N_21541,N_21761);
xnor U22308 (N_22308,N_21534,N_21847);
and U22309 (N_22309,N_21767,N_21687);
or U22310 (N_22310,N_21525,N_21899);
or U22311 (N_22311,N_21765,N_21779);
nor U22312 (N_22312,N_21886,N_21881);
nand U22313 (N_22313,N_21637,N_21613);
or U22314 (N_22314,N_21601,N_21985);
nand U22315 (N_22315,N_21569,N_21832);
nand U22316 (N_22316,N_21502,N_21955);
xor U22317 (N_22317,N_21753,N_21621);
and U22318 (N_22318,N_21861,N_21819);
xor U22319 (N_22319,N_21908,N_21807);
nor U22320 (N_22320,N_21895,N_21543);
nor U22321 (N_22321,N_21542,N_21733);
and U22322 (N_22322,N_21954,N_21847);
nor U22323 (N_22323,N_21751,N_21670);
nand U22324 (N_22324,N_21648,N_21780);
nand U22325 (N_22325,N_21949,N_21967);
or U22326 (N_22326,N_21820,N_21993);
xor U22327 (N_22327,N_21899,N_21698);
xor U22328 (N_22328,N_21537,N_21917);
xnor U22329 (N_22329,N_21773,N_21720);
and U22330 (N_22330,N_21858,N_21600);
or U22331 (N_22331,N_21613,N_21914);
nor U22332 (N_22332,N_21712,N_21511);
or U22333 (N_22333,N_21868,N_21908);
xor U22334 (N_22334,N_21868,N_21832);
or U22335 (N_22335,N_21643,N_21795);
and U22336 (N_22336,N_21714,N_21816);
nor U22337 (N_22337,N_21851,N_21854);
and U22338 (N_22338,N_21787,N_21954);
or U22339 (N_22339,N_21989,N_21764);
nand U22340 (N_22340,N_21761,N_21768);
and U22341 (N_22341,N_21645,N_21879);
nand U22342 (N_22342,N_21718,N_21683);
nor U22343 (N_22343,N_21589,N_21541);
nand U22344 (N_22344,N_21647,N_21558);
or U22345 (N_22345,N_21573,N_21629);
nor U22346 (N_22346,N_21643,N_21978);
xnor U22347 (N_22347,N_21795,N_21782);
nor U22348 (N_22348,N_21607,N_21653);
nor U22349 (N_22349,N_21565,N_21721);
nor U22350 (N_22350,N_21718,N_21598);
xor U22351 (N_22351,N_21775,N_21729);
or U22352 (N_22352,N_21697,N_21554);
and U22353 (N_22353,N_21628,N_21733);
or U22354 (N_22354,N_21535,N_21539);
nor U22355 (N_22355,N_21540,N_21647);
or U22356 (N_22356,N_21802,N_21904);
and U22357 (N_22357,N_21748,N_21887);
xor U22358 (N_22358,N_21916,N_21869);
nand U22359 (N_22359,N_21509,N_21850);
or U22360 (N_22360,N_21886,N_21664);
and U22361 (N_22361,N_21544,N_21968);
nor U22362 (N_22362,N_21597,N_21572);
and U22363 (N_22363,N_21953,N_21619);
and U22364 (N_22364,N_21648,N_21615);
or U22365 (N_22365,N_21623,N_21708);
and U22366 (N_22366,N_21753,N_21592);
xnor U22367 (N_22367,N_21525,N_21979);
xor U22368 (N_22368,N_21559,N_21528);
nor U22369 (N_22369,N_21817,N_21671);
nor U22370 (N_22370,N_21997,N_21906);
nor U22371 (N_22371,N_21691,N_21634);
and U22372 (N_22372,N_21679,N_21991);
nor U22373 (N_22373,N_21704,N_21858);
or U22374 (N_22374,N_21854,N_21573);
nand U22375 (N_22375,N_21916,N_21817);
nor U22376 (N_22376,N_21699,N_21708);
or U22377 (N_22377,N_21887,N_21655);
xor U22378 (N_22378,N_21959,N_21746);
xor U22379 (N_22379,N_21920,N_21767);
or U22380 (N_22380,N_21639,N_21888);
and U22381 (N_22381,N_21546,N_21929);
xnor U22382 (N_22382,N_21804,N_21696);
nor U22383 (N_22383,N_21593,N_21898);
or U22384 (N_22384,N_21627,N_21677);
nor U22385 (N_22385,N_21784,N_21979);
and U22386 (N_22386,N_21597,N_21688);
nand U22387 (N_22387,N_21734,N_21840);
nor U22388 (N_22388,N_21568,N_21522);
nand U22389 (N_22389,N_21537,N_21914);
xnor U22390 (N_22390,N_21708,N_21569);
and U22391 (N_22391,N_21647,N_21631);
and U22392 (N_22392,N_21641,N_21674);
nand U22393 (N_22393,N_21825,N_21858);
nand U22394 (N_22394,N_21904,N_21523);
and U22395 (N_22395,N_21546,N_21524);
nor U22396 (N_22396,N_21998,N_21994);
nor U22397 (N_22397,N_21731,N_21860);
xor U22398 (N_22398,N_21705,N_21584);
and U22399 (N_22399,N_21635,N_21572);
and U22400 (N_22400,N_21774,N_21536);
nor U22401 (N_22401,N_21990,N_21509);
or U22402 (N_22402,N_21685,N_21879);
nor U22403 (N_22403,N_21516,N_21724);
nand U22404 (N_22404,N_21845,N_21784);
and U22405 (N_22405,N_21735,N_21880);
and U22406 (N_22406,N_21587,N_21938);
xor U22407 (N_22407,N_21712,N_21810);
nor U22408 (N_22408,N_21992,N_21909);
xnor U22409 (N_22409,N_21561,N_21594);
nor U22410 (N_22410,N_21760,N_21978);
nor U22411 (N_22411,N_21605,N_21679);
or U22412 (N_22412,N_21666,N_21662);
nand U22413 (N_22413,N_21529,N_21591);
nand U22414 (N_22414,N_21776,N_21849);
and U22415 (N_22415,N_21618,N_21801);
and U22416 (N_22416,N_21836,N_21503);
nand U22417 (N_22417,N_21873,N_21654);
nand U22418 (N_22418,N_21971,N_21716);
and U22419 (N_22419,N_21799,N_21653);
or U22420 (N_22420,N_21570,N_21948);
and U22421 (N_22421,N_21834,N_21783);
and U22422 (N_22422,N_21578,N_21709);
nand U22423 (N_22423,N_21793,N_21833);
nand U22424 (N_22424,N_21582,N_21719);
xor U22425 (N_22425,N_21911,N_21714);
xor U22426 (N_22426,N_21558,N_21545);
or U22427 (N_22427,N_21893,N_21960);
xnor U22428 (N_22428,N_21639,N_21933);
nand U22429 (N_22429,N_21749,N_21573);
nand U22430 (N_22430,N_21718,N_21804);
xor U22431 (N_22431,N_21932,N_21921);
nor U22432 (N_22432,N_21841,N_21887);
nor U22433 (N_22433,N_21508,N_21690);
and U22434 (N_22434,N_21548,N_21536);
or U22435 (N_22435,N_21500,N_21958);
xor U22436 (N_22436,N_21926,N_21852);
nand U22437 (N_22437,N_21913,N_21727);
nand U22438 (N_22438,N_21984,N_21550);
or U22439 (N_22439,N_21725,N_21980);
or U22440 (N_22440,N_21915,N_21526);
nor U22441 (N_22441,N_21977,N_21728);
and U22442 (N_22442,N_21795,N_21822);
or U22443 (N_22443,N_21572,N_21708);
nand U22444 (N_22444,N_21941,N_21945);
nor U22445 (N_22445,N_21802,N_21571);
nand U22446 (N_22446,N_21507,N_21797);
nor U22447 (N_22447,N_21907,N_21710);
nor U22448 (N_22448,N_21616,N_21973);
nor U22449 (N_22449,N_21874,N_21943);
or U22450 (N_22450,N_21671,N_21541);
or U22451 (N_22451,N_21956,N_21864);
and U22452 (N_22452,N_21593,N_21699);
nor U22453 (N_22453,N_21585,N_21707);
and U22454 (N_22454,N_21802,N_21972);
nor U22455 (N_22455,N_21528,N_21982);
and U22456 (N_22456,N_21609,N_21642);
xnor U22457 (N_22457,N_21582,N_21983);
nand U22458 (N_22458,N_21713,N_21890);
or U22459 (N_22459,N_21794,N_21603);
or U22460 (N_22460,N_21801,N_21525);
and U22461 (N_22461,N_21544,N_21881);
or U22462 (N_22462,N_21622,N_21518);
nor U22463 (N_22463,N_21874,N_21618);
nand U22464 (N_22464,N_21804,N_21856);
and U22465 (N_22465,N_21756,N_21940);
or U22466 (N_22466,N_21996,N_21592);
xor U22467 (N_22467,N_21777,N_21522);
nor U22468 (N_22468,N_21884,N_21684);
and U22469 (N_22469,N_21844,N_21598);
nand U22470 (N_22470,N_21603,N_21645);
or U22471 (N_22471,N_21576,N_21698);
xnor U22472 (N_22472,N_21714,N_21896);
nand U22473 (N_22473,N_21859,N_21767);
and U22474 (N_22474,N_21931,N_21975);
xor U22475 (N_22475,N_21923,N_21843);
nand U22476 (N_22476,N_21874,N_21945);
and U22477 (N_22477,N_21870,N_21897);
xor U22478 (N_22478,N_21824,N_21967);
xor U22479 (N_22479,N_21519,N_21787);
nor U22480 (N_22480,N_21920,N_21750);
or U22481 (N_22481,N_21743,N_21721);
nor U22482 (N_22482,N_21761,N_21834);
nand U22483 (N_22483,N_21683,N_21785);
nor U22484 (N_22484,N_21642,N_21724);
or U22485 (N_22485,N_21526,N_21873);
nand U22486 (N_22486,N_21903,N_21883);
or U22487 (N_22487,N_21693,N_21899);
xor U22488 (N_22488,N_21706,N_21787);
nand U22489 (N_22489,N_21771,N_21542);
and U22490 (N_22490,N_21655,N_21653);
and U22491 (N_22491,N_21759,N_21863);
or U22492 (N_22492,N_21618,N_21746);
and U22493 (N_22493,N_21667,N_21703);
nand U22494 (N_22494,N_21910,N_21829);
nand U22495 (N_22495,N_21792,N_21709);
nand U22496 (N_22496,N_21764,N_21894);
nand U22497 (N_22497,N_21785,N_21626);
or U22498 (N_22498,N_21905,N_21600);
and U22499 (N_22499,N_21574,N_21543);
xnor U22500 (N_22500,N_22460,N_22031);
or U22501 (N_22501,N_22178,N_22052);
nand U22502 (N_22502,N_22427,N_22187);
xor U22503 (N_22503,N_22276,N_22199);
and U22504 (N_22504,N_22165,N_22195);
nor U22505 (N_22505,N_22074,N_22281);
nor U22506 (N_22506,N_22035,N_22134);
nand U22507 (N_22507,N_22216,N_22176);
nand U22508 (N_22508,N_22103,N_22426);
xnor U22509 (N_22509,N_22416,N_22497);
and U22510 (N_22510,N_22327,N_22136);
and U22511 (N_22511,N_22357,N_22262);
xnor U22512 (N_22512,N_22298,N_22405);
nand U22513 (N_22513,N_22459,N_22266);
or U22514 (N_22514,N_22450,N_22077);
nor U22515 (N_22515,N_22037,N_22108);
nand U22516 (N_22516,N_22062,N_22064);
or U22517 (N_22517,N_22294,N_22493);
or U22518 (N_22518,N_22182,N_22312);
nand U22519 (N_22519,N_22303,N_22481);
and U22520 (N_22520,N_22068,N_22209);
and U22521 (N_22521,N_22264,N_22353);
or U22522 (N_22522,N_22485,N_22058);
nand U22523 (N_22523,N_22235,N_22196);
xor U22524 (N_22524,N_22048,N_22275);
and U22525 (N_22525,N_22453,N_22192);
nor U22526 (N_22526,N_22226,N_22366);
or U22527 (N_22527,N_22398,N_22343);
and U22528 (N_22528,N_22401,N_22184);
xor U22529 (N_22529,N_22179,N_22468);
xnor U22530 (N_22530,N_22395,N_22040);
nor U22531 (N_22531,N_22297,N_22181);
nor U22532 (N_22532,N_22300,N_22149);
xnor U22533 (N_22533,N_22444,N_22081);
nor U22534 (N_22534,N_22095,N_22202);
or U22535 (N_22535,N_22307,N_22347);
and U22536 (N_22536,N_22162,N_22190);
xor U22537 (N_22537,N_22047,N_22364);
nand U22538 (N_22538,N_22396,N_22049);
and U22539 (N_22539,N_22213,N_22269);
or U22540 (N_22540,N_22145,N_22345);
xnor U22541 (N_22541,N_22334,N_22358);
xnor U22542 (N_22542,N_22492,N_22197);
nand U22543 (N_22543,N_22200,N_22194);
and U22544 (N_22544,N_22115,N_22311);
xor U22545 (N_22545,N_22024,N_22228);
and U22546 (N_22546,N_22191,N_22001);
xor U22547 (N_22547,N_22490,N_22105);
and U22548 (N_22548,N_22121,N_22158);
nand U22549 (N_22549,N_22137,N_22404);
nor U22550 (N_22550,N_22421,N_22154);
nor U22551 (N_22551,N_22270,N_22495);
nand U22552 (N_22552,N_22163,N_22113);
or U22553 (N_22553,N_22259,N_22032);
xnor U22554 (N_22554,N_22023,N_22221);
and U22555 (N_22555,N_22005,N_22310);
or U22556 (N_22556,N_22480,N_22333);
nor U22557 (N_22557,N_22377,N_22375);
nand U22558 (N_22558,N_22285,N_22146);
nand U22559 (N_22559,N_22189,N_22475);
and U22560 (N_22560,N_22484,N_22272);
or U22561 (N_22561,N_22252,N_22400);
xor U22562 (N_22562,N_22042,N_22373);
nor U22563 (N_22563,N_22329,N_22351);
xor U22564 (N_22564,N_22029,N_22284);
nor U22565 (N_22565,N_22044,N_22442);
xor U22566 (N_22566,N_22059,N_22314);
and U22567 (N_22567,N_22437,N_22063);
or U22568 (N_22568,N_22224,N_22286);
nor U22569 (N_22569,N_22099,N_22138);
nand U22570 (N_22570,N_22186,N_22390);
xor U22571 (N_22571,N_22229,N_22072);
nor U22572 (N_22572,N_22326,N_22458);
xnor U22573 (N_22573,N_22241,N_22243);
or U22574 (N_22574,N_22452,N_22087);
nand U22575 (N_22575,N_22340,N_22205);
xnor U22576 (N_22576,N_22466,N_22051);
or U22577 (N_22577,N_22217,N_22109);
and U22578 (N_22578,N_22467,N_22411);
and U22579 (N_22579,N_22282,N_22030);
and U22580 (N_22580,N_22443,N_22141);
xnor U22581 (N_22581,N_22096,N_22177);
nand U22582 (N_22582,N_22431,N_22295);
or U22583 (N_22583,N_22004,N_22389);
and U22584 (N_22584,N_22245,N_22370);
or U22585 (N_22585,N_22092,N_22082);
or U22586 (N_22586,N_22098,N_22006);
nand U22587 (N_22587,N_22150,N_22083);
and U22588 (N_22588,N_22265,N_22157);
nand U22589 (N_22589,N_22338,N_22362);
and U22590 (N_22590,N_22291,N_22316);
nor U22591 (N_22591,N_22139,N_22354);
nand U22592 (N_22592,N_22020,N_22382);
nand U22593 (N_22593,N_22477,N_22346);
and U22594 (N_22594,N_22323,N_22118);
and U22595 (N_22595,N_22449,N_22017);
or U22596 (N_22596,N_22424,N_22360);
xor U22597 (N_22597,N_22057,N_22003);
and U22598 (N_22598,N_22148,N_22432);
or U22599 (N_22599,N_22055,N_22361);
nor U22600 (N_22600,N_22129,N_22267);
xor U22601 (N_22601,N_22498,N_22408);
nand U22602 (N_22602,N_22188,N_22328);
or U22603 (N_22603,N_22406,N_22069);
nand U22604 (N_22604,N_22011,N_22412);
or U22605 (N_22605,N_22160,N_22420);
or U22606 (N_22606,N_22236,N_22341);
nand U22607 (N_22607,N_22487,N_22133);
xnor U22608 (N_22608,N_22026,N_22244);
or U22609 (N_22609,N_22293,N_22438);
nand U22610 (N_22610,N_22094,N_22218);
or U22611 (N_22611,N_22470,N_22451);
xnor U22612 (N_22612,N_22097,N_22014);
and U22613 (N_22613,N_22122,N_22039);
and U22614 (N_22614,N_22261,N_22463);
xor U22615 (N_22615,N_22240,N_22018);
nand U22616 (N_22616,N_22322,N_22385);
nor U22617 (N_22617,N_22499,N_22280);
nand U22618 (N_22618,N_22143,N_22309);
and U22619 (N_22619,N_22211,N_22397);
and U22620 (N_22620,N_22215,N_22388);
nor U22621 (N_22621,N_22394,N_22080);
and U22622 (N_22622,N_22234,N_22317);
nand U22623 (N_22623,N_22253,N_22491);
or U22624 (N_22624,N_22479,N_22016);
nand U22625 (N_22625,N_22287,N_22290);
and U22626 (N_22626,N_22367,N_22120);
or U22627 (N_22627,N_22066,N_22299);
nand U22628 (N_22628,N_22436,N_22445);
xnor U22629 (N_22629,N_22496,N_22379);
and U22630 (N_22630,N_22112,N_22075);
xor U22631 (N_22631,N_22156,N_22140);
xnor U22632 (N_22632,N_22000,N_22402);
nor U22633 (N_22633,N_22478,N_22247);
nor U22634 (N_22634,N_22117,N_22440);
or U22635 (N_22635,N_22413,N_22132);
xnor U22636 (N_22636,N_22337,N_22210);
nor U22637 (N_22637,N_22289,N_22170);
xnor U22638 (N_22638,N_22246,N_22474);
nor U22639 (N_22639,N_22387,N_22166);
nor U22640 (N_22640,N_22369,N_22242);
nor U22641 (N_22641,N_22447,N_22010);
or U22642 (N_22642,N_22230,N_22169);
nor U22643 (N_22643,N_22093,N_22255);
and U22644 (N_22644,N_22227,N_22473);
or U22645 (N_22645,N_22013,N_22414);
and U22646 (N_22646,N_22271,N_22292);
nor U22647 (N_22647,N_22464,N_22021);
nand U22648 (N_22648,N_22106,N_22356);
xor U22649 (N_22649,N_22116,N_22332);
nor U22650 (N_22650,N_22054,N_22482);
and U22651 (N_22651,N_22022,N_22283);
nor U22652 (N_22652,N_22131,N_22036);
or U22653 (N_22653,N_22012,N_22433);
xor U22654 (N_22654,N_22128,N_22041);
and U22655 (N_22655,N_22355,N_22315);
or U22656 (N_22656,N_22381,N_22008);
and U22657 (N_22657,N_22119,N_22212);
or U22658 (N_22658,N_22208,N_22203);
xnor U22659 (N_22659,N_22277,N_22324);
and U22660 (N_22660,N_22167,N_22256);
and U22661 (N_22661,N_22331,N_22350);
xnor U22662 (N_22662,N_22222,N_22248);
and U22663 (N_22663,N_22465,N_22104);
xnor U22664 (N_22664,N_22274,N_22476);
or U22665 (N_22665,N_22446,N_22147);
nor U22666 (N_22666,N_22231,N_22407);
or U22667 (N_22667,N_22045,N_22254);
xnor U22668 (N_22668,N_22151,N_22110);
xnor U22669 (N_22669,N_22296,N_22383);
nand U22670 (N_22670,N_22378,N_22304);
xnor U22671 (N_22671,N_22391,N_22114);
nand U22672 (N_22672,N_22100,N_22376);
or U22673 (N_22673,N_22457,N_22027);
nor U22674 (N_22674,N_22441,N_22273);
nor U22675 (N_22675,N_22174,N_22403);
xor U22676 (N_22676,N_22089,N_22085);
xor U22677 (N_22677,N_22219,N_22056);
and U22678 (N_22678,N_22380,N_22258);
or U22679 (N_22679,N_22251,N_22086);
and U22680 (N_22680,N_22288,N_22159);
nor U22681 (N_22681,N_22015,N_22155);
or U22682 (N_22682,N_22130,N_22019);
or U22683 (N_22683,N_22392,N_22126);
nor U22684 (N_22684,N_22090,N_22125);
nor U22685 (N_22685,N_22263,N_22193);
and U22686 (N_22686,N_22384,N_22180);
or U22687 (N_22687,N_22306,N_22279);
or U22688 (N_22688,N_22409,N_22363);
nor U22689 (N_22689,N_22305,N_22164);
and U22690 (N_22690,N_22061,N_22428);
nor U22691 (N_22691,N_22342,N_22065);
and U22692 (N_22692,N_22489,N_22127);
or U22693 (N_22693,N_22321,N_22483);
nor U22694 (N_22694,N_22425,N_22239);
nor U22695 (N_22695,N_22073,N_22050);
nand U22696 (N_22696,N_22301,N_22025);
or U22697 (N_22697,N_22336,N_22223);
nand U22698 (N_22698,N_22260,N_22423);
xor U22699 (N_22699,N_22101,N_22007);
xor U22700 (N_22700,N_22207,N_22472);
nand U22701 (N_22701,N_22175,N_22198);
and U22702 (N_22702,N_22325,N_22319);
nor U22703 (N_22703,N_22371,N_22454);
and U22704 (N_22704,N_22456,N_22429);
xnor U22705 (N_22705,N_22318,N_22461);
xor U22706 (N_22706,N_22469,N_22002);
nor U22707 (N_22707,N_22250,N_22201);
or U22708 (N_22708,N_22372,N_22349);
or U22709 (N_22709,N_22183,N_22335);
nor U22710 (N_22710,N_22034,N_22173);
xnor U22711 (N_22711,N_22455,N_22232);
nor U22712 (N_22712,N_22278,N_22009);
nor U22713 (N_22713,N_22204,N_22257);
or U22714 (N_22714,N_22418,N_22344);
xor U22715 (N_22715,N_22434,N_22399);
nand U22716 (N_22716,N_22494,N_22225);
nand U22717 (N_22717,N_22107,N_22206);
nor U22718 (N_22718,N_22320,N_22365);
nor U22719 (N_22719,N_22144,N_22070);
nand U22720 (N_22720,N_22471,N_22033);
xnor U22721 (N_22721,N_22417,N_22386);
nor U22722 (N_22722,N_22435,N_22268);
or U22723 (N_22723,N_22171,N_22043);
nor U22724 (N_22724,N_22168,N_22076);
and U22725 (N_22725,N_22102,N_22415);
nand U22726 (N_22726,N_22359,N_22124);
nand U22727 (N_22727,N_22462,N_22339);
nor U22728 (N_22728,N_22153,N_22123);
and U22729 (N_22729,N_22348,N_22308);
nand U22730 (N_22730,N_22046,N_22313);
nor U22731 (N_22731,N_22028,N_22053);
nor U22732 (N_22732,N_22060,N_22410);
or U22733 (N_22733,N_22368,N_22088);
nand U22734 (N_22734,N_22302,N_22185);
nand U22735 (N_22735,N_22038,N_22237);
xor U22736 (N_22736,N_22220,N_22152);
nand U22737 (N_22737,N_22439,N_22084);
xnor U22738 (N_22738,N_22172,N_22419);
or U22739 (N_22739,N_22422,N_22079);
xnor U22740 (N_22740,N_22161,N_22214);
or U22741 (N_22741,N_22078,N_22486);
and U22742 (N_22742,N_22067,N_22238);
nor U22743 (N_22743,N_22488,N_22448);
xor U22744 (N_22744,N_22142,N_22249);
or U22745 (N_22745,N_22135,N_22091);
or U22746 (N_22746,N_22374,N_22071);
nand U22747 (N_22747,N_22352,N_22330);
nand U22748 (N_22748,N_22430,N_22111);
nor U22749 (N_22749,N_22393,N_22233);
xnor U22750 (N_22750,N_22324,N_22304);
or U22751 (N_22751,N_22268,N_22337);
and U22752 (N_22752,N_22246,N_22168);
and U22753 (N_22753,N_22090,N_22193);
nor U22754 (N_22754,N_22262,N_22121);
nand U22755 (N_22755,N_22312,N_22369);
nor U22756 (N_22756,N_22185,N_22362);
nand U22757 (N_22757,N_22272,N_22394);
nand U22758 (N_22758,N_22036,N_22178);
and U22759 (N_22759,N_22296,N_22180);
or U22760 (N_22760,N_22056,N_22362);
nor U22761 (N_22761,N_22370,N_22263);
nor U22762 (N_22762,N_22339,N_22303);
or U22763 (N_22763,N_22094,N_22409);
xor U22764 (N_22764,N_22077,N_22499);
or U22765 (N_22765,N_22175,N_22007);
nand U22766 (N_22766,N_22093,N_22042);
nor U22767 (N_22767,N_22289,N_22238);
and U22768 (N_22768,N_22174,N_22486);
and U22769 (N_22769,N_22190,N_22375);
nor U22770 (N_22770,N_22006,N_22274);
and U22771 (N_22771,N_22181,N_22164);
and U22772 (N_22772,N_22261,N_22329);
nand U22773 (N_22773,N_22179,N_22243);
nor U22774 (N_22774,N_22191,N_22015);
and U22775 (N_22775,N_22159,N_22419);
nand U22776 (N_22776,N_22245,N_22236);
xor U22777 (N_22777,N_22177,N_22384);
xnor U22778 (N_22778,N_22272,N_22212);
nor U22779 (N_22779,N_22196,N_22127);
nand U22780 (N_22780,N_22328,N_22026);
nor U22781 (N_22781,N_22300,N_22271);
xnor U22782 (N_22782,N_22086,N_22394);
nor U22783 (N_22783,N_22250,N_22238);
and U22784 (N_22784,N_22271,N_22281);
nand U22785 (N_22785,N_22317,N_22402);
nor U22786 (N_22786,N_22197,N_22051);
or U22787 (N_22787,N_22007,N_22420);
or U22788 (N_22788,N_22304,N_22143);
nand U22789 (N_22789,N_22320,N_22035);
nand U22790 (N_22790,N_22369,N_22392);
nand U22791 (N_22791,N_22093,N_22214);
xor U22792 (N_22792,N_22078,N_22093);
nor U22793 (N_22793,N_22197,N_22373);
or U22794 (N_22794,N_22132,N_22170);
xor U22795 (N_22795,N_22217,N_22145);
nor U22796 (N_22796,N_22469,N_22400);
or U22797 (N_22797,N_22425,N_22144);
nand U22798 (N_22798,N_22169,N_22346);
and U22799 (N_22799,N_22129,N_22209);
nor U22800 (N_22800,N_22460,N_22418);
or U22801 (N_22801,N_22172,N_22313);
nor U22802 (N_22802,N_22179,N_22155);
nor U22803 (N_22803,N_22493,N_22243);
and U22804 (N_22804,N_22033,N_22066);
and U22805 (N_22805,N_22318,N_22247);
nand U22806 (N_22806,N_22303,N_22497);
and U22807 (N_22807,N_22240,N_22272);
xor U22808 (N_22808,N_22087,N_22055);
or U22809 (N_22809,N_22020,N_22168);
or U22810 (N_22810,N_22185,N_22162);
or U22811 (N_22811,N_22443,N_22451);
nand U22812 (N_22812,N_22487,N_22329);
nor U22813 (N_22813,N_22444,N_22489);
nor U22814 (N_22814,N_22205,N_22478);
and U22815 (N_22815,N_22344,N_22450);
nand U22816 (N_22816,N_22128,N_22203);
nand U22817 (N_22817,N_22207,N_22491);
nor U22818 (N_22818,N_22071,N_22171);
and U22819 (N_22819,N_22199,N_22092);
and U22820 (N_22820,N_22214,N_22353);
xor U22821 (N_22821,N_22222,N_22179);
or U22822 (N_22822,N_22060,N_22250);
nand U22823 (N_22823,N_22388,N_22223);
nor U22824 (N_22824,N_22160,N_22090);
nor U22825 (N_22825,N_22299,N_22256);
nor U22826 (N_22826,N_22044,N_22413);
and U22827 (N_22827,N_22249,N_22021);
xor U22828 (N_22828,N_22421,N_22160);
nor U22829 (N_22829,N_22093,N_22038);
or U22830 (N_22830,N_22092,N_22090);
and U22831 (N_22831,N_22346,N_22359);
or U22832 (N_22832,N_22154,N_22116);
nand U22833 (N_22833,N_22466,N_22141);
nor U22834 (N_22834,N_22322,N_22035);
or U22835 (N_22835,N_22135,N_22303);
or U22836 (N_22836,N_22283,N_22486);
nor U22837 (N_22837,N_22309,N_22130);
nand U22838 (N_22838,N_22407,N_22055);
or U22839 (N_22839,N_22387,N_22389);
xnor U22840 (N_22840,N_22398,N_22191);
or U22841 (N_22841,N_22301,N_22396);
or U22842 (N_22842,N_22382,N_22120);
nand U22843 (N_22843,N_22027,N_22489);
or U22844 (N_22844,N_22496,N_22348);
or U22845 (N_22845,N_22406,N_22015);
nor U22846 (N_22846,N_22360,N_22370);
and U22847 (N_22847,N_22412,N_22121);
nand U22848 (N_22848,N_22042,N_22036);
or U22849 (N_22849,N_22340,N_22075);
nor U22850 (N_22850,N_22491,N_22184);
nand U22851 (N_22851,N_22211,N_22258);
xor U22852 (N_22852,N_22001,N_22214);
xor U22853 (N_22853,N_22188,N_22210);
and U22854 (N_22854,N_22445,N_22143);
and U22855 (N_22855,N_22006,N_22324);
nor U22856 (N_22856,N_22427,N_22249);
xor U22857 (N_22857,N_22400,N_22056);
nand U22858 (N_22858,N_22260,N_22192);
nor U22859 (N_22859,N_22256,N_22099);
nor U22860 (N_22860,N_22357,N_22336);
and U22861 (N_22861,N_22141,N_22200);
xor U22862 (N_22862,N_22093,N_22013);
and U22863 (N_22863,N_22218,N_22329);
or U22864 (N_22864,N_22377,N_22137);
xor U22865 (N_22865,N_22368,N_22341);
xnor U22866 (N_22866,N_22204,N_22455);
xnor U22867 (N_22867,N_22183,N_22151);
nor U22868 (N_22868,N_22463,N_22336);
nand U22869 (N_22869,N_22286,N_22299);
or U22870 (N_22870,N_22059,N_22296);
or U22871 (N_22871,N_22159,N_22145);
nand U22872 (N_22872,N_22262,N_22489);
xor U22873 (N_22873,N_22272,N_22385);
nor U22874 (N_22874,N_22078,N_22437);
or U22875 (N_22875,N_22185,N_22229);
nor U22876 (N_22876,N_22257,N_22267);
or U22877 (N_22877,N_22145,N_22157);
or U22878 (N_22878,N_22100,N_22243);
and U22879 (N_22879,N_22114,N_22312);
and U22880 (N_22880,N_22109,N_22180);
and U22881 (N_22881,N_22481,N_22050);
or U22882 (N_22882,N_22493,N_22142);
or U22883 (N_22883,N_22468,N_22294);
and U22884 (N_22884,N_22485,N_22176);
xor U22885 (N_22885,N_22403,N_22123);
nor U22886 (N_22886,N_22029,N_22105);
nand U22887 (N_22887,N_22058,N_22115);
and U22888 (N_22888,N_22079,N_22242);
xnor U22889 (N_22889,N_22168,N_22207);
and U22890 (N_22890,N_22434,N_22068);
nor U22891 (N_22891,N_22299,N_22017);
and U22892 (N_22892,N_22029,N_22426);
or U22893 (N_22893,N_22315,N_22212);
xor U22894 (N_22894,N_22050,N_22231);
or U22895 (N_22895,N_22282,N_22062);
and U22896 (N_22896,N_22436,N_22363);
nor U22897 (N_22897,N_22192,N_22144);
xor U22898 (N_22898,N_22352,N_22338);
and U22899 (N_22899,N_22257,N_22036);
and U22900 (N_22900,N_22168,N_22196);
nor U22901 (N_22901,N_22011,N_22460);
and U22902 (N_22902,N_22438,N_22369);
xor U22903 (N_22903,N_22372,N_22454);
xnor U22904 (N_22904,N_22199,N_22465);
and U22905 (N_22905,N_22319,N_22214);
xor U22906 (N_22906,N_22147,N_22284);
and U22907 (N_22907,N_22089,N_22017);
and U22908 (N_22908,N_22270,N_22345);
xor U22909 (N_22909,N_22081,N_22184);
or U22910 (N_22910,N_22284,N_22205);
or U22911 (N_22911,N_22446,N_22120);
xnor U22912 (N_22912,N_22212,N_22038);
and U22913 (N_22913,N_22440,N_22004);
or U22914 (N_22914,N_22319,N_22060);
nor U22915 (N_22915,N_22368,N_22096);
xor U22916 (N_22916,N_22479,N_22070);
or U22917 (N_22917,N_22187,N_22191);
xnor U22918 (N_22918,N_22142,N_22122);
and U22919 (N_22919,N_22281,N_22401);
nor U22920 (N_22920,N_22204,N_22317);
or U22921 (N_22921,N_22304,N_22481);
nor U22922 (N_22922,N_22198,N_22153);
and U22923 (N_22923,N_22181,N_22109);
and U22924 (N_22924,N_22454,N_22424);
nand U22925 (N_22925,N_22408,N_22440);
xnor U22926 (N_22926,N_22302,N_22469);
nand U22927 (N_22927,N_22361,N_22168);
or U22928 (N_22928,N_22167,N_22186);
or U22929 (N_22929,N_22006,N_22317);
nand U22930 (N_22930,N_22479,N_22451);
and U22931 (N_22931,N_22436,N_22137);
and U22932 (N_22932,N_22256,N_22396);
xnor U22933 (N_22933,N_22416,N_22065);
nand U22934 (N_22934,N_22083,N_22311);
and U22935 (N_22935,N_22126,N_22025);
nor U22936 (N_22936,N_22414,N_22149);
xnor U22937 (N_22937,N_22116,N_22430);
xnor U22938 (N_22938,N_22249,N_22048);
nand U22939 (N_22939,N_22193,N_22473);
xor U22940 (N_22940,N_22236,N_22184);
xnor U22941 (N_22941,N_22115,N_22238);
nor U22942 (N_22942,N_22237,N_22311);
or U22943 (N_22943,N_22034,N_22005);
nand U22944 (N_22944,N_22420,N_22324);
and U22945 (N_22945,N_22458,N_22166);
and U22946 (N_22946,N_22120,N_22314);
or U22947 (N_22947,N_22185,N_22188);
and U22948 (N_22948,N_22471,N_22377);
nor U22949 (N_22949,N_22452,N_22167);
or U22950 (N_22950,N_22206,N_22373);
and U22951 (N_22951,N_22386,N_22083);
nor U22952 (N_22952,N_22357,N_22035);
or U22953 (N_22953,N_22298,N_22362);
or U22954 (N_22954,N_22334,N_22410);
nand U22955 (N_22955,N_22136,N_22337);
nand U22956 (N_22956,N_22099,N_22307);
or U22957 (N_22957,N_22387,N_22411);
nor U22958 (N_22958,N_22250,N_22326);
xnor U22959 (N_22959,N_22342,N_22315);
or U22960 (N_22960,N_22408,N_22396);
nand U22961 (N_22961,N_22157,N_22400);
or U22962 (N_22962,N_22054,N_22090);
xor U22963 (N_22963,N_22279,N_22061);
xnor U22964 (N_22964,N_22162,N_22266);
nor U22965 (N_22965,N_22268,N_22055);
nand U22966 (N_22966,N_22350,N_22319);
nand U22967 (N_22967,N_22029,N_22251);
nor U22968 (N_22968,N_22272,N_22291);
nor U22969 (N_22969,N_22209,N_22455);
nor U22970 (N_22970,N_22218,N_22115);
nand U22971 (N_22971,N_22050,N_22234);
or U22972 (N_22972,N_22004,N_22176);
or U22973 (N_22973,N_22424,N_22225);
nor U22974 (N_22974,N_22263,N_22319);
xor U22975 (N_22975,N_22263,N_22159);
or U22976 (N_22976,N_22482,N_22167);
and U22977 (N_22977,N_22481,N_22057);
nor U22978 (N_22978,N_22282,N_22089);
and U22979 (N_22979,N_22280,N_22041);
nand U22980 (N_22980,N_22397,N_22479);
nor U22981 (N_22981,N_22439,N_22112);
nand U22982 (N_22982,N_22342,N_22351);
or U22983 (N_22983,N_22018,N_22160);
nand U22984 (N_22984,N_22085,N_22330);
nand U22985 (N_22985,N_22461,N_22346);
or U22986 (N_22986,N_22303,N_22413);
or U22987 (N_22987,N_22016,N_22481);
or U22988 (N_22988,N_22235,N_22217);
nand U22989 (N_22989,N_22128,N_22210);
nand U22990 (N_22990,N_22481,N_22418);
nor U22991 (N_22991,N_22244,N_22072);
nor U22992 (N_22992,N_22126,N_22463);
nor U22993 (N_22993,N_22131,N_22156);
nand U22994 (N_22994,N_22384,N_22350);
and U22995 (N_22995,N_22351,N_22449);
nand U22996 (N_22996,N_22445,N_22338);
nand U22997 (N_22997,N_22206,N_22382);
nor U22998 (N_22998,N_22381,N_22470);
nor U22999 (N_22999,N_22282,N_22468);
nor U23000 (N_23000,N_22916,N_22931);
nor U23001 (N_23001,N_22977,N_22814);
xor U23002 (N_23002,N_22504,N_22670);
nand U23003 (N_23003,N_22922,N_22564);
nor U23004 (N_23004,N_22799,N_22585);
or U23005 (N_23005,N_22894,N_22573);
nand U23006 (N_23006,N_22740,N_22618);
or U23007 (N_23007,N_22508,N_22808);
or U23008 (N_23008,N_22907,N_22654);
xnor U23009 (N_23009,N_22739,N_22596);
nand U23010 (N_23010,N_22592,N_22721);
or U23011 (N_23011,N_22978,N_22662);
or U23012 (N_23012,N_22974,N_22823);
xnor U23013 (N_23013,N_22925,N_22617);
or U23014 (N_23014,N_22555,N_22559);
or U23015 (N_23015,N_22593,N_22944);
nor U23016 (N_23016,N_22581,N_22598);
nor U23017 (N_23017,N_22970,N_22834);
and U23018 (N_23018,N_22983,N_22909);
xnor U23019 (N_23019,N_22973,N_22883);
or U23020 (N_23020,N_22805,N_22603);
and U23021 (N_23021,N_22719,N_22787);
or U23022 (N_23022,N_22958,N_22841);
nor U23023 (N_23023,N_22996,N_22887);
nand U23024 (N_23024,N_22888,N_22891);
nor U23025 (N_23025,N_22949,N_22824);
xor U23026 (N_23026,N_22660,N_22623);
or U23027 (N_23027,N_22532,N_22992);
nand U23028 (N_23028,N_22928,N_22956);
nand U23029 (N_23029,N_22994,N_22524);
nor U23030 (N_23030,N_22519,N_22906);
nor U23031 (N_23031,N_22648,N_22857);
and U23032 (N_23032,N_22747,N_22801);
nor U23033 (N_23033,N_22501,N_22579);
nor U23034 (N_23034,N_22578,N_22625);
and U23035 (N_23035,N_22976,N_22753);
or U23036 (N_23036,N_22845,N_22547);
xnor U23037 (N_23037,N_22981,N_22993);
xnor U23038 (N_23038,N_22512,N_22927);
nor U23039 (N_23039,N_22785,N_22873);
xor U23040 (N_23040,N_22899,N_22766);
xor U23041 (N_23041,N_22803,N_22557);
xor U23042 (N_23042,N_22545,N_22954);
or U23043 (N_23043,N_22836,N_22505);
nor U23044 (N_23044,N_22597,N_22879);
xnor U23045 (N_23045,N_22699,N_22571);
or U23046 (N_23046,N_22502,N_22852);
nor U23047 (N_23047,N_22762,N_22975);
nand U23048 (N_23048,N_22631,N_22950);
or U23049 (N_23049,N_22535,N_22847);
nor U23050 (N_23050,N_22797,N_22500);
nand U23051 (N_23051,N_22902,N_22506);
xor U23052 (N_23052,N_22689,N_22685);
xor U23053 (N_23053,N_22754,N_22751);
and U23054 (N_23054,N_22565,N_22589);
or U23055 (N_23055,N_22517,N_22688);
and U23056 (N_23056,N_22724,N_22793);
nor U23057 (N_23057,N_22668,N_22948);
nor U23058 (N_23058,N_22653,N_22742);
or U23059 (N_23059,N_22672,N_22734);
and U23060 (N_23060,N_22686,N_22576);
nand U23061 (N_23061,N_22520,N_22582);
or U23062 (N_23062,N_22764,N_22586);
xor U23063 (N_23063,N_22613,N_22715);
and U23064 (N_23064,N_22548,N_22733);
nand U23065 (N_23065,N_22650,N_22725);
xor U23066 (N_23066,N_22886,N_22628);
and U23067 (N_23067,N_22651,N_22730);
or U23068 (N_23068,N_22904,N_22806);
or U23069 (N_23069,N_22854,N_22601);
nor U23070 (N_23070,N_22630,N_22966);
nand U23071 (N_23071,N_22741,N_22683);
nor U23072 (N_23072,N_22553,N_22702);
nor U23073 (N_23073,N_22998,N_22809);
xor U23074 (N_23074,N_22963,N_22930);
and U23075 (N_23075,N_22777,N_22861);
nand U23076 (N_23076,N_22935,N_22720);
or U23077 (N_23077,N_22965,N_22835);
xnor U23078 (N_23078,N_22611,N_22726);
nand U23079 (N_23079,N_22876,N_22679);
nor U23080 (N_23080,N_22594,N_22633);
nand U23081 (N_23081,N_22591,N_22892);
or U23082 (N_23082,N_22771,N_22637);
nor U23083 (N_23083,N_22772,N_22760);
xor U23084 (N_23084,N_22829,N_22914);
and U23085 (N_23085,N_22953,N_22599);
xnor U23086 (N_23086,N_22526,N_22657);
and U23087 (N_23087,N_22911,N_22819);
nand U23088 (N_23088,N_22813,N_22577);
and U23089 (N_23089,N_22758,N_22756);
xnor U23090 (N_23090,N_22972,N_22540);
xnor U23091 (N_23091,N_22893,N_22515);
nand U23092 (N_23092,N_22776,N_22775);
or U23093 (N_23093,N_22929,N_22749);
xnor U23094 (N_23094,N_22624,N_22616);
and U23095 (N_23095,N_22794,N_22622);
and U23096 (N_23096,N_22995,N_22716);
or U23097 (N_23097,N_22846,N_22516);
and U23098 (N_23098,N_22574,N_22800);
nand U23099 (N_23099,N_22642,N_22736);
and U23100 (N_23100,N_22527,N_22712);
nor U23101 (N_23101,N_22900,N_22746);
and U23102 (N_23102,N_22737,N_22643);
nor U23103 (N_23103,N_22536,N_22587);
nor U23104 (N_23104,N_22681,N_22588);
nor U23105 (N_23105,N_22752,N_22757);
xor U23106 (N_23106,N_22735,N_22853);
nand U23107 (N_23107,N_22684,N_22881);
and U23108 (N_23108,N_22696,N_22869);
xor U23109 (N_23109,N_22901,N_22868);
nand U23110 (N_23110,N_22666,N_22743);
and U23111 (N_23111,N_22945,N_22695);
nor U23112 (N_23112,N_22850,N_22678);
nor U23113 (N_23113,N_22838,N_22626);
or U23114 (N_23114,N_22882,N_22698);
nand U23115 (N_23115,N_22534,N_22822);
nand U23116 (N_23116,N_22700,N_22768);
nand U23117 (N_23117,N_22529,N_22862);
nor U23118 (N_23118,N_22844,N_22833);
xor U23119 (N_23119,N_22595,N_22513);
nand U23120 (N_23120,N_22874,N_22703);
xnor U23121 (N_23121,N_22788,N_22908);
nand U23122 (N_23122,N_22658,N_22632);
and U23123 (N_23123,N_22872,N_22986);
xnor U23124 (N_23124,N_22544,N_22912);
nor U23125 (N_23125,N_22647,N_22608);
nor U23126 (N_23126,N_22522,N_22665);
or U23127 (N_23127,N_22708,N_22942);
xnor U23128 (N_23128,N_22825,N_22773);
nor U23129 (N_23129,N_22732,N_22523);
nor U23130 (N_23130,N_22566,N_22980);
xor U23131 (N_23131,N_22820,N_22810);
and U23132 (N_23132,N_22690,N_22731);
and U23133 (N_23133,N_22755,N_22982);
or U23134 (N_23134,N_22895,N_22877);
xor U23135 (N_23135,N_22960,N_22843);
and U23136 (N_23136,N_22568,N_22584);
nand U23137 (N_23137,N_22832,N_22934);
and U23138 (N_23138,N_22604,N_22723);
or U23139 (N_23139,N_22811,N_22765);
nor U23140 (N_23140,N_22661,N_22827);
or U23141 (N_23141,N_22563,N_22514);
xnor U23142 (N_23142,N_22783,N_22807);
and U23143 (N_23143,N_22851,N_22826);
nand U23144 (N_23144,N_22656,N_22962);
nand U23145 (N_23145,N_22542,N_22669);
xor U23146 (N_23146,N_22748,N_22717);
nand U23147 (N_23147,N_22615,N_22667);
and U23148 (N_23148,N_22525,N_22614);
nand U23149 (N_23149,N_22511,N_22562);
and U23150 (N_23150,N_22636,N_22786);
nand U23151 (N_23151,N_22990,N_22521);
xnor U23152 (N_23152,N_22779,N_22884);
nor U23153 (N_23153,N_22691,N_22933);
nor U23154 (N_23154,N_22609,N_22959);
xor U23155 (N_23155,N_22984,N_22940);
nand U23156 (N_23156,N_22641,N_22759);
or U23157 (N_23157,N_22761,N_22727);
and U23158 (N_23158,N_22745,N_22898);
or U23159 (N_23159,N_22859,N_22664);
and U23160 (N_23160,N_22750,N_22946);
xnor U23161 (N_23161,N_22556,N_22644);
xor U23162 (N_23162,N_22863,N_22957);
and U23163 (N_23163,N_22640,N_22804);
and U23164 (N_23164,N_22921,N_22938);
nor U23165 (N_23165,N_22999,N_22896);
and U23166 (N_23166,N_22817,N_22952);
xnor U23167 (N_23167,N_22697,N_22509);
nor U23168 (N_23168,N_22989,N_22575);
nor U23169 (N_23169,N_22769,N_22780);
and U23170 (N_23170,N_22590,N_22729);
nor U23171 (N_23171,N_22791,N_22839);
xnor U23172 (N_23172,N_22570,N_22558);
and U23173 (N_23173,N_22913,N_22533);
and U23174 (N_23174,N_22692,N_22767);
nand U23175 (N_23175,N_22580,N_22530);
nand U23176 (N_23176,N_22627,N_22537);
and U23177 (N_23177,N_22890,N_22943);
nand U23178 (N_23178,N_22680,N_22828);
and U23179 (N_23179,N_22987,N_22655);
nor U23180 (N_23180,N_22812,N_22612);
nand U23181 (N_23181,N_22837,N_22961);
xnor U23182 (N_23182,N_22905,N_22889);
and U23183 (N_23183,N_22718,N_22583);
and U23184 (N_23184,N_22561,N_22936);
xor U23185 (N_23185,N_22560,N_22781);
xor U23186 (N_23186,N_22546,N_22967);
nand U23187 (N_23187,N_22802,N_22714);
and U23188 (N_23188,N_22864,N_22645);
nand U23189 (N_23189,N_22634,N_22652);
nand U23190 (N_23190,N_22503,N_22572);
or U23191 (N_23191,N_22932,N_22539);
or U23192 (N_23192,N_22855,N_22968);
xnor U23193 (N_23193,N_22705,N_22939);
or U23194 (N_23194,N_22738,N_22569);
or U23195 (N_23195,N_22620,N_22988);
or U23196 (N_23196,N_22635,N_22518);
xor U23197 (N_23197,N_22600,N_22870);
or U23198 (N_23198,N_22510,N_22885);
nor U23199 (N_23199,N_22763,N_22795);
nor U23200 (N_23200,N_22677,N_22774);
nor U23201 (N_23201,N_22639,N_22842);
nor U23202 (N_23202,N_22796,N_22709);
nand U23203 (N_23203,N_22673,N_22567);
xnor U23204 (N_23204,N_22675,N_22997);
nand U23205 (N_23205,N_22674,N_22964);
nor U23206 (N_23206,N_22713,N_22971);
nor U23207 (N_23207,N_22784,N_22897);
or U23208 (N_23208,N_22638,N_22818);
or U23209 (N_23209,N_22924,N_22878);
nand U23210 (N_23210,N_22865,N_22858);
or U23211 (N_23211,N_22693,N_22849);
nor U23212 (N_23212,N_22552,N_22815);
nor U23213 (N_23213,N_22621,N_22947);
and U23214 (N_23214,N_22770,N_22605);
nand U23215 (N_23215,N_22543,N_22646);
xor U23216 (N_23216,N_22607,N_22682);
nand U23217 (N_23217,N_22711,N_22816);
nor U23218 (N_23218,N_22649,N_22676);
or U23219 (N_23219,N_22926,N_22528);
or U23220 (N_23220,N_22728,N_22871);
or U23221 (N_23221,N_22551,N_22550);
nand U23222 (N_23222,N_22923,N_22782);
or U23223 (N_23223,N_22985,N_22744);
nor U23224 (N_23224,N_22917,N_22710);
nor U23225 (N_23225,N_22790,N_22821);
nor U23226 (N_23226,N_22778,N_22918);
and U23227 (N_23227,N_22722,N_22554);
nor U23228 (N_23228,N_22602,N_22991);
or U23229 (N_23229,N_22866,N_22941);
and U23230 (N_23230,N_22848,N_22840);
and U23231 (N_23231,N_22659,N_22694);
nand U23232 (N_23232,N_22831,N_22937);
or U23233 (N_23233,N_22860,N_22538);
xnor U23234 (N_23234,N_22955,N_22910);
or U23235 (N_23235,N_22507,N_22707);
and U23236 (N_23236,N_22606,N_22798);
xnor U23237 (N_23237,N_22687,N_22629);
and U23238 (N_23238,N_22619,N_22792);
xnor U23239 (N_23239,N_22880,N_22920);
or U23240 (N_23240,N_22706,N_22830);
nor U23241 (N_23241,N_22867,N_22671);
and U23242 (N_23242,N_22701,N_22915);
and U23243 (N_23243,N_22663,N_22903);
xor U23244 (N_23244,N_22875,N_22789);
and U23245 (N_23245,N_22856,N_22541);
nand U23246 (N_23246,N_22919,N_22969);
xnor U23247 (N_23247,N_22549,N_22704);
nand U23248 (N_23248,N_22610,N_22979);
nor U23249 (N_23249,N_22951,N_22531);
and U23250 (N_23250,N_22748,N_22781);
nand U23251 (N_23251,N_22643,N_22755);
nand U23252 (N_23252,N_22895,N_22503);
nand U23253 (N_23253,N_22886,N_22833);
and U23254 (N_23254,N_22670,N_22877);
and U23255 (N_23255,N_22740,N_22880);
xor U23256 (N_23256,N_22564,N_22868);
nor U23257 (N_23257,N_22902,N_22684);
xnor U23258 (N_23258,N_22621,N_22597);
or U23259 (N_23259,N_22888,N_22796);
nand U23260 (N_23260,N_22995,N_22933);
nand U23261 (N_23261,N_22828,N_22810);
or U23262 (N_23262,N_22978,N_22624);
xor U23263 (N_23263,N_22764,N_22515);
nand U23264 (N_23264,N_22697,N_22714);
xnor U23265 (N_23265,N_22852,N_22929);
xnor U23266 (N_23266,N_22913,N_22794);
and U23267 (N_23267,N_22885,N_22779);
nor U23268 (N_23268,N_22978,N_22814);
nand U23269 (N_23269,N_22738,N_22733);
xor U23270 (N_23270,N_22849,N_22975);
nor U23271 (N_23271,N_22628,N_22907);
nor U23272 (N_23272,N_22625,N_22772);
nor U23273 (N_23273,N_22916,N_22614);
and U23274 (N_23274,N_22658,N_22816);
xnor U23275 (N_23275,N_22675,N_22689);
or U23276 (N_23276,N_22512,N_22513);
or U23277 (N_23277,N_22880,N_22733);
nor U23278 (N_23278,N_22741,N_22930);
or U23279 (N_23279,N_22748,N_22831);
or U23280 (N_23280,N_22544,N_22901);
nand U23281 (N_23281,N_22981,N_22913);
nand U23282 (N_23282,N_22747,N_22696);
or U23283 (N_23283,N_22655,N_22679);
nand U23284 (N_23284,N_22852,N_22689);
and U23285 (N_23285,N_22965,N_22928);
nand U23286 (N_23286,N_22761,N_22542);
xnor U23287 (N_23287,N_22552,N_22534);
xor U23288 (N_23288,N_22555,N_22905);
and U23289 (N_23289,N_22987,N_22986);
nor U23290 (N_23290,N_22841,N_22592);
xnor U23291 (N_23291,N_22976,N_22785);
xnor U23292 (N_23292,N_22927,N_22970);
or U23293 (N_23293,N_22932,N_22863);
xnor U23294 (N_23294,N_22941,N_22653);
or U23295 (N_23295,N_22779,N_22558);
xnor U23296 (N_23296,N_22751,N_22808);
xor U23297 (N_23297,N_22816,N_22565);
nor U23298 (N_23298,N_22937,N_22645);
xnor U23299 (N_23299,N_22951,N_22546);
nor U23300 (N_23300,N_22543,N_22680);
xor U23301 (N_23301,N_22979,N_22793);
xor U23302 (N_23302,N_22547,N_22583);
nand U23303 (N_23303,N_22828,N_22720);
and U23304 (N_23304,N_22789,N_22865);
xnor U23305 (N_23305,N_22613,N_22698);
xor U23306 (N_23306,N_22823,N_22772);
nor U23307 (N_23307,N_22513,N_22741);
or U23308 (N_23308,N_22917,N_22932);
and U23309 (N_23309,N_22513,N_22506);
and U23310 (N_23310,N_22948,N_22998);
nand U23311 (N_23311,N_22615,N_22751);
and U23312 (N_23312,N_22680,N_22970);
nor U23313 (N_23313,N_22514,N_22760);
nand U23314 (N_23314,N_22538,N_22810);
or U23315 (N_23315,N_22883,N_22684);
or U23316 (N_23316,N_22538,N_22691);
nand U23317 (N_23317,N_22632,N_22875);
or U23318 (N_23318,N_22693,N_22723);
nand U23319 (N_23319,N_22576,N_22642);
and U23320 (N_23320,N_22726,N_22505);
nor U23321 (N_23321,N_22990,N_22524);
nor U23322 (N_23322,N_22665,N_22919);
xnor U23323 (N_23323,N_22623,N_22679);
nand U23324 (N_23324,N_22678,N_22635);
nand U23325 (N_23325,N_22868,N_22591);
nor U23326 (N_23326,N_22858,N_22976);
nand U23327 (N_23327,N_22780,N_22574);
nand U23328 (N_23328,N_22621,N_22632);
nand U23329 (N_23329,N_22809,N_22660);
and U23330 (N_23330,N_22635,N_22655);
or U23331 (N_23331,N_22890,N_22871);
nor U23332 (N_23332,N_22937,N_22540);
nand U23333 (N_23333,N_22929,N_22635);
xnor U23334 (N_23334,N_22544,N_22888);
nand U23335 (N_23335,N_22960,N_22846);
and U23336 (N_23336,N_22731,N_22717);
nand U23337 (N_23337,N_22908,N_22563);
and U23338 (N_23338,N_22675,N_22938);
xnor U23339 (N_23339,N_22976,N_22834);
nand U23340 (N_23340,N_22817,N_22947);
nor U23341 (N_23341,N_22861,N_22782);
xor U23342 (N_23342,N_22780,N_22508);
and U23343 (N_23343,N_22832,N_22879);
nand U23344 (N_23344,N_22510,N_22508);
or U23345 (N_23345,N_22699,N_22634);
nor U23346 (N_23346,N_22694,N_22517);
nand U23347 (N_23347,N_22872,N_22530);
or U23348 (N_23348,N_22650,N_22538);
nand U23349 (N_23349,N_22642,N_22755);
xnor U23350 (N_23350,N_22740,N_22847);
nor U23351 (N_23351,N_22772,N_22789);
nand U23352 (N_23352,N_22541,N_22779);
nand U23353 (N_23353,N_22777,N_22638);
nor U23354 (N_23354,N_22930,N_22947);
or U23355 (N_23355,N_22777,N_22801);
nand U23356 (N_23356,N_22754,N_22933);
and U23357 (N_23357,N_22696,N_22691);
nor U23358 (N_23358,N_22843,N_22869);
nand U23359 (N_23359,N_22772,N_22906);
xor U23360 (N_23360,N_22551,N_22832);
xor U23361 (N_23361,N_22872,N_22949);
xor U23362 (N_23362,N_22992,N_22738);
xor U23363 (N_23363,N_22590,N_22993);
xnor U23364 (N_23364,N_22874,N_22810);
nand U23365 (N_23365,N_22722,N_22751);
and U23366 (N_23366,N_22589,N_22734);
xor U23367 (N_23367,N_22653,N_22566);
xor U23368 (N_23368,N_22776,N_22623);
or U23369 (N_23369,N_22763,N_22759);
nor U23370 (N_23370,N_22720,N_22577);
nand U23371 (N_23371,N_22757,N_22936);
nand U23372 (N_23372,N_22677,N_22771);
and U23373 (N_23373,N_22627,N_22799);
xor U23374 (N_23374,N_22713,N_22530);
nand U23375 (N_23375,N_22832,N_22725);
or U23376 (N_23376,N_22986,N_22781);
xor U23377 (N_23377,N_22726,N_22656);
and U23378 (N_23378,N_22626,N_22907);
or U23379 (N_23379,N_22553,N_22692);
nor U23380 (N_23380,N_22863,N_22980);
xor U23381 (N_23381,N_22541,N_22718);
or U23382 (N_23382,N_22927,N_22609);
and U23383 (N_23383,N_22763,N_22628);
nor U23384 (N_23384,N_22586,N_22961);
nand U23385 (N_23385,N_22740,N_22539);
nor U23386 (N_23386,N_22938,N_22995);
and U23387 (N_23387,N_22989,N_22828);
and U23388 (N_23388,N_22623,N_22692);
or U23389 (N_23389,N_22935,N_22703);
xor U23390 (N_23390,N_22598,N_22999);
or U23391 (N_23391,N_22878,N_22997);
or U23392 (N_23392,N_22503,N_22614);
nor U23393 (N_23393,N_22523,N_22718);
nand U23394 (N_23394,N_22589,N_22686);
nand U23395 (N_23395,N_22742,N_22667);
xor U23396 (N_23396,N_22532,N_22548);
nor U23397 (N_23397,N_22753,N_22692);
and U23398 (N_23398,N_22821,N_22686);
or U23399 (N_23399,N_22885,N_22636);
nor U23400 (N_23400,N_22710,N_22558);
and U23401 (N_23401,N_22771,N_22571);
nor U23402 (N_23402,N_22598,N_22514);
nor U23403 (N_23403,N_22899,N_22668);
or U23404 (N_23404,N_22737,N_22971);
and U23405 (N_23405,N_22570,N_22676);
nor U23406 (N_23406,N_22888,N_22929);
or U23407 (N_23407,N_22834,N_22722);
and U23408 (N_23408,N_22983,N_22518);
and U23409 (N_23409,N_22880,N_22689);
nand U23410 (N_23410,N_22770,N_22608);
nor U23411 (N_23411,N_22845,N_22576);
xor U23412 (N_23412,N_22717,N_22934);
nor U23413 (N_23413,N_22931,N_22848);
or U23414 (N_23414,N_22722,N_22985);
nor U23415 (N_23415,N_22860,N_22985);
xnor U23416 (N_23416,N_22590,N_22685);
xnor U23417 (N_23417,N_22824,N_22731);
and U23418 (N_23418,N_22517,N_22511);
nand U23419 (N_23419,N_22793,N_22541);
nor U23420 (N_23420,N_22643,N_22760);
xor U23421 (N_23421,N_22626,N_22503);
nor U23422 (N_23422,N_22745,N_22813);
or U23423 (N_23423,N_22532,N_22723);
and U23424 (N_23424,N_22601,N_22657);
xor U23425 (N_23425,N_22768,N_22608);
nor U23426 (N_23426,N_22938,N_22504);
xnor U23427 (N_23427,N_22683,N_22721);
or U23428 (N_23428,N_22821,N_22793);
or U23429 (N_23429,N_22806,N_22696);
or U23430 (N_23430,N_22520,N_22613);
or U23431 (N_23431,N_22640,N_22746);
or U23432 (N_23432,N_22753,N_22543);
and U23433 (N_23433,N_22597,N_22559);
nor U23434 (N_23434,N_22728,N_22536);
nand U23435 (N_23435,N_22588,N_22954);
and U23436 (N_23436,N_22592,N_22794);
xnor U23437 (N_23437,N_22945,N_22614);
or U23438 (N_23438,N_22608,N_22784);
xor U23439 (N_23439,N_22525,N_22596);
nand U23440 (N_23440,N_22986,N_22571);
nor U23441 (N_23441,N_22536,N_22746);
xnor U23442 (N_23442,N_22646,N_22619);
or U23443 (N_23443,N_22672,N_22881);
and U23444 (N_23444,N_22548,N_22895);
and U23445 (N_23445,N_22975,N_22946);
nor U23446 (N_23446,N_22671,N_22612);
and U23447 (N_23447,N_22679,N_22828);
or U23448 (N_23448,N_22674,N_22914);
nand U23449 (N_23449,N_22660,N_22931);
nor U23450 (N_23450,N_22798,N_22592);
and U23451 (N_23451,N_22724,N_22731);
xor U23452 (N_23452,N_22659,N_22538);
or U23453 (N_23453,N_22734,N_22632);
nand U23454 (N_23454,N_22519,N_22898);
nor U23455 (N_23455,N_22607,N_22654);
xnor U23456 (N_23456,N_22733,N_22796);
or U23457 (N_23457,N_22875,N_22716);
xnor U23458 (N_23458,N_22563,N_22990);
nand U23459 (N_23459,N_22548,N_22770);
and U23460 (N_23460,N_22613,N_22790);
nor U23461 (N_23461,N_22948,N_22766);
nand U23462 (N_23462,N_22629,N_22895);
nor U23463 (N_23463,N_22715,N_22824);
and U23464 (N_23464,N_22710,N_22789);
and U23465 (N_23465,N_22726,N_22755);
nand U23466 (N_23466,N_22695,N_22677);
xnor U23467 (N_23467,N_22850,N_22853);
nor U23468 (N_23468,N_22808,N_22602);
nand U23469 (N_23469,N_22646,N_22928);
xnor U23470 (N_23470,N_22911,N_22981);
xor U23471 (N_23471,N_22878,N_22934);
or U23472 (N_23472,N_22702,N_22776);
xor U23473 (N_23473,N_22990,N_22532);
nand U23474 (N_23474,N_22804,N_22974);
nor U23475 (N_23475,N_22934,N_22527);
nand U23476 (N_23476,N_22680,N_22749);
nand U23477 (N_23477,N_22702,N_22810);
and U23478 (N_23478,N_22785,N_22922);
and U23479 (N_23479,N_22648,N_22807);
xor U23480 (N_23480,N_22994,N_22860);
nor U23481 (N_23481,N_22594,N_22682);
nand U23482 (N_23482,N_22747,N_22554);
or U23483 (N_23483,N_22989,N_22592);
nand U23484 (N_23484,N_22646,N_22934);
and U23485 (N_23485,N_22637,N_22544);
or U23486 (N_23486,N_22979,N_22983);
nor U23487 (N_23487,N_22641,N_22655);
nand U23488 (N_23488,N_22640,N_22599);
xor U23489 (N_23489,N_22956,N_22896);
and U23490 (N_23490,N_22830,N_22723);
or U23491 (N_23491,N_22964,N_22734);
nand U23492 (N_23492,N_22891,N_22916);
and U23493 (N_23493,N_22865,N_22726);
and U23494 (N_23494,N_22749,N_22807);
or U23495 (N_23495,N_22550,N_22834);
or U23496 (N_23496,N_22905,N_22759);
nand U23497 (N_23497,N_22783,N_22718);
nor U23498 (N_23498,N_22718,N_22988);
and U23499 (N_23499,N_22700,N_22603);
or U23500 (N_23500,N_23109,N_23225);
xnor U23501 (N_23501,N_23024,N_23220);
or U23502 (N_23502,N_23296,N_23104);
xor U23503 (N_23503,N_23288,N_23447);
nor U23504 (N_23504,N_23073,N_23187);
nor U23505 (N_23505,N_23402,N_23097);
nor U23506 (N_23506,N_23072,N_23283);
xnor U23507 (N_23507,N_23486,N_23054);
or U23508 (N_23508,N_23184,N_23491);
and U23509 (N_23509,N_23102,N_23190);
nand U23510 (N_23510,N_23356,N_23274);
nor U23511 (N_23511,N_23131,N_23299);
nor U23512 (N_23512,N_23162,N_23132);
nor U23513 (N_23513,N_23223,N_23487);
nand U23514 (N_23514,N_23313,N_23485);
and U23515 (N_23515,N_23352,N_23361);
nor U23516 (N_23516,N_23284,N_23429);
nand U23517 (N_23517,N_23256,N_23069);
and U23518 (N_23518,N_23456,N_23366);
nor U23519 (N_23519,N_23037,N_23320);
and U23520 (N_23520,N_23202,N_23259);
and U23521 (N_23521,N_23114,N_23362);
nand U23522 (N_23522,N_23473,N_23492);
xnor U23523 (N_23523,N_23247,N_23345);
nand U23524 (N_23524,N_23413,N_23075);
nand U23525 (N_23525,N_23330,N_23423);
nor U23526 (N_23526,N_23198,N_23360);
and U23527 (N_23527,N_23390,N_23373);
and U23528 (N_23528,N_23101,N_23196);
nand U23529 (N_23529,N_23208,N_23448);
and U23530 (N_23530,N_23233,N_23269);
or U23531 (N_23531,N_23185,N_23482);
xnor U23532 (N_23532,N_23086,N_23125);
xor U23533 (N_23533,N_23410,N_23497);
nor U23534 (N_23534,N_23004,N_23213);
xor U23535 (N_23535,N_23389,N_23437);
and U23536 (N_23536,N_23239,N_23059);
nor U23537 (N_23537,N_23412,N_23050);
nor U23538 (N_23538,N_23401,N_23346);
and U23539 (N_23539,N_23297,N_23419);
nor U23540 (N_23540,N_23121,N_23280);
nand U23541 (N_23541,N_23182,N_23153);
nand U23542 (N_23542,N_23295,N_23078);
or U23543 (N_23543,N_23260,N_23065);
and U23544 (N_23544,N_23219,N_23234);
nand U23545 (N_23545,N_23082,N_23192);
xor U23546 (N_23546,N_23014,N_23355);
nor U23547 (N_23547,N_23146,N_23112);
or U23548 (N_23548,N_23304,N_23191);
or U23549 (N_23549,N_23285,N_23479);
nand U23550 (N_23550,N_23427,N_23206);
nand U23551 (N_23551,N_23480,N_23438);
xor U23552 (N_23552,N_23032,N_23110);
xnor U23553 (N_23553,N_23309,N_23431);
and U23554 (N_23554,N_23230,N_23221);
and U23555 (N_23555,N_23314,N_23042);
or U23556 (N_23556,N_23255,N_23106);
nor U23557 (N_23557,N_23012,N_23026);
or U23558 (N_23558,N_23426,N_23077);
nor U23559 (N_23559,N_23444,N_23264);
nand U23560 (N_23560,N_23216,N_23029);
or U23561 (N_23561,N_23325,N_23249);
nand U23562 (N_23562,N_23128,N_23009);
xor U23563 (N_23563,N_23094,N_23041);
and U23564 (N_23564,N_23393,N_23034);
nand U23565 (N_23565,N_23120,N_23115);
xor U23566 (N_23566,N_23087,N_23186);
xor U23567 (N_23567,N_23158,N_23375);
or U23568 (N_23568,N_23273,N_23167);
nor U23569 (N_23569,N_23489,N_23181);
nand U23570 (N_23570,N_23027,N_23145);
and U23571 (N_23571,N_23062,N_23048);
nand U23572 (N_23572,N_23481,N_23136);
nor U23573 (N_23573,N_23342,N_23380);
xnor U23574 (N_23574,N_23395,N_23416);
xnor U23575 (N_23575,N_23396,N_23047);
or U23576 (N_23576,N_23160,N_23147);
xnor U23577 (N_23577,N_23166,N_23323);
and U23578 (N_23578,N_23488,N_23333);
xor U23579 (N_23579,N_23460,N_23116);
and U23580 (N_23580,N_23122,N_23322);
or U23581 (N_23581,N_23270,N_23175);
xor U23582 (N_23582,N_23275,N_23326);
nor U23583 (N_23583,N_23250,N_23392);
nor U23584 (N_23584,N_23176,N_23040);
nand U23585 (N_23585,N_23126,N_23183);
nor U23586 (N_23586,N_23254,N_23263);
and U23587 (N_23587,N_23006,N_23081);
xor U23588 (N_23588,N_23237,N_23155);
nand U23589 (N_23589,N_23177,N_23033);
nor U23590 (N_23590,N_23312,N_23031);
or U23591 (N_23591,N_23432,N_23405);
xnor U23592 (N_23592,N_23007,N_23089);
nor U23593 (N_23593,N_23357,N_23408);
nand U23594 (N_23594,N_23088,N_23468);
nand U23595 (N_23595,N_23466,N_23194);
and U23596 (N_23596,N_23113,N_23002);
or U23597 (N_23597,N_23334,N_23134);
and U23598 (N_23598,N_23257,N_23303);
nand U23599 (N_23599,N_23052,N_23400);
and U23600 (N_23600,N_23328,N_23496);
nand U23601 (N_23601,N_23420,N_23241);
nor U23602 (N_23602,N_23246,N_23471);
nor U23603 (N_23603,N_23163,N_23058);
nor U23604 (N_23604,N_23051,N_23472);
xnor U23605 (N_23605,N_23200,N_23318);
nand U23606 (N_23606,N_23148,N_23119);
xor U23607 (N_23607,N_23368,N_23045);
and U23608 (N_23608,N_23203,N_23484);
or U23609 (N_23609,N_23080,N_23035);
nor U23610 (N_23610,N_23016,N_23343);
or U23611 (N_23611,N_23272,N_23067);
and U23612 (N_23612,N_23071,N_23316);
nand U23613 (N_23613,N_23229,N_23271);
or U23614 (N_23614,N_23324,N_23397);
xor U23615 (N_23615,N_23470,N_23238);
and U23616 (N_23616,N_23404,N_23363);
nor U23617 (N_23617,N_23372,N_23076);
nor U23618 (N_23618,N_23144,N_23474);
nand U23619 (N_23619,N_23387,N_23278);
and U23620 (N_23620,N_23302,N_23277);
or U23621 (N_23621,N_23476,N_23337);
nor U23622 (N_23622,N_23245,N_23243);
or U23623 (N_23623,N_23378,N_23056);
and U23624 (N_23624,N_23188,N_23382);
xor U23625 (N_23625,N_23193,N_23055);
and U23626 (N_23626,N_23399,N_23098);
nand U23627 (N_23627,N_23418,N_23061);
nor U23628 (N_23628,N_23025,N_23493);
nand U23629 (N_23629,N_23276,N_23150);
or U23630 (N_23630,N_23358,N_23329);
nand U23631 (N_23631,N_23411,N_23053);
or U23632 (N_23632,N_23107,N_23212);
xnor U23633 (N_23633,N_23123,N_23139);
nand U23634 (N_23634,N_23242,N_23178);
or U23635 (N_23635,N_23459,N_23317);
and U23636 (N_23636,N_23172,N_23407);
nand U23637 (N_23637,N_23261,N_23301);
and U23638 (N_23638,N_23453,N_23443);
nand U23639 (N_23639,N_23038,N_23279);
nor U23640 (N_23640,N_23371,N_23018);
nor U23641 (N_23641,N_23100,N_23341);
or U23642 (N_23642,N_23354,N_23209);
and U23643 (N_23643,N_23010,N_23044);
and U23644 (N_23644,N_23422,N_23462);
nor U23645 (N_23645,N_23290,N_23450);
and U23646 (N_23646,N_23099,N_23091);
xnor U23647 (N_23647,N_23461,N_23003);
or U23648 (N_23648,N_23327,N_23311);
nor U23649 (N_23649,N_23074,N_23282);
or U23650 (N_23650,N_23377,N_23335);
or U23651 (N_23651,N_23210,N_23036);
and U23652 (N_23652,N_23452,N_23179);
nor U23653 (N_23653,N_23173,N_23433);
xor U23654 (N_23654,N_23451,N_23068);
xnor U23655 (N_23655,N_23321,N_23490);
nand U23656 (N_23656,N_23300,N_23454);
and U23657 (N_23657,N_23103,N_23289);
xor U23658 (N_23658,N_23351,N_23201);
nor U23659 (N_23659,N_23475,N_23394);
nand U23660 (N_23660,N_23286,N_23359);
xnor U23661 (N_23661,N_23319,N_23463);
and U23662 (N_23662,N_23305,N_23469);
or U23663 (N_23663,N_23157,N_23159);
or U23664 (N_23664,N_23133,N_23066);
or U23665 (N_23665,N_23294,N_23298);
or U23666 (N_23666,N_23174,N_23215);
nand U23667 (N_23667,N_23436,N_23140);
or U23668 (N_23668,N_23046,N_23171);
and U23669 (N_23669,N_23258,N_23118);
xnor U23670 (N_23670,N_23268,N_23030);
and U23671 (N_23671,N_23434,N_23379);
or U23672 (N_23672,N_23374,N_23008);
xnor U23673 (N_23673,N_23415,N_23370);
or U23674 (N_23674,N_23070,N_23364);
and U23675 (N_23675,N_23265,N_23039);
xnor U23676 (N_23676,N_23331,N_23079);
nand U23677 (N_23677,N_23227,N_23266);
nand U23678 (N_23678,N_23465,N_23308);
and U23679 (N_23679,N_23214,N_23170);
nand U23680 (N_23680,N_23011,N_23442);
xnor U23681 (N_23681,N_23236,N_23001);
nor U23682 (N_23682,N_23483,N_23424);
nand U23683 (N_23683,N_23409,N_23154);
nand U23684 (N_23684,N_23398,N_23262);
and U23685 (N_23685,N_23307,N_23156);
xor U23686 (N_23686,N_23494,N_23083);
nand U23687 (N_23687,N_23127,N_23092);
nand U23688 (N_23688,N_23498,N_23417);
nor U23689 (N_23689,N_23207,N_23267);
nor U23690 (N_23690,N_23129,N_23152);
or U23691 (N_23691,N_23063,N_23199);
nor U23692 (N_23692,N_23446,N_23085);
nor U23693 (N_23693,N_23135,N_23478);
xnor U23694 (N_23694,N_23464,N_23332);
xnor U23695 (N_23695,N_23224,N_23228);
nand U23696 (N_23696,N_23151,N_23439);
nand U23697 (N_23697,N_23222,N_23365);
and U23698 (N_23698,N_23111,N_23391);
xor U23699 (N_23699,N_23138,N_23165);
and U23700 (N_23700,N_23414,N_23403);
and U23701 (N_23701,N_23457,N_23244);
and U23702 (N_23702,N_23441,N_23385);
nor U23703 (N_23703,N_23495,N_23093);
or U23704 (N_23704,N_23445,N_23381);
or U23705 (N_23705,N_23369,N_23240);
nand U23706 (N_23706,N_23435,N_23336);
xnor U23707 (N_23707,N_23440,N_23340);
or U23708 (N_23708,N_23353,N_23021);
or U23709 (N_23709,N_23057,N_23310);
or U23710 (N_23710,N_23020,N_23000);
xnor U23711 (N_23711,N_23350,N_23306);
and U23712 (N_23712,N_23291,N_23023);
nor U23713 (N_23713,N_23455,N_23060);
and U23714 (N_23714,N_23049,N_23384);
or U23715 (N_23715,N_23232,N_23425);
or U23716 (N_23716,N_23211,N_23252);
nand U23717 (N_23717,N_23204,N_23499);
and U23718 (N_23718,N_23137,N_23235);
nand U23719 (N_23719,N_23084,N_23281);
nor U23720 (N_23720,N_23458,N_23349);
nand U23721 (N_23721,N_23019,N_23164);
xnor U23722 (N_23722,N_23005,N_23406);
xnor U23723 (N_23723,N_23231,N_23217);
nand U23724 (N_23724,N_23017,N_23467);
nor U23725 (N_23725,N_23205,N_23130);
xnor U23726 (N_23726,N_23141,N_23095);
xnor U23727 (N_23727,N_23169,N_23226);
or U23728 (N_23728,N_23248,N_23108);
and U23729 (N_23729,N_23367,N_23388);
xor U23730 (N_23730,N_23096,N_23292);
nand U23731 (N_23731,N_23253,N_23043);
and U23732 (N_23732,N_23143,N_23477);
and U23733 (N_23733,N_23197,N_23218);
nor U23734 (N_23734,N_23347,N_23105);
nor U23735 (N_23735,N_23124,N_23428);
xor U23736 (N_23736,N_23090,N_23168);
nor U23737 (N_23737,N_23022,N_23195);
and U23738 (N_23738,N_23180,N_23142);
nand U23739 (N_23739,N_23287,N_23421);
and U23740 (N_23740,N_23251,N_23348);
and U23741 (N_23741,N_23339,N_23161);
and U23742 (N_23742,N_23064,N_23338);
or U23743 (N_23743,N_23383,N_23015);
xnor U23744 (N_23744,N_23117,N_23344);
nand U23745 (N_23745,N_23430,N_23149);
or U23746 (N_23746,N_23386,N_23013);
or U23747 (N_23747,N_23376,N_23028);
or U23748 (N_23748,N_23293,N_23315);
xnor U23749 (N_23749,N_23189,N_23449);
xor U23750 (N_23750,N_23079,N_23403);
or U23751 (N_23751,N_23242,N_23076);
or U23752 (N_23752,N_23142,N_23103);
or U23753 (N_23753,N_23397,N_23304);
or U23754 (N_23754,N_23068,N_23222);
or U23755 (N_23755,N_23112,N_23348);
nand U23756 (N_23756,N_23482,N_23476);
and U23757 (N_23757,N_23313,N_23387);
nor U23758 (N_23758,N_23285,N_23300);
nand U23759 (N_23759,N_23278,N_23330);
xor U23760 (N_23760,N_23431,N_23100);
xor U23761 (N_23761,N_23286,N_23422);
nor U23762 (N_23762,N_23084,N_23329);
nor U23763 (N_23763,N_23291,N_23246);
or U23764 (N_23764,N_23169,N_23222);
xor U23765 (N_23765,N_23121,N_23259);
or U23766 (N_23766,N_23413,N_23186);
xor U23767 (N_23767,N_23476,N_23166);
or U23768 (N_23768,N_23170,N_23105);
nor U23769 (N_23769,N_23489,N_23197);
nor U23770 (N_23770,N_23371,N_23281);
and U23771 (N_23771,N_23488,N_23167);
or U23772 (N_23772,N_23171,N_23376);
and U23773 (N_23773,N_23308,N_23491);
xor U23774 (N_23774,N_23230,N_23234);
nand U23775 (N_23775,N_23349,N_23006);
or U23776 (N_23776,N_23042,N_23423);
nor U23777 (N_23777,N_23042,N_23383);
xnor U23778 (N_23778,N_23384,N_23048);
and U23779 (N_23779,N_23488,N_23104);
and U23780 (N_23780,N_23255,N_23096);
nand U23781 (N_23781,N_23283,N_23015);
nor U23782 (N_23782,N_23488,N_23031);
nand U23783 (N_23783,N_23164,N_23313);
xnor U23784 (N_23784,N_23315,N_23335);
xor U23785 (N_23785,N_23358,N_23281);
nor U23786 (N_23786,N_23101,N_23329);
or U23787 (N_23787,N_23077,N_23261);
xor U23788 (N_23788,N_23369,N_23478);
nand U23789 (N_23789,N_23344,N_23318);
nor U23790 (N_23790,N_23014,N_23210);
or U23791 (N_23791,N_23361,N_23090);
nand U23792 (N_23792,N_23497,N_23031);
and U23793 (N_23793,N_23188,N_23402);
xnor U23794 (N_23794,N_23312,N_23051);
nand U23795 (N_23795,N_23438,N_23412);
nand U23796 (N_23796,N_23220,N_23463);
nor U23797 (N_23797,N_23129,N_23407);
or U23798 (N_23798,N_23331,N_23171);
xor U23799 (N_23799,N_23117,N_23047);
xor U23800 (N_23800,N_23003,N_23395);
or U23801 (N_23801,N_23062,N_23309);
nand U23802 (N_23802,N_23079,N_23064);
nand U23803 (N_23803,N_23057,N_23096);
xnor U23804 (N_23804,N_23421,N_23370);
and U23805 (N_23805,N_23310,N_23378);
nor U23806 (N_23806,N_23364,N_23462);
xnor U23807 (N_23807,N_23431,N_23274);
xnor U23808 (N_23808,N_23085,N_23498);
nor U23809 (N_23809,N_23358,N_23121);
xnor U23810 (N_23810,N_23223,N_23206);
or U23811 (N_23811,N_23254,N_23114);
and U23812 (N_23812,N_23172,N_23224);
nor U23813 (N_23813,N_23065,N_23436);
nand U23814 (N_23814,N_23029,N_23403);
nand U23815 (N_23815,N_23070,N_23202);
nand U23816 (N_23816,N_23047,N_23366);
or U23817 (N_23817,N_23357,N_23452);
xnor U23818 (N_23818,N_23312,N_23127);
and U23819 (N_23819,N_23408,N_23137);
and U23820 (N_23820,N_23119,N_23123);
nand U23821 (N_23821,N_23041,N_23301);
or U23822 (N_23822,N_23233,N_23496);
or U23823 (N_23823,N_23166,N_23295);
nor U23824 (N_23824,N_23261,N_23210);
nor U23825 (N_23825,N_23151,N_23488);
nand U23826 (N_23826,N_23146,N_23180);
and U23827 (N_23827,N_23474,N_23204);
nor U23828 (N_23828,N_23045,N_23003);
xnor U23829 (N_23829,N_23090,N_23212);
or U23830 (N_23830,N_23182,N_23253);
or U23831 (N_23831,N_23010,N_23401);
nor U23832 (N_23832,N_23310,N_23093);
xnor U23833 (N_23833,N_23304,N_23394);
xnor U23834 (N_23834,N_23032,N_23024);
and U23835 (N_23835,N_23085,N_23186);
nor U23836 (N_23836,N_23162,N_23464);
xnor U23837 (N_23837,N_23347,N_23206);
or U23838 (N_23838,N_23032,N_23066);
nor U23839 (N_23839,N_23070,N_23173);
xor U23840 (N_23840,N_23112,N_23310);
nand U23841 (N_23841,N_23022,N_23242);
nand U23842 (N_23842,N_23040,N_23057);
nor U23843 (N_23843,N_23010,N_23166);
xnor U23844 (N_23844,N_23159,N_23235);
nor U23845 (N_23845,N_23408,N_23199);
and U23846 (N_23846,N_23298,N_23096);
and U23847 (N_23847,N_23004,N_23173);
xor U23848 (N_23848,N_23282,N_23362);
and U23849 (N_23849,N_23458,N_23264);
or U23850 (N_23850,N_23193,N_23134);
or U23851 (N_23851,N_23248,N_23137);
and U23852 (N_23852,N_23382,N_23309);
nor U23853 (N_23853,N_23256,N_23272);
or U23854 (N_23854,N_23498,N_23375);
or U23855 (N_23855,N_23090,N_23281);
xor U23856 (N_23856,N_23121,N_23200);
nor U23857 (N_23857,N_23097,N_23404);
nand U23858 (N_23858,N_23325,N_23071);
xnor U23859 (N_23859,N_23257,N_23187);
and U23860 (N_23860,N_23226,N_23212);
and U23861 (N_23861,N_23227,N_23086);
xor U23862 (N_23862,N_23189,N_23284);
nand U23863 (N_23863,N_23307,N_23153);
xor U23864 (N_23864,N_23098,N_23349);
nand U23865 (N_23865,N_23133,N_23100);
nand U23866 (N_23866,N_23192,N_23123);
and U23867 (N_23867,N_23257,N_23217);
nor U23868 (N_23868,N_23063,N_23118);
or U23869 (N_23869,N_23366,N_23051);
xor U23870 (N_23870,N_23281,N_23470);
nand U23871 (N_23871,N_23093,N_23342);
nor U23872 (N_23872,N_23072,N_23354);
or U23873 (N_23873,N_23057,N_23371);
nor U23874 (N_23874,N_23345,N_23436);
xor U23875 (N_23875,N_23013,N_23168);
nand U23876 (N_23876,N_23415,N_23283);
xnor U23877 (N_23877,N_23139,N_23246);
or U23878 (N_23878,N_23039,N_23447);
nor U23879 (N_23879,N_23473,N_23124);
and U23880 (N_23880,N_23460,N_23440);
or U23881 (N_23881,N_23336,N_23495);
nor U23882 (N_23882,N_23486,N_23045);
and U23883 (N_23883,N_23137,N_23210);
and U23884 (N_23884,N_23471,N_23253);
and U23885 (N_23885,N_23167,N_23483);
and U23886 (N_23886,N_23324,N_23444);
xor U23887 (N_23887,N_23315,N_23032);
nand U23888 (N_23888,N_23230,N_23437);
nand U23889 (N_23889,N_23424,N_23201);
or U23890 (N_23890,N_23423,N_23202);
or U23891 (N_23891,N_23144,N_23422);
xnor U23892 (N_23892,N_23191,N_23342);
nand U23893 (N_23893,N_23462,N_23213);
and U23894 (N_23894,N_23056,N_23437);
and U23895 (N_23895,N_23483,N_23406);
or U23896 (N_23896,N_23449,N_23170);
and U23897 (N_23897,N_23192,N_23197);
xnor U23898 (N_23898,N_23393,N_23008);
xor U23899 (N_23899,N_23162,N_23253);
and U23900 (N_23900,N_23273,N_23109);
xor U23901 (N_23901,N_23044,N_23207);
nor U23902 (N_23902,N_23478,N_23448);
xor U23903 (N_23903,N_23168,N_23020);
and U23904 (N_23904,N_23198,N_23359);
nor U23905 (N_23905,N_23113,N_23164);
nor U23906 (N_23906,N_23283,N_23419);
and U23907 (N_23907,N_23104,N_23420);
and U23908 (N_23908,N_23384,N_23444);
or U23909 (N_23909,N_23221,N_23415);
or U23910 (N_23910,N_23342,N_23330);
xor U23911 (N_23911,N_23187,N_23371);
nand U23912 (N_23912,N_23182,N_23438);
or U23913 (N_23913,N_23464,N_23494);
nor U23914 (N_23914,N_23195,N_23475);
xnor U23915 (N_23915,N_23196,N_23245);
nor U23916 (N_23916,N_23230,N_23075);
xnor U23917 (N_23917,N_23194,N_23115);
xnor U23918 (N_23918,N_23209,N_23017);
nand U23919 (N_23919,N_23251,N_23318);
nor U23920 (N_23920,N_23353,N_23498);
or U23921 (N_23921,N_23372,N_23018);
or U23922 (N_23922,N_23261,N_23384);
and U23923 (N_23923,N_23317,N_23337);
and U23924 (N_23924,N_23476,N_23387);
xnor U23925 (N_23925,N_23080,N_23292);
or U23926 (N_23926,N_23352,N_23324);
or U23927 (N_23927,N_23469,N_23471);
or U23928 (N_23928,N_23166,N_23217);
nand U23929 (N_23929,N_23135,N_23233);
or U23930 (N_23930,N_23410,N_23419);
or U23931 (N_23931,N_23156,N_23414);
nand U23932 (N_23932,N_23433,N_23277);
nand U23933 (N_23933,N_23054,N_23296);
nor U23934 (N_23934,N_23076,N_23353);
xnor U23935 (N_23935,N_23314,N_23327);
nand U23936 (N_23936,N_23232,N_23402);
xor U23937 (N_23937,N_23211,N_23180);
nor U23938 (N_23938,N_23366,N_23314);
nor U23939 (N_23939,N_23271,N_23465);
nor U23940 (N_23940,N_23144,N_23473);
and U23941 (N_23941,N_23194,N_23028);
xor U23942 (N_23942,N_23448,N_23290);
xor U23943 (N_23943,N_23360,N_23340);
nand U23944 (N_23944,N_23294,N_23094);
xor U23945 (N_23945,N_23096,N_23243);
xor U23946 (N_23946,N_23332,N_23258);
nor U23947 (N_23947,N_23264,N_23450);
or U23948 (N_23948,N_23240,N_23487);
nor U23949 (N_23949,N_23083,N_23385);
nand U23950 (N_23950,N_23202,N_23067);
xnor U23951 (N_23951,N_23357,N_23100);
and U23952 (N_23952,N_23147,N_23081);
nand U23953 (N_23953,N_23432,N_23250);
or U23954 (N_23954,N_23308,N_23095);
nand U23955 (N_23955,N_23306,N_23144);
or U23956 (N_23956,N_23008,N_23014);
nand U23957 (N_23957,N_23197,N_23204);
nand U23958 (N_23958,N_23312,N_23039);
xor U23959 (N_23959,N_23270,N_23260);
nor U23960 (N_23960,N_23261,N_23457);
nand U23961 (N_23961,N_23039,N_23063);
nand U23962 (N_23962,N_23039,N_23419);
and U23963 (N_23963,N_23320,N_23030);
or U23964 (N_23964,N_23348,N_23497);
xnor U23965 (N_23965,N_23008,N_23076);
nand U23966 (N_23966,N_23218,N_23302);
nor U23967 (N_23967,N_23025,N_23115);
and U23968 (N_23968,N_23020,N_23455);
nand U23969 (N_23969,N_23463,N_23342);
or U23970 (N_23970,N_23342,N_23393);
nor U23971 (N_23971,N_23435,N_23137);
or U23972 (N_23972,N_23386,N_23104);
or U23973 (N_23973,N_23489,N_23461);
or U23974 (N_23974,N_23286,N_23063);
xnor U23975 (N_23975,N_23023,N_23216);
and U23976 (N_23976,N_23002,N_23326);
nand U23977 (N_23977,N_23303,N_23380);
xor U23978 (N_23978,N_23192,N_23201);
xor U23979 (N_23979,N_23117,N_23418);
and U23980 (N_23980,N_23422,N_23082);
nand U23981 (N_23981,N_23168,N_23014);
nand U23982 (N_23982,N_23218,N_23018);
or U23983 (N_23983,N_23373,N_23462);
nor U23984 (N_23984,N_23394,N_23087);
xor U23985 (N_23985,N_23142,N_23442);
nor U23986 (N_23986,N_23362,N_23107);
nor U23987 (N_23987,N_23331,N_23187);
xnor U23988 (N_23988,N_23245,N_23304);
nand U23989 (N_23989,N_23332,N_23090);
or U23990 (N_23990,N_23300,N_23135);
nor U23991 (N_23991,N_23125,N_23026);
or U23992 (N_23992,N_23126,N_23462);
nor U23993 (N_23993,N_23210,N_23414);
nor U23994 (N_23994,N_23399,N_23263);
or U23995 (N_23995,N_23002,N_23129);
xor U23996 (N_23996,N_23478,N_23205);
or U23997 (N_23997,N_23263,N_23325);
or U23998 (N_23998,N_23452,N_23037);
and U23999 (N_23999,N_23220,N_23312);
and U24000 (N_24000,N_23711,N_23900);
and U24001 (N_24001,N_23644,N_23662);
and U24002 (N_24002,N_23555,N_23932);
and U24003 (N_24003,N_23746,N_23905);
nand U24004 (N_24004,N_23933,N_23643);
nand U24005 (N_24005,N_23604,N_23530);
and U24006 (N_24006,N_23612,N_23901);
nor U24007 (N_24007,N_23969,N_23944);
nand U24008 (N_24008,N_23584,N_23910);
nand U24009 (N_24009,N_23947,N_23741);
or U24010 (N_24010,N_23852,N_23693);
and U24011 (N_24011,N_23809,N_23542);
nand U24012 (N_24012,N_23760,N_23864);
and U24013 (N_24013,N_23758,N_23548);
nand U24014 (N_24014,N_23841,N_23569);
or U24015 (N_24015,N_23583,N_23502);
nor U24016 (N_24016,N_23768,N_23810);
nor U24017 (N_24017,N_23788,N_23615);
nor U24018 (N_24018,N_23750,N_23642);
and U24019 (N_24019,N_23889,N_23505);
or U24020 (N_24020,N_23596,N_23704);
and U24021 (N_24021,N_23909,N_23576);
and U24022 (N_24022,N_23707,N_23560);
xor U24023 (N_24023,N_23582,N_23722);
or U24024 (N_24024,N_23580,N_23877);
or U24025 (N_24025,N_23970,N_23546);
nand U24026 (N_24026,N_23938,N_23949);
nand U24027 (N_24027,N_23640,N_23518);
nor U24028 (N_24028,N_23531,N_23708);
nor U24029 (N_24029,N_23975,N_23958);
and U24030 (N_24030,N_23766,N_23813);
nand U24031 (N_24031,N_23617,N_23748);
and U24032 (N_24032,N_23936,N_23562);
and U24033 (N_24033,N_23775,N_23902);
and U24034 (N_24034,N_23781,N_23802);
nand U24035 (N_24035,N_23669,N_23821);
xor U24036 (N_24036,N_23737,N_23656);
or U24037 (N_24037,N_23501,N_23872);
and U24038 (N_24038,N_23827,N_23745);
xnor U24039 (N_24039,N_23607,N_23687);
or U24040 (N_24040,N_23744,N_23719);
nand U24041 (N_24041,N_23620,N_23660);
and U24042 (N_24042,N_23538,N_23839);
nand U24043 (N_24043,N_23886,N_23843);
and U24044 (N_24044,N_23525,N_23913);
or U24045 (N_24045,N_23962,N_23982);
nor U24046 (N_24046,N_23819,N_23539);
nor U24047 (N_24047,N_23876,N_23753);
xnor U24048 (N_24048,N_23757,N_23606);
and U24049 (N_24049,N_23875,N_23641);
or U24050 (N_24050,N_23570,N_23694);
xnor U24051 (N_24051,N_23511,N_23890);
nand U24052 (N_24052,N_23684,N_23920);
or U24053 (N_24053,N_23586,N_23591);
and U24054 (N_24054,N_23808,N_23811);
xor U24055 (N_24055,N_23628,N_23903);
nor U24056 (N_24056,N_23537,N_23956);
nand U24057 (N_24057,N_23953,N_23714);
or U24058 (N_24058,N_23602,N_23697);
or U24059 (N_24059,N_23820,N_23510);
and U24060 (N_24060,N_23790,N_23836);
or U24061 (N_24061,N_23554,N_23850);
nand U24062 (N_24062,N_23859,N_23792);
xor U24063 (N_24063,N_23611,N_23624);
or U24064 (N_24064,N_23659,N_23838);
nor U24065 (N_24065,N_23559,N_23671);
nor U24066 (N_24066,N_23964,N_23732);
xor U24067 (N_24067,N_23655,N_23651);
or U24068 (N_24068,N_23565,N_23989);
nand U24069 (N_24069,N_23873,N_23908);
or U24070 (N_24070,N_23550,N_23778);
and U24071 (N_24071,N_23513,N_23921);
and U24072 (N_24072,N_23618,N_23541);
xnor U24073 (N_24073,N_23812,N_23817);
nor U24074 (N_24074,N_23833,N_23965);
xor U24075 (N_24075,N_23557,N_23725);
nand U24076 (N_24076,N_23540,N_23919);
nor U24077 (N_24077,N_23941,N_23828);
nand U24078 (N_24078,N_23629,N_23855);
nand U24079 (N_24079,N_23796,N_23634);
and U24080 (N_24080,N_23881,N_23930);
and U24081 (N_24081,N_23755,N_23705);
and U24082 (N_24082,N_23592,N_23623);
nor U24083 (N_24083,N_23619,N_23863);
or U24084 (N_24084,N_23912,N_23966);
nor U24085 (N_24085,N_23504,N_23779);
nand U24086 (N_24086,N_23625,N_23682);
or U24087 (N_24087,N_23955,N_23840);
and U24088 (N_24088,N_23514,N_23950);
nand U24089 (N_24089,N_23506,N_23916);
nor U24090 (N_24090,N_23922,N_23699);
and U24091 (N_24091,N_23545,N_23519);
xnor U24092 (N_24092,N_23782,N_23742);
or U24093 (N_24093,N_23767,N_23885);
nand U24094 (N_24094,N_23512,N_23552);
nor U24095 (N_24095,N_23971,N_23579);
or U24096 (N_24096,N_23526,N_23700);
xnor U24097 (N_24097,N_23516,N_23658);
xor U24098 (N_24098,N_23721,N_23581);
or U24099 (N_24099,N_23589,N_23981);
nand U24100 (N_24100,N_23603,N_23804);
xnor U24101 (N_24101,N_23897,N_23702);
or U24102 (N_24102,N_23980,N_23578);
nand U24103 (N_24103,N_23712,N_23977);
nor U24104 (N_24104,N_23769,N_23547);
and U24105 (N_24105,N_23923,N_23717);
or U24106 (N_24106,N_23567,N_23871);
nor U24107 (N_24107,N_23899,N_23785);
nor U24108 (N_24108,N_23799,N_23638);
nand U24109 (N_24109,N_23738,N_23904);
and U24110 (N_24110,N_23621,N_23993);
and U24111 (N_24111,N_23528,N_23880);
or U24112 (N_24112,N_23743,N_23637);
nand U24113 (N_24113,N_23566,N_23847);
nor U24114 (N_24114,N_23887,N_23690);
nor U24115 (N_24115,N_23544,N_23527);
and U24116 (N_24116,N_23730,N_23952);
and U24117 (N_24117,N_23801,N_23780);
nor U24118 (N_24118,N_23650,N_23927);
and U24119 (N_24119,N_23549,N_23984);
or U24120 (N_24120,N_23532,N_23815);
nand U24121 (N_24121,N_23853,N_23703);
or U24122 (N_24122,N_23696,N_23568);
nand U24123 (N_24123,N_23613,N_23600);
nand U24124 (N_24124,N_23635,N_23830);
xnor U24125 (N_24125,N_23798,N_23867);
nor U24126 (N_24126,N_23507,N_23595);
and U24127 (N_24127,N_23882,N_23848);
nor U24128 (N_24128,N_23729,N_23915);
nor U24129 (N_24129,N_23892,N_23879);
nor U24130 (N_24130,N_23783,N_23657);
nor U24131 (N_24131,N_23960,N_23670);
nand U24132 (N_24132,N_23898,N_23533);
nor U24133 (N_24133,N_23534,N_23961);
xnor U24134 (N_24134,N_23574,N_23990);
nor U24135 (N_24135,N_23529,N_23816);
or U24136 (N_24136,N_23866,N_23724);
xor U24137 (N_24137,N_23661,N_23939);
and U24138 (N_24138,N_23829,N_23503);
or U24139 (N_24139,N_23870,N_23926);
and U24140 (N_24140,N_23973,N_23771);
or U24141 (N_24141,N_23883,N_23614);
nand U24142 (N_24142,N_23807,N_23786);
xnor U24143 (N_24143,N_23972,N_23633);
nand U24144 (N_24144,N_23713,N_23826);
nor U24145 (N_24145,N_23718,N_23987);
and U24146 (N_24146,N_23665,N_23851);
and U24147 (N_24147,N_23627,N_23911);
xnor U24148 (N_24148,N_23951,N_23673);
nand U24149 (N_24149,N_23789,N_23692);
and U24150 (N_24150,N_23685,N_23677);
and U24151 (N_24151,N_23734,N_23945);
nor U24152 (N_24152,N_23543,N_23777);
and U24153 (N_24153,N_23608,N_23698);
xor U24154 (N_24154,N_23551,N_23998);
nand U24155 (N_24155,N_23822,N_23996);
nand U24156 (N_24156,N_23942,N_23818);
nor U24157 (N_24157,N_23861,N_23772);
xnor U24158 (N_24158,N_23649,N_23832);
nand U24159 (N_24159,N_23854,N_23935);
and U24160 (N_24160,N_23963,N_23868);
xnor U24161 (N_24161,N_23858,N_23636);
or U24162 (N_24162,N_23645,N_23837);
xnor U24163 (N_24163,N_23740,N_23934);
or U24164 (N_24164,N_23835,N_23857);
nand U24165 (N_24165,N_23598,N_23918);
xnor U24166 (N_24166,N_23917,N_23884);
xor U24167 (N_24167,N_23862,N_23577);
nor U24168 (N_24168,N_23731,N_23759);
and U24169 (N_24169,N_23986,N_23773);
nor U24170 (N_24170,N_23680,N_23626);
nor U24171 (N_24171,N_23794,N_23710);
xnor U24172 (N_24172,N_23701,N_23517);
and U24173 (N_24173,N_23594,N_23940);
nor U24174 (N_24174,N_23795,N_23959);
nor U24175 (N_24175,N_23667,N_23823);
xor U24176 (N_24176,N_23564,N_23834);
nand U24177 (N_24177,N_23558,N_23895);
and U24178 (N_24178,N_23985,N_23679);
nand U24179 (N_24179,N_23509,N_23686);
nor U24180 (N_24180,N_23522,N_23845);
and U24181 (N_24181,N_23979,N_23995);
and U24182 (N_24182,N_23556,N_23590);
nand U24183 (N_24183,N_23747,N_23695);
nor U24184 (N_24184,N_23846,N_23597);
or U24185 (N_24185,N_23793,N_23683);
or U24186 (N_24186,N_23653,N_23946);
nand U24187 (N_24187,N_23770,N_23508);
or U24188 (N_24188,N_23978,N_23948);
nand U24189 (N_24189,N_23844,N_23787);
or U24190 (N_24190,N_23865,N_23925);
nor U24191 (N_24191,N_23791,N_23761);
and U24192 (N_24192,N_23736,N_23929);
nand U24193 (N_24193,N_23974,N_23675);
nand U24194 (N_24194,N_23616,N_23756);
nor U24195 (N_24195,N_23869,N_23520);
and U24196 (N_24196,N_23954,N_23874);
or U24197 (N_24197,N_23575,N_23894);
or U24198 (N_24198,N_23733,N_23587);
and U24199 (N_24199,N_23924,N_23751);
or U24200 (N_24200,N_23967,N_23878);
nor U24201 (N_24201,N_23893,N_23535);
nor U24202 (N_24202,N_23776,N_23856);
nor U24203 (N_24203,N_23928,N_23676);
xnor U24204 (N_24204,N_23983,N_23739);
nand U24205 (N_24205,N_23914,N_23931);
xor U24206 (N_24206,N_23896,N_23521);
nor U24207 (N_24207,N_23639,N_23715);
xnor U24208 (N_24208,N_23968,N_23824);
nand U24209 (N_24209,N_23654,N_23803);
xor U24210 (N_24210,N_23601,N_23814);
and U24211 (N_24211,N_23999,N_23666);
nand U24212 (N_24212,N_23588,N_23500);
nand U24213 (N_24213,N_23716,N_23524);
nand U24214 (N_24214,N_23515,N_23907);
nand U24215 (N_24215,N_23727,N_23605);
nor U24216 (N_24216,N_23691,N_23891);
nor U24217 (N_24217,N_23764,N_23765);
and U24218 (N_24218,N_23709,N_23585);
xnor U24219 (N_24219,N_23664,N_23797);
xor U24220 (N_24220,N_23805,N_23735);
xor U24221 (N_24221,N_23663,N_23752);
xor U24222 (N_24222,N_23622,N_23723);
nand U24223 (N_24223,N_23672,N_23726);
and U24224 (N_24224,N_23957,N_23572);
nand U24225 (N_24225,N_23647,N_23860);
and U24226 (N_24226,N_23609,N_23610);
xor U24227 (N_24227,N_23991,N_23831);
nand U24228 (N_24228,N_23749,N_23688);
or U24229 (N_24229,N_23561,N_23800);
xnor U24230 (N_24230,N_23536,N_23976);
xnor U24231 (N_24231,N_23668,N_23646);
and U24232 (N_24232,N_23888,N_23648);
xnor U24233 (N_24233,N_23806,N_23706);
or U24234 (N_24234,N_23754,N_23631);
nor U24235 (N_24235,N_23992,N_23728);
nor U24236 (N_24236,N_23720,N_23678);
and U24237 (N_24237,N_23988,N_23937);
or U24238 (N_24238,N_23763,N_23762);
nor U24239 (N_24239,N_23774,N_23563);
and U24240 (N_24240,N_23842,N_23681);
nor U24241 (N_24241,N_23630,N_23571);
or U24242 (N_24242,N_23599,N_23523);
or U24243 (N_24243,N_23943,N_23997);
xor U24244 (N_24244,N_23573,N_23906);
xor U24245 (N_24245,N_23689,N_23784);
and U24246 (N_24246,N_23674,N_23849);
and U24247 (N_24247,N_23632,N_23994);
and U24248 (N_24248,N_23593,N_23553);
and U24249 (N_24249,N_23652,N_23825);
or U24250 (N_24250,N_23732,N_23927);
nand U24251 (N_24251,N_23698,N_23954);
and U24252 (N_24252,N_23946,N_23659);
and U24253 (N_24253,N_23933,N_23641);
nor U24254 (N_24254,N_23569,N_23807);
or U24255 (N_24255,N_23894,N_23605);
or U24256 (N_24256,N_23665,N_23613);
xnor U24257 (N_24257,N_23678,N_23559);
and U24258 (N_24258,N_23618,N_23646);
and U24259 (N_24259,N_23841,N_23675);
xor U24260 (N_24260,N_23685,N_23844);
and U24261 (N_24261,N_23845,N_23658);
nand U24262 (N_24262,N_23812,N_23921);
and U24263 (N_24263,N_23598,N_23814);
or U24264 (N_24264,N_23934,N_23770);
nand U24265 (N_24265,N_23783,N_23945);
nor U24266 (N_24266,N_23855,N_23538);
or U24267 (N_24267,N_23768,N_23730);
nor U24268 (N_24268,N_23600,N_23711);
nand U24269 (N_24269,N_23945,N_23988);
or U24270 (N_24270,N_23840,N_23841);
and U24271 (N_24271,N_23962,N_23521);
and U24272 (N_24272,N_23698,N_23900);
xnor U24273 (N_24273,N_23705,N_23526);
and U24274 (N_24274,N_23957,N_23853);
nor U24275 (N_24275,N_23880,N_23891);
xor U24276 (N_24276,N_23712,N_23757);
or U24277 (N_24277,N_23690,N_23615);
and U24278 (N_24278,N_23547,N_23892);
xnor U24279 (N_24279,N_23666,N_23852);
nand U24280 (N_24280,N_23510,N_23869);
and U24281 (N_24281,N_23531,N_23706);
nand U24282 (N_24282,N_23714,N_23721);
and U24283 (N_24283,N_23871,N_23930);
nor U24284 (N_24284,N_23695,N_23539);
or U24285 (N_24285,N_23590,N_23920);
and U24286 (N_24286,N_23818,N_23577);
nor U24287 (N_24287,N_23971,N_23539);
xnor U24288 (N_24288,N_23505,N_23584);
xnor U24289 (N_24289,N_23828,N_23903);
xnor U24290 (N_24290,N_23923,N_23932);
or U24291 (N_24291,N_23995,N_23516);
xnor U24292 (N_24292,N_23610,N_23672);
and U24293 (N_24293,N_23856,N_23686);
nor U24294 (N_24294,N_23603,N_23904);
and U24295 (N_24295,N_23557,N_23912);
xnor U24296 (N_24296,N_23563,N_23966);
or U24297 (N_24297,N_23819,N_23934);
xnor U24298 (N_24298,N_23505,N_23840);
xnor U24299 (N_24299,N_23662,N_23577);
nand U24300 (N_24300,N_23916,N_23613);
nand U24301 (N_24301,N_23508,N_23875);
nand U24302 (N_24302,N_23878,N_23930);
or U24303 (N_24303,N_23613,N_23674);
and U24304 (N_24304,N_23545,N_23914);
xor U24305 (N_24305,N_23998,N_23676);
nor U24306 (N_24306,N_23807,N_23648);
nand U24307 (N_24307,N_23936,N_23941);
xor U24308 (N_24308,N_23770,N_23698);
and U24309 (N_24309,N_23829,N_23953);
and U24310 (N_24310,N_23605,N_23802);
xnor U24311 (N_24311,N_23929,N_23880);
and U24312 (N_24312,N_23720,N_23725);
or U24313 (N_24313,N_23888,N_23949);
or U24314 (N_24314,N_23993,N_23942);
nand U24315 (N_24315,N_23576,N_23571);
or U24316 (N_24316,N_23985,N_23508);
or U24317 (N_24317,N_23785,N_23634);
xnor U24318 (N_24318,N_23559,N_23638);
nor U24319 (N_24319,N_23901,N_23955);
or U24320 (N_24320,N_23928,N_23705);
or U24321 (N_24321,N_23724,N_23553);
or U24322 (N_24322,N_23997,N_23915);
nand U24323 (N_24323,N_23990,N_23910);
and U24324 (N_24324,N_23583,N_23906);
nor U24325 (N_24325,N_23866,N_23717);
nor U24326 (N_24326,N_23832,N_23565);
nand U24327 (N_24327,N_23600,N_23912);
or U24328 (N_24328,N_23547,N_23567);
and U24329 (N_24329,N_23670,N_23625);
nor U24330 (N_24330,N_23532,N_23675);
or U24331 (N_24331,N_23891,N_23701);
or U24332 (N_24332,N_23650,N_23826);
xnor U24333 (N_24333,N_23887,N_23821);
and U24334 (N_24334,N_23901,N_23862);
or U24335 (N_24335,N_23707,N_23722);
nand U24336 (N_24336,N_23797,N_23942);
xnor U24337 (N_24337,N_23507,N_23537);
nor U24338 (N_24338,N_23823,N_23754);
nor U24339 (N_24339,N_23590,N_23968);
and U24340 (N_24340,N_23885,N_23844);
nor U24341 (N_24341,N_23758,N_23915);
nand U24342 (N_24342,N_23883,N_23513);
nor U24343 (N_24343,N_23589,N_23690);
nand U24344 (N_24344,N_23670,N_23907);
nand U24345 (N_24345,N_23519,N_23529);
nand U24346 (N_24346,N_23925,N_23575);
or U24347 (N_24347,N_23571,N_23915);
xnor U24348 (N_24348,N_23780,N_23731);
nand U24349 (N_24349,N_23989,N_23542);
xor U24350 (N_24350,N_23918,N_23711);
and U24351 (N_24351,N_23606,N_23843);
nand U24352 (N_24352,N_23812,N_23940);
or U24353 (N_24353,N_23688,N_23634);
xor U24354 (N_24354,N_23691,N_23841);
nand U24355 (N_24355,N_23761,N_23756);
or U24356 (N_24356,N_23805,N_23768);
nor U24357 (N_24357,N_23603,N_23565);
nor U24358 (N_24358,N_23824,N_23893);
nor U24359 (N_24359,N_23842,N_23912);
nor U24360 (N_24360,N_23911,N_23803);
nor U24361 (N_24361,N_23917,N_23531);
xnor U24362 (N_24362,N_23734,N_23709);
xor U24363 (N_24363,N_23881,N_23547);
xor U24364 (N_24364,N_23513,N_23946);
nand U24365 (N_24365,N_23848,N_23515);
nand U24366 (N_24366,N_23605,N_23678);
nor U24367 (N_24367,N_23902,N_23545);
and U24368 (N_24368,N_23933,N_23652);
xor U24369 (N_24369,N_23721,N_23882);
xor U24370 (N_24370,N_23841,N_23663);
xor U24371 (N_24371,N_23723,N_23808);
nor U24372 (N_24372,N_23878,N_23786);
nand U24373 (N_24373,N_23958,N_23844);
xor U24374 (N_24374,N_23833,N_23688);
and U24375 (N_24375,N_23683,N_23680);
or U24376 (N_24376,N_23577,N_23866);
xor U24377 (N_24377,N_23827,N_23915);
nor U24378 (N_24378,N_23563,N_23726);
nor U24379 (N_24379,N_23783,N_23505);
nor U24380 (N_24380,N_23821,N_23912);
or U24381 (N_24381,N_23994,N_23812);
or U24382 (N_24382,N_23551,N_23868);
and U24383 (N_24383,N_23574,N_23788);
and U24384 (N_24384,N_23633,N_23666);
and U24385 (N_24385,N_23755,N_23617);
or U24386 (N_24386,N_23993,N_23971);
xnor U24387 (N_24387,N_23826,N_23797);
xor U24388 (N_24388,N_23899,N_23864);
nor U24389 (N_24389,N_23809,N_23795);
and U24390 (N_24390,N_23736,N_23649);
nand U24391 (N_24391,N_23750,N_23984);
nand U24392 (N_24392,N_23918,N_23793);
xor U24393 (N_24393,N_23849,N_23633);
and U24394 (N_24394,N_23945,N_23758);
nor U24395 (N_24395,N_23837,N_23586);
or U24396 (N_24396,N_23624,N_23986);
or U24397 (N_24397,N_23841,N_23782);
nor U24398 (N_24398,N_23667,N_23575);
nand U24399 (N_24399,N_23983,N_23764);
and U24400 (N_24400,N_23815,N_23975);
nor U24401 (N_24401,N_23760,N_23641);
nor U24402 (N_24402,N_23960,N_23767);
and U24403 (N_24403,N_23661,N_23666);
or U24404 (N_24404,N_23763,N_23894);
or U24405 (N_24405,N_23972,N_23688);
and U24406 (N_24406,N_23979,N_23946);
or U24407 (N_24407,N_23721,N_23688);
xnor U24408 (N_24408,N_23675,N_23907);
xnor U24409 (N_24409,N_23897,N_23662);
xor U24410 (N_24410,N_23812,N_23865);
or U24411 (N_24411,N_23733,N_23633);
nand U24412 (N_24412,N_23771,N_23839);
nor U24413 (N_24413,N_23683,N_23837);
or U24414 (N_24414,N_23735,N_23862);
nand U24415 (N_24415,N_23698,N_23989);
and U24416 (N_24416,N_23808,N_23580);
nand U24417 (N_24417,N_23961,N_23510);
or U24418 (N_24418,N_23778,N_23868);
xnor U24419 (N_24419,N_23769,N_23581);
xnor U24420 (N_24420,N_23680,N_23711);
and U24421 (N_24421,N_23631,N_23705);
nor U24422 (N_24422,N_23818,N_23753);
or U24423 (N_24423,N_23880,N_23791);
and U24424 (N_24424,N_23873,N_23772);
or U24425 (N_24425,N_23922,N_23935);
nor U24426 (N_24426,N_23541,N_23815);
xor U24427 (N_24427,N_23566,N_23824);
or U24428 (N_24428,N_23673,N_23752);
nor U24429 (N_24429,N_23995,N_23544);
or U24430 (N_24430,N_23658,N_23804);
and U24431 (N_24431,N_23739,N_23679);
or U24432 (N_24432,N_23871,N_23901);
xnor U24433 (N_24433,N_23623,N_23551);
or U24434 (N_24434,N_23549,N_23949);
xnor U24435 (N_24435,N_23907,N_23567);
nor U24436 (N_24436,N_23713,N_23870);
xor U24437 (N_24437,N_23580,N_23870);
xnor U24438 (N_24438,N_23948,N_23713);
and U24439 (N_24439,N_23540,N_23735);
or U24440 (N_24440,N_23567,N_23803);
xor U24441 (N_24441,N_23661,N_23783);
or U24442 (N_24442,N_23585,N_23682);
nor U24443 (N_24443,N_23518,N_23994);
nor U24444 (N_24444,N_23642,N_23530);
nand U24445 (N_24445,N_23809,N_23792);
and U24446 (N_24446,N_23724,N_23619);
or U24447 (N_24447,N_23700,N_23518);
or U24448 (N_24448,N_23826,N_23510);
nand U24449 (N_24449,N_23920,N_23901);
xor U24450 (N_24450,N_23750,N_23910);
nand U24451 (N_24451,N_23854,N_23924);
nor U24452 (N_24452,N_23675,N_23701);
xnor U24453 (N_24453,N_23938,N_23595);
and U24454 (N_24454,N_23584,N_23537);
nand U24455 (N_24455,N_23749,N_23914);
xnor U24456 (N_24456,N_23872,N_23889);
nor U24457 (N_24457,N_23651,N_23744);
or U24458 (N_24458,N_23960,N_23592);
xnor U24459 (N_24459,N_23573,N_23590);
nand U24460 (N_24460,N_23722,N_23615);
or U24461 (N_24461,N_23564,N_23554);
or U24462 (N_24462,N_23675,N_23670);
and U24463 (N_24463,N_23948,N_23926);
nand U24464 (N_24464,N_23825,N_23846);
or U24465 (N_24465,N_23528,N_23792);
nor U24466 (N_24466,N_23881,N_23710);
nand U24467 (N_24467,N_23759,N_23718);
or U24468 (N_24468,N_23568,N_23706);
nor U24469 (N_24469,N_23875,N_23543);
xnor U24470 (N_24470,N_23856,N_23533);
nor U24471 (N_24471,N_23553,N_23862);
and U24472 (N_24472,N_23817,N_23907);
or U24473 (N_24473,N_23652,N_23894);
or U24474 (N_24474,N_23629,N_23519);
nand U24475 (N_24475,N_23844,N_23877);
or U24476 (N_24476,N_23622,N_23839);
xor U24477 (N_24477,N_23608,N_23720);
xor U24478 (N_24478,N_23776,N_23546);
and U24479 (N_24479,N_23843,N_23750);
and U24480 (N_24480,N_23782,N_23619);
or U24481 (N_24481,N_23891,N_23835);
and U24482 (N_24482,N_23825,N_23649);
or U24483 (N_24483,N_23550,N_23633);
or U24484 (N_24484,N_23622,N_23931);
or U24485 (N_24485,N_23784,N_23619);
nand U24486 (N_24486,N_23724,N_23689);
xor U24487 (N_24487,N_23945,N_23887);
xor U24488 (N_24488,N_23758,N_23870);
and U24489 (N_24489,N_23856,N_23940);
or U24490 (N_24490,N_23870,N_23632);
and U24491 (N_24491,N_23505,N_23717);
or U24492 (N_24492,N_23848,N_23517);
nand U24493 (N_24493,N_23699,N_23633);
xor U24494 (N_24494,N_23635,N_23938);
nor U24495 (N_24495,N_23849,N_23597);
nor U24496 (N_24496,N_23685,N_23674);
nor U24497 (N_24497,N_23688,N_23912);
nor U24498 (N_24498,N_23996,N_23683);
nand U24499 (N_24499,N_23602,N_23523);
xnor U24500 (N_24500,N_24252,N_24335);
xor U24501 (N_24501,N_24237,N_24355);
nor U24502 (N_24502,N_24090,N_24127);
or U24503 (N_24503,N_24100,N_24381);
xor U24504 (N_24504,N_24314,N_24091);
nand U24505 (N_24505,N_24162,N_24138);
nand U24506 (N_24506,N_24329,N_24227);
and U24507 (N_24507,N_24185,N_24034);
nand U24508 (N_24508,N_24461,N_24083);
or U24509 (N_24509,N_24099,N_24240);
nor U24510 (N_24510,N_24277,N_24315);
nor U24511 (N_24511,N_24089,N_24125);
nand U24512 (N_24512,N_24268,N_24232);
nor U24513 (N_24513,N_24128,N_24476);
nand U24514 (N_24514,N_24215,N_24046);
nand U24515 (N_24515,N_24163,N_24003);
xnor U24516 (N_24516,N_24343,N_24475);
nand U24517 (N_24517,N_24195,N_24431);
xnor U24518 (N_24518,N_24312,N_24327);
or U24519 (N_24519,N_24360,N_24486);
nand U24520 (N_24520,N_24256,N_24351);
and U24521 (N_24521,N_24228,N_24129);
nand U24522 (N_24522,N_24258,N_24285);
or U24523 (N_24523,N_24344,N_24160);
xor U24524 (N_24524,N_24141,N_24088);
and U24525 (N_24525,N_24177,N_24297);
or U24526 (N_24526,N_24147,N_24331);
nor U24527 (N_24527,N_24325,N_24173);
and U24528 (N_24528,N_24121,N_24487);
xnor U24529 (N_24529,N_24316,N_24328);
or U24530 (N_24530,N_24114,N_24432);
and U24531 (N_24531,N_24133,N_24483);
and U24532 (N_24532,N_24056,N_24479);
nand U24533 (N_24533,N_24363,N_24382);
xnor U24534 (N_24534,N_24282,N_24451);
nand U24535 (N_24535,N_24218,N_24288);
or U24536 (N_24536,N_24037,N_24437);
nand U24537 (N_24537,N_24322,N_24212);
nand U24538 (N_24538,N_24337,N_24208);
or U24539 (N_24539,N_24107,N_24404);
or U24540 (N_24540,N_24048,N_24217);
and U24541 (N_24541,N_24006,N_24278);
xnor U24542 (N_24542,N_24478,N_24402);
and U24543 (N_24543,N_24324,N_24093);
and U24544 (N_24544,N_24482,N_24293);
and U24545 (N_24545,N_24059,N_24167);
or U24546 (N_24546,N_24233,N_24098);
xor U24547 (N_24547,N_24462,N_24384);
or U24548 (N_24548,N_24452,N_24105);
or U24549 (N_24549,N_24375,N_24072);
nor U24550 (N_24550,N_24029,N_24126);
nor U24551 (N_24551,N_24349,N_24092);
nor U24552 (N_24552,N_24300,N_24436);
and U24553 (N_24553,N_24455,N_24317);
xnor U24554 (N_24554,N_24248,N_24229);
nand U24555 (N_24555,N_24145,N_24313);
nor U24556 (N_24556,N_24387,N_24320);
nor U24557 (N_24557,N_24020,N_24017);
xor U24558 (N_24558,N_24231,N_24249);
or U24559 (N_24559,N_24050,N_24019);
or U24560 (N_24560,N_24397,N_24250);
xnor U24561 (N_24561,N_24388,N_24203);
or U24562 (N_24562,N_24257,N_24193);
nor U24563 (N_24563,N_24018,N_24309);
and U24564 (N_24564,N_24008,N_24415);
xor U24565 (N_24565,N_24354,N_24175);
nand U24566 (N_24566,N_24043,N_24152);
and U24567 (N_24567,N_24409,N_24025);
and U24568 (N_24568,N_24362,N_24253);
or U24569 (N_24569,N_24368,N_24084);
nor U24570 (N_24570,N_24047,N_24271);
nand U24571 (N_24571,N_24036,N_24400);
and U24572 (N_24572,N_24396,N_24033);
and U24573 (N_24573,N_24184,N_24474);
nor U24574 (N_24574,N_24393,N_24200);
nand U24575 (N_24575,N_24374,N_24022);
and U24576 (N_24576,N_24281,N_24266);
xnor U24577 (N_24577,N_24367,N_24273);
or U24578 (N_24578,N_24446,N_24246);
nor U24579 (N_24579,N_24210,N_24305);
nor U24580 (N_24580,N_24183,N_24386);
xor U24581 (N_24581,N_24011,N_24028);
nand U24582 (N_24582,N_24139,N_24222);
xnor U24583 (N_24583,N_24440,N_24395);
xor U24584 (N_24584,N_24377,N_24352);
and U24585 (N_24585,N_24135,N_24295);
xnor U24586 (N_24586,N_24361,N_24369);
nand U24587 (N_24587,N_24169,N_24030);
and U24588 (N_24588,N_24366,N_24074);
and U24589 (N_24589,N_24284,N_24408);
xnor U24590 (N_24590,N_24079,N_24272);
and U24591 (N_24591,N_24182,N_24421);
xnor U24592 (N_24592,N_24241,N_24111);
xor U24593 (N_24593,N_24294,N_24132);
nand U24594 (N_24594,N_24379,N_24358);
xor U24595 (N_24595,N_24154,N_24004);
and U24596 (N_24596,N_24380,N_24264);
xnor U24597 (N_24597,N_24498,N_24353);
nand U24598 (N_24598,N_24181,N_24109);
xor U24599 (N_24599,N_24097,N_24291);
xnor U24600 (N_24600,N_24443,N_24458);
nor U24601 (N_24601,N_24494,N_24174);
nand U24602 (N_24602,N_24411,N_24283);
xnor U24603 (N_24603,N_24051,N_24308);
or U24604 (N_24604,N_24336,N_24130);
or U24605 (N_24605,N_24045,N_24068);
or U24606 (N_24606,N_24450,N_24287);
xor U24607 (N_24607,N_24430,N_24077);
and U24608 (N_24608,N_24364,N_24274);
xnor U24609 (N_24609,N_24301,N_24170);
nor U24610 (N_24610,N_24131,N_24269);
nor U24611 (N_24611,N_24065,N_24262);
nand U24612 (N_24612,N_24340,N_24307);
nand U24613 (N_24613,N_24075,N_24027);
or U24614 (N_24614,N_24279,N_24464);
xnor U24615 (N_24615,N_24267,N_24326);
xnor U24616 (N_24616,N_24497,N_24457);
xor U24617 (N_24617,N_24347,N_24157);
xnor U24618 (N_24618,N_24164,N_24302);
xnor U24619 (N_24619,N_24081,N_24063);
nand U24620 (N_24620,N_24298,N_24255);
or U24621 (N_24621,N_24191,N_24166);
or U24622 (N_24622,N_24251,N_24234);
nor U24623 (N_24623,N_24254,N_24338);
nand U24624 (N_24624,N_24124,N_24192);
and U24625 (N_24625,N_24001,N_24123);
nand U24626 (N_24626,N_24206,N_24319);
and U24627 (N_24627,N_24263,N_24194);
nor U24628 (N_24628,N_24010,N_24078);
or U24629 (N_24629,N_24031,N_24055);
and U24630 (N_24630,N_24376,N_24244);
or U24631 (N_24631,N_24219,N_24221);
nor U24632 (N_24632,N_24496,N_24242);
xor U24633 (N_24633,N_24463,N_24188);
nor U24634 (N_24634,N_24239,N_24243);
nor U24635 (N_24635,N_24172,N_24371);
nand U24636 (N_24636,N_24425,N_24468);
nand U24637 (N_24637,N_24005,N_24424);
and U24638 (N_24638,N_24113,N_24062);
or U24639 (N_24639,N_24009,N_24158);
nand U24640 (N_24640,N_24197,N_24439);
and U24641 (N_24641,N_24477,N_24067);
nor U24642 (N_24642,N_24000,N_24426);
nor U24643 (N_24643,N_24303,N_24357);
xor U24644 (N_24644,N_24042,N_24394);
nor U24645 (N_24645,N_24339,N_24418);
nor U24646 (N_24646,N_24275,N_24176);
and U24647 (N_24647,N_24416,N_24235);
nor U24648 (N_24648,N_24155,N_24398);
nor U24649 (N_24649,N_24086,N_24156);
xnor U24650 (N_24650,N_24087,N_24481);
and U24651 (N_24651,N_24015,N_24417);
nor U24652 (N_24652,N_24286,N_24103);
xnor U24653 (N_24653,N_24104,N_24151);
xnor U24654 (N_24654,N_24201,N_24310);
or U24655 (N_24655,N_24153,N_24070);
or U24656 (N_24656,N_24306,N_24460);
or U24657 (N_24657,N_24054,N_24341);
or U24658 (N_24658,N_24171,N_24423);
xor U24659 (N_24659,N_24061,N_24044);
nor U24660 (N_24660,N_24385,N_24134);
nand U24661 (N_24661,N_24204,N_24187);
nand U24662 (N_24662,N_24444,N_24230);
or U24663 (N_24663,N_24220,N_24378);
nor U24664 (N_24664,N_24429,N_24345);
nor U24665 (N_24665,N_24356,N_24467);
xnor U24666 (N_24666,N_24115,N_24459);
xnor U24667 (N_24667,N_24292,N_24270);
and U24668 (N_24668,N_24214,N_24112);
xnor U24669 (N_24669,N_24276,N_24441);
xor U24670 (N_24670,N_24346,N_24499);
nor U24671 (N_24671,N_24280,N_24236);
and U24672 (N_24672,N_24304,N_24140);
nand U24673 (N_24673,N_24420,N_24108);
and U24674 (N_24674,N_24096,N_24122);
or U24675 (N_24675,N_24106,N_24066);
nor U24676 (N_24676,N_24143,N_24101);
nor U24677 (N_24677,N_24120,N_24007);
xnor U24678 (N_24678,N_24383,N_24202);
nand U24679 (N_24679,N_24410,N_24198);
xnor U24680 (N_24680,N_24290,N_24161);
xnor U24681 (N_24681,N_24469,N_24073);
nor U24682 (N_24682,N_24032,N_24442);
nand U24683 (N_24683,N_24095,N_24053);
or U24684 (N_24684,N_24060,N_24413);
or U24685 (N_24685,N_24216,N_24348);
nand U24686 (N_24686,N_24449,N_24247);
or U24687 (N_24687,N_24412,N_24076);
nand U24688 (N_24688,N_24488,N_24406);
and U24689 (N_24689,N_24265,N_24480);
or U24690 (N_24690,N_24144,N_24082);
xor U24691 (N_24691,N_24052,N_24058);
and U24692 (N_24692,N_24419,N_24350);
nor U24693 (N_24693,N_24039,N_24165);
xnor U24694 (N_24694,N_24370,N_24071);
xnor U24695 (N_24695,N_24493,N_24489);
nand U24696 (N_24696,N_24407,N_24445);
and U24697 (N_24697,N_24405,N_24289);
nand U24698 (N_24698,N_24433,N_24168);
and U24699 (N_24699,N_24148,N_24372);
and U24700 (N_24700,N_24453,N_24323);
nand U24701 (N_24701,N_24490,N_24041);
and U24702 (N_24702,N_24110,N_24466);
xnor U24703 (N_24703,N_24142,N_24146);
nor U24704 (N_24704,N_24318,N_24150);
xor U24705 (N_24705,N_24472,N_24064);
nor U24706 (N_24706,N_24403,N_24137);
or U24707 (N_24707,N_24392,N_24399);
nand U24708 (N_24708,N_24069,N_24334);
or U24709 (N_24709,N_24434,N_24473);
xnor U24710 (N_24710,N_24149,N_24332);
xnor U24711 (N_24711,N_24016,N_24190);
nand U24712 (N_24712,N_24199,N_24085);
nand U24713 (N_24713,N_24080,N_24021);
nand U24714 (N_24714,N_24209,N_24422);
or U24715 (N_24715,N_24189,N_24495);
nor U24716 (N_24716,N_24186,N_24035);
and U24717 (N_24717,N_24238,N_24296);
nand U24718 (N_24718,N_24428,N_24485);
and U24719 (N_24719,N_24102,N_24117);
xor U24720 (N_24720,N_24225,N_24213);
and U24721 (N_24721,N_24401,N_24435);
nor U24722 (N_24722,N_24471,N_24456);
nor U24723 (N_24723,N_24260,N_24330);
and U24724 (N_24724,N_24492,N_24012);
nand U24725 (N_24725,N_24196,N_24359);
and U24726 (N_24726,N_24484,N_24119);
xor U24727 (N_24727,N_24365,N_24211);
xnor U24728 (N_24728,N_24470,N_24259);
nor U24729 (N_24729,N_24178,N_24049);
xnor U24730 (N_24730,N_24261,N_24118);
and U24731 (N_24731,N_24224,N_24207);
nor U24732 (N_24732,N_24094,N_24179);
and U24733 (N_24733,N_24024,N_24389);
and U24734 (N_24734,N_24454,N_24205);
xor U24735 (N_24735,N_24448,N_24491);
nand U24736 (N_24736,N_24427,N_24465);
nor U24737 (N_24737,N_24373,N_24038);
nand U24738 (N_24738,N_24002,N_24414);
or U24739 (N_24739,N_24223,N_24342);
or U24740 (N_24740,N_24333,N_24299);
and U24741 (N_24741,N_24321,N_24026);
nor U24742 (N_24742,N_24159,N_24226);
nand U24743 (N_24743,N_24438,N_24447);
xor U24744 (N_24744,N_24245,N_24390);
and U24745 (N_24745,N_24116,N_24311);
xor U24746 (N_24746,N_24057,N_24023);
and U24747 (N_24747,N_24013,N_24180);
and U24748 (N_24748,N_24136,N_24014);
or U24749 (N_24749,N_24391,N_24040);
nor U24750 (N_24750,N_24379,N_24151);
and U24751 (N_24751,N_24272,N_24498);
nand U24752 (N_24752,N_24159,N_24346);
and U24753 (N_24753,N_24295,N_24220);
or U24754 (N_24754,N_24138,N_24027);
nor U24755 (N_24755,N_24419,N_24163);
xor U24756 (N_24756,N_24278,N_24481);
or U24757 (N_24757,N_24212,N_24471);
nor U24758 (N_24758,N_24257,N_24130);
or U24759 (N_24759,N_24436,N_24355);
xor U24760 (N_24760,N_24035,N_24008);
and U24761 (N_24761,N_24444,N_24301);
nor U24762 (N_24762,N_24341,N_24330);
xor U24763 (N_24763,N_24184,N_24300);
and U24764 (N_24764,N_24379,N_24020);
nor U24765 (N_24765,N_24130,N_24228);
xnor U24766 (N_24766,N_24153,N_24327);
nor U24767 (N_24767,N_24184,N_24264);
and U24768 (N_24768,N_24083,N_24459);
xnor U24769 (N_24769,N_24241,N_24444);
nor U24770 (N_24770,N_24030,N_24443);
xor U24771 (N_24771,N_24387,N_24041);
and U24772 (N_24772,N_24249,N_24081);
xor U24773 (N_24773,N_24497,N_24083);
and U24774 (N_24774,N_24078,N_24139);
xnor U24775 (N_24775,N_24042,N_24103);
nand U24776 (N_24776,N_24085,N_24120);
xnor U24777 (N_24777,N_24332,N_24183);
or U24778 (N_24778,N_24041,N_24007);
and U24779 (N_24779,N_24441,N_24109);
nand U24780 (N_24780,N_24010,N_24034);
nor U24781 (N_24781,N_24116,N_24473);
nor U24782 (N_24782,N_24159,N_24194);
xnor U24783 (N_24783,N_24441,N_24389);
and U24784 (N_24784,N_24342,N_24072);
and U24785 (N_24785,N_24350,N_24150);
and U24786 (N_24786,N_24337,N_24229);
nor U24787 (N_24787,N_24457,N_24022);
nor U24788 (N_24788,N_24423,N_24363);
xnor U24789 (N_24789,N_24440,N_24120);
nand U24790 (N_24790,N_24217,N_24317);
xnor U24791 (N_24791,N_24285,N_24220);
nand U24792 (N_24792,N_24336,N_24053);
and U24793 (N_24793,N_24356,N_24121);
nand U24794 (N_24794,N_24354,N_24343);
or U24795 (N_24795,N_24285,N_24404);
nand U24796 (N_24796,N_24337,N_24148);
xnor U24797 (N_24797,N_24182,N_24267);
or U24798 (N_24798,N_24301,N_24162);
xor U24799 (N_24799,N_24403,N_24181);
and U24800 (N_24800,N_24208,N_24292);
nor U24801 (N_24801,N_24496,N_24265);
nor U24802 (N_24802,N_24206,N_24426);
nor U24803 (N_24803,N_24277,N_24472);
nand U24804 (N_24804,N_24448,N_24353);
nor U24805 (N_24805,N_24124,N_24105);
or U24806 (N_24806,N_24465,N_24061);
or U24807 (N_24807,N_24192,N_24183);
xor U24808 (N_24808,N_24378,N_24199);
nand U24809 (N_24809,N_24495,N_24354);
nor U24810 (N_24810,N_24212,N_24010);
nand U24811 (N_24811,N_24114,N_24002);
nand U24812 (N_24812,N_24071,N_24097);
nor U24813 (N_24813,N_24306,N_24200);
and U24814 (N_24814,N_24452,N_24322);
nand U24815 (N_24815,N_24349,N_24237);
nand U24816 (N_24816,N_24462,N_24351);
and U24817 (N_24817,N_24172,N_24497);
xnor U24818 (N_24818,N_24376,N_24449);
xor U24819 (N_24819,N_24048,N_24067);
xor U24820 (N_24820,N_24118,N_24401);
and U24821 (N_24821,N_24252,N_24166);
or U24822 (N_24822,N_24468,N_24304);
xor U24823 (N_24823,N_24276,N_24128);
and U24824 (N_24824,N_24271,N_24280);
nand U24825 (N_24825,N_24157,N_24305);
nand U24826 (N_24826,N_24368,N_24279);
or U24827 (N_24827,N_24239,N_24297);
xor U24828 (N_24828,N_24248,N_24260);
nor U24829 (N_24829,N_24017,N_24296);
nor U24830 (N_24830,N_24490,N_24050);
nand U24831 (N_24831,N_24068,N_24122);
and U24832 (N_24832,N_24327,N_24365);
nor U24833 (N_24833,N_24406,N_24451);
xnor U24834 (N_24834,N_24287,N_24058);
and U24835 (N_24835,N_24185,N_24406);
nand U24836 (N_24836,N_24237,N_24064);
nor U24837 (N_24837,N_24186,N_24109);
and U24838 (N_24838,N_24083,N_24149);
nor U24839 (N_24839,N_24070,N_24315);
and U24840 (N_24840,N_24246,N_24383);
xnor U24841 (N_24841,N_24059,N_24041);
nor U24842 (N_24842,N_24064,N_24261);
and U24843 (N_24843,N_24279,N_24156);
xnor U24844 (N_24844,N_24102,N_24100);
or U24845 (N_24845,N_24005,N_24253);
nor U24846 (N_24846,N_24210,N_24264);
xnor U24847 (N_24847,N_24480,N_24094);
nand U24848 (N_24848,N_24445,N_24002);
xor U24849 (N_24849,N_24203,N_24177);
nand U24850 (N_24850,N_24164,N_24367);
or U24851 (N_24851,N_24165,N_24433);
nor U24852 (N_24852,N_24276,N_24222);
xor U24853 (N_24853,N_24466,N_24123);
or U24854 (N_24854,N_24246,N_24276);
nand U24855 (N_24855,N_24009,N_24077);
or U24856 (N_24856,N_24316,N_24288);
and U24857 (N_24857,N_24104,N_24222);
and U24858 (N_24858,N_24334,N_24440);
xnor U24859 (N_24859,N_24028,N_24418);
nor U24860 (N_24860,N_24446,N_24232);
nand U24861 (N_24861,N_24472,N_24068);
and U24862 (N_24862,N_24296,N_24207);
nand U24863 (N_24863,N_24291,N_24488);
nor U24864 (N_24864,N_24391,N_24314);
and U24865 (N_24865,N_24250,N_24363);
nor U24866 (N_24866,N_24175,N_24160);
and U24867 (N_24867,N_24369,N_24046);
and U24868 (N_24868,N_24003,N_24160);
xor U24869 (N_24869,N_24348,N_24185);
nor U24870 (N_24870,N_24279,N_24114);
nand U24871 (N_24871,N_24228,N_24492);
nand U24872 (N_24872,N_24029,N_24065);
or U24873 (N_24873,N_24402,N_24099);
and U24874 (N_24874,N_24488,N_24224);
nand U24875 (N_24875,N_24063,N_24234);
nor U24876 (N_24876,N_24018,N_24340);
xor U24877 (N_24877,N_24014,N_24012);
or U24878 (N_24878,N_24234,N_24483);
nand U24879 (N_24879,N_24487,N_24039);
xor U24880 (N_24880,N_24192,N_24379);
or U24881 (N_24881,N_24223,N_24417);
xnor U24882 (N_24882,N_24293,N_24211);
nor U24883 (N_24883,N_24176,N_24336);
and U24884 (N_24884,N_24100,N_24098);
nor U24885 (N_24885,N_24358,N_24254);
xor U24886 (N_24886,N_24382,N_24392);
or U24887 (N_24887,N_24295,N_24008);
nor U24888 (N_24888,N_24041,N_24331);
and U24889 (N_24889,N_24376,N_24298);
nand U24890 (N_24890,N_24204,N_24022);
and U24891 (N_24891,N_24306,N_24280);
or U24892 (N_24892,N_24451,N_24045);
or U24893 (N_24893,N_24131,N_24415);
nand U24894 (N_24894,N_24006,N_24381);
nor U24895 (N_24895,N_24445,N_24017);
nand U24896 (N_24896,N_24047,N_24429);
xnor U24897 (N_24897,N_24218,N_24309);
xor U24898 (N_24898,N_24232,N_24299);
and U24899 (N_24899,N_24137,N_24356);
nor U24900 (N_24900,N_24332,N_24349);
nand U24901 (N_24901,N_24498,N_24468);
and U24902 (N_24902,N_24314,N_24318);
and U24903 (N_24903,N_24250,N_24082);
nand U24904 (N_24904,N_24214,N_24303);
and U24905 (N_24905,N_24266,N_24445);
and U24906 (N_24906,N_24218,N_24399);
or U24907 (N_24907,N_24120,N_24051);
nand U24908 (N_24908,N_24056,N_24136);
or U24909 (N_24909,N_24396,N_24323);
and U24910 (N_24910,N_24486,N_24284);
nand U24911 (N_24911,N_24173,N_24443);
nor U24912 (N_24912,N_24393,N_24381);
nor U24913 (N_24913,N_24335,N_24153);
xor U24914 (N_24914,N_24162,N_24430);
nand U24915 (N_24915,N_24043,N_24061);
or U24916 (N_24916,N_24479,N_24463);
and U24917 (N_24917,N_24088,N_24055);
nor U24918 (N_24918,N_24055,N_24306);
nand U24919 (N_24919,N_24383,N_24297);
nand U24920 (N_24920,N_24458,N_24354);
xor U24921 (N_24921,N_24329,N_24139);
nor U24922 (N_24922,N_24270,N_24355);
or U24923 (N_24923,N_24405,N_24286);
and U24924 (N_24924,N_24272,N_24439);
and U24925 (N_24925,N_24127,N_24200);
nand U24926 (N_24926,N_24429,N_24045);
nor U24927 (N_24927,N_24147,N_24225);
nand U24928 (N_24928,N_24265,N_24335);
nor U24929 (N_24929,N_24476,N_24390);
nor U24930 (N_24930,N_24079,N_24240);
nor U24931 (N_24931,N_24287,N_24331);
nand U24932 (N_24932,N_24149,N_24169);
nand U24933 (N_24933,N_24381,N_24358);
nand U24934 (N_24934,N_24068,N_24429);
nand U24935 (N_24935,N_24385,N_24189);
nand U24936 (N_24936,N_24122,N_24383);
xnor U24937 (N_24937,N_24014,N_24040);
and U24938 (N_24938,N_24284,N_24296);
xor U24939 (N_24939,N_24344,N_24009);
xor U24940 (N_24940,N_24279,N_24113);
and U24941 (N_24941,N_24269,N_24086);
nand U24942 (N_24942,N_24044,N_24051);
nor U24943 (N_24943,N_24107,N_24240);
and U24944 (N_24944,N_24496,N_24348);
and U24945 (N_24945,N_24137,N_24211);
nand U24946 (N_24946,N_24292,N_24305);
and U24947 (N_24947,N_24126,N_24083);
xnor U24948 (N_24948,N_24356,N_24116);
and U24949 (N_24949,N_24046,N_24475);
nor U24950 (N_24950,N_24059,N_24250);
nand U24951 (N_24951,N_24100,N_24338);
and U24952 (N_24952,N_24083,N_24016);
xnor U24953 (N_24953,N_24252,N_24324);
and U24954 (N_24954,N_24351,N_24212);
nand U24955 (N_24955,N_24301,N_24446);
nor U24956 (N_24956,N_24095,N_24319);
and U24957 (N_24957,N_24341,N_24178);
nand U24958 (N_24958,N_24015,N_24149);
xor U24959 (N_24959,N_24269,N_24160);
and U24960 (N_24960,N_24021,N_24131);
or U24961 (N_24961,N_24182,N_24088);
nor U24962 (N_24962,N_24058,N_24337);
or U24963 (N_24963,N_24139,N_24463);
or U24964 (N_24964,N_24057,N_24148);
xnor U24965 (N_24965,N_24212,N_24377);
and U24966 (N_24966,N_24125,N_24083);
xor U24967 (N_24967,N_24012,N_24404);
or U24968 (N_24968,N_24490,N_24093);
xnor U24969 (N_24969,N_24391,N_24063);
nand U24970 (N_24970,N_24037,N_24420);
and U24971 (N_24971,N_24492,N_24079);
xor U24972 (N_24972,N_24007,N_24299);
nor U24973 (N_24973,N_24223,N_24480);
or U24974 (N_24974,N_24120,N_24248);
or U24975 (N_24975,N_24182,N_24394);
xnor U24976 (N_24976,N_24023,N_24233);
and U24977 (N_24977,N_24166,N_24046);
or U24978 (N_24978,N_24367,N_24025);
and U24979 (N_24979,N_24114,N_24149);
and U24980 (N_24980,N_24258,N_24419);
or U24981 (N_24981,N_24060,N_24102);
and U24982 (N_24982,N_24457,N_24260);
and U24983 (N_24983,N_24012,N_24231);
or U24984 (N_24984,N_24368,N_24183);
xor U24985 (N_24985,N_24054,N_24422);
nand U24986 (N_24986,N_24289,N_24212);
nor U24987 (N_24987,N_24499,N_24212);
nand U24988 (N_24988,N_24136,N_24103);
and U24989 (N_24989,N_24124,N_24423);
and U24990 (N_24990,N_24060,N_24340);
nor U24991 (N_24991,N_24149,N_24495);
or U24992 (N_24992,N_24338,N_24189);
nand U24993 (N_24993,N_24047,N_24396);
nand U24994 (N_24994,N_24332,N_24305);
xor U24995 (N_24995,N_24127,N_24468);
xor U24996 (N_24996,N_24378,N_24466);
xnor U24997 (N_24997,N_24182,N_24448);
nor U24998 (N_24998,N_24245,N_24087);
nor U24999 (N_24999,N_24305,N_24082);
or UO_0 (O_0,N_24906,N_24934);
xnor UO_1 (O_1,N_24570,N_24712);
nor UO_2 (O_2,N_24855,N_24775);
and UO_3 (O_3,N_24814,N_24820);
nand UO_4 (O_4,N_24549,N_24778);
nand UO_5 (O_5,N_24543,N_24900);
nor UO_6 (O_6,N_24637,N_24800);
and UO_7 (O_7,N_24657,N_24614);
nand UO_8 (O_8,N_24997,N_24667);
nand UO_9 (O_9,N_24733,N_24786);
nor UO_10 (O_10,N_24604,N_24884);
nand UO_11 (O_11,N_24694,N_24904);
nand UO_12 (O_12,N_24548,N_24795);
and UO_13 (O_13,N_24647,N_24984);
and UO_14 (O_14,N_24518,N_24522);
nor UO_15 (O_15,N_24933,N_24501);
xnor UO_16 (O_16,N_24837,N_24737);
xnor UO_17 (O_17,N_24994,N_24920);
nand UO_18 (O_18,N_24658,N_24698);
nand UO_19 (O_19,N_24690,N_24895);
nand UO_20 (O_20,N_24661,N_24921);
and UO_21 (O_21,N_24845,N_24515);
or UO_22 (O_22,N_24819,N_24953);
xor UO_23 (O_23,N_24665,N_24640);
xnor UO_24 (O_24,N_24623,N_24909);
or UO_25 (O_25,N_24977,N_24727);
nor UO_26 (O_26,N_24776,N_24966);
xor UO_27 (O_27,N_24551,N_24681);
nand UO_28 (O_28,N_24868,N_24982);
nand UO_29 (O_29,N_24958,N_24862);
nor UO_30 (O_30,N_24738,N_24622);
or UO_31 (O_31,N_24618,N_24908);
xnor UO_32 (O_32,N_24724,N_24575);
and UO_33 (O_33,N_24603,N_24630);
xnor UO_34 (O_34,N_24610,N_24705);
xnor UO_35 (O_35,N_24502,N_24653);
xor UO_36 (O_36,N_24644,N_24968);
or UO_37 (O_37,N_24767,N_24582);
xor UO_38 (O_38,N_24898,N_24936);
or UO_39 (O_39,N_24663,N_24863);
xor UO_40 (O_40,N_24545,N_24726);
nand UO_41 (O_41,N_24883,N_24973);
nand UO_42 (O_42,N_24537,N_24815);
or UO_43 (O_43,N_24998,N_24826);
or UO_44 (O_44,N_24676,N_24860);
nand UO_45 (O_45,N_24505,N_24834);
and UO_46 (O_46,N_24817,N_24987);
or UO_47 (O_47,N_24593,N_24873);
or UO_48 (O_48,N_24695,N_24613);
and UO_49 (O_49,N_24639,N_24509);
and UO_50 (O_50,N_24580,N_24880);
or UO_51 (O_51,N_24824,N_24939);
and UO_52 (O_52,N_24739,N_24704);
nand UO_53 (O_53,N_24650,N_24875);
nor UO_54 (O_54,N_24943,N_24867);
xor UO_55 (O_55,N_24774,N_24882);
xnor UO_56 (O_56,N_24682,N_24876);
xnor UO_57 (O_57,N_24595,N_24986);
nor UO_58 (O_58,N_24835,N_24975);
nor UO_59 (O_59,N_24707,N_24631);
and UO_60 (O_60,N_24568,N_24999);
nor UO_61 (O_61,N_24662,N_24585);
nand UO_62 (O_62,N_24757,N_24716);
xor UO_63 (O_63,N_24976,N_24664);
or UO_64 (O_64,N_24576,N_24679);
or UO_65 (O_65,N_24821,N_24890);
nor UO_66 (O_66,N_24621,N_24980);
or UO_67 (O_67,N_24500,N_24762);
xor UO_68 (O_68,N_24523,N_24572);
nor UO_69 (O_69,N_24857,N_24912);
nand UO_70 (O_70,N_24856,N_24945);
xnor UO_71 (O_71,N_24683,N_24581);
nand UO_72 (O_72,N_24590,N_24625);
and UO_73 (O_73,N_24810,N_24638);
nor UO_74 (O_74,N_24748,N_24780);
and UO_75 (O_75,N_24669,N_24678);
xor UO_76 (O_76,N_24632,N_24811);
nand UO_77 (O_77,N_24554,N_24988);
nor UO_78 (O_78,N_24872,N_24965);
xor UO_79 (O_79,N_24563,N_24889);
nand UO_80 (O_80,N_24583,N_24866);
nand UO_81 (O_81,N_24544,N_24660);
and UO_82 (O_82,N_24927,N_24619);
nor UO_83 (O_83,N_24722,N_24938);
or UO_84 (O_84,N_24513,N_24928);
nand UO_85 (O_85,N_24859,N_24533);
or UO_86 (O_86,N_24552,N_24879);
or UO_87 (O_87,N_24615,N_24559);
xor UO_88 (O_88,N_24910,N_24950);
nor UO_89 (O_89,N_24643,N_24808);
xor UO_90 (O_90,N_24700,N_24736);
or UO_91 (O_91,N_24874,N_24753);
nand UO_92 (O_92,N_24978,N_24840);
xnor UO_93 (O_93,N_24635,N_24526);
nor UO_94 (O_94,N_24508,N_24573);
or UO_95 (O_95,N_24797,N_24981);
nand UO_96 (O_96,N_24806,N_24801);
or UO_97 (O_97,N_24930,N_24751);
or UO_98 (O_98,N_24729,N_24961);
nor UO_99 (O_99,N_24914,N_24848);
nor UO_100 (O_100,N_24510,N_24577);
and UO_101 (O_101,N_24948,N_24645);
nor UO_102 (O_102,N_24701,N_24956);
or UO_103 (O_103,N_24746,N_24536);
xor UO_104 (O_104,N_24611,N_24646);
nand UO_105 (O_105,N_24560,N_24864);
and UO_106 (O_106,N_24571,N_24606);
xor UO_107 (O_107,N_24829,N_24564);
xnor UO_108 (O_108,N_24957,N_24745);
nor UO_109 (O_109,N_24807,N_24711);
nand UO_110 (O_110,N_24922,N_24550);
and UO_111 (O_111,N_24507,N_24962);
xor UO_112 (O_112,N_24932,N_24574);
and UO_113 (O_113,N_24731,N_24885);
nand UO_114 (O_114,N_24633,N_24990);
nor UO_115 (O_115,N_24717,N_24556);
and UO_116 (O_116,N_24967,N_24626);
xor UO_117 (O_117,N_24854,N_24607);
nor UO_118 (O_118,N_24747,N_24937);
xor UO_119 (O_119,N_24963,N_24710);
nor UO_120 (O_120,N_24760,N_24796);
or UO_121 (O_121,N_24771,N_24805);
nand UO_122 (O_122,N_24628,N_24627);
and UO_123 (O_123,N_24519,N_24531);
nand UO_124 (O_124,N_24787,N_24702);
nand UO_125 (O_125,N_24735,N_24851);
xnor UO_126 (O_126,N_24569,N_24617);
xor UO_127 (O_127,N_24598,N_24899);
nand UO_128 (O_128,N_24752,N_24878);
nor UO_129 (O_129,N_24743,N_24608);
and UO_130 (O_130,N_24793,N_24916);
and UO_131 (O_131,N_24947,N_24955);
xnor UO_132 (O_132,N_24750,N_24557);
or UO_133 (O_133,N_24517,N_24991);
xor UO_134 (O_134,N_24901,N_24685);
xor UO_135 (O_135,N_24656,N_24865);
xnor UO_136 (O_136,N_24706,N_24589);
or UO_137 (O_137,N_24539,N_24915);
and UO_138 (O_138,N_24555,N_24730);
or UO_139 (O_139,N_24566,N_24830);
nor UO_140 (O_140,N_24983,N_24512);
nand UO_141 (O_141,N_24668,N_24514);
or UO_142 (O_142,N_24527,N_24770);
xnor UO_143 (O_143,N_24913,N_24675);
and UO_144 (O_144,N_24940,N_24680);
nand UO_145 (O_145,N_24734,N_24942);
xor UO_146 (O_146,N_24849,N_24652);
or UO_147 (O_147,N_24684,N_24929);
or UO_148 (O_148,N_24979,N_24709);
nand UO_149 (O_149,N_24594,N_24789);
and UO_150 (O_150,N_24782,N_24558);
and UO_151 (O_151,N_24996,N_24565);
or UO_152 (O_152,N_24798,N_24586);
xor UO_153 (O_153,N_24597,N_24959);
or UO_154 (O_154,N_24538,N_24532);
or UO_155 (O_155,N_24763,N_24813);
nand UO_156 (O_156,N_24740,N_24567);
xnor UO_157 (O_157,N_24624,N_24905);
nor UO_158 (O_158,N_24870,N_24516);
nor UO_159 (O_159,N_24839,N_24699);
or UO_160 (O_160,N_24941,N_24654);
and UO_161 (O_161,N_24827,N_24842);
and UO_162 (O_162,N_24641,N_24954);
nand UO_163 (O_163,N_24535,N_24836);
nand UO_164 (O_164,N_24755,N_24969);
nand UO_165 (O_165,N_24917,N_24773);
and UO_166 (O_166,N_24732,N_24769);
nor UO_167 (O_167,N_24850,N_24911);
nor UO_168 (O_168,N_24708,N_24579);
xor UO_169 (O_169,N_24651,N_24749);
nand UO_170 (O_170,N_24688,N_24765);
xor UO_171 (O_171,N_24891,N_24553);
or UO_172 (O_172,N_24541,N_24525);
nor UO_173 (O_173,N_24670,N_24689);
xor UO_174 (O_174,N_24612,N_24718);
nor UO_175 (O_175,N_24561,N_24768);
nor UO_176 (O_176,N_24600,N_24728);
nor UO_177 (O_177,N_24674,N_24723);
or UO_178 (O_178,N_24601,N_24926);
xnor UO_179 (O_179,N_24721,N_24951);
nand UO_180 (O_180,N_24791,N_24799);
or UO_181 (O_181,N_24822,N_24742);
or UO_182 (O_182,N_24972,N_24599);
nor UO_183 (O_183,N_24992,N_24605);
or UO_184 (O_184,N_24825,N_24852);
and UO_185 (O_185,N_24672,N_24964);
and UO_186 (O_186,N_24671,N_24844);
nor UO_187 (O_187,N_24693,N_24602);
nor UO_188 (O_188,N_24673,N_24578);
or UO_189 (O_189,N_24703,N_24714);
nand UO_190 (O_190,N_24903,N_24785);
xnor UO_191 (O_191,N_24893,N_24833);
nand UO_192 (O_192,N_24636,N_24896);
nand UO_193 (O_193,N_24790,N_24907);
xor UO_194 (O_194,N_24846,N_24562);
xnor UO_195 (O_195,N_24783,N_24741);
nand UO_196 (O_196,N_24788,N_24588);
and UO_197 (O_197,N_24779,N_24547);
nand UO_198 (O_198,N_24871,N_24823);
nand UO_199 (O_199,N_24935,N_24616);
nor UO_200 (O_200,N_24858,N_24534);
xor UO_201 (O_201,N_24843,N_24620);
or UO_202 (O_202,N_24596,N_24521);
nor UO_203 (O_203,N_24715,N_24696);
or UO_204 (O_204,N_24960,N_24892);
nor UO_205 (O_205,N_24832,N_24949);
xor UO_206 (O_206,N_24520,N_24974);
xnor UO_207 (O_207,N_24506,N_24503);
nor UO_208 (O_208,N_24802,N_24528);
nand UO_209 (O_209,N_24888,N_24924);
xnor UO_210 (O_210,N_24902,N_24591);
xnor UO_211 (O_211,N_24925,N_24659);
xnor UO_212 (O_212,N_24759,N_24803);
and UO_213 (O_213,N_24919,N_24792);
and UO_214 (O_214,N_24542,N_24540);
xor UO_215 (O_215,N_24692,N_24781);
xor UO_216 (O_216,N_24887,N_24546);
xor UO_217 (O_217,N_24869,N_24530);
or UO_218 (O_218,N_24853,N_24995);
xnor UO_219 (O_219,N_24764,N_24841);
or UO_220 (O_220,N_24894,N_24529);
or UO_221 (O_221,N_24609,N_24861);
nand UO_222 (O_222,N_24809,N_24587);
nor UO_223 (O_223,N_24818,N_24993);
and UO_224 (O_224,N_24944,N_24648);
nand UO_225 (O_225,N_24923,N_24766);
xor UO_226 (O_226,N_24918,N_24720);
xnor UO_227 (O_227,N_24649,N_24666);
xor UO_228 (O_228,N_24634,N_24719);
or UO_229 (O_229,N_24524,N_24772);
or UO_230 (O_230,N_24897,N_24831);
or UO_231 (O_231,N_24754,N_24970);
nand UO_232 (O_232,N_24804,N_24828);
xor UO_233 (O_233,N_24952,N_24584);
nand UO_234 (O_234,N_24886,N_24816);
nand UO_235 (O_235,N_24655,N_24847);
nand UO_236 (O_236,N_24629,N_24677);
and UO_237 (O_237,N_24794,N_24971);
and UO_238 (O_238,N_24697,N_24713);
xor UO_239 (O_239,N_24687,N_24777);
or UO_240 (O_240,N_24989,N_24931);
or UO_241 (O_241,N_24877,N_24756);
xor UO_242 (O_242,N_24758,N_24686);
nand UO_243 (O_243,N_24744,N_24985);
xnor UO_244 (O_244,N_24946,N_24812);
and UO_245 (O_245,N_24511,N_24725);
xnor UO_246 (O_246,N_24838,N_24784);
nand UO_247 (O_247,N_24504,N_24691);
and UO_248 (O_248,N_24761,N_24881);
nand UO_249 (O_249,N_24592,N_24642);
and UO_250 (O_250,N_24521,N_24590);
or UO_251 (O_251,N_24863,N_24635);
and UO_252 (O_252,N_24539,N_24719);
or UO_253 (O_253,N_24877,N_24600);
and UO_254 (O_254,N_24500,N_24642);
xnor UO_255 (O_255,N_24660,N_24667);
or UO_256 (O_256,N_24557,N_24671);
or UO_257 (O_257,N_24814,N_24997);
nand UO_258 (O_258,N_24531,N_24922);
nor UO_259 (O_259,N_24502,N_24835);
or UO_260 (O_260,N_24511,N_24963);
nor UO_261 (O_261,N_24876,N_24888);
nand UO_262 (O_262,N_24594,N_24953);
nand UO_263 (O_263,N_24947,N_24815);
nor UO_264 (O_264,N_24665,N_24602);
nand UO_265 (O_265,N_24748,N_24869);
xor UO_266 (O_266,N_24550,N_24825);
nor UO_267 (O_267,N_24833,N_24954);
and UO_268 (O_268,N_24941,N_24550);
nor UO_269 (O_269,N_24992,N_24884);
or UO_270 (O_270,N_24973,N_24830);
and UO_271 (O_271,N_24534,N_24897);
nand UO_272 (O_272,N_24735,N_24896);
xor UO_273 (O_273,N_24747,N_24869);
xor UO_274 (O_274,N_24505,N_24930);
nor UO_275 (O_275,N_24556,N_24814);
nor UO_276 (O_276,N_24530,N_24680);
or UO_277 (O_277,N_24615,N_24997);
xor UO_278 (O_278,N_24508,N_24933);
and UO_279 (O_279,N_24643,N_24759);
xor UO_280 (O_280,N_24704,N_24978);
and UO_281 (O_281,N_24938,N_24631);
or UO_282 (O_282,N_24809,N_24990);
nand UO_283 (O_283,N_24855,N_24664);
or UO_284 (O_284,N_24932,N_24656);
nor UO_285 (O_285,N_24919,N_24503);
nor UO_286 (O_286,N_24989,N_24618);
and UO_287 (O_287,N_24508,N_24572);
or UO_288 (O_288,N_24888,N_24889);
and UO_289 (O_289,N_24568,N_24839);
nand UO_290 (O_290,N_24789,N_24767);
nor UO_291 (O_291,N_24791,N_24852);
and UO_292 (O_292,N_24605,N_24826);
nand UO_293 (O_293,N_24915,N_24626);
nand UO_294 (O_294,N_24791,N_24797);
xor UO_295 (O_295,N_24982,N_24935);
and UO_296 (O_296,N_24791,N_24864);
or UO_297 (O_297,N_24813,N_24829);
nand UO_298 (O_298,N_24521,N_24850);
or UO_299 (O_299,N_24768,N_24886);
nand UO_300 (O_300,N_24857,N_24948);
nor UO_301 (O_301,N_24841,N_24718);
or UO_302 (O_302,N_24997,N_24666);
nor UO_303 (O_303,N_24735,N_24651);
nand UO_304 (O_304,N_24801,N_24615);
nor UO_305 (O_305,N_24747,N_24613);
nand UO_306 (O_306,N_24928,N_24771);
nand UO_307 (O_307,N_24826,N_24727);
xor UO_308 (O_308,N_24872,N_24791);
and UO_309 (O_309,N_24650,N_24641);
and UO_310 (O_310,N_24542,N_24829);
or UO_311 (O_311,N_24746,N_24921);
nand UO_312 (O_312,N_24708,N_24613);
nand UO_313 (O_313,N_24668,N_24641);
or UO_314 (O_314,N_24669,N_24758);
nor UO_315 (O_315,N_24640,N_24928);
and UO_316 (O_316,N_24981,N_24905);
nand UO_317 (O_317,N_24941,N_24689);
nand UO_318 (O_318,N_24858,N_24632);
nor UO_319 (O_319,N_24653,N_24500);
nand UO_320 (O_320,N_24762,N_24590);
xnor UO_321 (O_321,N_24900,N_24786);
xnor UO_322 (O_322,N_24652,N_24552);
xnor UO_323 (O_323,N_24534,N_24915);
and UO_324 (O_324,N_24923,N_24991);
xor UO_325 (O_325,N_24845,N_24643);
and UO_326 (O_326,N_24725,N_24910);
or UO_327 (O_327,N_24909,N_24976);
nand UO_328 (O_328,N_24987,N_24755);
nor UO_329 (O_329,N_24788,N_24998);
or UO_330 (O_330,N_24505,N_24793);
nor UO_331 (O_331,N_24624,N_24629);
nand UO_332 (O_332,N_24745,N_24758);
and UO_333 (O_333,N_24982,N_24615);
nand UO_334 (O_334,N_24747,N_24667);
or UO_335 (O_335,N_24631,N_24564);
nor UO_336 (O_336,N_24978,N_24532);
and UO_337 (O_337,N_24897,N_24693);
or UO_338 (O_338,N_24547,N_24676);
or UO_339 (O_339,N_24752,N_24593);
nor UO_340 (O_340,N_24846,N_24620);
or UO_341 (O_341,N_24950,N_24547);
or UO_342 (O_342,N_24745,N_24517);
or UO_343 (O_343,N_24561,N_24778);
or UO_344 (O_344,N_24738,N_24696);
or UO_345 (O_345,N_24770,N_24947);
or UO_346 (O_346,N_24773,N_24923);
and UO_347 (O_347,N_24892,N_24536);
xnor UO_348 (O_348,N_24981,N_24735);
nor UO_349 (O_349,N_24625,N_24704);
xnor UO_350 (O_350,N_24611,N_24908);
and UO_351 (O_351,N_24838,N_24975);
nand UO_352 (O_352,N_24674,N_24784);
or UO_353 (O_353,N_24884,N_24993);
or UO_354 (O_354,N_24506,N_24964);
or UO_355 (O_355,N_24663,N_24936);
xnor UO_356 (O_356,N_24523,N_24566);
and UO_357 (O_357,N_24613,N_24674);
and UO_358 (O_358,N_24827,N_24939);
nor UO_359 (O_359,N_24712,N_24679);
xnor UO_360 (O_360,N_24715,N_24990);
nor UO_361 (O_361,N_24660,N_24790);
xor UO_362 (O_362,N_24572,N_24813);
nand UO_363 (O_363,N_24624,N_24711);
nand UO_364 (O_364,N_24691,N_24596);
xnor UO_365 (O_365,N_24737,N_24833);
nand UO_366 (O_366,N_24822,N_24976);
nor UO_367 (O_367,N_24627,N_24814);
xor UO_368 (O_368,N_24959,N_24701);
xnor UO_369 (O_369,N_24597,N_24553);
and UO_370 (O_370,N_24970,N_24875);
and UO_371 (O_371,N_24639,N_24580);
and UO_372 (O_372,N_24934,N_24858);
and UO_373 (O_373,N_24931,N_24589);
or UO_374 (O_374,N_24946,N_24757);
nand UO_375 (O_375,N_24824,N_24975);
or UO_376 (O_376,N_24984,N_24959);
nor UO_377 (O_377,N_24818,N_24537);
and UO_378 (O_378,N_24597,N_24775);
xor UO_379 (O_379,N_24513,N_24525);
nor UO_380 (O_380,N_24762,N_24595);
xor UO_381 (O_381,N_24801,N_24944);
xnor UO_382 (O_382,N_24568,N_24643);
and UO_383 (O_383,N_24616,N_24790);
and UO_384 (O_384,N_24795,N_24609);
and UO_385 (O_385,N_24780,N_24740);
and UO_386 (O_386,N_24530,N_24517);
nor UO_387 (O_387,N_24736,N_24703);
xor UO_388 (O_388,N_24577,N_24580);
or UO_389 (O_389,N_24540,N_24632);
xnor UO_390 (O_390,N_24720,N_24814);
or UO_391 (O_391,N_24840,N_24710);
xnor UO_392 (O_392,N_24963,N_24774);
or UO_393 (O_393,N_24671,N_24942);
nor UO_394 (O_394,N_24612,N_24990);
xnor UO_395 (O_395,N_24679,N_24768);
nor UO_396 (O_396,N_24932,N_24808);
nor UO_397 (O_397,N_24829,N_24687);
or UO_398 (O_398,N_24974,N_24652);
nand UO_399 (O_399,N_24508,N_24564);
nor UO_400 (O_400,N_24664,N_24615);
or UO_401 (O_401,N_24818,N_24849);
xor UO_402 (O_402,N_24925,N_24785);
nor UO_403 (O_403,N_24690,N_24646);
nor UO_404 (O_404,N_24753,N_24745);
nand UO_405 (O_405,N_24894,N_24742);
or UO_406 (O_406,N_24624,N_24888);
nand UO_407 (O_407,N_24852,N_24614);
and UO_408 (O_408,N_24896,N_24664);
nand UO_409 (O_409,N_24831,N_24520);
nor UO_410 (O_410,N_24566,N_24776);
xnor UO_411 (O_411,N_24724,N_24707);
and UO_412 (O_412,N_24624,N_24519);
and UO_413 (O_413,N_24785,N_24915);
nor UO_414 (O_414,N_24562,N_24892);
or UO_415 (O_415,N_24636,N_24906);
xor UO_416 (O_416,N_24939,N_24847);
and UO_417 (O_417,N_24840,N_24547);
nand UO_418 (O_418,N_24973,N_24903);
nor UO_419 (O_419,N_24640,N_24557);
and UO_420 (O_420,N_24537,N_24720);
nand UO_421 (O_421,N_24782,N_24569);
nor UO_422 (O_422,N_24907,N_24973);
nor UO_423 (O_423,N_24596,N_24945);
and UO_424 (O_424,N_24562,N_24521);
xnor UO_425 (O_425,N_24922,N_24783);
and UO_426 (O_426,N_24635,N_24885);
xnor UO_427 (O_427,N_24814,N_24955);
nor UO_428 (O_428,N_24702,N_24603);
xnor UO_429 (O_429,N_24961,N_24770);
nand UO_430 (O_430,N_24564,N_24955);
and UO_431 (O_431,N_24587,N_24695);
or UO_432 (O_432,N_24901,N_24933);
nand UO_433 (O_433,N_24667,N_24852);
nand UO_434 (O_434,N_24977,N_24873);
and UO_435 (O_435,N_24738,N_24771);
or UO_436 (O_436,N_24593,N_24762);
xnor UO_437 (O_437,N_24736,N_24997);
nor UO_438 (O_438,N_24736,N_24964);
and UO_439 (O_439,N_24645,N_24796);
or UO_440 (O_440,N_24919,N_24506);
nand UO_441 (O_441,N_24745,N_24829);
nand UO_442 (O_442,N_24741,N_24860);
and UO_443 (O_443,N_24568,N_24699);
xor UO_444 (O_444,N_24862,N_24947);
and UO_445 (O_445,N_24666,N_24884);
nand UO_446 (O_446,N_24627,N_24792);
or UO_447 (O_447,N_24951,N_24502);
or UO_448 (O_448,N_24570,N_24710);
xor UO_449 (O_449,N_24902,N_24911);
nand UO_450 (O_450,N_24695,N_24785);
or UO_451 (O_451,N_24763,N_24761);
nor UO_452 (O_452,N_24929,N_24816);
xnor UO_453 (O_453,N_24718,N_24687);
xor UO_454 (O_454,N_24669,N_24833);
nand UO_455 (O_455,N_24935,N_24521);
nand UO_456 (O_456,N_24618,N_24566);
or UO_457 (O_457,N_24782,N_24953);
xor UO_458 (O_458,N_24566,N_24937);
nor UO_459 (O_459,N_24619,N_24990);
nand UO_460 (O_460,N_24904,N_24631);
xor UO_461 (O_461,N_24964,N_24850);
xor UO_462 (O_462,N_24632,N_24776);
xor UO_463 (O_463,N_24657,N_24634);
or UO_464 (O_464,N_24925,N_24702);
xor UO_465 (O_465,N_24550,N_24944);
xnor UO_466 (O_466,N_24588,N_24595);
or UO_467 (O_467,N_24643,N_24884);
nand UO_468 (O_468,N_24524,N_24847);
nand UO_469 (O_469,N_24620,N_24632);
or UO_470 (O_470,N_24951,N_24679);
nor UO_471 (O_471,N_24799,N_24609);
xnor UO_472 (O_472,N_24874,N_24895);
xor UO_473 (O_473,N_24855,N_24919);
nand UO_474 (O_474,N_24688,N_24656);
xnor UO_475 (O_475,N_24864,N_24610);
or UO_476 (O_476,N_24586,N_24957);
xnor UO_477 (O_477,N_24747,N_24998);
nand UO_478 (O_478,N_24871,N_24947);
nand UO_479 (O_479,N_24778,N_24819);
and UO_480 (O_480,N_24575,N_24604);
nor UO_481 (O_481,N_24978,N_24719);
and UO_482 (O_482,N_24970,N_24716);
and UO_483 (O_483,N_24546,N_24733);
or UO_484 (O_484,N_24652,N_24906);
nand UO_485 (O_485,N_24537,N_24723);
or UO_486 (O_486,N_24729,N_24906);
and UO_487 (O_487,N_24900,N_24583);
nand UO_488 (O_488,N_24568,N_24767);
nor UO_489 (O_489,N_24531,N_24581);
nand UO_490 (O_490,N_24825,N_24897);
xor UO_491 (O_491,N_24562,N_24730);
or UO_492 (O_492,N_24942,N_24958);
nor UO_493 (O_493,N_24953,N_24915);
xnor UO_494 (O_494,N_24997,N_24795);
xnor UO_495 (O_495,N_24970,N_24565);
nor UO_496 (O_496,N_24829,N_24936);
and UO_497 (O_497,N_24720,N_24928);
nand UO_498 (O_498,N_24893,N_24895);
and UO_499 (O_499,N_24934,N_24515);
xor UO_500 (O_500,N_24504,N_24817);
and UO_501 (O_501,N_24662,N_24518);
nand UO_502 (O_502,N_24812,N_24648);
xnor UO_503 (O_503,N_24788,N_24617);
and UO_504 (O_504,N_24585,N_24925);
nor UO_505 (O_505,N_24817,N_24849);
xnor UO_506 (O_506,N_24675,N_24627);
or UO_507 (O_507,N_24744,N_24505);
and UO_508 (O_508,N_24505,N_24970);
and UO_509 (O_509,N_24763,N_24531);
xnor UO_510 (O_510,N_24587,N_24665);
nand UO_511 (O_511,N_24632,N_24838);
and UO_512 (O_512,N_24728,N_24516);
nand UO_513 (O_513,N_24695,N_24898);
nor UO_514 (O_514,N_24588,N_24962);
xor UO_515 (O_515,N_24629,N_24751);
xor UO_516 (O_516,N_24731,N_24509);
nand UO_517 (O_517,N_24606,N_24628);
and UO_518 (O_518,N_24831,N_24696);
nand UO_519 (O_519,N_24612,N_24864);
nor UO_520 (O_520,N_24513,N_24870);
or UO_521 (O_521,N_24736,N_24837);
xnor UO_522 (O_522,N_24785,N_24653);
nand UO_523 (O_523,N_24967,N_24603);
or UO_524 (O_524,N_24948,N_24843);
and UO_525 (O_525,N_24879,N_24636);
xor UO_526 (O_526,N_24728,N_24843);
xor UO_527 (O_527,N_24570,N_24896);
or UO_528 (O_528,N_24664,N_24645);
nor UO_529 (O_529,N_24768,N_24552);
xor UO_530 (O_530,N_24562,N_24859);
xor UO_531 (O_531,N_24754,N_24509);
and UO_532 (O_532,N_24534,N_24950);
nand UO_533 (O_533,N_24639,N_24934);
or UO_534 (O_534,N_24504,N_24820);
and UO_535 (O_535,N_24856,N_24985);
or UO_536 (O_536,N_24812,N_24983);
xor UO_537 (O_537,N_24799,N_24984);
and UO_538 (O_538,N_24836,N_24684);
nor UO_539 (O_539,N_24973,N_24880);
or UO_540 (O_540,N_24731,N_24838);
xnor UO_541 (O_541,N_24905,N_24527);
nor UO_542 (O_542,N_24934,N_24580);
nand UO_543 (O_543,N_24913,N_24543);
nand UO_544 (O_544,N_24755,N_24924);
and UO_545 (O_545,N_24643,N_24666);
and UO_546 (O_546,N_24860,N_24584);
xnor UO_547 (O_547,N_24945,N_24527);
and UO_548 (O_548,N_24854,N_24777);
xnor UO_549 (O_549,N_24620,N_24744);
or UO_550 (O_550,N_24547,N_24681);
or UO_551 (O_551,N_24546,N_24611);
nand UO_552 (O_552,N_24546,N_24594);
or UO_553 (O_553,N_24784,N_24743);
xor UO_554 (O_554,N_24895,N_24791);
nand UO_555 (O_555,N_24696,N_24655);
nor UO_556 (O_556,N_24578,N_24906);
and UO_557 (O_557,N_24647,N_24709);
or UO_558 (O_558,N_24528,N_24968);
nand UO_559 (O_559,N_24971,N_24833);
xor UO_560 (O_560,N_24948,N_24707);
nand UO_561 (O_561,N_24848,N_24862);
xor UO_562 (O_562,N_24993,N_24725);
nor UO_563 (O_563,N_24634,N_24885);
nor UO_564 (O_564,N_24632,N_24893);
and UO_565 (O_565,N_24834,N_24741);
or UO_566 (O_566,N_24506,N_24864);
nor UO_567 (O_567,N_24886,N_24555);
and UO_568 (O_568,N_24673,N_24761);
or UO_569 (O_569,N_24967,N_24792);
and UO_570 (O_570,N_24769,N_24723);
xnor UO_571 (O_571,N_24619,N_24950);
xnor UO_572 (O_572,N_24875,N_24889);
xnor UO_573 (O_573,N_24502,N_24917);
and UO_574 (O_574,N_24790,N_24561);
and UO_575 (O_575,N_24594,N_24584);
nor UO_576 (O_576,N_24775,N_24732);
nor UO_577 (O_577,N_24903,N_24545);
xnor UO_578 (O_578,N_24683,N_24580);
nand UO_579 (O_579,N_24681,N_24924);
nand UO_580 (O_580,N_24643,N_24502);
nor UO_581 (O_581,N_24705,N_24584);
and UO_582 (O_582,N_24998,N_24534);
and UO_583 (O_583,N_24667,N_24664);
or UO_584 (O_584,N_24710,N_24805);
nand UO_585 (O_585,N_24528,N_24597);
nor UO_586 (O_586,N_24926,N_24680);
nand UO_587 (O_587,N_24936,N_24852);
xnor UO_588 (O_588,N_24508,N_24506);
xor UO_589 (O_589,N_24654,N_24946);
nor UO_590 (O_590,N_24545,N_24806);
nand UO_591 (O_591,N_24802,N_24578);
nand UO_592 (O_592,N_24841,N_24723);
nor UO_593 (O_593,N_24873,N_24783);
and UO_594 (O_594,N_24519,N_24796);
nor UO_595 (O_595,N_24643,N_24861);
and UO_596 (O_596,N_24902,N_24890);
nor UO_597 (O_597,N_24880,N_24824);
and UO_598 (O_598,N_24781,N_24829);
nand UO_599 (O_599,N_24890,N_24681);
or UO_600 (O_600,N_24826,N_24709);
and UO_601 (O_601,N_24925,N_24870);
nor UO_602 (O_602,N_24971,N_24548);
nor UO_603 (O_603,N_24615,N_24582);
xor UO_604 (O_604,N_24994,N_24821);
nor UO_605 (O_605,N_24653,N_24613);
nand UO_606 (O_606,N_24835,N_24570);
xnor UO_607 (O_607,N_24806,N_24677);
or UO_608 (O_608,N_24508,N_24693);
xnor UO_609 (O_609,N_24644,N_24568);
nand UO_610 (O_610,N_24828,N_24618);
nand UO_611 (O_611,N_24982,N_24917);
nor UO_612 (O_612,N_24887,N_24571);
nor UO_613 (O_613,N_24916,N_24622);
xor UO_614 (O_614,N_24546,N_24725);
xnor UO_615 (O_615,N_24657,N_24703);
and UO_616 (O_616,N_24741,N_24510);
nor UO_617 (O_617,N_24961,N_24859);
nor UO_618 (O_618,N_24681,N_24680);
nand UO_619 (O_619,N_24568,N_24883);
and UO_620 (O_620,N_24817,N_24548);
nor UO_621 (O_621,N_24615,N_24785);
xor UO_622 (O_622,N_24884,N_24567);
and UO_623 (O_623,N_24872,N_24849);
nor UO_624 (O_624,N_24679,N_24968);
nor UO_625 (O_625,N_24681,N_24925);
nor UO_626 (O_626,N_24540,N_24956);
and UO_627 (O_627,N_24967,N_24673);
and UO_628 (O_628,N_24731,N_24524);
nand UO_629 (O_629,N_24867,N_24709);
xnor UO_630 (O_630,N_24569,N_24965);
and UO_631 (O_631,N_24574,N_24822);
nor UO_632 (O_632,N_24634,N_24802);
xnor UO_633 (O_633,N_24618,N_24627);
or UO_634 (O_634,N_24661,N_24618);
nor UO_635 (O_635,N_24972,N_24936);
and UO_636 (O_636,N_24650,N_24974);
and UO_637 (O_637,N_24645,N_24521);
nor UO_638 (O_638,N_24715,N_24764);
xnor UO_639 (O_639,N_24894,N_24521);
nand UO_640 (O_640,N_24682,N_24542);
nor UO_641 (O_641,N_24811,N_24750);
or UO_642 (O_642,N_24558,N_24710);
and UO_643 (O_643,N_24646,N_24506);
or UO_644 (O_644,N_24703,N_24788);
nand UO_645 (O_645,N_24806,N_24922);
or UO_646 (O_646,N_24883,N_24708);
nand UO_647 (O_647,N_24780,N_24988);
nand UO_648 (O_648,N_24872,N_24556);
nand UO_649 (O_649,N_24925,N_24783);
or UO_650 (O_650,N_24721,N_24892);
nor UO_651 (O_651,N_24597,N_24661);
nand UO_652 (O_652,N_24501,N_24504);
and UO_653 (O_653,N_24794,N_24711);
or UO_654 (O_654,N_24888,N_24591);
nand UO_655 (O_655,N_24771,N_24865);
nor UO_656 (O_656,N_24897,N_24889);
or UO_657 (O_657,N_24723,N_24504);
nor UO_658 (O_658,N_24518,N_24956);
xor UO_659 (O_659,N_24801,N_24985);
or UO_660 (O_660,N_24648,N_24842);
nand UO_661 (O_661,N_24580,N_24789);
or UO_662 (O_662,N_24991,N_24752);
nand UO_663 (O_663,N_24941,N_24965);
and UO_664 (O_664,N_24920,N_24823);
nor UO_665 (O_665,N_24572,N_24544);
nand UO_666 (O_666,N_24801,N_24599);
nor UO_667 (O_667,N_24772,N_24659);
xor UO_668 (O_668,N_24700,N_24801);
and UO_669 (O_669,N_24594,N_24797);
or UO_670 (O_670,N_24888,N_24849);
or UO_671 (O_671,N_24863,N_24571);
and UO_672 (O_672,N_24683,N_24992);
and UO_673 (O_673,N_24655,N_24557);
nor UO_674 (O_674,N_24800,N_24710);
xor UO_675 (O_675,N_24654,N_24601);
or UO_676 (O_676,N_24839,N_24734);
or UO_677 (O_677,N_24899,N_24974);
nor UO_678 (O_678,N_24733,N_24657);
or UO_679 (O_679,N_24980,N_24991);
or UO_680 (O_680,N_24699,N_24604);
and UO_681 (O_681,N_24570,N_24909);
xnor UO_682 (O_682,N_24666,N_24545);
and UO_683 (O_683,N_24864,N_24965);
xnor UO_684 (O_684,N_24757,N_24659);
xor UO_685 (O_685,N_24507,N_24968);
or UO_686 (O_686,N_24890,N_24796);
or UO_687 (O_687,N_24912,N_24749);
or UO_688 (O_688,N_24858,N_24615);
xnor UO_689 (O_689,N_24832,N_24527);
xor UO_690 (O_690,N_24723,N_24706);
nor UO_691 (O_691,N_24981,N_24796);
xor UO_692 (O_692,N_24777,N_24920);
and UO_693 (O_693,N_24878,N_24561);
and UO_694 (O_694,N_24893,N_24802);
nor UO_695 (O_695,N_24764,N_24960);
nand UO_696 (O_696,N_24528,N_24904);
nand UO_697 (O_697,N_24812,N_24956);
xor UO_698 (O_698,N_24796,N_24921);
or UO_699 (O_699,N_24548,N_24777);
nor UO_700 (O_700,N_24898,N_24614);
nor UO_701 (O_701,N_24794,N_24723);
and UO_702 (O_702,N_24811,N_24581);
or UO_703 (O_703,N_24502,N_24719);
nor UO_704 (O_704,N_24604,N_24616);
or UO_705 (O_705,N_24664,N_24770);
or UO_706 (O_706,N_24628,N_24514);
nand UO_707 (O_707,N_24664,N_24905);
nand UO_708 (O_708,N_24956,N_24550);
nand UO_709 (O_709,N_24742,N_24688);
and UO_710 (O_710,N_24733,N_24717);
or UO_711 (O_711,N_24544,N_24831);
xnor UO_712 (O_712,N_24954,N_24976);
and UO_713 (O_713,N_24641,N_24673);
xnor UO_714 (O_714,N_24817,N_24834);
nand UO_715 (O_715,N_24706,N_24566);
nor UO_716 (O_716,N_24590,N_24859);
and UO_717 (O_717,N_24530,N_24614);
and UO_718 (O_718,N_24823,N_24878);
and UO_719 (O_719,N_24922,N_24604);
xnor UO_720 (O_720,N_24743,N_24718);
or UO_721 (O_721,N_24588,N_24635);
nor UO_722 (O_722,N_24974,N_24798);
or UO_723 (O_723,N_24629,N_24823);
and UO_724 (O_724,N_24539,N_24717);
nor UO_725 (O_725,N_24958,N_24519);
xnor UO_726 (O_726,N_24678,N_24934);
or UO_727 (O_727,N_24844,N_24812);
nand UO_728 (O_728,N_24713,N_24645);
xor UO_729 (O_729,N_24713,N_24716);
nor UO_730 (O_730,N_24990,N_24650);
xor UO_731 (O_731,N_24901,N_24890);
nor UO_732 (O_732,N_24816,N_24869);
or UO_733 (O_733,N_24927,N_24805);
or UO_734 (O_734,N_24564,N_24795);
xor UO_735 (O_735,N_24885,N_24984);
xor UO_736 (O_736,N_24518,N_24862);
xor UO_737 (O_737,N_24695,N_24921);
nor UO_738 (O_738,N_24736,N_24731);
xor UO_739 (O_739,N_24539,N_24726);
nand UO_740 (O_740,N_24694,N_24847);
nand UO_741 (O_741,N_24599,N_24826);
and UO_742 (O_742,N_24584,N_24738);
or UO_743 (O_743,N_24892,N_24927);
or UO_744 (O_744,N_24682,N_24649);
nor UO_745 (O_745,N_24555,N_24557);
xnor UO_746 (O_746,N_24530,N_24862);
and UO_747 (O_747,N_24533,N_24658);
nor UO_748 (O_748,N_24877,N_24809);
xor UO_749 (O_749,N_24509,N_24608);
xnor UO_750 (O_750,N_24580,N_24927);
nand UO_751 (O_751,N_24663,N_24792);
or UO_752 (O_752,N_24983,N_24829);
or UO_753 (O_753,N_24593,N_24528);
nand UO_754 (O_754,N_24862,N_24580);
xnor UO_755 (O_755,N_24739,N_24754);
or UO_756 (O_756,N_24944,N_24750);
nand UO_757 (O_757,N_24660,N_24571);
xor UO_758 (O_758,N_24664,N_24957);
or UO_759 (O_759,N_24592,N_24536);
nand UO_760 (O_760,N_24890,N_24764);
nor UO_761 (O_761,N_24907,N_24609);
or UO_762 (O_762,N_24923,N_24622);
nor UO_763 (O_763,N_24532,N_24592);
or UO_764 (O_764,N_24948,N_24957);
xnor UO_765 (O_765,N_24744,N_24773);
nor UO_766 (O_766,N_24821,N_24596);
or UO_767 (O_767,N_24773,N_24504);
xor UO_768 (O_768,N_24714,N_24781);
nand UO_769 (O_769,N_24723,N_24959);
nand UO_770 (O_770,N_24757,N_24959);
xnor UO_771 (O_771,N_24541,N_24631);
and UO_772 (O_772,N_24973,N_24711);
or UO_773 (O_773,N_24803,N_24999);
nand UO_774 (O_774,N_24909,N_24807);
nand UO_775 (O_775,N_24729,N_24891);
xnor UO_776 (O_776,N_24843,N_24733);
xnor UO_777 (O_777,N_24973,N_24788);
xor UO_778 (O_778,N_24729,N_24697);
nand UO_779 (O_779,N_24853,N_24705);
or UO_780 (O_780,N_24589,N_24729);
xnor UO_781 (O_781,N_24620,N_24723);
nand UO_782 (O_782,N_24846,N_24791);
and UO_783 (O_783,N_24630,N_24586);
and UO_784 (O_784,N_24525,N_24919);
xor UO_785 (O_785,N_24901,N_24976);
xor UO_786 (O_786,N_24900,N_24763);
nand UO_787 (O_787,N_24559,N_24912);
nand UO_788 (O_788,N_24724,N_24771);
or UO_789 (O_789,N_24966,N_24516);
or UO_790 (O_790,N_24810,N_24711);
nor UO_791 (O_791,N_24583,N_24994);
or UO_792 (O_792,N_24555,N_24836);
or UO_793 (O_793,N_24535,N_24532);
nand UO_794 (O_794,N_24855,N_24515);
nor UO_795 (O_795,N_24711,N_24580);
or UO_796 (O_796,N_24543,N_24961);
and UO_797 (O_797,N_24934,N_24632);
nand UO_798 (O_798,N_24740,N_24659);
xnor UO_799 (O_799,N_24824,N_24527);
nor UO_800 (O_800,N_24610,N_24572);
and UO_801 (O_801,N_24676,N_24507);
or UO_802 (O_802,N_24833,N_24810);
and UO_803 (O_803,N_24592,N_24843);
nor UO_804 (O_804,N_24505,N_24678);
and UO_805 (O_805,N_24744,N_24925);
or UO_806 (O_806,N_24750,N_24562);
nor UO_807 (O_807,N_24732,N_24514);
and UO_808 (O_808,N_24506,N_24519);
nor UO_809 (O_809,N_24566,N_24718);
and UO_810 (O_810,N_24649,N_24763);
xor UO_811 (O_811,N_24540,N_24570);
xnor UO_812 (O_812,N_24877,N_24989);
nand UO_813 (O_813,N_24585,N_24517);
xor UO_814 (O_814,N_24974,N_24814);
or UO_815 (O_815,N_24530,N_24542);
nand UO_816 (O_816,N_24939,N_24539);
nand UO_817 (O_817,N_24677,N_24994);
nand UO_818 (O_818,N_24957,N_24718);
xnor UO_819 (O_819,N_24876,N_24997);
nor UO_820 (O_820,N_24892,N_24549);
nand UO_821 (O_821,N_24907,N_24872);
nand UO_822 (O_822,N_24894,N_24842);
nand UO_823 (O_823,N_24951,N_24638);
xor UO_824 (O_824,N_24627,N_24645);
nand UO_825 (O_825,N_24896,N_24644);
and UO_826 (O_826,N_24921,N_24698);
nand UO_827 (O_827,N_24817,N_24616);
nor UO_828 (O_828,N_24853,N_24554);
xnor UO_829 (O_829,N_24914,N_24699);
nand UO_830 (O_830,N_24711,N_24964);
nand UO_831 (O_831,N_24913,N_24563);
or UO_832 (O_832,N_24597,N_24514);
xnor UO_833 (O_833,N_24787,N_24694);
and UO_834 (O_834,N_24565,N_24710);
nand UO_835 (O_835,N_24534,N_24884);
and UO_836 (O_836,N_24776,N_24917);
nor UO_837 (O_837,N_24717,N_24601);
and UO_838 (O_838,N_24754,N_24821);
or UO_839 (O_839,N_24507,N_24795);
and UO_840 (O_840,N_24974,N_24808);
xor UO_841 (O_841,N_24882,N_24742);
nor UO_842 (O_842,N_24784,N_24580);
nor UO_843 (O_843,N_24863,N_24702);
nand UO_844 (O_844,N_24592,N_24679);
or UO_845 (O_845,N_24656,N_24824);
nor UO_846 (O_846,N_24529,N_24560);
xor UO_847 (O_847,N_24553,N_24547);
nand UO_848 (O_848,N_24848,N_24521);
and UO_849 (O_849,N_24522,N_24546);
nand UO_850 (O_850,N_24887,N_24987);
nor UO_851 (O_851,N_24812,N_24980);
xor UO_852 (O_852,N_24719,N_24803);
and UO_853 (O_853,N_24969,N_24940);
and UO_854 (O_854,N_24502,N_24863);
or UO_855 (O_855,N_24652,N_24934);
nand UO_856 (O_856,N_24792,N_24767);
and UO_857 (O_857,N_24747,N_24804);
nor UO_858 (O_858,N_24674,N_24823);
nand UO_859 (O_859,N_24675,N_24710);
or UO_860 (O_860,N_24685,N_24908);
xor UO_861 (O_861,N_24808,N_24746);
nand UO_862 (O_862,N_24703,N_24602);
or UO_863 (O_863,N_24647,N_24985);
and UO_864 (O_864,N_24827,N_24698);
or UO_865 (O_865,N_24894,N_24712);
and UO_866 (O_866,N_24636,N_24869);
nand UO_867 (O_867,N_24764,N_24550);
or UO_868 (O_868,N_24710,N_24922);
nand UO_869 (O_869,N_24696,N_24993);
or UO_870 (O_870,N_24980,N_24721);
nand UO_871 (O_871,N_24536,N_24822);
or UO_872 (O_872,N_24564,N_24685);
xnor UO_873 (O_873,N_24506,N_24766);
nor UO_874 (O_874,N_24964,N_24854);
nor UO_875 (O_875,N_24919,N_24529);
nor UO_876 (O_876,N_24983,N_24769);
or UO_877 (O_877,N_24785,N_24756);
xor UO_878 (O_878,N_24877,N_24647);
and UO_879 (O_879,N_24730,N_24936);
xnor UO_880 (O_880,N_24613,N_24889);
or UO_881 (O_881,N_24913,N_24559);
nor UO_882 (O_882,N_24799,N_24516);
xnor UO_883 (O_883,N_24611,N_24571);
nand UO_884 (O_884,N_24541,N_24570);
and UO_885 (O_885,N_24995,N_24998);
or UO_886 (O_886,N_24758,N_24677);
or UO_887 (O_887,N_24503,N_24816);
nand UO_888 (O_888,N_24663,N_24623);
or UO_889 (O_889,N_24594,N_24730);
nand UO_890 (O_890,N_24686,N_24805);
nor UO_891 (O_891,N_24805,N_24533);
and UO_892 (O_892,N_24767,N_24864);
and UO_893 (O_893,N_24679,N_24959);
nor UO_894 (O_894,N_24972,N_24725);
and UO_895 (O_895,N_24844,N_24919);
xnor UO_896 (O_896,N_24946,N_24971);
and UO_897 (O_897,N_24942,N_24935);
xor UO_898 (O_898,N_24560,N_24933);
nand UO_899 (O_899,N_24615,N_24782);
nor UO_900 (O_900,N_24579,N_24776);
nor UO_901 (O_901,N_24685,N_24889);
and UO_902 (O_902,N_24936,N_24658);
or UO_903 (O_903,N_24565,N_24652);
nand UO_904 (O_904,N_24588,N_24578);
nor UO_905 (O_905,N_24859,N_24500);
or UO_906 (O_906,N_24717,N_24607);
nand UO_907 (O_907,N_24507,N_24567);
xnor UO_908 (O_908,N_24775,N_24773);
xor UO_909 (O_909,N_24808,N_24773);
nand UO_910 (O_910,N_24831,N_24723);
xor UO_911 (O_911,N_24714,N_24628);
nand UO_912 (O_912,N_24637,N_24834);
xnor UO_913 (O_913,N_24612,N_24989);
xnor UO_914 (O_914,N_24940,N_24912);
nand UO_915 (O_915,N_24836,N_24818);
xor UO_916 (O_916,N_24593,N_24707);
xnor UO_917 (O_917,N_24654,N_24757);
or UO_918 (O_918,N_24670,N_24663);
nor UO_919 (O_919,N_24796,N_24658);
nand UO_920 (O_920,N_24965,N_24744);
and UO_921 (O_921,N_24531,N_24937);
xor UO_922 (O_922,N_24511,N_24632);
nand UO_923 (O_923,N_24637,N_24887);
nand UO_924 (O_924,N_24581,N_24656);
xnor UO_925 (O_925,N_24511,N_24985);
and UO_926 (O_926,N_24508,N_24754);
nor UO_927 (O_927,N_24562,N_24752);
nand UO_928 (O_928,N_24817,N_24756);
nor UO_929 (O_929,N_24823,N_24538);
xor UO_930 (O_930,N_24881,N_24867);
nand UO_931 (O_931,N_24654,N_24862);
and UO_932 (O_932,N_24985,N_24996);
nor UO_933 (O_933,N_24529,N_24540);
nor UO_934 (O_934,N_24834,N_24691);
and UO_935 (O_935,N_24911,N_24950);
xnor UO_936 (O_936,N_24640,N_24874);
or UO_937 (O_937,N_24969,N_24728);
or UO_938 (O_938,N_24935,N_24592);
nand UO_939 (O_939,N_24828,N_24899);
nand UO_940 (O_940,N_24527,N_24719);
nor UO_941 (O_941,N_24995,N_24514);
nand UO_942 (O_942,N_24530,N_24647);
or UO_943 (O_943,N_24945,N_24791);
and UO_944 (O_944,N_24911,N_24718);
or UO_945 (O_945,N_24929,N_24692);
or UO_946 (O_946,N_24821,N_24567);
or UO_947 (O_947,N_24844,N_24796);
nor UO_948 (O_948,N_24613,N_24911);
and UO_949 (O_949,N_24602,N_24901);
nand UO_950 (O_950,N_24509,N_24700);
nand UO_951 (O_951,N_24569,N_24999);
nand UO_952 (O_952,N_24519,N_24916);
xor UO_953 (O_953,N_24513,N_24894);
xor UO_954 (O_954,N_24782,N_24780);
xor UO_955 (O_955,N_24853,N_24803);
and UO_956 (O_956,N_24701,N_24999);
and UO_957 (O_957,N_24659,N_24530);
and UO_958 (O_958,N_24736,N_24749);
or UO_959 (O_959,N_24786,N_24791);
xnor UO_960 (O_960,N_24710,N_24775);
nand UO_961 (O_961,N_24961,N_24692);
or UO_962 (O_962,N_24670,N_24774);
nand UO_963 (O_963,N_24939,N_24535);
nor UO_964 (O_964,N_24965,N_24591);
xnor UO_965 (O_965,N_24748,N_24593);
nor UO_966 (O_966,N_24767,N_24695);
nand UO_967 (O_967,N_24766,N_24891);
or UO_968 (O_968,N_24544,N_24511);
and UO_969 (O_969,N_24740,N_24841);
xnor UO_970 (O_970,N_24537,N_24972);
xor UO_971 (O_971,N_24909,N_24795);
and UO_972 (O_972,N_24594,N_24611);
nor UO_973 (O_973,N_24964,N_24825);
xnor UO_974 (O_974,N_24595,N_24503);
xnor UO_975 (O_975,N_24639,N_24706);
or UO_976 (O_976,N_24947,N_24521);
xor UO_977 (O_977,N_24548,N_24541);
or UO_978 (O_978,N_24632,N_24503);
xnor UO_979 (O_979,N_24920,N_24883);
nor UO_980 (O_980,N_24968,N_24590);
nor UO_981 (O_981,N_24894,N_24967);
nor UO_982 (O_982,N_24688,N_24519);
nor UO_983 (O_983,N_24789,N_24699);
and UO_984 (O_984,N_24758,N_24780);
xor UO_985 (O_985,N_24967,N_24800);
or UO_986 (O_986,N_24857,N_24544);
and UO_987 (O_987,N_24655,N_24863);
nand UO_988 (O_988,N_24861,N_24631);
or UO_989 (O_989,N_24784,N_24993);
nand UO_990 (O_990,N_24945,N_24963);
nand UO_991 (O_991,N_24955,N_24790);
xnor UO_992 (O_992,N_24931,N_24592);
nor UO_993 (O_993,N_24648,N_24731);
or UO_994 (O_994,N_24632,N_24557);
or UO_995 (O_995,N_24946,N_24914);
xnor UO_996 (O_996,N_24794,N_24789);
or UO_997 (O_997,N_24530,N_24536);
nand UO_998 (O_998,N_24903,N_24806);
nor UO_999 (O_999,N_24936,N_24509);
and UO_1000 (O_1000,N_24669,N_24622);
xnor UO_1001 (O_1001,N_24690,N_24574);
or UO_1002 (O_1002,N_24698,N_24542);
xnor UO_1003 (O_1003,N_24783,N_24716);
nor UO_1004 (O_1004,N_24796,N_24653);
xnor UO_1005 (O_1005,N_24999,N_24506);
and UO_1006 (O_1006,N_24808,N_24750);
nand UO_1007 (O_1007,N_24511,N_24715);
nor UO_1008 (O_1008,N_24868,N_24790);
and UO_1009 (O_1009,N_24762,N_24973);
xor UO_1010 (O_1010,N_24863,N_24617);
or UO_1011 (O_1011,N_24839,N_24604);
xnor UO_1012 (O_1012,N_24815,N_24675);
and UO_1013 (O_1013,N_24772,N_24511);
and UO_1014 (O_1014,N_24957,N_24829);
nor UO_1015 (O_1015,N_24594,N_24802);
nand UO_1016 (O_1016,N_24629,N_24683);
or UO_1017 (O_1017,N_24969,N_24650);
nand UO_1018 (O_1018,N_24967,N_24852);
and UO_1019 (O_1019,N_24517,N_24802);
or UO_1020 (O_1020,N_24795,N_24901);
xor UO_1021 (O_1021,N_24616,N_24816);
nand UO_1022 (O_1022,N_24889,N_24957);
or UO_1023 (O_1023,N_24535,N_24912);
and UO_1024 (O_1024,N_24628,N_24795);
and UO_1025 (O_1025,N_24628,N_24639);
nand UO_1026 (O_1026,N_24794,N_24504);
or UO_1027 (O_1027,N_24609,N_24562);
nor UO_1028 (O_1028,N_24626,N_24996);
and UO_1029 (O_1029,N_24776,N_24763);
xnor UO_1030 (O_1030,N_24696,N_24960);
xnor UO_1031 (O_1031,N_24571,N_24804);
or UO_1032 (O_1032,N_24565,N_24837);
or UO_1033 (O_1033,N_24643,N_24769);
and UO_1034 (O_1034,N_24709,N_24900);
and UO_1035 (O_1035,N_24676,N_24862);
nor UO_1036 (O_1036,N_24534,N_24944);
nor UO_1037 (O_1037,N_24865,N_24827);
nor UO_1038 (O_1038,N_24704,N_24856);
nor UO_1039 (O_1039,N_24563,N_24893);
nand UO_1040 (O_1040,N_24577,N_24820);
xnor UO_1041 (O_1041,N_24694,N_24817);
nor UO_1042 (O_1042,N_24531,N_24806);
or UO_1043 (O_1043,N_24859,N_24724);
xnor UO_1044 (O_1044,N_24608,N_24728);
nand UO_1045 (O_1045,N_24923,N_24891);
xor UO_1046 (O_1046,N_24535,N_24878);
or UO_1047 (O_1047,N_24852,N_24506);
xor UO_1048 (O_1048,N_24583,N_24787);
nand UO_1049 (O_1049,N_24874,N_24594);
and UO_1050 (O_1050,N_24600,N_24860);
and UO_1051 (O_1051,N_24708,N_24561);
nand UO_1052 (O_1052,N_24960,N_24575);
and UO_1053 (O_1053,N_24557,N_24881);
nand UO_1054 (O_1054,N_24747,N_24566);
nand UO_1055 (O_1055,N_24940,N_24918);
nand UO_1056 (O_1056,N_24972,N_24524);
and UO_1057 (O_1057,N_24904,N_24589);
and UO_1058 (O_1058,N_24691,N_24995);
nand UO_1059 (O_1059,N_24966,N_24747);
xnor UO_1060 (O_1060,N_24838,N_24792);
or UO_1061 (O_1061,N_24624,N_24786);
or UO_1062 (O_1062,N_24501,N_24938);
or UO_1063 (O_1063,N_24665,N_24672);
xnor UO_1064 (O_1064,N_24646,N_24696);
nand UO_1065 (O_1065,N_24704,N_24716);
nand UO_1066 (O_1066,N_24664,N_24708);
nor UO_1067 (O_1067,N_24671,N_24637);
nand UO_1068 (O_1068,N_24640,N_24881);
and UO_1069 (O_1069,N_24576,N_24849);
nor UO_1070 (O_1070,N_24520,N_24786);
nor UO_1071 (O_1071,N_24727,N_24616);
or UO_1072 (O_1072,N_24756,N_24806);
nor UO_1073 (O_1073,N_24626,N_24920);
and UO_1074 (O_1074,N_24548,N_24505);
and UO_1075 (O_1075,N_24785,N_24827);
nand UO_1076 (O_1076,N_24778,N_24555);
nand UO_1077 (O_1077,N_24904,N_24501);
nand UO_1078 (O_1078,N_24502,N_24749);
and UO_1079 (O_1079,N_24913,N_24631);
xor UO_1080 (O_1080,N_24706,N_24684);
or UO_1081 (O_1081,N_24782,N_24872);
nand UO_1082 (O_1082,N_24669,N_24522);
and UO_1083 (O_1083,N_24620,N_24862);
nor UO_1084 (O_1084,N_24687,N_24925);
and UO_1085 (O_1085,N_24894,N_24637);
xnor UO_1086 (O_1086,N_24853,N_24585);
and UO_1087 (O_1087,N_24938,N_24981);
nand UO_1088 (O_1088,N_24867,N_24566);
and UO_1089 (O_1089,N_24530,N_24580);
or UO_1090 (O_1090,N_24925,N_24874);
and UO_1091 (O_1091,N_24886,N_24934);
nor UO_1092 (O_1092,N_24737,N_24562);
xor UO_1093 (O_1093,N_24750,N_24910);
or UO_1094 (O_1094,N_24985,N_24948);
and UO_1095 (O_1095,N_24958,N_24815);
nor UO_1096 (O_1096,N_24808,N_24961);
xor UO_1097 (O_1097,N_24840,N_24791);
xnor UO_1098 (O_1098,N_24847,N_24695);
and UO_1099 (O_1099,N_24745,N_24846);
xor UO_1100 (O_1100,N_24943,N_24690);
or UO_1101 (O_1101,N_24612,N_24862);
and UO_1102 (O_1102,N_24988,N_24860);
or UO_1103 (O_1103,N_24787,N_24839);
nor UO_1104 (O_1104,N_24562,N_24781);
nor UO_1105 (O_1105,N_24770,N_24919);
nor UO_1106 (O_1106,N_24871,N_24563);
xnor UO_1107 (O_1107,N_24899,N_24508);
nand UO_1108 (O_1108,N_24987,N_24502);
nand UO_1109 (O_1109,N_24551,N_24770);
xor UO_1110 (O_1110,N_24930,N_24775);
or UO_1111 (O_1111,N_24515,N_24930);
xnor UO_1112 (O_1112,N_24940,N_24788);
and UO_1113 (O_1113,N_24898,N_24827);
nor UO_1114 (O_1114,N_24894,N_24715);
nor UO_1115 (O_1115,N_24541,N_24831);
or UO_1116 (O_1116,N_24936,N_24968);
nor UO_1117 (O_1117,N_24895,N_24619);
nor UO_1118 (O_1118,N_24592,N_24638);
nor UO_1119 (O_1119,N_24659,N_24759);
or UO_1120 (O_1120,N_24662,N_24583);
nor UO_1121 (O_1121,N_24725,N_24955);
nor UO_1122 (O_1122,N_24774,N_24934);
or UO_1123 (O_1123,N_24909,N_24962);
nor UO_1124 (O_1124,N_24936,N_24915);
nor UO_1125 (O_1125,N_24502,N_24608);
nand UO_1126 (O_1126,N_24556,N_24938);
nand UO_1127 (O_1127,N_24843,N_24820);
xor UO_1128 (O_1128,N_24954,N_24771);
or UO_1129 (O_1129,N_24971,N_24725);
or UO_1130 (O_1130,N_24846,N_24708);
nor UO_1131 (O_1131,N_24580,N_24609);
and UO_1132 (O_1132,N_24615,N_24791);
nor UO_1133 (O_1133,N_24798,N_24941);
nand UO_1134 (O_1134,N_24774,N_24519);
nand UO_1135 (O_1135,N_24618,N_24526);
xor UO_1136 (O_1136,N_24769,N_24902);
and UO_1137 (O_1137,N_24605,N_24828);
nor UO_1138 (O_1138,N_24503,N_24778);
xor UO_1139 (O_1139,N_24799,N_24668);
xnor UO_1140 (O_1140,N_24588,N_24711);
nor UO_1141 (O_1141,N_24965,N_24783);
and UO_1142 (O_1142,N_24647,N_24660);
xnor UO_1143 (O_1143,N_24585,N_24897);
xor UO_1144 (O_1144,N_24988,N_24513);
nand UO_1145 (O_1145,N_24530,N_24800);
and UO_1146 (O_1146,N_24953,N_24713);
or UO_1147 (O_1147,N_24991,N_24677);
or UO_1148 (O_1148,N_24777,N_24636);
nand UO_1149 (O_1149,N_24669,N_24642);
xnor UO_1150 (O_1150,N_24922,N_24503);
nand UO_1151 (O_1151,N_24506,N_24538);
and UO_1152 (O_1152,N_24973,N_24895);
or UO_1153 (O_1153,N_24522,N_24945);
nand UO_1154 (O_1154,N_24631,N_24884);
nand UO_1155 (O_1155,N_24531,N_24953);
nand UO_1156 (O_1156,N_24743,N_24550);
and UO_1157 (O_1157,N_24891,N_24742);
and UO_1158 (O_1158,N_24840,N_24919);
xor UO_1159 (O_1159,N_24510,N_24669);
and UO_1160 (O_1160,N_24759,N_24738);
or UO_1161 (O_1161,N_24904,N_24657);
nand UO_1162 (O_1162,N_24511,N_24863);
xnor UO_1163 (O_1163,N_24559,N_24767);
xnor UO_1164 (O_1164,N_24931,N_24549);
nand UO_1165 (O_1165,N_24866,N_24725);
and UO_1166 (O_1166,N_24514,N_24897);
nor UO_1167 (O_1167,N_24894,N_24796);
xnor UO_1168 (O_1168,N_24843,N_24583);
nand UO_1169 (O_1169,N_24733,N_24541);
or UO_1170 (O_1170,N_24856,N_24586);
xnor UO_1171 (O_1171,N_24609,N_24572);
or UO_1172 (O_1172,N_24879,N_24688);
and UO_1173 (O_1173,N_24883,N_24562);
and UO_1174 (O_1174,N_24761,N_24638);
nor UO_1175 (O_1175,N_24756,N_24839);
nand UO_1176 (O_1176,N_24930,N_24858);
and UO_1177 (O_1177,N_24513,N_24502);
nor UO_1178 (O_1178,N_24719,N_24545);
nand UO_1179 (O_1179,N_24542,N_24840);
xnor UO_1180 (O_1180,N_24875,N_24846);
nor UO_1181 (O_1181,N_24897,N_24518);
nor UO_1182 (O_1182,N_24777,N_24621);
nand UO_1183 (O_1183,N_24869,N_24501);
and UO_1184 (O_1184,N_24703,N_24802);
or UO_1185 (O_1185,N_24866,N_24931);
and UO_1186 (O_1186,N_24941,N_24603);
nor UO_1187 (O_1187,N_24780,N_24645);
or UO_1188 (O_1188,N_24526,N_24807);
or UO_1189 (O_1189,N_24657,N_24694);
nand UO_1190 (O_1190,N_24645,N_24673);
nor UO_1191 (O_1191,N_24582,N_24624);
xor UO_1192 (O_1192,N_24615,N_24701);
xnor UO_1193 (O_1193,N_24768,N_24614);
and UO_1194 (O_1194,N_24549,N_24709);
xor UO_1195 (O_1195,N_24718,N_24739);
or UO_1196 (O_1196,N_24624,N_24558);
xor UO_1197 (O_1197,N_24642,N_24574);
or UO_1198 (O_1198,N_24985,N_24821);
xor UO_1199 (O_1199,N_24870,N_24621);
and UO_1200 (O_1200,N_24814,N_24584);
xnor UO_1201 (O_1201,N_24624,N_24611);
or UO_1202 (O_1202,N_24583,N_24649);
and UO_1203 (O_1203,N_24879,N_24686);
or UO_1204 (O_1204,N_24563,N_24622);
nor UO_1205 (O_1205,N_24751,N_24924);
and UO_1206 (O_1206,N_24590,N_24811);
nand UO_1207 (O_1207,N_24970,N_24558);
or UO_1208 (O_1208,N_24693,N_24661);
nor UO_1209 (O_1209,N_24877,N_24613);
nand UO_1210 (O_1210,N_24825,N_24729);
nand UO_1211 (O_1211,N_24875,N_24533);
and UO_1212 (O_1212,N_24889,N_24610);
xor UO_1213 (O_1213,N_24815,N_24588);
and UO_1214 (O_1214,N_24926,N_24817);
and UO_1215 (O_1215,N_24784,N_24902);
nor UO_1216 (O_1216,N_24686,N_24898);
or UO_1217 (O_1217,N_24582,N_24962);
and UO_1218 (O_1218,N_24548,N_24850);
or UO_1219 (O_1219,N_24545,N_24525);
nor UO_1220 (O_1220,N_24688,N_24912);
or UO_1221 (O_1221,N_24849,N_24529);
or UO_1222 (O_1222,N_24759,N_24665);
nor UO_1223 (O_1223,N_24842,N_24834);
or UO_1224 (O_1224,N_24526,N_24729);
or UO_1225 (O_1225,N_24680,N_24679);
nor UO_1226 (O_1226,N_24806,N_24703);
or UO_1227 (O_1227,N_24870,N_24725);
xnor UO_1228 (O_1228,N_24525,N_24705);
or UO_1229 (O_1229,N_24925,N_24605);
or UO_1230 (O_1230,N_24883,N_24862);
or UO_1231 (O_1231,N_24970,N_24735);
or UO_1232 (O_1232,N_24656,N_24583);
nor UO_1233 (O_1233,N_24502,N_24836);
and UO_1234 (O_1234,N_24555,N_24754);
xnor UO_1235 (O_1235,N_24860,N_24631);
xor UO_1236 (O_1236,N_24532,N_24632);
nand UO_1237 (O_1237,N_24980,N_24907);
and UO_1238 (O_1238,N_24938,N_24700);
xnor UO_1239 (O_1239,N_24777,N_24580);
nand UO_1240 (O_1240,N_24576,N_24583);
nor UO_1241 (O_1241,N_24706,N_24794);
nand UO_1242 (O_1242,N_24615,N_24868);
and UO_1243 (O_1243,N_24971,N_24607);
xor UO_1244 (O_1244,N_24919,N_24724);
and UO_1245 (O_1245,N_24597,N_24580);
nor UO_1246 (O_1246,N_24880,N_24536);
or UO_1247 (O_1247,N_24668,N_24878);
and UO_1248 (O_1248,N_24500,N_24541);
and UO_1249 (O_1249,N_24878,N_24819);
nand UO_1250 (O_1250,N_24980,N_24818);
nor UO_1251 (O_1251,N_24553,N_24806);
and UO_1252 (O_1252,N_24866,N_24580);
or UO_1253 (O_1253,N_24662,N_24921);
or UO_1254 (O_1254,N_24555,N_24508);
nand UO_1255 (O_1255,N_24904,N_24542);
nor UO_1256 (O_1256,N_24815,N_24877);
xor UO_1257 (O_1257,N_24900,N_24916);
nor UO_1258 (O_1258,N_24859,N_24629);
nor UO_1259 (O_1259,N_24653,N_24867);
nand UO_1260 (O_1260,N_24628,N_24581);
and UO_1261 (O_1261,N_24734,N_24800);
nor UO_1262 (O_1262,N_24822,N_24561);
and UO_1263 (O_1263,N_24788,N_24724);
and UO_1264 (O_1264,N_24754,N_24613);
nor UO_1265 (O_1265,N_24990,N_24572);
or UO_1266 (O_1266,N_24719,N_24958);
xor UO_1267 (O_1267,N_24581,N_24987);
or UO_1268 (O_1268,N_24928,N_24569);
nor UO_1269 (O_1269,N_24927,N_24818);
nand UO_1270 (O_1270,N_24744,N_24644);
and UO_1271 (O_1271,N_24691,N_24564);
nor UO_1272 (O_1272,N_24552,N_24829);
or UO_1273 (O_1273,N_24983,N_24694);
nand UO_1274 (O_1274,N_24594,N_24516);
xnor UO_1275 (O_1275,N_24835,N_24992);
xnor UO_1276 (O_1276,N_24601,N_24862);
or UO_1277 (O_1277,N_24995,N_24801);
nor UO_1278 (O_1278,N_24589,N_24533);
nor UO_1279 (O_1279,N_24988,N_24850);
xnor UO_1280 (O_1280,N_24958,N_24573);
xnor UO_1281 (O_1281,N_24876,N_24825);
xor UO_1282 (O_1282,N_24531,N_24671);
nor UO_1283 (O_1283,N_24769,N_24704);
xor UO_1284 (O_1284,N_24539,N_24881);
and UO_1285 (O_1285,N_24677,N_24862);
xor UO_1286 (O_1286,N_24806,N_24763);
xnor UO_1287 (O_1287,N_24692,N_24785);
xnor UO_1288 (O_1288,N_24672,N_24644);
or UO_1289 (O_1289,N_24778,N_24929);
nand UO_1290 (O_1290,N_24704,N_24653);
nor UO_1291 (O_1291,N_24580,N_24875);
nand UO_1292 (O_1292,N_24734,N_24903);
or UO_1293 (O_1293,N_24651,N_24580);
xor UO_1294 (O_1294,N_24880,N_24928);
nor UO_1295 (O_1295,N_24715,N_24655);
nor UO_1296 (O_1296,N_24666,N_24550);
nand UO_1297 (O_1297,N_24665,N_24775);
nor UO_1298 (O_1298,N_24739,N_24579);
xnor UO_1299 (O_1299,N_24990,N_24776);
or UO_1300 (O_1300,N_24881,N_24783);
nand UO_1301 (O_1301,N_24514,N_24947);
or UO_1302 (O_1302,N_24695,N_24978);
nand UO_1303 (O_1303,N_24722,N_24735);
nor UO_1304 (O_1304,N_24770,N_24785);
nor UO_1305 (O_1305,N_24957,N_24823);
or UO_1306 (O_1306,N_24957,N_24593);
or UO_1307 (O_1307,N_24797,N_24833);
nor UO_1308 (O_1308,N_24828,N_24710);
xnor UO_1309 (O_1309,N_24731,N_24915);
nand UO_1310 (O_1310,N_24628,N_24541);
and UO_1311 (O_1311,N_24924,N_24948);
or UO_1312 (O_1312,N_24635,N_24559);
and UO_1313 (O_1313,N_24882,N_24917);
or UO_1314 (O_1314,N_24944,N_24690);
and UO_1315 (O_1315,N_24852,N_24981);
nand UO_1316 (O_1316,N_24883,N_24680);
or UO_1317 (O_1317,N_24954,N_24894);
nand UO_1318 (O_1318,N_24840,N_24988);
or UO_1319 (O_1319,N_24937,N_24691);
xor UO_1320 (O_1320,N_24536,N_24507);
xor UO_1321 (O_1321,N_24636,N_24671);
and UO_1322 (O_1322,N_24657,N_24776);
nor UO_1323 (O_1323,N_24754,N_24662);
or UO_1324 (O_1324,N_24818,N_24535);
xnor UO_1325 (O_1325,N_24950,N_24649);
and UO_1326 (O_1326,N_24946,N_24630);
and UO_1327 (O_1327,N_24989,N_24571);
and UO_1328 (O_1328,N_24597,N_24686);
nor UO_1329 (O_1329,N_24516,N_24583);
xnor UO_1330 (O_1330,N_24717,N_24595);
xnor UO_1331 (O_1331,N_24795,N_24946);
or UO_1332 (O_1332,N_24704,N_24965);
nor UO_1333 (O_1333,N_24689,N_24792);
nand UO_1334 (O_1334,N_24955,N_24533);
xnor UO_1335 (O_1335,N_24743,N_24927);
and UO_1336 (O_1336,N_24951,N_24746);
nor UO_1337 (O_1337,N_24506,N_24582);
xnor UO_1338 (O_1338,N_24947,N_24881);
and UO_1339 (O_1339,N_24807,N_24543);
or UO_1340 (O_1340,N_24799,N_24560);
or UO_1341 (O_1341,N_24596,N_24911);
nand UO_1342 (O_1342,N_24611,N_24917);
xnor UO_1343 (O_1343,N_24643,N_24817);
xnor UO_1344 (O_1344,N_24950,N_24729);
xor UO_1345 (O_1345,N_24773,N_24793);
and UO_1346 (O_1346,N_24825,N_24669);
and UO_1347 (O_1347,N_24972,N_24530);
xnor UO_1348 (O_1348,N_24951,N_24982);
and UO_1349 (O_1349,N_24911,N_24914);
or UO_1350 (O_1350,N_24644,N_24772);
nand UO_1351 (O_1351,N_24921,N_24940);
xnor UO_1352 (O_1352,N_24993,N_24573);
xor UO_1353 (O_1353,N_24637,N_24621);
xnor UO_1354 (O_1354,N_24810,N_24659);
nand UO_1355 (O_1355,N_24903,N_24817);
nor UO_1356 (O_1356,N_24996,N_24718);
nor UO_1357 (O_1357,N_24812,N_24997);
nand UO_1358 (O_1358,N_24966,N_24810);
or UO_1359 (O_1359,N_24921,N_24590);
and UO_1360 (O_1360,N_24860,N_24594);
nand UO_1361 (O_1361,N_24779,N_24728);
nand UO_1362 (O_1362,N_24937,N_24742);
nor UO_1363 (O_1363,N_24526,N_24614);
nor UO_1364 (O_1364,N_24568,N_24841);
nor UO_1365 (O_1365,N_24785,N_24779);
xor UO_1366 (O_1366,N_24579,N_24767);
nand UO_1367 (O_1367,N_24522,N_24919);
or UO_1368 (O_1368,N_24627,N_24679);
nor UO_1369 (O_1369,N_24558,N_24658);
xor UO_1370 (O_1370,N_24603,N_24979);
nand UO_1371 (O_1371,N_24935,N_24636);
nand UO_1372 (O_1372,N_24666,N_24989);
nand UO_1373 (O_1373,N_24627,N_24565);
nor UO_1374 (O_1374,N_24511,N_24859);
or UO_1375 (O_1375,N_24935,N_24704);
xor UO_1376 (O_1376,N_24948,N_24516);
or UO_1377 (O_1377,N_24981,N_24575);
xor UO_1378 (O_1378,N_24864,N_24844);
and UO_1379 (O_1379,N_24802,N_24581);
nor UO_1380 (O_1380,N_24763,N_24829);
xnor UO_1381 (O_1381,N_24842,N_24985);
nor UO_1382 (O_1382,N_24685,N_24983);
nor UO_1383 (O_1383,N_24504,N_24572);
and UO_1384 (O_1384,N_24791,N_24726);
and UO_1385 (O_1385,N_24609,N_24697);
xor UO_1386 (O_1386,N_24672,N_24527);
nand UO_1387 (O_1387,N_24642,N_24613);
xnor UO_1388 (O_1388,N_24669,N_24729);
xor UO_1389 (O_1389,N_24617,N_24514);
nor UO_1390 (O_1390,N_24730,N_24718);
nor UO_1391 (O_1391,N_24689,N_24760);
or UO_1392 (O_1392,N_24689,N_24865);
xor UO_1393 (O_1393,N_24903,N_24500);
and UO_1394 (O_1394,N_24605,N_24633);
or UO_1395 (O_1395,N_24846,N_24506);
xnor UO_1396 (O_1396,N_24768,N_24883);
and UO_1397 (O_1397,N_24529,N_24866);
nor UO_1398 (O_1398,N_24824,N_24613);
xor UO_1399 (O_1399,N_24839,N_24509);
nand UO_1400 (O_1400,N_24536,N_24727);
nand UO_1401 (O_1401,N_24638,N_24566);
or UO_1402 (O_1402,N_24618,N_24633);
xnor UO_1403 (O_1403,N_24694,N_24556);
and UO_1404 (O_1404,N_24825,N_24745);
xor UO_1405 (O_1405,N_24585,N_24703);
xor UO_1406 (O_1406,N_24802,N_24589);
or UO_1407 (O_1407,N_24772,N_24767);
nand UO_1408 (O_1408,N_24600,N_24947);
nand UO_1409 (O_1409,N_24619,N_24965);
nand UO_1410 (O_1410,N_24726,N_24740);
xnor UO_1411 (O_1411,N_24854,N_24512);
and UO_1412 (O_1412,N_24629,N_24577);
xnor UO_1413 (O_1413,N_24505,N_24616);
xnor UO_1414 (O_1414,N_24950,N_24560);
xnor UO_1415 (O_1415,N_24780,N_24989);
xor UO_1416 (O_1416,N_24867,N_24888);
nor UO_1417 (O_1417,N_24758,N_24667);
or UO_1418 (O_1418,N_24612,N_24819);
xnor UO_1419 (O_1419,N_24918,N_24631);
nand UO_1420 (O_1420,N_24524,N_24926);
nand UO_1421 (O_1421,N_24519,N_24959);
xnor UO_1422 (O_1422,N_24986,N_24998);
nand UO_1423 (O_1423,N_24832,N_24799);
nor UO_1424 (O_1424,N_24735,N_24942);
nor UO_1425 (O_1425,N_24861,N_24865);
and UO_1426 (O_1426,N_24563,N_24592);
and UO_1427 (O_1427,N_24822,N_24583);
and UO_1428 (O_1428,N_24995,N_24582);
xnor UO_1429 (O_1429,N_24515,N_24635);
nand UO_1430 (O_1430,N_24608,N_24786);
xor UO_1431 (O_1431,N_24776,N_24882);
nand UO_1432 (O_1432,N_24603,N_24800);
and UO_1433 (O_1433,N_24944,N_24879);
xor UO_1434 (O_1434,N_24586,N_24551);
or UO_1435 (O_1435,N_24547,N_24688);
or UO_1436 (O_1436,N_24812,N_24649);
xor UO_1437 (O_1437,N_24736,N_24572);
xor UO_1438 (O_1438,N_24904,N_24834);
nor UO_1439 (O_1439,N_24536,N_24523);
and UO_1440 (O_1440,N_24724,N_24708);
nand UO_1441 (O_1441,N_24788,N_24927);
nand UO_1442 (O_1442,N_24637,N_24594);
nor UO_1443 (O_1443,N_24534,N_24663);
or UO_1444 (O_1444,N_24944,N_24564);
xnor UO_1445 (O_1445,N_24551,N_24793);
xor UO_1446 (O_1446,N_24621,N_24612);
or UO_1447 (O_1447,N_24734,N_24921);
xnor UO_1448 (O_1448,N_24962,N_24719);
nor UO_1449 (O_1449,N_24826,N_24900);
nor UO_1450 (O_1450,N_24664,N_24801);
xor UO_1451 (O_1451,N_24632,N_24660);
or UO_1452 (O_1452,N_24998,N_24520);
or UO_1453 (O_1453,N_24517,N_24631);
or UO_1454 (O_1454,N_24671,N_24928);
nand UO_1455 (O_1455,N_24916,N_24699);
and UO_1456 (O_1456,N_24684,N_24938);
and UO_1457 (O_1457,N_24717,N_24897);
xor UO_1458 (O_1458,N_24858,N_24607);
and UO_1459 (O_1459,N_24951,N_24578);
nor UO_1460 (O_1460,N_24706,N_24740);
nand UO_1461 (O_1461,N_24789,N_24527);
nor UO_1462 (O_1462,N_24677,N_24645);
nand UO_1463 (O_1463,N_24690,N_24691);
nor UO_1464 (O_1464,N_24799,N_24585);
nand UO_1465 (O_1465,N_24998,N_24848);
xor UO_1466 (O_1466,N_24726,N_24708);
or UO_1467 (O_1467,N_24761,N_24910);
or UO_1468 (O_1468,N_24803,N_24651);
nand UO_1469 (O_1469,N_24893,N_24714);
or UO_1470 (O_1470,N_24966,N_24700);
or UO_1471 (O_1471,N_24763,N_24716);
nor UO_1472 (O_1472,N_24722,N_24998);
nor UO_1473 (O_1473,N_24583,N_24547);
and UO_1474 (O_1474,N_24929,N_24899);
and UO_1475 (O_1475,N_24910,N_24826);
or UO_1476 (O_1476,N_24698,N_24738);
nand UO_1477 (O_1477,N_24581,N_24641);
nand UO_1478 (O_1478,N_24997,N_24791);
or UO_1479 (O_1479,N_24995,N_24816);
and UO_1480 (O_1480,N_24884,N_24619);
and UO_1481 (O_1481,N_24917,N_24928);
nand UO_1482 (O_1482,N_24911,N_24546);
nand UO_1483 (O_1483,N_24979,N_24738);
and UO_1484 (O_1484,N_24672,N_24575);
and UO_1485 (O_1485,N_24547,N_24618);
nor UO_1486 (O_1486,N_24714,N_24634);
nand UO_1487 (O_1487,N_24818,N_24954);
xnor UO_1488 (O_1488,N_24599,N_24750);
and UO_1489 (O_1489,N_24798,N_24965);
nor UO_1490 (O_1490,N_24878,N_24908);
or UO_1491 (O_1491,N_24756,N_24981);
and UO_1492 (O_1492,N_24910,N_24640);
xnor UO_1493 (O_1493,N_24871,N_24644);
or UO_1494 (O_1494,N_24884,N_24613);
and UO_1495 (O_1495,N_24837,N_24918);
xor UO_1496 (O_1496,N_24797,N_24587);
nor UO_1497 (O_1497,N_24842,N_24969);
and UO_1498 (O_1498,N_24976,N_24640);
nand UO_1499 (O_1499,N_24698,N_24801);
nand UO_1500 (O_1500,N_24646,N_24988);
nor UO_1501 (O_1501,N_24568,N_24664);
or UO_1502 (O_1502,N_24720,N_24731);
xnor UO_1503 (O_1503,N_24849,N_24575);
or UO_1504 (O_1504,N_24507,N_24704);
nor UO_1505 (O_1505,N_24739,N_24875);
and UO_1506 (O_1506,N_24601,N_24903);
and UO_1507 (O_1507,N_24690,N_24726);
nand UO_1508 (O_1508,N_24642,N_24753);
xnor UO_1509 (O_1509,N_24730,N_24865);
xnor UO_1510 (O_1510,N_24914,N_24690);
nor UO_1511 (O_1511,N_24997,N_24850);
or UO_1512 (O_1512,N_24744,N_24684);
or UO_1513 (O_1513,N_24949,N_24659);
nor UO_1514 (O_1514,N_24686,N_24828);
nand UO_1515 (O_1515,N_24709,N_24927);
and UO_1516 (O_1516,N_24950,N_24929);
or UO_1517 (O_1517,N_24530,N_24834);
and UO_1518 (O_1518,N_24625,N_24782);
xnor UO_1519 (O_1519,N_24659,N_24696);
or UO_1520 (O_1520,N_24749,N_24812);
and UO_1521 (O_1521,N_24901,N_24951);
xor UO_1522 (O_1522,N_24636,N_24533);
and UO_1523 (O_1523,N_24583,N_24683);
and UO_1524 (O_1524,N_24795,N_24871);
xnor UO_1525 (O_1525,N_24645,N_24905);
nor UO_1526 (O_1526,N_24951,N_24728);
or UO_1527 (O_1527,N_24782,N_24748);
nor UO_1528 (O_1528,N_24716,N_24854);
nor UO_1529 (O_1529,N_24755,N_24715);
or UO_1530 (O_1530,N_24685,N_24524);
and UO_1531 (O_1531,N_24595,N_24973);
and UO_1532 (O_1532,N_24808,N_24655);
nand UO_1533 (O_1533,N_24938,N_24613);
nor UO_1534 (O_1534,N_24869,N_24645);
xor UO_1535 (O_1535,N_24986,N_24712);
xor UO_1536 (O_1536,N_24763,N_24648);
xnor UO_1537 (O_1537,N_24974,N_24818);
or UO_1538 (O_1538,N_24804,N_24522);
xor UO_1539 (O_1539,N_24776,N_24609);
xor UO_1540 (O_1540,N_24541,N_24774);
and UO_1541 (O_1541,N_24520,N_24769);
or UO_1542 (O_1542,N_24968,N_24827);
and UO_1543 (O_1543,N_24806,N_24582);
or UO_1544 (O_1544,N_24543,N_24692);
xnor UO_1545 (O_1545,N_24943,N_24555);
or UO_1546 (O_1546,N_24993,N_24769);
nor UO_1547 (O_1547,N_24594,N_24852);
xnor UO_1548 (O_1548,N_24764,N_24717);
nand UO_1549 (O_1549,N_24548,N_24893);
and UO_1550 (O_1550,N_24553,N_24514);
nand UO_1551 (O_1551,N_24506,N_24574);
and UO_1552 (O_1552,N_24843,N_24628);
and UO_1553 (O_1553,N_24742,N_24523);
or UO_1554 (O_1554,N_24578,N_24813);
xnor UO_1555 (O_1555,N_24897,N_24709);
nand UO_1556 (O_1556,N_24871,N_24901);
and UO_1557 (O_1557,N_24934,N_24581);
nor UO_1558 (O_1558,N_24922,N_24924);
or UO_1559 (O_1559,N_24774,N_24940);
and UO_1560 (O_1560,N_24750,N_24662);
or UO_1561 (O_1561,N_24590,N_24591);
or UO_1562 (O_1562,N_24992,N_24682);
nor UO_1563 (O_1563,N_24912,N_24826);
nand UO_1564 (O_1564,N_24538,N_24608);
xnor UO_1565 (O_1565,N_24699,N_24586);
nand UO_1566 (O_1566,N_24521,N_24685);
xor UO_1567 (O_1567,N_24619,N_24818);
nor UO_1568 (O_1568,N_24732,N_24842);
nand UO_1569 (O_1569,N_24549,N_24518);
nor UO_1570 (O_1570,N_24707,N_24585);
and UO_1571 (O_1571,N_24850,N_24832);
nor UO_1572 (O_1572,N_24747,N_24785);
xnor UO_1573 (O_1573,N_24982,N_24625);
or UO_1574 (O_1574,N_24676,N_24771);
xnor UO_1575 (O_1575,N_24693,N_24850);
nor UO_1576 (O_1576,N_24760,N_24601);
nor UO_1577 (O_1577,N_24542,N_24699);
nor UO_1578 (O_1578,N_24743,N_24843);
nor UO_1579 (O_1579,N_24679,N_24971);
nor UO_1580 (O_1580,N_24702,N_24512);
or UO_1581 (O_1581,N_24520,N_24697);
xnor UO_1582 (O_1582,N_24912,N_24691);
nand UO_1583 (O_1583,N_24622,N_24831);
or UO_1584 (O_1584,N_24638,N_24532);
xnor UO_1585 (O_1585,N_24895,N_24775);
or UO_1586 (O_1586,N_24856,N_24640);
nand UO_1587 (O_1587,N_24883,N_24647);
xor UO_1588 (O_1588,N_24549,N_24776);
nor UO_1589 (O_1589,N_24709,N_24788);
or UO_1590 (O_1590,N_24814,N_24841);
and UO_1591 (O_1591,N_24869,N_24586);
nand UO_1592 (O_1592,N_24810,N_24741);
and UO_1593 (O_1593,N_24763,N_24869);
or UO_1594 (O_1594,N_24507,N_24738);
nor UO_1595 (O_1595,N_24976,N_24554);
nand UO_1596 (O_1596,N_24564,N_24525);
nand UO_1597 (O_1597,N_24958,N_24578);
nor UO_1598 (O_1598,N_24582,N_24943);
or UO_1599 (O_1599,N_24885,N_24958);
nor UO_1600 (O_1600,N_24852,N_24745);
or UO_1601 (O_1601,N_24869,N_24912);
or UO_1602 (O_1602,N_24558,N_24818);
xnor UO_1603 (O_1603,N_24873,N_24696);
nand UO_1604 (O_1604,N_24590,N_24536);
nor UO_1605 (O_1605,N_24502,N_24875);
nor UO_1606 (O_1606,N_24618,N_24551);
nor UO_1607 (O_1607,N_24554,N_24909);
xnor UO_1608 (O_1608,N_24636,N_24863);
xor UO_1609 (O_1609,N_24543,N_24672);
nor UO_1610 (O_1610,N_24814,N_24780);
xnor UO_1611 (O_1611,N_24528,N_24755);
or UO_1612 (O_1612,N_24585,N_24928);
and UO_1613 (O_1613,N_24752,N_24771);
nor UO_1614 (O_1614,N_24531,N_24878);
and UO_1615 (O_1615,N_24651,N_24754);
and UO_1616 (O_1616,N_24571,N_24536);
or UO_1617 (O_1617,N_24914,N_24550);
xnor UO_1618 (O_1618,N_24937,N_24570);
nand UO_1619 (O_1619,N_24606,N_24703);
nor UO_1620 (O_1620,N_24584,N_24916);
xnor UO_1621 (O_1621,N_24698,N_24644);
nor UO_1622 (O_1622,N_24777,N_24831);
nor UO_1623 (O_1623,N_24827,N_24915);
and UO_1624 (O_1624,N_24631,N_24691);
nand UO_1625 (O_1625,N_24657,N_24519);
xnor UO_1626 (O_1626,N_24593,N_24854);
nor UO_1627 (O_1627,N_24801,N_24585);
nor UO_1628 (O_1628,N_24918,N_24539);
or UO_1629 (O_1629,N_24784,N_24732);
xor UO_1630 (O_1630,N_24537,N_24529);
or UO_1631 (O_1631,N_24700,N_24703);
or UO_1632 (O_1632,N_24764,N_24745);
xor UO_1633 (O_1633,N_24903,N_24642);
nor UO_1634 (O_1634,N_24683,N_24578);
nor UO_1635 (O_1635,N_24825,N_24836);
nand UO_1636 (O_1636,N_24651,N_24799);
nor UO_1637 (O_1637,N_24978,N_24917);
or UO_1638 (O_1638,N_24905,N_24893);
and UO_1639 (O_1639,N_24617,N_24605);
and UO_1640 (O_1640,N_24761,N_24890);
xor UO_1641 (O_1641,N_24509,N_24539);
nor UO_1642 (O_1642,N_24780,N_24828);
nor UO_1643 (O_1643,N_24670,N_24516);
nand UO_1644 (O_1644,N_24545,N_24635);
nor UO_1645 (O_1645,N_24638,N_24560);
and UO_1646 (O_1646,N_24888,N_24979);
nand UO_1647 (O_1647,N_24652,N_24618);
xor UO_1648 (O_1648,N_24796,N_24606);
nor UO_1649 (O_1649,N_24823,N_24870);
nor UO_1650 (O_1650,N_24923,N_24965);
and UO_1651 (O_1651,N_24899,N_24735);
or UO_1652 (O_1652,N_24697,N_24830);
xor UO_1653 (O_1653,N_24985,N_24918);
xnor UO_1654 (O_1654,N_24883,N_24629);
xor UO_1655 (O_1655,N_24787,N_24738);
nand UO_1656 (O_1656,N_24747,N_24546);
nand UO_1657 (O_1657,N_24843,N_24863);
nand UO_1658 (O_1658,N_24781,N_24570);
xor UO_1659 (O_1659,N_24904,N_24933);
and UO_1660 (O_1660,N_24760,N_24786);
nand UO_1661 (O_1661,N_24752,N_24866);
and UO_1662 (O_1662,N_24721,N_24584);
nand UO_1663 (O_1663,N_24687,N_24948);
or UO_1664 (O_1664,N_24610,N_24842);
xor UO_1665 (O_1665,N_24990,N_24598);
xnor UO_1666 (O_1666,N_24945,N_24656);
or UO_1667 (O_1667,N_24871,N_24595);
nand UO_1668 (O_1668,N_24563,N_24800);
or UO_1669 (O_1669,N_24870,N_24815);
nand UO_1670 (O_1670,N_24631,N_24596);
or UO_1671 (O_1671,N_24932,N_24591);
and UO_1672 (O_1672,N_24711,N_24789);
and UO_1673 (O_1673,N_24686,N_24972);
xnor UO_1674 (O_1674,N_24770,N_24556);
and UO_1675 (O_1675,N_24690,N_24776);
nor UO_1676 (O_1676,N_24535,N_24764);
and UO_1677 (O_1677,N_24572,N_24579);
and UO_1678 (O_1678,N_24594,N_24944);
or UO_1679 (O_1679,N_24829,N_24568);
nand UO_1680 (O_1680,N_24849,N_24670);
nor UO_1681 (O_1681,N_24650,N_24918);
and UO_1682 (O_1682,N_24685,N_24916);
or UO_1683 (O_1683,N_24535,N_24506);
xnor UO_1684 (O_1684,N_24974,N_24515);
xor UO_1685 (O_1685,N_24885,N_24949);
xor UO_1686 (O_1686,N_24990,N_24761);
nand UO_1687 (O_1687,N_24849,N_24681);
and UO_1688 (O_1688,N_24570,N_24950);
and UO_1689 (O_1689,N_24516,N_24849);
nor UO_1690 (O_1690,N_24930,N_24665);
nand UO_1691 (O_1691,N_24761,N_24766);
nand UO_1692 (O_1692,N_24812,N_24695);
nand UO_1693 (O_1693,N_24576,N_24828);
and UO_1694 (O_1694,N_24850,N_24998);
xor UO_1695 (O_1695,N_24680,N_24651);
xnor UO_1696 (O_1696,N_24945,N_24605);
or UO_1697 (O_1697,N_24591,N_24754);
or UO_1698 (O_1698,N_24846,N_24520);
xor UO_1699 (O_1699,N_24997,N_24707);
nor UO_1700 (O_1700,N_24950,N_24643);
and UO_1701 (O_1701,N_24770,N_24667);
and UO_1702 (O_1702,N_24750,N_24896);
and UO_1703 (O_1703,N_24845,N_24604);
xnor UO_1704 (O_1704,N_24963,N_24697);
nor UO_1705 (O_1705,N_24588,N_24931);
and UO_1706 (O_1706,N_24814,N_24748);
or UO_1707 (O_1707,N_24825,N_24547);
xnor UO_1708 (O_1708,N_24674,N_24609);
nand UO_1709 (O_1709,N_24515,N_24604);
nand UO_1710 (O_1710,N_24768,N_24751);
nor UO_1711 (O_1711,N_24898,N_24967);
or UO_1712 (O_1712,N_24949,N_24549);
or UO_1713 (O_1713,N_24911,N_24716);
xor UO_1714 (O_1714,N_24573,N_24770);
or UO_1715 (O_1715,N_24837,N_24648);
and UO_1716 (O_1716,N_24521,N_24543);
and UO_1717 (O_1717,N_24603,N_24507);
nand UO_1718 (O_1718,N_24610,N_24600);
nor UO_1719 (O_1719,N_24537,N_24706);
or UO_1720 (O_1720,N_24542,N_24922);
or UO_1721 (O_1721,N_24922,N_24989);
xnor UO_1722 (O_1722,N_24793,N_24564);
or UO_1723 (O_1723,N_24841,N_24937);
xnor UO_1724 (O_1724,N_24561,N_24696);
nor UO_1725 (O_1725,N_24614,N_24866);
nand UO_1726 (O_1726,N_24779,N_24816);
xor UO_1727 (O_1727,N_24714,N_24542);
xor UO_1728 (O_1728,N_24582,N_24988);
nor UO_1729 (O_1729,N_24895,N_24965);
nand UO_1730 (O_1730,N_24814,N_24761);
nand UO_1731 (O_1731,N_24534,N_24520);
xor UO_1732 (O_1732,N_24691,N_24752);
and UO_1733 (O_1733,N_24769,N_24793);
nor UO_1734 (O_1734,N_24989,N_24905);
and UO_1735 (O_1735,N_24853,N_24547);
and UO_1736 (O_1736,N_24520,N_24834);
and UO_1737 (O_1737,N_24516,N_24765);
or UO_1738 (O_1738,N_24982,N_24839);
nand UO_1739 (O_1739,N_24631,N_24637);
nor UO_1740 (O_1740,N_24709,N_24551);
and UO_1741 (O_1741,N_24590,N_24633);
xnor UO_1742 (O_1742,N_24556,N_24816);
nand UO_1743 (O_1743,N_24832,N_24875);
and UO_1744 (O_1744,N_24516,N_24866);
xnor UO_1745 (O_1745,N_24601,N_24618);
or UO_1746 (O_1746,N_24735,N_24690);
or UO_1747 (O_1747,N_24723,N_24788);
xnor UO_1748 (O_1748,N_24687,N_24582);
xnor UO_1749 (O_1749,N_24975,N_24597);
nand UO_1750 (O_1750,N_24863,N_24664);
nand UO_1751 (O_1751,N_24584,N_24996);
and UO_1752 (O_1752,N_24644,N_24860);
nand UO_1753 (O_1753,N_24736,N_24581);
and UO_1754 (O_1754,N_24927,N_24971);
nor UO_1755 (O_1755,N_24542,N_24661);
xnor UO_1756 (O_1756,N_24658,N_24784);
xnor UO_1757 (O_1757,N_24904,N_24752);
nand UO_1758 (O_1758,N_24978,N_24893);
and UO_1759 (O_1759,N_24665,N_24825);
or UO_1760 (O_1760,N_24943,N_24639);
and UO_1761 (O_1761,N_24765,N_24708);
nor UO_1762 (O_1762,N_24619,N_24539);
and UO_1763 (O_1763,N_24819,N_24619);
nor UO_1764 (O_1764,N_24779,N_24801);
xor UO_1765 (O_1765,N_24570,N_24568);
nor UO_1766 (O_1766,N_24830,N_24614);
and UO_1767 (O_1767,N_24622,N_24644);
xnor UO_1768 (O_1768,N_24908,N_24997);
and UO_1769 (O_1769,N_24658,N_24638);
nor UO_1770 (O_1770,N_24530,N_24898);
nand UO_1771 (O_1771,N_24838,N_24847);
nor UO_1772 (O_1772,N_24807,N_24529);
and UO_1773 (O_1773,N_24845,N_24621);
and UO_1774 (O_1774,N_24737,N_24962);
or UO_1775 (O_1775,N_24782,N_24966);
xor UO_1776 (O_1776,N_24710,N_24612);
or UO_1777 (O_1777,N_24841,N_24990);
or UO_1778 (O_1778,N_24612,N_24978);
nand UO_1779 (O_1779,N_24748,N_24984);
xor UO_1780 (O_1780,N_24743,N_24948);
xnor UO_1781 (O_1781,N_24829,N_24625);
xor UO_1782 (O_1782,N_24985,N_24787);
nand UO_1783 (O_1783,N_24787,N_24845);
xnor UO_1784 (O_1784,N_24898,N_24789);
nand UO_1785 (O_1785,N_24784,N_24816);
or UO_1786 (O_1786,N_24887,N_24584);
xnor UO_1787 (O_1787,N_24763,N_24847);
and UO_1788 (O_1788,N_24663,N_24886);
and UO_1789 (O_1789,N_24963,N_24900);
xnor UO_1790 (O_1790,N_24610,N_24752);
and UO_1791 (O_1791,N_24764,N_24706);
nor UO_1792 (O_1792,N_24988,N_24929);
xor UO_1793 (O_1793,N_24883,N_24665);
nand UO_1794 (O_1794,N_24724,N_24609);
nor UO_1795 (O_1795,N_24648,N_24512);
nor UO_1796 (O_1796,N_24962,N_24802);
and UO_1797 (O_1797,N_24578,N_24619);
nor UO_1798 (O_1798,N_24715,N_24629);
and UO_1799 (O_1799,N_24769,N_24984);
xnor UO_1800 (O_1800,N_24883,N_24725);
nor UO_1801 (O_1801,N_24555,N_24944);
nand UO_1802 (O_1802,N_24645,N_24851);
nor UO_1803 (O_1803,N_24881,N_24988);
xnor UO_1804 (O_1804,N_24929,N_24771);
nor UO_1805 (O_1805,N_24637,N_24842);
xnor UO_1806 (O_1806,N_24649,N_24817);
xnor UO_1807 (O_1807,N_24883,N_24690);
and UO_1808 (O_1808,N_24957,N_24702);
xor UO_1809 (O_1809,N_24705,N_24949);
or UO_1810 (O_1810,N_24639,N_24616);
xor UO_1811 (O_1811,N_24518,N_24749);
xnor UO_1812 (O_1812,N_24954,N_24885);
and UO_1813 (O_1813,N_24703,N_24953);
and UO_1814 (O_1814,N_24835,N_24804);
and UO_1815 (O_1815,N_24986,N_24881);
xor UO_1816 (O_1816,N_24830,N_24940);
or UO_1817 (O_1817,N_24512,N_24681);
or UO_1818 (O_1818,N_24827,N_24700);
and UO_1819 (O_1819,N_24913,N_24699);
xnor UO_1820 (O_1820,N_24804,N_24599);
or UO_1821 (O_1821,N_24983,N_24870);
and UO_1822 (O_1822,N_24610,N_24719);
and UO_1823 (O_1823,N_24775,N_24934);
or UO_1824 (O_1824,N_24912,N_24703);
and UO_1825 (O_1825,N_24618,N_24784);
or UO_1826 (O_1826,N_24856,N_24733);
nand UO_1827 (O_1827,N_24680,N_24736);
xor UO_1828 (O_1828,N_24872,N_24971);
xnor UO_1829 (O_1829,N_24559,N_24682);
or UO_1830 (O_1830,N_24542,N_24934);
or UO_1831 (O_1831,N_24788,N_24785);
or UO_1832 (O_1832,N_24518,N_24571);
nor UO_1833 (O_1833,N_24721,N_24974);
nand UO_1834 (O_1834,N_24590,N_24594);
xnor UO_1835 (O_1835,N_24932,N_24522);
nand UO_1836 (O_1836,N_24886,N_24889);
xor UO_1837 (O_1837,N_24521,N_24959);
nor UO_1838 (O_1838,N_24687,N_24695);
nand UO_1839 (O_1839,N_24964,N_24934);
and UO_1840 (O_1840,N_24680,N_24887);
nor UO_1841 (O_1841,N_24714,N_24749);
nand UO_1842 (O_1842,N_24500,N_24730);
nand UO_1843 (O_1843,N_24604,N_24935);
xnor UO_1844 (O_1844,N_24583,N_24771);
nor UO_1845 (O_1845,N_24808,N_24583);
or UO_1846 (O_1846,N_24871,N_24910);
nor UO_1847 (O_1847,N_24965,N_24903);
or UO_1848 (O_1848,N_24999,N_24959);
or UO_1849 (O_1849,N_24734,N_24601);
and UO_1850 (O_1850,N_24623,N_24502);
xnor UO_1851 (O_1851,N_24582,N_24557);
nand UO_1852 (O_1852,N_24708,N_24675);
nand UO_1853 (O_1853,N_24664,N_24983);
or UO_1854 (O_1854,N_24634,N_24684);
or UO_1855 (O_1855,N_24848,N_24777);
nand UO_1856 (O_1856,N_24740,N_24521);
and UO_1857 (O_1857,N_24699,N_24578);
and UO_1858 (O_1858,N_24574,N_24805);
and UO_1859 (O_1859,N_24889,N_24857);
nor UO_1860 (O_1860,N_24905,N_24914);
and UO_1861 (O_1861,N_24660,N_24510);
or UO_1862 (O_1862,N_24969,N_24587);
or UO_1863 (O_1863,N_24791,N_24783);
xor UO_1864 (O_1864,N_24657,N_24889);
and UO_1865 (O_1865,N_24574,N_24857);
nand UO_1866 (O_1866,N_24891,N_24903);
and UO_1867 (O_1867,N_24732,N_24559);
or UO_1868 (O_1868,N_24697,N_24836);
or UO_1869 (O_1869,N_24943,N_24928);
nand UO_1870 (O_1870,N_24764,N_24643);
xnor UO_1871 (O_1871,N_24861,N_24737);
and UO_1872 (O_1872,N_24937,N_24875);
and UO_1873 (O_1873,N_24833,N_24801);
or UO_1874 (O_1874,N_24709,N_24737);
nor UO_1875 (O_1875,N_24518,N_24506);
nor UO_1876 (O_1876,N_24926,N_24765);
or UO_1877 (O_1877,N_24601,N_24940);
xor UO_1878 (O_1878,N_24993,N_24531);
and UO_1879 (O_1879,N_24721,N_24557);
nor UO_1880 (O_1880,N_24888,N_24532);
or UO_1881 (O_1881,N_24754,N_24645);
or UO_1882 (O_1882,N_24818,N_24988);
nand UO_1883 (O_1883,N_24869,N_24706);
nand UO_1884 (O_1884,N_24658,N_24749);
nand UO_1885 (O_1885,N_24615,N_24879);
nor UO_1886 (O_1886,N_24716,N_24759);
or UO_1887 (O_1887,N_24952,N_24757);
xor UO_1888 (O_1888,N_24811,N_24538);
and UO_1889 (O_1889,N_24849,N_24583);
or UO_1890 (O_1890,N_24909,N_24531);
or UO_1891 (O_1891,N_24976,N_24924);
xnor UO_1892 (O_1892,N_24922,N_24929);
xnor UO_1893 (O_1893,N_24617,N_24635);
or UO_1894 (O_1894,N_24634,N_24605);
nand UO_1895 (O_1895,N_24797,N_24935);
nor UO_1896 (O_1896,N_24792,N_24887);
nor UO_1897 (O_1897,N_24883,N_24893);
and UO_1898 (O_1898,N_24637,N_24670);
and UO_1899 (O_1899,N_24717,N_24757);
and UO_1900 (O_1900,N_24990,N_24768);
and UO_1901 (O_1901,N_24730,N_24510);
nor UO_1902 (O_1902,N_24629,N_24953);
or UO_1903 (O_1903,N_24968,N_24813);
and UO_1904 (O_1904,N_24591,N_24828);
nand UO_1905 (O_1905,N_24650,N_24596);
nand UO_1906 (O_1906,N_24959,N_24751);
xnor UO_1907 (O_1907,N_24801,N_24579);
xnor UO_1908 (O_1908,N_24606,N_24883);
and UO_1909 (O_1909,N_24704,N_24753);
xnor UO_1910 (O_1910,N_24585,N_24810);
or UO_1911 (O_1911,N_24593,N_24577);
nand UO_1912 (O_1912,N_24954,N_24883);
nor UO_1913 (O_1913,N_24592,N_24739);
nor UO_1914 (O_1914,N_24531,N_24810);
nand UO_1915 (O_1915,N_24814,N_24732);
or UO_1916 (O_1916,N_24984,N_24938);
nand UO_1917 (O_1917,N_24778,N_24974);
nor UO_1918 (O_1918,N_24842,N_24813);
nor UO_1919 (O_1919,N_24956,N_24809);
or UO_1920 (O_1920,N_24602,N_24658);
xnor UO_1921 (O_1921,N_24877,N_24968);
and UO_1922 (O_1922,N_24611,N_24592);
nand UO_1923 (O_1923,N_24880,N_24683);
xnor UO_1924 (O_1924,N_24569,N_24868);
nor UO_1925 (O_1925,N_24530,N_24544);
nand UO_1926 (O_1926,N_24783,N_24964);
xor UO_1927 (O_1927,N_24599,N_24879);
nor UO_1928 (O_1928,N_24707,N_24521);
and UO_1929 (O_1929,N_24962,N_24769);
xnor UO_1930 (O_1930,N_24915,N_24769);
nor UO_1931 (O_1931,N_24505,N_24923);
and UO_1932 (O_1932,N_24707,N_24786);
nand UO_1933 (O_1933,N_24722,N_24649);
xor UO_1934 (O_1934,N_24601,N_24913);
xnor UO_1935 (O_1935,N_24864,N_24531);
nand UO_1936 (O_1936,N_24874,N_24541);
xor UO_1937 (O_1937,N_24665,N_24772);
nand UO_1938 (O_1938,N_24805,N_24626);
nand UO_1939 (O_1939,N_24750,N_24939);
and UO_1940 (O_1940,N_24737,N_24593);
xnor UO_1941 (O_1941,N_24755,N_24915);
or UO_1942 (O_1942,N_24912,N_24761);
and UO_1943 (O_1943,N_24633,N_24725);
and UO_1944 (O_1944,N_24943,N_24742);
xnor UO_1945 (O_1945,N_24950,N_24702);
or UO_1946 (O_1946,N_24991,N_24963);
and UO_1947 (O_1947,N_24557,N_24543);
nand UO_1948 (O_1948,N_24839,N_24746);
xor UO_1949 (O_1949,N_24622,N_24509);
nor UO_1950 (O_1950,N_24541,N_24924);
and UO_1951 (O_1951,N_24701,N_24791);
and UO_1952 (O_1952,N_24785,N_24860);
nor UO_1953 (O_1953,N_24729,N_24609);
or UO_1954 (O_1954,N_24650,N_24881);
xor UO_1955 (O_1955,N_24568,N_24519);
and UO_1956 (O_1956,N_24763,N_24821);
xnor UO_1957 (O_1957,N_24865,N_24588);
and UO_1958 (O_1958,N_24613,N_24667);
xnor UO_1959 (O_1959,N_24996,N_24968);
or UO_1960 (O_1960,N_24549,N_24540);
nand UO_1961 (O_1961,N_24943,N_24812);
nor UO_1962 (O_1962,N_24954,N_24963);
nor UO_1963 (O_1963,N_24738,N_24959);
xnor UO_1964 (O_1964,N_24692,N_24753);
nor UO_1965 (O_1965,N_24967,N_24777);
xnor UO_1966 (O_1966,N_24688,N_24843);
or UO_1967 (O_1967,N_24722,N_24835);
or UO_1968 (O_1968,N_24685,N_24760);
or UO_1969 (O_1969,N_24713,N_24837);
or UO_1970 (O_1970,N_24582,N_24520);
xor UO_1971 (O_1971,N_24915,N_24542);
nor UO_1972 (O_1972,N_24992,N_24588);
or UO_1973 (O_1973,N_24807,N_24694);
and UO_1974 (O_1974,N_24728,N_24719);
xor UO_1975 (O_1975,N_24578,N_24525);
nand UO_1976 (O_1976,N_24577,N_24574);
xnor UO_1977 (O_1977,N_24861,N_24926);
and UO_1978 (O_1978,N_24579,N_24700);
and UO_1979 (O_1979,N_24779,N_24984);
xnor UO_1980 (O_1980,N_24713,N_24714);
nor UO_1981 (O_1981,N_24775,N_24532);
xor UO_1982 (O_1982,N_24880,N_24700);
xnor UO_1983 (O_1983,N_24708,N_24819);
and UO_1984 (O_1984,N_24880,N_24749);
and UO_1985 (O_1985,N_24529,N_24908);
nor UO_1986 (O_1986,N_24634,N_24915);
nor UO_1987 (O_1987,N_24968,N_24603);
nor UO_1988 (O_1988,N_24984,N_24652);
xnor UO_1989 (O_1989,N_24515,N_24612);
and UO_1990 (O_1990,N_24656,N_24761);
nor UO_1991 (O_1991,N_24552,N_24868);
nor UO_1992 (O_1992,N_24520,N_24622);
nand UO_1993 (O_1993,N_24958,N_24513);
nand UO_1994 (O_1994,N_24558,N_24874);
xnor UO_1995 (O_1995,N_24950,N_24689);
xnor UO_1996 (O_1996,N_24819,N_24701);
or UO_1997 (O_1997,N_24801,N_24880);
xnor UO_1998 (O_1998,N_24654,N_24892);
xnor UO_1999 (O_1999,N_24956,N_24593);
nand UO_2000 (O_2000,N_24988,N_24856);
or UO_2001 (O_2001,N_24805,N_24779);
nor UO_2002 (O_2002,N_24864,N_24584);
nand UO_2003 (O_2003,N_24967,N_24849);
or UO_2004 (O_2004,N_24665,N_24948);
or UO_2005 (O_2005,N_24925,N_24522);
and UO_2006 (O_2006,N_24550,N_24578);
and UO_2007 (O_2007,N_24584,N_24516);
nand UO_2008 (O_2008,N_24909,N_24696);
nand UO_2009 (O_2009,N_24592,N_24956);
or UO_2010 (O_2010,N_24834,N_24539);
xnor UO_2011 (O_2011,N_24799,N_24744);
xnor UO_2012 (O_2012,N_24593,N_24920);
and UO_2013 (O_2013,N_24766,N_24705);
and UO_2014 (O_2014,N_24696,N_24711);
nor UO_2015 (O_2015,N_24889,N_24644);
nor UO_2016 (O_2016,N_24867,N_24944);
nand UO_2017 (O_2017,N_24611,N_24664);
nor UO_2018 (O_2018,N_24538,N_24881);
nand UO_2019 (O_2019,N_24923,N_24952);
and UO_2020 (O_2020,N_24814,N_24816);
nor UO_2021 (O_2021,N_24549,N_24874);
xnor UO_2022 (O_2022,N_24990,N_24505);
xor UO_2023 (O_2023,N_24875,N_24874);
and UO_2024 (O_2024,N_24727,N_24514);
nand UO_2025 (O_2025,N_24792,N_24645);
and UO_2026 (O_2026,N_24652,N_24732);
or UO_2027 (O_2027,N_24912,N_24607);
and UO_2028 (O_2028,N_24597,N_24816);
xnor UO_2029 (O_2029,N_24864,N_24740);
xor UO_2030 (O_2030,N_24660,N_24904);
or UO_2031 (O_2031,N_24794,N_24791);
or UO_2032 (O_2032,N_24741,N_24892);
or UO_2033 (O_2033,N_24986,N_24709);
xor UO_2034 (O_2034,N_24841,N_24601);
or UO_2035 (O_2035,N_24957,N_24747);
or UO_2036 (O_2036,N_24871,N_24688);
nand UO_2037 (O_2037,N_24973,N_24780);
nor UO_2038 (O_2038,N_24724,N_24657);
xor UO_2039 (O_2039,N_24930,N_24754);
and UO_2040 (O_2040,N_24944,N_24862);
xor UO_2041 (O_2041,N_24507,N_24885);
nor UO_2042 (O_2042,N_24546,N_24838);
nor UO_2043 (O_2043,N_24541,N_24522);
and UO_2044 (O_2044,N_24576,N_24665);
nor UO_2045 (O_2045,N_24938,N_24957);
nand UO_2046 (O_2046,N_24815,N_24796);
or UO_2047 (O_2047,N_24644,N_24767);
or UO_2048 (O_2048,N_24601,N_24797);
xor UO_2049 (O_2049,N_24546,N_24643);
xor UO_2050 (O_2050,N_24681,N_24847);
nor UO_2051 (O_2051,N_24950,N_24974);
xor UO_2052 (O_2052,N_24843,N_24524);
and UO_2053 (O_2053,N_24886,N_24641);
nor UO_2054 (O_2054,N_24510,N_24674);
nor UO_2055 (O_2055,N_24670,N_24582);
or UO_2056 (O_2056,N_24924,N_24661);
xnor UO_2057 (O_2057,N_24521,N_24866);
or UO_2058 (O_2058,N_24855,N_24731);
or UO_2059 (O_2059,N_24644,N_24770);
and UO_2060 (O_2060,N_24587,N_24661);
nor UO_2061 (O_2061,N_24861,N_24804);
nor UO_2062 (O_2062,N_24851,N_24596);
nand UO_2063 (O_2063,N_24598,N_24658);
and UO_2064 (O_2064,N_24874,N_24570);
or UO_2065 (O_2065,N_24986,N_24868);
nor UO_2066 (O_2066,N_24869,N_24615);
or UO_2067 (O_2067,N_24559,N_24764);
xnor UO_2068 (O_2068,N_24959,N_24733);
xor UO_2069 (O_2069,N_24901,N_24826);
nor UO_2070 (O_2070,N_24935,N_24847);
or UO_2071 (O_2071,N_24624,N_24983);
xnor UO_2072 (O_2072,N_24721,N_24940);
nor UO_2073 (O_2073,N_24707,N_24992);
xor UO_2074 (O_2074,N_24684,N_24920);
nor UO_2075 (O_2075,N_24994,N_24972);
or UO_2076 (O_2076,N_24996,N_24932);
or UO_2077 (O_2077,N_24611,N_24692);
or UO_2078 (O_2078,N_24595,N_24890);
nand UO_2079 (O_2079,N_24872,N_24842);
and UO_2080 (O_2080,N_24933,N_24876);
and UO_2081 (O_2081,N_24801,N_24797);
xor UO_2082 (O_2082,N_24573,N_24820);
or UO_2083 (O_2083,N_24527,N_24942);
and UO_2084 (O_2084,N_24880,N_24943);
nand UO_2085 (O_2085,N_24837,N_24827);
and UO_2086 (O_2086,N_24785,N_24764);
nand UO_2087 (O_2087,N_24529,N_24584);
or UO_2088 (O_2088,N_24781,N_24689);
and UO_2089 (O_2089,N_24731,N_24842);
nand UO_2090 (O_2090,N_24731,N_24806);
nor UO_2091 (O_2091,N_24818,N_24521);
or UO_2092 (O_2092,N_24986,N_24544);
or UO_2093 (O_2093,N_24979,N_24661);
and UO_2094 (O_2094,N_24854,N_24709);
and UO_2095 (O_2095,N_24917,N_24927);
xnor UO_2096 (O_2096,N_24918,N_24994);
or UO_2097 (O_2097,N_24882,N_24547);
or UO_2098 (O_2098,N_24957,N_24946);
nor UO_2099 (O_2099,N_24775,N_24990);
nand UO_2100 (O_2100,N_24765,N_24532);
nand UO_2101 (O_2101,N_24803,N_24676);
xor UO_2102 (O_2102,N_24545,N_24942);
or UO_2103 (O_2103,N_24881,N_24792);
or UO_2104 (O_2104,N_24974,N_24672);
nand UO_2105 (O_2105,N_24632,N_24844);
and UO_2106 (O_2106,N_24727,N_24781);
xnor UO_2107 (O_2107,N_24800,N_24765);
or UO_2108 (O_2108,N_24929,N_24658);
xor UO_2109 (O_2109,N_24777,N_24605);
nor UO_2110 (O_2110,N_24728,N_24641);
or UO_2111 (O_2111,N_24805,N_24509);
and UO_2112 (O_2112,N_24770,N_24748);
or UO_2113 (O_2113,N_24578,N_24910);
or UO_2114 (O_2114,N_24558,N_24585);
nand UO_2115 (O_2115,N_24966,N_24541);
nor UO_2116 (O_2116,N_24772,N_24572);
or UO_2117 (O_2117,N_24698,N_24888);
xor UO_2118 (O_2118,N_24626,N_24644);
and UO_2119 (O_2119,N_24567,N_24606);
xor UO_2120 (O_2120,N_24838,N_24670);
xor UO_2121 (O_2121,N_24847,N_24881);
and UO_2122 (O_2122,N_24911,N_24994);
nand UO_2123 (O_2123,N_24745,N_24747);
and UO_2124 (O_2124,N_24899,N_24552);
and UO_2125 (O_2125,N_24676,N_24891);
nor UO_2126 (O_2126,N_24630,N_24618);
nand UO_2127 (O_2127,N_24648,N_24749);
and UO_2128 (O_2128,N_24819,N_24967);
nand UO_2129 (O_2129,N_24673,N_24687);
or UO_2130 (O_2130,N_24788,N_24778);
nor UO_2131 (O_2131,N_24609,N_24909);
xnor UO_2132 (O_2132,N_24843,N_24998);
xor UO_2133 (O_2133,N_24934,N_24952);
nor UO_2134 (O_2134,N_24789,N_24985);
or UO_2135 (O_2135,N_24620,N_24687);
or UO_2136 (O_2136,N_24698,N_24756);
or UO_2137 (O_2137,N_24687,N_24874);
nand UO_2138 (O_2138,N_24912,N_24871);
and UO_2139 (O_2139,N_24533,N_24987);
nor UO_2140 (O_2140,N_24970,N_24847);
nor UO_2141 (O_2141,N_24926,N_24619);
or UO_2142 (O_2142,N_24688,N_24836);
or UO_2143 (O_2143,N_24614,N_24639);
and UO_2144 (O_2144,N_24982,N_24661);
and UO_2145 (O_2145,N_24563,N_24679);
and UO_2146 (O_2146,N_24719,N_24643);
xor UO_2147 (O_2147,N_24868,N_24565);
and UO_2148 (O_2148,N_24615,N_24968);
nand UO_2149 (O_2149,N_24819,N_24527);
or UO_2150 (O_2150,N_24981,N_24541);
xnor UO_2151 (O_2151,N_24907,N_24739);
nand UO_2152 (O_2152,N_24755,N_24948);
nand UO_2153 (O_2153,N_24808,N_24973);
nand UO_2154 (O_2154,N_24995,N_24526);
nor UO_2155 (O_2155,N_24862,N_24984);
and UO_2156 (O_2156,N_24670,N_24619);
xor UO_2157 (O_2157,N_24772,N_24504);
or UO_2158 (O_2158,N_24572,N_24509);
and UO_2159 (O_2159,N_24567,N_24506);
or UO_2160 (O_2160,N_24976,N_24996);
and UO_2161 (O_2161,N_24593,N_24773);
and UO_2162 (O_2162,N_24687,N_24548);
or UO_2163 (O_2163,N_24960,N_24918);
nand UO_2164 (O_2164,N_24935,N_24983);
nor UO_2165 (O_2165,N_24564,N_24714);
or UO_2166 (O_2166,N_24982,N_24611);
xor UO_2167 (O_2167,N_24538,N_24531);
nor UO_2168 (O_2168,N_24759,N_24839);
nor UO_2169 (O_2169,N_24554,N_24533);
xnor UO_2170 (O_2170,N_24986,N_24731);
nand UO_2171 (O_2171,N_24924,N_24699);
nor UO_2172 (O_2172,N_24909,N_24997);
and UO_2173 (O_2173,N_24763,N_24841);
nor UO_2174 (O_2174,N_24874,N_24653);
nand UO_2175 (O_2175,N_24645,N_24669);
and UO_2176 (O_2176,N_24937,N_24591);
xor UO_2177 (O_2177,N_24594,N_24657);
nand UO_2178 (O_2178,N_24543,N_24711);
nor UO_2179 (O_2179,N_24667,N_24915);
or UO_2180 (O_2180,N_24715,N_24753);
nor UO_2181 (O_2181,N_24531,N_24759);
and UO_2182 (O_2182,N_24926,N_24518);
nor UO_2183 (O_2183,N_24751,N_24789);
xnor UO_2184 (O_2184,N_24931,N_24952);
and UO_2185 (O_2185,N_24710,N_24724);
and UO_2186 (O_2186,N_24925,N_24893);
nand UO_2187 (O_2187,N_24567,N_24786);
nand UO_2188 (O_2188,N_24537,N_24546);
nor UO_2189 (O_2189,N_24674,N_24564);
and UO_2190 (O_2190,N_24747,N_24687);
xnor UO_2191 (O_2191,N_24997,N_24999);
nor UO_2192 (O_2192,N_24941,N_24588);
nand UO_2193 (O_2193,N_24667,N_24665);
xnor UO_2194 (O_2194,N_24571,N_24551);
xnor UO_2195 (O_2195,N_24975,N_24744);
nand UO_2196 (O_2196,N_24568,N_24957);
nand UO_2197 (O_2197,N_24744,N_24665);
and UO_2198 (O_2198,N_24880,N_24771);
nor UO_2199 (O_2199,N_24716,N_24645);
xor UO_2200 (O_2200,N_24597,N_24979);
nor UO_2201 (O_2201,N_24903,N_24643);
xor UO_2202 (O_2202,N_24756,N_24808);
xnor UO_2203 (O_2203,N_24986,N_24645);
nor UO_2204 (O_2204,N_24511,N_24646);
or UO_2205 (O_2205,N_24570,N_24522);
and UO_2206 (O_2206,N_24860,N_24707);
and UO_2207 (O_2207,N_24560,N_24669);
nor UO_2208 (O_2208,N_24899,N_24674);
and UO_2209 (O_2209,N_24574,N_24643);
or UO_2210 (O_2210,N_24771,N_24949);
xor UO_2211 (O_2211,N_24972,N_24744);
or UO_2212 (O_2212,N_24900,N_24707);
and UO_2213 (O_2213,N_24782,N_24754);
xor UO_2214 (O_2214,N_24679,N_24717);
nand UO_2215 (O_2215,N_24881,N_24642);
xnor UO_2216 (O_2216,N_24918,N_24789);
or UO_2217 (O_2217,N_24602,N_24591);
and UO_2218 (O_2218,N_24727,N_24730);
nand UO_2219 (O_2219,N_24510,N_24827);
nor UO_2220 (O_2220,N_24753,N_24932);
xor UO_2221 (O_2221,N_24532,N_24755);
nor UO_2222 (O_2222,N_24517,N_24831);
xnor UO_2223 (O_2223,N_24541,N_24753);
nor UO_2224 (O_2224,N_24693,N_24942);
nand UO_2225 (O_2225,N_24865,N_24657);
xnor UO_2226 (O_2226,N_24833,N_24513);
or UO_2227 (O_2227,N_24530,N_24718);
nand UO_2228 (O_2228,N_24886,N_24873);
and UO_2229 (O_2229,N_24517,N_24922);
xor UO_2230 (O_2230,N_24547,N_24590);
nor UO_2231 (O_2231,N_24690,N_24602);
nand UO_2232 (O_2232,N_24583,N_24545);
and UO_2233 (O_2233,N_24844,N_24587);
xor UO_2234 (O_2234,N_24901,N_24622);
nor UO_2235 (O_2235,N_24606,N_24882);
nand UO_2236 (O_2236,N_24985,N_24531);
nand UO_2237 (O_2237,N_24546,N_24649);
or UO_2238 (O_2238,N_24554,N_24503);
and UO_2239 (O_2239,N_24723,N_24570);
or UO_2240 (O_2240,N_24900,N_24682);
nor UO_2241 (O_2241,N_24562,N_24525);
nand UO_2242 (O_2242,N_24646,N_24806);
nand UO_2243 (O_2243,N_24570,N_24659);
nand UO_2244 (O_2244,N_24857,N_24872);
and UO_2245 (O_2245,N_24678,N_24648);
nor UO_2246 (O_2246,N_24549,N_24795);
and UO_2247 (O_2247,N_24912,N_24650);
nor UO_2248 (O_2248,N_24625,N_24608);
nand UO_2249 (O_2249,N_24635,N_24998);
xor UO_2250 (O_2250,N_24997,N_24524);
nor UO_2251 (O_2251,N_24669,N_24978);
and UO_2252 (O_2252,N_24856,N_24795);
or UO_2253 (O_2253,N_24826,N_24939);
nand UO_2254 (O_2254,N_24995,N_24994);
nand UO_2255 (O_2255,N_24708,N_24875);
xor UO_2256 (O_2256,N_24811,N_24964);
or UO_2257 (O_2257,N_24592,N_24826);
and UO_2258 (O_2258,N_24871,N_24968);
and UO_2259 (O_2259,N_24722,N_24555);
or UO_2260 (O_2260,N_24545,N_24521);
nor UO_2261 (O_2261,N_24846,N_24947);
xor UO_2262 (O_2262,N_24901,N_24917);
or UO_2263 (O_2263,N_24540,N_24716);
xor UO_2264 (O_2264,N_24616,N_24787);
xor UO_2265 (O_2265,N_24845,N_24751);
nand UO_2266 (O_2266,N_24651,N_24796);
nor UO_2267 (O_2267,N_24717,N_24806);
or UO_2268 (O_2268,N_24789,N_24664);
nor UO_2269 (O_2269,N_24998,N_24671);
and UO_2270 (O_2270,N_24666,N_24685);
and UO_2271 (O_2271,N_24581,N_24914);
or UO_2272 (O_2272,N_24869,N_24986);
and UO_2273 (O_2273,N_24856,N_24929);
nand UO_2274 (O_2274,N_24859,N_24957);
nor UO_2275 (O_2275,N_24967,N_24984);
nand UO_2276 (O_2276,N_24575,N_24668);
or UO_2277 (O_2277,N_24696,N_24851);
or UO_2278 (O_2278,N_24640,N_24858);
nand UO_2279 (O_2279,N_24861,N_24719);
or UO_2280 (O_2280,N_24960,N_24589);
and UO_2281 (O_2281,N_24872,N_24802);
nand UO_2282 (O_2282,N_24795,N_24554);
or UO_2283 (O_2283,N_24806,N_24720);
nand UO_2284 (O_2284,N_24938,N_24711);
or UO_2285 (O_2285,N_24665,N_24643);
and UO_2286 (O_2286,N_24622,N_24718);
nor UO_2287 (O_2287,N_24574,N_24796);
nor UO_2288 (O_2288,N_24713,N_24538);
xor UO_2289 (O_2289,N_24707,N_24616);
and UO_2290 (O_2290,N_24993,N_24525);
xor UO_2291 (O_2291,N_24676,N_24572);
nor UO_2292 (O_2292,N_24604,N_24821);
nand UO_2293 (O_2293,N_24517,N_24923);
xor UO_2294 (O_2294,N_24732,N_24752);
or UO_2295 (O_2295,N_24693,N_24649);
nand UO_2296 (O_2296,N_24604,N_24678);
or UO_2297 (O_2297,N_24923,N_24926);
nor UO_2298 (O_2298,N_24584,N_24773);
nor UO_2299 (O_2299,N_24684,N_24978);
nor UO_2300 (O_2300,N_24529,N_24690);
nand UO_2301 (O_2301,N_24836,N_24874);
and UO_2302 (O_2302,N_24589,N_24514);
nand UO_2303 (O_2303,N_24780,N_24503);
nand UO_2304 (O_2304,N_24956,N_24942);
nor UO_2305 (O_2305,N_24514,N_24924);
nand UO_2306 (O_2306,N_24805,N_24965);
xnor UO_2307 (O_2307,N_24606,N_24946);
or UO_2308 (O_2308,N_24531,N_24693);
and UO_2309 (O_2309,N_24861,N_24644);
nand UO_2310 (O_2310,N_24777,N_24739);
nand UO_2311 (O_2311,N_24753,N_24911);
nor UO_2312 (O_2312,N_24588,N_24721);
and UO_2313 (O_2313,N_24611,N_24742);
xnor UO_2314 (O_2314,N_24840,N_24989);
and UO_2315 (O_2315,N_24807,N_24927);
and UO_2316 (O_2316,N_24821,N_24855);
or UO_2317 (O_2317,N_24631,N_24640);
nor UO_2318 (O_2318,N_24744,N_24776);
nor UO_2319 (O_2319,N_24961,N_24801);
and UO_2320 (O_2320,N_24820,N_24693);
xnor UO_2321 (O_2321,N_24599,N_24655);
xnor UO_2322 (O_2322,N_24681,N_24959);
xor UO_2323 (O_2323,N_24945,N_24696);
nor UO_2324 (O_2324,N_24834,N_24812);
and UO_2325 (O_2325,N_24576,N_24797);
xnor UO_2326 (O_2326,N_24722,N_24783);
and UO_2327 (O_2327,N_24757,N_24961);
nand UO_2328 (O_2328,N_24658,N_24554);
xor UO_2329 (O_2329,N_24538,N_24956);
xor UO_2330 (O_2330,N_24738,N_24587);
xor UO_2331 (O_2331,N_24757,N_24653);
xor UO_2332 (O_2332,N_24670,N_24599);
and UO_2333 (O_2333,N_24502,N_24582);
nor UO_2334 (O_2334,N_24534,N_24717);
nand UO_2335 (O_2335,N_24549,N_24747);
xor UO_2336 (O_2336,N_24526,N_24849);
and UO_2337 (O_2337,N_24566,N_24759);
xnor UO_2338 (O_2338,N_24628,N_24850);
and UO_2339 (O_2339,N_24873,N_24861);
or UO_2340 (O_2340,N_24898,N_24836);
xnor UO_2341 (O_2341,N_24806,N_24696);
nand UO_2342 (O_2342,N_24750,N_24994);
xor UO_2343 (O_2343,N_24773,N_24546);
nor UO_2344 (O_2344,N_24841,N_24634);
nor UO_2345 (O_2345,N_24700,N_24940);
nor UO_2346 (O_2346,N_24649,N_24890);
nand UO_2347 (O_2347,N_24614,N_24590);
nor UO_2348 (O_2348,N_24548,N_24866);
xor UO_2349 (O_2349,N_24697,N_24620);
nand UO_2350 (O_2350,N_24533,N_24665);
and UO_2351 (O_2351,N_24620,N_24845);
nand UO_2352 (O_2352,N_24595,N_24926);
nand UO_2353 (O_2353,N_24842,N_24501);
nand UO_2354 (O_2354,N_24594,N_24971);
xnor UO_2355 (O_2355,N_24526,N_24609);
nand UO_2356 (O_2356,N_24761,N_24892);
xnor UO_2357 (O_2357,N_24955,N_24628);
nand UO_2358 (O_2358,N_24687,N_24931);
xor UO_2359 (O_2359,N_24658,N_24939);
xor UO_2360 (O_2360,N_24909,N_24726);
nand UO_2361 (O_2361,N_24997,N_24893);
and UO_2362 (O_2362,N_24671,N_24907);
nand UO_2363 (O_2363,N_24664,N_24627);
and UO_2364 (O_2364,N_24679,N_24700);
nand UO_2365 (O_2365,N_24666,N_24912);
or UO_2366 (O_2366,N_24781,N_24541);
nand UO_2367 (O_2367,N_24994,N_24503);
xnor UO_2368 (O_2368,N_24710,N_24743);
nand UO_2369 (O_2369,N_24954,N_24614);
or UO_2370 (O_2370,N_24819,N_24566);
or UO_2371 (O_2371,N_24923,N_24704);
nor UO_2372 (O_2372,N_24613,N_24573);
xnor UO_2373 (O_2373,N_24953,N_24717);
and UO_2374 (O_2374,N_24585,N_24950);
nor UO_2375 (O_2375,N_24673,N_24722);
xor UO_2376 (O_2376,N_24953,N_24583);
or UO_2377 (O_2377,N_24720,N_24809);
xnor UO_2378 (O_2378,N_24582,N_24911);
nand UO_2379 (O_2379,N_24767,N_24987);
or UO_2380 (O_2380,N_24571,N_24509);
or UO_2381 (O_2381,N_24695,N_24699);
nor UO_2382 (O_2382,N_24601,N_24794);
nor UO_2383 (O_2383,N_24802,N_24894);
or UO_2384 (O_2384,N_24923,N_24746);
nor UO_2385 (O_2385,N_24986,N_24534);
nor UO_2386 (O_2386,N_24900,N_24934);
nand UO_2387 (O_2387,N_24963,N_24597);
nor UO_2388 (O_2388,N_24620,N_24705);
and UO_2389 (O_2389,N_24729,N_24699);
nor UO_2390 (O_2390,N_24733,N_24878);
nand UO_2391 (O_2391,N_24889,N_24919);
and UO_2392 (O_2392,N_24740,N_24919);
and UO_2393 (O_2393,N_24941,N_24914);
nor UO_2394 (O_2394,N_24959,N_24868);
nand UO_2395 (O_2395,N_24577,N_24775);
xnor UO_2396 (O_2396,N_24833,N_24636);
and UO_2397 (O_2397,N_24857,N_24720);
xor UO_2398 (O_2398,N_24931,N_24860);
nor UO_2399 (O_2399,N_24760,N_24888);
xnor UO_2400 (O_2400,N_24845,N_24565);
nor UO_2401 (O_2401,N_24687,N_24520);
nand UO_2402 (O_2402,N_24543,N_24637);
nor UO_2403 (O_2403,N_24612,N_24756);
and UO_2404 (O_2404,N_24966,N_24910);
nand UO_2405 (O_2405,N_24672,N_24893);
and UO_2406 (O_2406,N_24980,N_24546);
or UO_2407 (O_2407,N_24926,N_24568);
nor UO_2408 (O_2408,N_24924,N_24964);
nor UO_2409 (O_2409,N_24775,N_24743);
nor UO_2410 (O_2410,N_24628,N_24880);
nor UO_2411 (O_2411,N_24567,N_24634);
or UO_2412 (O_2412,N_24776,N_24928);
or UO_2413 (O_2413,N_24783,N_24805);
xor UO_2414 (O_2414,N_24989,N_24548);
nand UO_2415 (O_2415,N_24813,N_24770);
xor UO_2416 (O_2416,N_24889,N_24842);
nor UO_2417 (O_2417,N_24675,N_24511);
nor UO_2418 (O_2418,N_24695,N_24888);
nand UO_2419 (O_2419,N_24825,N_24702);
or UO_2420 (O_2420,N_24825,N_24596);
xnor UO_2421 (O_2421,N_24600,N_24988);
nand UO_2422 (O_2422,N_24673,N_24741);
nand UO_2423 (O_2423,N_24909,N_24677);
xor UO_2424 (O_2424,N_24520,N_24863);
and UO_2425 (O_2425,N_24936,N_24600);
and UO_2426 (O_2426,N_24583,N_24938);
or UO_2427 (O_2427,N_24800,N_24593);
xnor UO_2428 (O_2428,N_24929,N_24790);
xnor UO_2429 (O_2429,N_24555,N_24763);
nor UO_2430 (O_2430,N_24562,N_24643);
or UO_2431 (O_2431,N_24789,N_24820);
xor UO_2432 (O_2432,N_24751,N_24603);
nor UO_2433 (O_2433,N_24919,N_24604);
and UO_2434 (O_2434,N_24860,N_24641);
or UO_2435 (O_2435,N_24937,N_24872);
nor UO_2436 (O_2436,N_24760,N_24823);
nor UO_2437 (O_2437,N_24747,N_24706);
or UO_2438 (O_2438,N_24659,N_24918);
nand UO_2439 (O_2439,N_24681,N_24918);
and UO_2440 (O_2440,N_24657,N_24799);
xor UO_2441 (O_2441,N_24849,N_24639);
or UO_2442 (O_2442,N_24790,N_24538);
nand UO_2443 (O_2443,N_24534,N_24631);
nand UO_2444 (O_2444,N_24953,N_24789);
nand UO_2445 (O_2445,N_24708,N_24655);
nand UO_2446 (O_2446,N_24900,N_24894);
nand UO_2447 (O_2447,N_24592,N_24839);
nor UO_2448 (O_2448,N_24966,N_24804);
nand UO_2449 (O_2449,N_24677,N_24765);
and UO_2450 (O_2450,N_24826,N_24762);
xnor UO_2451 (O_2451,N_24902,N_24679);
nand UO_2452 (O_2452,N_24941,N_24841);
or UO_2453 (O_2453,N_24944,N_24905);
nor UO_2454 (O_2454,N_24735,N_24983);
and UO_2455 (O_2455,N_24515,N_24848);
nor UO_2456 (O_2456,N_24795,N_24761);
nor UO_2457 (O_2457,N_24947,N_24611);
nand UO_2458 (O_2458,N_24882,N_24596);
nor UO_2459 (O_2459,N_24602,N_24635);
or UO_2460 (O_2460,N_24833,N_24780);
nor UO_2461 (O_2461,N_24807,N_24771);
nand UO_2462 (O_2462,N_24870,N_24995);
or UO_2463 (O_2463,N_24629,N_24685);
and UO_2464 (O_2464,N_24740,N_24675);
and UO_2465 (O_2465,N_24802,N_24878);
and UO_2466 (O_2466,N_24660,N_24952);
nor UO_2467 (O_2467,N_24771,N_24745);
or UO_2468 (O_2468,N_24933,N_24511);
or UO_2469 (O_2469,N_24614,N_24680);
nand UO_2470 (O_2470,N_24942,N_24978);
and UO_2471 (O_2471,N_24656,N_24631);
or UO_2472 (O_2472,N_24724,N_24789);
xor UO_2473 (O_2473,N_24847,N_24856);
or UO_2474 (O_2474,N_24735,N_24724);
and UO_2475 (O_2475,N_24562,N_24564);
and UO_2476 (O_2476,N_24835,N_24655);
nor UO_2477 (O_2477,N_24981,N_24950);
nor UO_2478 (O_2478,N_24772,N_24964);
nand UO_2479 (O_2479,N_24552,N_24631);
xor UO_2480 (O_2480,N_24897,N_24914);
or UO_2481 (O_2481,N_24651,N_24733);
xor UO_2482 (O_2482,N_24571,N_24524);
xnor UO_2483 (O_2483,N_24519,N_24640);
nand UO_2484 (O_2484,N_24824,N_24990);
or UO_2485 (O_2485,N_24730,N_24772);
or UO_2486 (O_2486,N_24513,N_24573);
and UO_2487 (O_2487,N_24779,N_24520);
and UO_2488 (O_2488,N_24882,N_24854);
nand UO_2489 (O_2489,N_24765,N_24630);
and UO_2490 (O_2490,N_24969,N_24581);
xor UO_2491 (O_2491,N_24619,N_24796);
nor UO_2492 (O_2492,N_24581,N_24521);
nor UO_2493 (O_2493,N_24694,N_24856);
nand UO_2494 (O_2494,N_24561,N_24866);
xnor UO_2495 (O_2495,N_24665,N_24720);
or UO_2496 (O_2496,N_24833,N_24524);
nor UO_2497 (O_2497,N_24880,N_24650);
or UO_2498 (O_2498,N_24608,N_24572);
and UO_2499 (O_2499,N_24712,N_24946);
or UO_2500 (O_2500,N_24807,N_24992);
nand UO_2501 (O_2501,N_24784,N_24701);
nand UO_2502 (O_2502,N_24535,N_24894);
nand UO_2503 (O_2503,N_24966,N_24973);
and UO_2504 (O_2504,N_24756,N_24791);
nand UO_2505 (O_2505,N_24932,N_24874);
or UO_2506 (O_2506,N_24752,N_24607);
or UO_2507 (O_2507,N_24723,N_24774);
and UO_2508 (O_2508,N_24833,N_24985);
nand UO_2509 (O_2509,N_24917,N_24871);
xnor UO_2510 (O_2510,N_24864,N_24959);
and UO_2511 (O_2511,N_24746,N_24724);
and UO_2512 (O_2512,N_24671,N_24900);
or UO_2513 (O_2513,N_24920,N_24660);
xor UO_2514 (O_2514,N_24692,N_24552);
nor UO_2515 (O_2515,N_24783,N_24941);
nand UO_2516 (O_2516,N_24744,N_24535);
xnor UO_2517 (O_2517,N_24702,N_24628);
nand UO_2518 (O_2518,N_24877,N_24908);
and UO_2519 (O_2519,N_24713,N_24738);
nor UO_2520 (O_2520,N_24968,N_24921);
or UO_2521 (O_2521,N_24990,N_24540);
xor UO_2522 (O_2522,N_24866,N_24940);
or UO_2523 (O_2523,N_24902,N_24500);
or UO_2524 (O_2524,N_24852,N_24596);
xnor UO_2525 (O_2525,N_24636,N_24646);
and UO_2526 (O_2526,N_24775,N_24564);
nand UO_2527 (O_2527,N_24685,N_24870);
or UO_2528 (O_2528,N_24912,N_24637);
nand UO_2529 (O_2529,N_24534,N_24886);
nor UO_2530 (O_2530,N_24595,N_24833);
or UO_2531 (O_2531,N_24592,N_24731);
and UO_2532 (O_2532,N_24590,N_24681);
or UO_2533 (O_2533,N_24646,N_24569);
xor UO_2534 (O_2534,N_24754,N_24547);
xor UO_2535 (O_2535,N_24526,N_24961);
nand UO_2536 (O_2536,N_24808,N_24908);
xor UO_2537 (O_2537,N_24967,N_24689);
and UO_2538 (O_2538,N_24923,N_24693);
nand UO_2539 (O_2539,N_24630,N_24957);
or UO_2540 (O_2540,N_24635,N_24865);
nor UO_2541 (O_2541,N_24701,N_24520);
and UO_2542 (O_2542,N_24617,N_24828);
and UO_2543 (O_2543,N_24973,N_24814);
and UO_2544 (O_2544,N_24954,N_24970);
and UO_2545 (O_2545,N_24930,N_24866);
or UO_2546 (O_2546,N_24642,N_24544);
or UO_2547 (O_2547,N_24775,N_24696);
or UO_2548 (O_2548,N_24685,N_24582);
nand UO_2549 (O_2549,N_24865,N_24682);
xnor UO_2550 (O_2550,N_24812,N_24696);
or UO_2551 (O_2551,N_24758,N_24820);
xor UO_2552 (O_2552,N_24710,N_24902);
nor UO_2553 (O_2553,N_24897,N_24662);
xor UO_2554 (O_2554,N_24579,N_24546);
nor UO_2555 (O_2555,N_24652,N_24877);
nor UO_2556 (O_2556,N_24524,N_24557);
nor UO_2557 (O_2557,N_24827,N_24905);
or UO_2558 (O_2558,N_24574,N_24746);
and UO_2559 (O_2559,N_24630,N_24635);
nand UO_2560 (O_2560,N_24901,N_24916);
and UO_2561 (O_2561,N_24798,N_24942);
nor UO_2562 (O_2562,N_24889,N_24514);
nand UO_2563 (O_2563,N_24620,N_24689);
nor UO_2564 (O_2564,N_24805,N_24612);
and UO_2565 (O_2565,N_24962,N_24658);
nor UO_2566 (O_2566,N_24798,N_24519);
and UO_2567 (O_2567,N_24528,N_24717);
xnor UO_2568 (O_2568,N_24675,N_24819);
and UO_2569 (O_2569,N_24969,N_24697);
or UO_2570 (O_2570,N_24645,N_24749);
and UO_2571 (O_2571,N_24909,N_24565);
nand UO_2572 (O_2572,N_24699,N_24936);
nand UO_2573 (O_2573,N_24810,N_24541);
and UO_2574 (O_2574,N_24998,N_24744);
and UO_2575 (O_2575,N_24688,N_24963);
nor UO_2576 (O_2576,N_24548,N_24869);
nor UO_2577 (O_2577,N_24596,N_24671);
or UO_2578 (O_2578,N_24804,N_24812);
nand UO_2579 (O_2579,N_24709,N_24815);
xnor UO_2580 (O_2580,N_24774,N_24638);
xor UO_2581 (O_2581,N_24654,N_24994);
xnor UO_2582 (O_2582,N_24863,N_24630);
nor UO_2583 (O_2583,N_24902,N_24642);
nand UO_2584 (O_2584,N_24741,N_24717);
nand UO_2585 (O_2585,N_24644,N_24833);
xor UO_2586 (O_2586,N_24872,N_24818);
xor UO_2587 (O_2587,N_24609,N_24686);
and UO_2588 (O_2588,N_24671,N_24768);
nor UO_2589 (O_2589,N_24591,N_24758);
or UO_2590 (O_2590,N_24931,N_24674);
nor UO_2591 (O_2591,N_24755,N_24699);
and UO_2592 (O_2592,N_24640,N_24753);
or UO_2593 (O_2593,N_24621,N_24698);
nor UO_2594 (O_2594,N_24509,N_24783);
or UO_2595 (O_2595,N_24531,N_24578);
xor UO_2596 (O_2596,N_24924,N_24894);
nand UO_2597 (O_2597,N_24827,N_24836);
nand UO_2598 (O_2598,N_24552,N_24525);
and UO_2599 (O_2599,N_24709,N_24963);
and UO_2600 (O_2600,N_24962,N_24774);
xnor UO_2601 (O_2601,N_24861,N_24575);
and UO_2602 (O_2602,N_24722,N_24750);
nor UO_2603 (O_2603,N_24887,N_24724);
xor UO_2604 (O_2604,N_24966,N_24717);
or UO_2605 (O_2605,N_24603,N_24647);
xor UO_2606 (O_2606,N_24929,N_24653);
nor UO_2607 (O_2607,N_24664,N_24806);
or UO_2608 (O_2608,N_24897,N_24699);
or UO_2609 (O_2609,N_24736,N_24910);
nor UO_2610 (O_2610,N_24608,N_24993);
or UO_2611 (O_2611,N_24625,N_24618);
nor UO_2612 (O_2612,N_24660,N_24803);
and UO_2613 (O_2613,N_24587,N_24554);
nand UO_2614 (O_2614,N_24855,N_24574);
nand UO_2615 (O_2615,N_24541,N_24712);
nor UO_2616 (O_2616,N_24527,N_24534);
or UO_2617 (O_2617,N_24707,N_24976);
nor UO_2618 (O_2618,N_24797,N_24802);
nor UO_2619 (O_2619,N_24859,N_24544);
and UO_2620 (O_2620,N_24768,N_24697);
and UO_2621 (O_2621,N_24829,N_24589);
nand UO_2622 (O_2622,N_24587,N_24837);
nand UO_2623 (O_2623,N_24910,N_24635);
nor UO_2624 (O_2624,N_24936,N_24649);
and UO_2625 (O_2625,N_24941,N_24695);
and UO_2626 (O_2626,N_24600,N_24802);
nand UO_2627 (O_2627,N_24520,N_24715);
and UO_2628 (O_2628,N_24943,N_24595);
or UO_2629 (O_2629,N_24689,N_24955);
xor UO_2630 (O_2630,N_24981,N_24989);
nand UO_2631 (O_2631,N_24999,N_24523);
and UO_2632 (O_2632,N_24592,N_24654);
and UO_2633 (O_2633,N_24960,N_24541);
nor UO_2634 (O_2634,N_24676,N_24518);
xor UO_2635 (O_2635,N_24905,N_24505);
nor UO_2636 (O_2636,N_24917,N_24935);
nand UO_2637 (O_2637,N_24839,N_24624);
nand UO_2638 (O_2638,N_24557,N_24875);
or UO_2639 (O_2639,N_24541,N_24614);
xnor UO_2640 (O_2640,N_24939,N_24968);
xnor UO_2641 (O_2641,N_24805,N_24562);
nor UO_2642 (O_2642,N_24663,N_24751);
or UO_2643 (O_2643,N_24872,N_24607);
and UO_2644 (O_2644,N_24650,N_24562);
nand UO_2645 (O_2645,N_24864,N_24628);
nor UO_2646 (O_2646,N_24758,N_24789);
and UO_2647 (O_2647,N_24500,N_24679);
nand UO_2648 (O_2648,N_24941,N_24915);
xor UO_2649 (O_2649,N_24748,N_24956);
nor UO_2650 (O_2650,N_24506,N_24711);
and UO_2651 (O_2651,N_24652,N_24617);
nor UO_2652 (O_2652,N_24508,N_24761);
or UO_2653 (O_2653,N_24936,N_24919);
or UO_2654 (O_2654,N_24572,N_24592);
xor UO_2655 (O_2655,N_24806,N_24726);
xnor UO_2656 (O_2656,N_24833,N_24685);
or UO_2657 (O_2657,N_24509,N_24892);
or UO_2658 (O_2658,N_24614,N_24528);
xor UO_2659 (O_2659,N_24976,N_24872);
xor UO_2660 (O_2660,N_24958,N_24919);
and UO_2661 (O_2661,N_24919,N_24820);
nand UO_2662 (O_2662,N_24989,N_24557);
and UO_2663 (O_2663,N_24599,N_24799);
or UO_2664 (O_2664,N_24911,N_24893);
xor UO_2665 (O_2665,N_24546,N_24825);
nand UO_2666 (O_2666,N_24673,N_24828);
and UO_2667 (O_2667,N_24930,N_24948);
or UO_2668 (O_2668,N_24602,N_24799);
nor UO_2669 (O_2669,N_24916,N_24999);
nand UO_2670 (O_2670,N_24695,N_24972);
and UO_2671 (O_2671,N_24689,N_24678);
or UO_2672 (O_2672,N_24564,N_24885);
xor UO_2673 (O_2673,N_24684,N_24788);
or UO_2674 (O_2674,N_24506,N_24635);
nor UO_2675 (O_2675,N_24667,N_24850);
nor UO_2676 (O_2676,N_24525,N_24799);
nor UO_2677 (O_2677,N_24964,N_24714);
nand UO_2678 (O_2678,N_24841,N_24577);
nor UO_2679 (O_2679,N_24636,N_24604);
nor UO_2680 (O_2680,N_24760,N_24657);
and UO_2681 (O_2681,N_24641,N_24823);
nor UO_2682 (O_2682,N_24997,N_24849);
nor UO_2683 (O_2683,N_24992,N_24697);
and UO_2684 (O_2684,N_24681,N_24806);
and UO_2685 (O_2685,N_24968,N_24699);
xnor UO_2686 (O_2686,N_24935,N_24709);
and UO_2687 (O_2687,N_24561,N_24814);
nand UO_2688 (O_2688,N_24598,N_24806);
nand UO_2689 (O_2689,N_24571,N_24882);
nand UO_2690 (O_2690,N_24625,N_24910);
xor UO_2691 (O_2691,N_24839,N_24860);
or UO_2692 (O_2692,N_24974,N_24706);
and UO_2693 (O_2693,N_24818,N_24790);
xor UO_2694 (O_2694,N_24703,N_24914);
nand UO_2695 (O_2695,N_24509,N_24880);
nor UO_2696 (O_2696,N_24726,N_24668);
xor UO_2697 (O_2697,N_24981,N_24633);
and UO_2698 (O_2698,N_24842,N_24907);
xor UO_2699 (O_2699,N_24614,N_24563);
xnor UO_2700 (O_2700,N_24567,N_24964);
nand UO_2701 (O_2701,N_24631,N_24522);
nand UO_2702 (O_2702,N_24962,N_24530);
xnor UO_2703 (O_2703,N_24567,N_24503);
or UO_2704 (O_2704,N_24553,N_24696);
nand UO_2705 (O_2705,N_24805,N_24665);
xor UO_2706 (O_2706,N_24993,N_24686);
or UO_2707 (O_2707,N_24939,N_24707);
or UO_2708 (O_2708,N_24905,N_24594);
nor UO_2709 (O_2709,N_24759,N_24831);
nor UO_2710 (O_2710,N_24623,N_24618);
xor UO_2711 (O_2711,N_24692,N_24639);
and UO_2712 (O_2712,N_24547,N_24778);
nand UO_2713 (O_2713,N_24627,N_24641);
or UO_2714 (O_2714,N_24976,N_24879);
xor UO_2715 (O_2715,N_24616,N_24586);
xor UO_2716 (O_2716,N_24963,N_24516);
nor UO_2717 (O_2717,N_24564,N_24963);
and UO_2718 (O_2718,N_24608,N_24616);
nor UO_2719 (O_2719,N_24546,N_24792);
xor UO_2720 (O_2720,N_24534,N_24939);
nor UO_2721 (O_2721,N_24953,N_24604);
xnor UO_2722 (O_2722,N_24884,N_24755);
nor UO_2723 (O_2723,N_24827,N_24901);
nand UO_2724 (O_2724,N_24694,N_24557);
and UO_2725 (O_2725,N_24602,N_24628);
xnor UO_2726 (O_2726,N_24884,N_24596);
and UO_2727 (O_2727,N_24691,N_24584);
xor UO_2728 (O_2728,N_24537,N_24895);
nor UO_2729 (O_2729,N_24693,N_24877);
and UO_2730 (O_2730,N_24732,N_24654);
or UO_2731 (O_2731,N_24622,N_24801);
and UO_2732 (O_2732,N_24626,N_24923);
nor UO_2733 (O_2733,N_24606,N_24997);
and UO_2734 (O_2734,N_24779,N_24542);
nand UO_2735 (O_2735,N_24965,N_24611);
xnor UO_2736 (O_2736,N_24671,N_24816);
xor UO_2737 (O_2737,N_24658,N_24887);
or UO_2738 (O_2738,N_24567,N_24807);
and UO_2739 (O_2739,N_24678,N_24627);
nor UO_2740 (O_2740,N_24913,N_24604);
or UO_2741 (O_2741,N_24827,N_24889);
xor UO_2742 (O_2742,N_24697,N_24536);
nor UO_2743 (O_2743,N_24992,N_24832);
and UO_2744 (O_2744,N_24657,N_24539);
and UO_2745 (O_2745,N_24734,N_24742);
and UO_2746 (O_2746,N_24865,N_24688);
xnor UO_2747 (O_2747,N_24730,N_24861);
or UO_2748 (O_2748,N_24805,N_24644);
xnor UO_2749 (O_2749,N_24612,N_24762);
nand UO_2750 (O_2750,N_24609,N_24841);
nor UO_2751 (O_2751,N_24938,N_24525);
xnor UO_2752 (O_2752,N_24530,N_24809);
or UO_2753 (O_2753,N_24789,N_24652);
xnor UO_2754 (O_2754,N_24743,N_24553);
nand UO_2755 (O_2755,N_24538,N_24997);
or UO_2756 (O_2756,N_24729,N_24534);
nor UO_2757 (O_2757,N_24846,N_24782);
nand UO_2758 (O_2758,N_24611,N_24699);
nand UO_2759 (O_2759,N_24784,N_24908);
and UO_2760 (O_2760,N_24525,N_24727);
and UO_2761 (O_2761,N_24734,N_24863);
nand UO_2762 (O_2762,N_24811,N_24809);
xnor UO_2763 (O_2763,N_24893,N_24816);
nand UO_2764 (O_2764,N_24580,N_24919);
or UO_2765 (O_2765,N_24641,N_24928);
nor UO_2766 (O_2766,N_24717,N_24879);
and UO_2767 (O_2767,N_24836,N_24973);
or UO_2768 (O_2768,N_24728,N_24882);
and UO_2769 (O_2769,N_24729,N_24803);
nor UO_2770 (O_2770,N_24978,N_24903);
nor UO_2771 (O_2771,N_24978,N_24933);
nand UO_2772 (O_2772,N_24605,N_24871);
and UO_2773 (O_2773,N_24567,N_24581);
and UO_2774 (O_2774,N_24632,N_24640);
or UO_2775 (O_2775,N_24535,N_24659);
or UO_2776 (O_2776,N_24880,N_24516);
and UO_2777 (O_2777,N_24872,N_24982);
and UO_2778 (O_2778,N_24828,N_24956);
xor UO_2779 (O_2779,N_24595,N_24975);
xor UO_2780 (O_2780,N_24689,N_24694);
nor UO_2781 (O_2781,N_24922,N_24561);
or UO_2782 (O_2782,N_24990,N_24996);
xnor UO_2783 (O_2783,N_24757,N_24529);
nor UO_2784 (O_2784,N_24620,N_24546);
xnor UO_2785 (O_2785,N_24950,N_24823);
xor UO_2786 (O_2786,N_24582,N_24665);
or UO_2787 (O_2787,N_24820,N_24968);
xor UO_2788 (O_2788,N_24628,N_24861);
xnor UO_2789 (O_2789,N_24878,N_24998);
and UO_2790 (O_2790,N_24913,N_24918);
nand UO_2791 (O_2791,N_24861,N_24738);
and UO_2792 (O_2792,N_24856,N_24605);
or UO_2793 (O_2793,N_24937,N_24640);
nor UO_2794 (O_2794,N_24667,N_24952);
and UO_2795 (O_2795,N_24946,N_24707);
xnor UO_2796 (O_2796,N_24589,N_24522);
and UO_2797 (O_2797,N_24836,N_24830);
xor UO_2798 (O_2798,N_24510,N_24890);
nor UO_2799 (O_2799,N_24791,N_24693);
xor UO_2800 (O_2800,N_24535,N_24520);
nor UO_2801 (O_2801,N_24803,N_24666);
xor UO_2802 (O_2802,N_24587,N_24677);
and UO_2803 (O_2803,N_24575,N_24691);
or UO_2804 (O_2804,N_24794,N_24870);
nand UO_2805 (O_2805,N_24923,N_24515);
xnor UO_2806 (O_2806,N_24615,N_24813);
xnor UO_2807 (O_2807,N_24907,N_24991);
nand UO_2808 (O_2808,N_24846,N_24615);
xnor UO_2809 (O_2809,N_24624,N_24593);
nor UO_2810 (O_2810,N_24562,N_24878);
nand UO_2811 (O_2811,N_24961,N_24872);
nor UO_2812 (O_2812,N_24528,N_24924);
and UO_2813 (O_2813,N_24647,N_24768);
nor UO_2814 (O_2814,N_24896,N_24972);
or UO_2815 (O_2815,N_24714,N_24504);
nand UO_2816 (O_2816,N_24765,N_24758);
or UO_2817 (O_2817,N_24648,N_24977);
xnor UO_2818 (O_2818,N_24645,N_24763);
xor UO_2819 (O_2819,N_24823,N_24649);
and UO_2820 (O_2820,N_24676,N_24917);
nand UO_2821 (O_2821,N_24703,N_24508);
nand UO_2822 (O_2822,N_24647,N_24838);
nand UO_2823 (O_2823,N_24759,N_24819);
nand UO_2824 (O_2824,N_24783,N_24620);
xnor UO_2825 (O_2825,N_24632,N_24972);
nor UO_2826 (O_2826,N_24866,N_24907);
xor UO_2827 (O_2827,N_24871,N_24833);
or UO_2828 (O_2828,N_24568,N_24953);
or UO_2829 (O_2829,N_24896,N_24746);
nor UO_2830 (O_2830,N_24699,N_24808);
nor UO_2831 (O_2831,N_24898,N_24762);
and UO_2832 (O_2832,N_24786,N_24860);
nor UO_2833 (O_2833,N_24629,N_24851);
nor UO_2834 (O_2834,N_24987,N_24902);
nand UO_2835 (O_2835,N_24927,N_24939);
xnor UO_2836 (O_2836,N_24714,N_24798);
xnor UO_2837 (O_2837,N_24957,N_24895);
and UO_2838 (O_2838,N_24867,N_24649);
and UO_2839 (O_2839,N_24934,N_24822);
and UO_2840 (O_2840,N_24755,N_24742);
nor UO_2841 (O_2841,N_24982,N_24539);
nand UO_2842 (O_2842,N_24544,N_24645);
nand UO_2843 (O_2843,N_24984,N_24796);
nor UO_2844 (O_2844,N_24925,N_24621);
xnor UO_2845 (O_2845,N_24662,N_24850);
or UO_2846 (O_2846,N_24639,N_24883);
and UO_2847 (O_2847,N_24544,N_24678);
nor UO_2848 (O_2848,N_24658,N_24537);
nand UO_2849 (O_2849,N_24728,N_24621);
and UO_2850 (O_2850,N_24981,N_24794);
nor UO_2851 (O_2851,N_24988,N_24653);
nand UO_2852 (O_2852,N_24660,N_24708);
or UO_2853 (O_2853,N_24923,N_24886);
or UO_2854 (O_2854,N_24516,N_24602);
nor UO_2855 (O_2855,N_24604,N_24920);
xnor UO_2856 (O_2856,N_24591,N_24796);
or UO_2857 (O_2857,N_24620,N_24544);
or UO_2858 (O_2858,N_24780,N_24511);
nand UO_2859 (O_2859,N_24857,N_24621);
nor UO_2860 (O_2860,N_24925,N_24746);
nand UO_2861 (O_2861,N_24933,N_24738);
or UO_2862 (O_2862,N_24891,N_24825);
or UO_2863 (O_2863,N_24706,N_24881);
xnor UO_2864 (O_2864,N_24594,N_24801);
nor UO_2865 (O_2865,N_24805,N_24793);
or UO_2866 (O_2866,N_24892,N_24764);
xor UO_2867 (O_2867,N_24629,N_24664);
and UO_2868 (O_2868,N_24991,N_24860);
nor UO_2869 (O_2869,N_24911,N_24928);
or UO_2870 (O_2870,N_24869,N_24661);
nand UO_2871 (O_2871,N_24992,N_24804);
nand UO_2872 (O_2872,N_24519,N_24766);
or UO_2873 (O_2873,N_24923,N_24727);
or UO_2874 (O_2874,N_24889,N_24998);
nand UO_2875 (O_2875,N_24766,N_24731);
xor UO_2876 (O_2876,N_24885,N_24502);
or UO_2877 (O_2877,N_24511,N_24606);
nor UO_2878 (O_2878,N_24518,N_24689);
nand UO_2879 (O_2879,N_24773,N_24829);
and UO_2880 (O_2880,N_24704,N_24741);
and UO_2881 (O_2881,N_24832,N_24913);
xor UO_2882 (O_2882,N_24630,N_24681);
xor UO_2883 (O_2883,N_24552,N_24869);
nor UO_2884 (O_2884,N_24926,N_24657);
xor UO_2885 (O_2885,N_24610,N_24779);
xnor UO_2886 (O_2886,N_24746,N_24857);
xor UO_2887 (O_2887,N_24577,N_24774);
nand UO_2888 (O_2888,N_24841,N_24824);
nand UO_2889 (O_2889,N_24593,N_24765);
nor UO_2890 (O_2890,N_24609,N_24702);
xnor UO_2891 (O_2891,N_24520,N_24625);
nor UO_2892 (O_2892,N_24939,N_24891);
and UO_2893 (O_2893,N_24659,N_24978);
or UO_2894 (O_2894,N_24812,N_24937);
or UO_2895 (O_2895,N_24699,N_24521);
nor UO_2896 (O_2896,N_24591,N_24866);
and UO_2897 (O_2897,N_24856,N_24560);
nand UO_2898 (O_2898,N_24834,N_24532);
and UO_2899 (O_2899,N_24954,N_24511);
and UO_2900 (O_2900,N_24598,N_24840);
nand UO_2901 (O_2901,N_24846,N_24970);
nand UO_2902 (O_2902,N_24740,N_24583);
or UO_2903 (O_2903,N_24614,N_24889);
nand UO_2904 (O_2904,N_24999,N_24979);
or UO_2905 (O_2905,N_24713,N_24985);
nor UO_2906 (O_2906,N_24806,N_24810);
xnor UO_2907 (O_2907,N_24882,N_24731);
or UO_2908 (O_2908,N_24738,N_24712);
xnor UO_2909 (O_2909,N_24695,N_24884);
nand UO_2910 (O_2910,N_24932,N_24898);
or UO_2911 (O_2911,N_24701,N_24975);
nor UO_2912 (O_2912,N_24865,N_24994);
xor UO_2913 (O_2913,N_24953,N_24569);
or UO_2914 (O_2914,N_24924,N_24606);
nand UO_2915 (O_2915,N_24659,N_24800);
nand UO_2916 (O_2916,N_24619,N_24868);
xnor UO_2917 (O_2917,N_24555,N_24827);
or UO_2918 (O_2918,N_24687,N_24564);
nor UO_2919 (O_2919,N_24904,N_24969);
nor UO_2920 (O_2920,N_24777,N_24817);
nor UO_2921 (O_2921,N_24543,N_24677);
nor UO_2922 (O_2922,N_24932,N_24669);
and UO_2923 (O_2923,N_24852,N_24702);
and UO_2924 (O_2924,N_24819,N_24995);
and UO_2925 (O_2925,N_24781,N_24623);
and UO_2926 (O_2926,N_24659,N_24790);
nand UO_2927 (O_2927,N_24975,N_24596);
and UO_2928 (O_2928,N_24894,N_24554);
nand UO_2929 (O_2929,N_24942,N_24756);
xor UO_2930 (O_2930,N_24571,N_24908);
or UO_2931 (O_2931,N_24958,N_24554);
nor UO_2932 (O_2932,N_24953,N_24917);
or UO_2933 (O_2933,N_24525,N_24781);
nor UO_2934 (O_2934,N_24854,N_24822);
nand UO_2935 (O_2935,N_24643,N_24856);
and UO_2936 (O_2936,N_24502,N_24681);
and UO_2937 (O_2937,N_24960,N_24733);
and UO_2938 (O_2938,N_24516,N_24558);
nor UO_2939 (O_2939,N_24837,N_24728);
and UO_2940 (O_2940,N_24553,N_24724);
xor UO_2941 (O_2941,N_24575,N_24552);
or UO_2942 (O_2942,N_24612,N_24655);
xor UO_2943 (O_2943,N_24938,N_24622);
nand UO_2944 (O_2944,N_24876,N_24556);
xor UO_2945 (O_2945,N_24997,N_24778);
nor UO_2946 (O_2946,N_24575,N_24894);
nor UO_2947 (O_2947,N_24889,N_24895);
nand UO_2948 (O_2948,N_24604,N_24671);
xnor UO_2949 (O_2949,N_24742,N_24786);
nand UO_2950 (O_2950,N_24712,N_24613);
nand UO_2951 (O_2951,N_24552,N_24779);
xnor UO_2952 (O_2952,N_24789,N_24995);
or UO_2953 (O_2953,N_24832,N_24668);
or UO_2954 (O_2954,N_24599,N_24683);
and UO_2955 (O_2955,N_24662,N_24573);
nor UO_2956 (O_2956,N_24954,N_24870);
nand UO_2957 (O_2957,N_24609,N_24748);
nand UO_2958 (O_2958,N_24696,N_24685);
xnor UO_2959 (O_2959,N_24525,N_24788);
and UO_2960 (O_2960,N_24697,N_24622);
nand UO_2961 (O_2961,N_24531,N_24831);
nand UO_2962 (O_2962,N_24982,N_24788);
and UO_2963 (O_2963,N_24593,N_24898);
nand UO_2964 (O_2964,N_24652,N_24504);
nand UO_2965 (O_2965,N_24751,N_24601);
or UO_2966 (O_2966,N_24770,N_24501);
nand UO_2967 (O_2967,N_24563,N_24682);
xnor UO_2968 (O_2968,N_24723,N_24685);
xor UO_2969 (O_2969,N_24928,N_24518);
and UO_2970 (O_2970,N_24840,N_24528);
nand UO_2971 (O_2971,N_24881,N_24896);
or UO_2972 (O_2972,N_24809,N_24605);
and UO_2973 (O_2973,N_24541,N_24948);
xnor UO_2974 (O_2974,N_24998,N_24759);
xor UO_2975 (O_2975,N_24919,N_24882);
nand UO_2976 (O_2976,N_24878,N_24617);
nand UO_2977 (O_2977,N_24618,N_24531);
or UO_2978 (O_2978,N_24759,N_24583);
and UO_2979 (O_2979,N_24930,N_24661);
nand UO_2980 (O_2980,N_24717,N_24683);
xnor UO_2981 (O_2981,N_24503,N_24578);
and UO_2982 (O_2982,N_24530,N_24876);
and UO_2983 (O_2983,N_24683,N_24764);
or UO_2984 (O_2984,N_24717,N_24604);
or UO_2985 (O_2985,N_24938,N_24812);
and UO_2986 (O_2986,N_24899,N_24903);
or UO_2987 (O_2987,N_24870,N_24922);
xor UO_2988 (O_2988,N_24619,N_24892);
xor UO_2989 (O_2989,N_24876,N_24903);
xor UO_2990 (O_2990,N_24526,N_24594);
nor UO_2991 (O_2991,N_24562,N_24800);
or UO_2992 (O_2992,N_24928,N_24997);
xor UO_2993 (O_2993,N_24513,N_24799);
or UO_2994 (O_2994,N_24927,N_24570);
xor UO_2995 (O_2995,N_24774,N_24893);
nand UO_2996 (O_2996,N_24534,N_24518);
nor UO_2997 (O_2997,N_24870,N_24761);
nor UO_2998 (O_2998,N_24819,N_24761);
and UO_2999 (O_2999,N_24804,N_24859);
endmodule