module basic_1000_10000_1500_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_77,In_674);
xnor U1 (N_1,In_503,In_297);
or U2 (N_2,In_409,In_425);
nor U3 (N_3,In_890,In_858);
nor U4 (N_4,In_311,In_208);
xnor U5 (N_5,In_748,In_967);
nor U6 (N_6,In_542,In_44);
xor U7 (N_7,In_371,In_68);
and U8 (N_8,In_463,In_288);
and U9 (N_9,In_79,In_388);
nand U10 (N_10,In_85,In_113);
nand U11 (N_11,In_485,In_57);
or U12 (N_12,In_680,In_339);
nand U13 (N_13,In_779,In_508);
or U14 (N_14,In_277,In_211);
or U15 (N_15,In_49,In_134);
and U16 (N_16,In_133,In_222);
and U17 (N_17,In_185,In_873);
nor U18 (N_18,In_290,In_27);
nor U19 (N_19,In_661,In_794);
xnor U20 (N_20,In_156,In_189);
and U21 (N_21,In_422,In_381);
nor U22 (N_22,In_7,In_796);
and U23 (N_23,In_398,In_0);
and U24 (N_24,In_584,In_480);
or U25 (N_25,In_482,In_833);
or U26 (N_26,In_334,In_497);
xor U27 (N_27,In_86,In_565);
xor U28 (N_28,In_617,In_214);
and U29 (N_29,In_338,In_636);
nor U30 (N_30,In_15,In_708);
and U31 (N_31,In_595,In_778);
nand U32 (N_32,In_275,In_696);
nand U33 (N_33,In_712,In_135);
nand U34 (N_34,In_915,In_406);
and U35 (N_35,In_386,In_457);
nor U36 (N_36,In_357,In_535);
nor U37 (N_37,In_854,In_511);
nor U38 (N_38,In_885,In_435);
nor U39 (N_39,In_193,In_744);
or U40 (N_40,In_307,In_969);
or U41 (N_41,In_194,In_775);
nor U42 (N_42,In_152,In_175);
nand U43 (N_43,In_606,In_760);
nor U44 (N_44,In_167,In_881);
and U45 (N_45,In_530,In_981);
nand U46 (N_46,In_559,In_868);
or U47 (N_47,In_627,In_819);
nor U48 (N_48,In_160,In_898);
nor U49 (N_49,In_414,In_434);
and U50 (N_50,In_822,In_355);
nand U51 (N_51,In_412,In_618);
nor U52 (N_52,In_766,In_418);
nand U53 (N_53,In_459,In_830);
and U54 (N_54,In_863,In_241);
nand U55 (N_55,In_592,In_664);
or U56 (N_56,In_536,In_832);
xnor U57 (N_57,In_367,In_954);
nand U58 (N_58,In_207,In_839);
or U59 (N_59,In_337,In_4);
nand U60 (N_60,In_147,In_601);
nor U61 (N_61,In_816,In_526);
nand U62 (N_62,In_173,In_332);
nand U63 (N_63,In_267,In_590);
or U64 (N_64,In_893,In_174);
or U65 (N_65,In_46,In_23);
and U66 (N_66,In_827,In_797);
and U67 (N_67,In_493,In_95);
and U68 (N_68,In_293,In_187);
nor U69 (N_69,In_629,In_181);
or U70 (N_70,In_652,In_91);
nand U71 (N_71,In_116,In_826);
nor U72 (N_72,In_573,In_271);
and U73 (N_73,In_413,In_487);
and U74 (N_74,In_453,In_424);
and U75 (N_75,In_249,In_335);
and U76 (N_76,In_206,In_410);
and U77 (N_77,In_221,In_694);
nand U78 (N_78,In_824,In_204);
and U79 (N_79,In_648,In_103);
nor U80 (N_80,In_917,In_679);
or U81 (N_81,In_12,In_415);
and U82 (N_82,In_707,In_743);
and U83 (N_83,In_663,In_318);
and U84 (N_84,In_727,In_899);
nand U85 (N_85,In_693,In_660);
nor U86 (N_86,In_562,In_940);
or U87 (N_87,In_382,In_118);
or U88 (N_88,In_162,In_5);
and U89 (N_89,In_80,In_54);
nor U90 (N_90,In_745,In_846);
xor U91 (N_91,In_923,In_336);
or U92 (N_92,In_352,In_87);
or U93 (N_93,In_729,In_150);
and U94 (N_94,In_914,In_948);
or U95 (N_95,In_452,In_490);
and U96 (N_96,In_228,In_588);
nor U97 (N_97,In_884,In_3);
nand U98 (N_98,In_951,In_281);
and U99 (N_99,In_484,In_986);
or U100 (N_100,In_356,In_427);
nor U101 (N_101,In_966,In_583);
nand U102 (N_102,In_810,In_548);
nand U103 (N_103,In_200,In_780);
and U104 (N_104,In_887,In_419);
or U105 (N_105,In_843,In_107);
nand U106 (N_106,In_404,In_359);
nor U107 (N_107,In_531,In_396);
nor U108 (N_108,In_73,In_402);
xnor U109 (N_109,In_937,In_781);
nor U110 (N_110,In_443,In_544);
nand U111 (N_111,In_977,In_861);
or U112 (N_112,In_31,In_261);
or U113 (N_113,In_84,In_309);
and U114 (N_114,In_755,In_279);
nand U115 (N_115,In_445,In_978);
nor U116 (N_116,In_869,In_945);
nand U117 (N_117,In_697,In_762);
nand U118 (N_118,In_849,In_537);
and U119 (N_119,In_64,In_676);
nor U120 (N_120,In_649,In_34);
or U121 (N_121,In_327,In_580);
nand U122 (N_122,In_539,In_625);
nor U123 (N_123,In_268,In_245);
and U124 (N_124,In_782,In_946);
xnor U125 (N_125,In_972,In_768);
nand U126 (N_126,In_691,In_60);
nand U127 (N_127,In_866,In_577);
nor U128 (N_128,In_259,In_574);
nor U129 (N_129,In_933,In_958);
or U130 (N_130,In_557,In_795);
nor U131 (N_131,In_26,In_837);
nand U132 (N_132,In_812,In_913);
and U133 (N_133,In_353,In_820);
nand U134 (N_134,In_872,In_515);
xnor U135 (N_135,In_883,In_244);
and U136 (N_136,In_231,In_860);
or U137 (N_137,In_274,In_792);
and U138 (N_138,In_513,In_975);
nor U139 (N_139,In_262,In_528);
nor U140 (N_140,In_420,In_551);
nor U141 (N_141,In_13,In_669);
and U142 (N_142,In_767,In_300);
xnor U143 (N_143,In_151,In_599);
or U144 (N_144,In_670,In_989);
nor U145 (N_145,In_753,In_608);
xnor U146 (N_146,In_844,In_876);
nor U147 (N_147,In_104,In_98);
and U148 (N_148,In_329,In_918);
and U149 (N_149,In_639,In_75);
nand U150 (N_150,In_19,In_128);
nor U151 (N_151,In_234,In_489);
nor U152 (N_152,In_260,In_454);
xnor U153 (N_153,In_560,In_704);
or U154 (N_154,In_806,In_289);
nor U155 (N_155,In_864,In_465);
nor U156 (N_156,In_90,In_751);
or U157 (N_157,In_730,In_436);
nand U158 (N_158,In_93,In_344);
nor U159 (N_159,In_610,In_518);
or U160 (N_160,In_350,In_879);
nand U161 (N_161,In_106,In_581);
xor U162 (N_162,In_379,In_220);
xnor U163 (N_163,In_524,In_659);
nand U164 (N_164,In_600,In_127);
and U165 (N_165,In_81,In_437);
nand U166 (N_166,In_593,In_502);
or U167 (N_167,In_397,In_613);
and U168 (N_168,In_455,In_591);
and U169 (N_169,In_125,In_247);
and U170 (N_170,In_121,In_21);
xnor U171 (N_171,In_351,In_813);
nand U172 (N_172,In_891,In_364);
or U173 (N_173,In_165,In_145);
and U174 (N_174,In_146,In_793);
nor U175 (N_175,In_2,In_102);
or U176 (N_176,In_195,In_24);
and U177 (N_177,In_874,In_186);
or U178 (N_178,In_769,In_942);
or U179 (N_179,In_30,In_305);
and U180 (N_180,In_633,In_667);
nand U181 (N_181,In_495,In_51);
nand U182 (N_182,In_752,In_862);
nor U183 (N_183,In_69,In_225);
nor U184 (N_184,In_678,In_505);
or U185 (N_185,In_199,In_934);
nand U186 (N_186,In_809,In_94);
or U187 (N_187,In_110,In_354);
and U188 (N_188,In_473,In_994);
nand U189 (N_189,In_324,In_431);
and U190 (N_190,In_283,In_714);
nor U191 (N_191,In_159,In_142);
nor U192 (N_192,In_988,In_39);
nor U193 (N_193,In_735,In_377);
or U194 (N_194,In_984,In_76);
nand U195 (N_195,In_461,In_925);
nand U196 (N_196,In_963,In_799);
nor U197 (N_197,In_525,In_257);
xnor U198 (N_198,In_558,In_37);
or U199 (N_199,In_728,In_428);
or U200 (N_200,In_850,In_657);
or U201 (N_201,In_952,In_423);
nand U202 (N_202,In_673,In_519);
or U203 (N_203,In_197,In_835);
and U204 (N_204,In_772,In_22);
xor U205 (N_205,In_690,In_201);
and U206 (N_206,In_349,In_492);
and U207 (N_207,In_999,In_276);
nand U208 (N_208,In_790,In_615);
nor U209 (N_209,In_70,In_761);
or U210 (N_210,In_89,In_582);
nor U211 (N_211,In_702,In_469);
nor U212 (N_212,In_153,In_255);
nor U213 (N_213,In_552,In_654);
or U214 (N_214,In_366,In_805);
nor U215 (N_215,In_58,In_213);
nor U216 (N_216,In_677,In_32);
or U217 (N_217,In_916,In_976);
or U218 (N_218,In_734,In_789);
nand U219 (N_219,In_756,In_330);
xnor U220 (N_220,In_739,In_446);
and U221 (N_221,In_96,In_266);
nand U222 (N_222,In_814,In_196);
and U223 (N_223,In_429,In_987);
nand U224 (N_224,In_741,In_785);
xnor U225 (N_225,In_836,In_626);
or U226 (N_226,In_763,In_631);
and U227 (N_227,In_912,In_112);
nor U228 (N_228,In_251,In_853);
nand U229 (N_229,In_383,In_348);
and U230 (N_230,In_645,In_962);
xor U231 (N_231,In_227,In_757);
and U232 (N_232,In_229,In_687);
nor U233 (N_233,In_233,In_807);
and U234 (N_234,In_650,In_296);
or U235 (N_235,In_564,In_10);
nand U236 (N_236,In_571,In_928);
and U237 (N_237,In_272,In_802);
nor U238 (N_238,In_252,In_341);
nand U239 (N_239,In_968,In_541);
or U240 (N_240,In_665,In_164);
xnor U241 (N_241,In_685,In_961);
or U242 (N_242,In_630,In_852);
nor U243 (N_243,In_566,In_360);
nand U244 (N_244,In_749,In_53);
and U245 (N_245,In_910,In_897);
or U246 (N_246,In_139,In_363);
or U247 (N_247,In_131,In_389);
or U248 (N_248,In_859,In_280);
nand U249 (N_249,In_892,In_343);
nand U250 (N_250,In_273,In_500);
and U251 (N_251,In_787,In_433);
or U252 (N_252,In_88,In_394);
or U253 (N_253,In_698,In_479);
and U254 (N_254,In_686,In_907);
nor U255 (N_255,In_403,In_731);
xnor U256 (N_256,In_587,In_243);
nand U257 (N_257,In_370,In_672);
or U258 (N_258,In_450,In_67);
or U259 (N_259,In_902,In_522);
nor U260 (N_260,In_949,In_701);
or U261 (N_261,In_263,In_292);
nor U262 (N_262,In_927,In_115);
nor U263 (N_263,In_20,In_230);
or U264 (N_264,In_765,In_284);
or U265 (N_265,In_959,In_303);
and U266 (N_266,In_579,In_442);
nand U267 (N_267,In_432,In_798);
nand U268 (N_268,In_250,In_725);
xor U269 (N_269,In_170,In_521);
nor U270 (N_270,In_59,In_373);
and U271 (N_271,In_746,In_632);
and U272 (N_272,In_737,In_460);
nor U273 (N_273,In_317,In_998);
nor U274 (N_274,In_66,In_732);
xor U275 (N_275,In_742,In_378);
and U276 (N_276,In_689,In_320);
nand U277 (N_277,In_140,In_821);
nor U278 (N_278,In_563,In_865);
or U279 (N_279,In_101,In_333);
or U280 (N_280,In_705,In_831);
nand U281 (N_281,In_190,In_609);
xor U282 (N_282,In_567,In_527);
nor U283 (N_283,In_662,In_471);
nand U284 (N_284,In_904,In_776);
nand U285 (N_285,In_417,In_240);
and U286 (N_286,In_561,In_903);
or U287 (N_287,In_611,In_711);
nor U288 (N_288,In_997,In_323);
or U289 (N_289,In_971,In_294);
nor U290 (N_290,In_543,In_517);
nor U291 (N_291,In_188,In_920);
nand U292 (N_292,In_720,In_834);
or U293 (N_293,In_804,In_168);
and U294 (N_294,In_264,In_786);
and U295 (N_295,In_520,In_498);
nand U296 (N_296,In_950,In_395);
nand U297 (N_297,In_614,In_651);
and U298 (N_298,In_299,In_439);
or U299 (N_299,In_331,In_61);
nand U300 (N_300,In_808,In_970);
and U301 (N_301,In_235,In_304);
or U302 (N_302,In_342,In_390);
nand U303 (N_303,In_236,In_932);
nand U304 (N_304,In_965,In_387);
nor U305 (N_305,In_124,In_688);
nor U306 (N_306,In_120,In_210);
xor U307 (N_307,In_468,In_212);
and U308 (N_308,In_671,In_620);
nor U309 (N_309,In_393,In_472);
and U310 (N_310,In_921,In_576);
nand U311 (N_311,In_100,In_656);
nor U312 (N_312,In_215,In_33);
and U313 (N_313,In_895,In_623);
nor U314 (N_314,In_646,In_25);
nand U315 (N_315,In_486,In_365);
and U316 (N_316,In_510,In_216);
or U317 (N_317,In_960,In_842);
nor U318 (N_318,In_622,In_132);
and U319 (N_319,In_1,In_555);
and U320 (N_320,In_313,In_713);
nand U321 (N_321,In_302,In_644);
or U322 (N_322,In_924,In_384);
or U323 (N_323,In_758,In_628);
nand U324 (N_324,In_218,In_483);
nor U325 (N_325,In_62,In_990);
nand U326 (N_326,In_78,In_771);
and U327 (N_327,In_974,In_889);
nand U328 (N_328,In_178,In_594);
or U329 (N_329,In_385,In_163);
and U330 (N_330,In_941,In_438);
xnor U331 (N_331,In_641,In_14);
or U332 (N_332,In_901,In_870);
and U333 (N_333,In_703,In_791);
and U334 (N_334,In_896,In_991);
nor U335 (N_335,In_532,In_71);
nor U336 (N_336,In_538,In_391);
and U337 (N_337,In_295,In_724);
nand U338 (N_338,In_65,In_788);
nor U339 (N_339,In_926,In_695);
and U340 (N_340,In_143,In_871);
or U341 (N_341,In_491,In_494);
nand U342 (N_342,In_621,In_717);
and U343 (N_343,In_955,In_176);
or U344 (N_344,In_43,In_957);
nor U345 (N_345,In_298,In_774);
nor U346 (N_346,In_444,In_604);
nor U347 (N_347,In_306,In_578);
nand U348 (N_348,In_764,In_985);
xor U349 (N_349,In_715,In_516);
nand U350 (N_350,In_840,In_52);
nand U351 (N_351,In_709,In_137);
and U352 (N_352,In_750,In_825);
and U353 (N_353,In_253,In_488);
and U354 (N_354,In_637,In_326);
nand U355 (N_355,In_114,In_42);
nor U356 (N_356,In_922,In_655);
or U357 (N_357,In_722,In_909);
or U358 (N_358,In_880,In_346);
nor U359 (N_359,In_286,In_523);
nand U360 (N_360,In_700,In_938);
nand U361 (N_361,In_278,In_270);
or U362 (N_362,In_647,In_108);
or U363 (N_363,In_144,In_449);
and U364 (N_364,In_801,In_224);
nor U365 (N_365,In_166,In_258);
xnor U366 (N_366,In_282,In_408);
or U367 (N_367,In_29,In_347);
or U368 (N_368,In_17,In_556);
and U369 (N_369,In_803,In_710);
nor U370 (N_370,In_223,In_640);
nor U371 (N_371,In_930,In_507);
nand U372 (N_372,In_553,In_470);
or U373 (N_373,In_63,In_856);
nand U374 (N_374,In_18,In_919);
and U375 (N_375,In_619,In_514);
nand U376 (N_376,In_867,In_456);
or U377 (N_377,In_589,In_586);
nand U378 (N_378,In_602,In_105);
xor U379 (N_379,In_430,In_192);
or U380 (N_380,In_754,In_154);
and U381 (N_381,In_109,In_130);
or U382 (N_382,In_369,In_111);
nand U383 (N_383,In_180,In_447);
nand U384 (N_384,In_9,In_421);
or U385 (N_385,In_939,In_183);
and U386 (N_386,In_770,In_56);
xnor U387 (N_387,In_28,In_900);
or U388 (N_388,In_345,In_35);
nor U389 (N_389,In_911,In_248);
or U390 (N_390,In_41,In_426);
or U391 (N_391,In_478,In_740);
nand U392 (N_392,In_980,In_401);
nand U393 (N_393,In_529,In_845);
nand U394 (N_394,In_8,In_596);
nand U395 (N_395,In_179,In_198);
nor U396 (N_396,In_585,In_226);
nor U397 (N_397,In_848,In_291);
xor U398 (N_398,In_405,In_607);
nor U399 (N_399,In_238,In_6);
and U400 (N_400,In_747,In_82);
xor U401 (N_401,In_316,In_718);
nor U402 (N_402,In_310,In_182);
nor U403 (N_403,In_314,In_256);
nor U404 (N_404,In_45,In_123);
nand U405 (N_405,In_375,In_823);
or U406 (N_406,In_504,In_285);
nor U407 (N_407,In_466,In_547);
and U408 (N_408,In_501,In_237);
nand U409 (N_409,In_119,In_572);
nor U410 (N_410,In_141,In_815);
or U411 (N_411,In_246,In_308);
or U412 (N_412,In_828,In_759);
nand U413 (N_413,In_47,In_545);
nor U414 (N_414,In_161,In_400);
or U415 (N_415,In_624,In_973);
or U416 (N_416,In_362,In_157);
nor U417 (N_417,In_777,In_875);
xnor U418 (N_418,In_706,In_947);
nand U419 (N_419,In_612,In_851);
nand U420 (N_420,In_155,In_817);
or U421 (N_421,In_169,In_117);
nor U422 (N_422,In_841,In_506);
nor U423 (N_423,In_953,In_509);
nor U424 (N_424,In_499,In_605);
nand U425 (N_425,In_800,In_462);
nand U426 (N_426,In_996,In_982);
nor U427 (N_427,In_983,In_908);
and U428 (N_428,In_368,In_943);
xor U429 (N_429,In_638,In_719);
or U430 (N_430,In_16,In_857);
nor U431 (N_431,In_40,In_675);
or U432 (N_432,In_138,In_217);
nand U433 (N_433,In_315,In_684);
or U434 (N_434,In_392,In_936);
nand U435 (N_435,In_411,In_126);
nand U436 (N_436,In_242,In_97);
nor U437 (N_437,In_886,In_407);
nor U438 (N_438,In_549,In_50);
nand U439 (N_439,In_733,In_888);
nor U440 (N_440,In_209,In_475);
or U441 (N_441,In_603,In_546);
or U442 (N_442,In_668,In_340);
nor U443 (N_443,In_653,In_441);
or U444 (N_444,In_301,In_992);
or U445 (N_445,In_328,In_935);
or U446 (N_446,In_597,In_550);
nand U447 (N_447,In_534,In_172);
and U448 (N_448,In_321,In_682);
and U449 (N_449,In_372,In_205);
nor U450 (N_450,In_122,In_554);
and U451 (N_451,In_906,In_905);
nor U452 (N_452,In_616,In_634);
nor U453 (N_453,In_993,In_964);
or U454 (N_454,In_956,In_995);
nor U455 (N_455,In_540,In_148);
xor U456 (N_456,In_721,In_448);
or U457 (N_457,In_979,In_72);
nor U458 (N_458,In_882,In_319);
xnor U459 (N_459,In_36,In_877);
nand U460 (N_460,In_136,In_931);
nand U461 (N_461,In_699,In_202);
nand U462 (N_462,In_48,In_773);
nor U463 (N_463,In_451,In_738);
or U464 (N_464,In_726,In_658);
nor U465 (N_465,In_784,In_254);
xnor U466 (N_466,In_361,In_598);
nand U467 (N_467,In_74,In_380);
nor U468 (N_468,In_149,In_736);
nand U469 (N_469,In_440,In_692);
or U470 (N_470,In_239,In_467);
or U471 (N_471,In_838,In_184);
nand U472 (N_472,In_496,In_158);
and U473 (N_473,In_878,In_575);
nand U474 (N_474,In_512,In_269);
or U475 (N_475,In_265,In_458);
nor U476 (N_476,In_219,In_399);
and U477 (N_477,In_635,In_177);
nand U478 (N_478,In_666,In_464);
xnor U479 (N_479,In_312,In_374);
xor U480 (N_480,In_929,In_783);
and U481 (N_481,In_847,In_83);
nor U482 (N_482,In_129,In_643);
nand U483 (N_483,In_481,In_829);
nand U484 (N_484,In_55,In_894);
nor U485 (N_485,In_358,In_322);
xnor U486 (N_486,In_232,In_944);
xor U487 (N_487,In_38,In_11);
nor U488 (N_488,In_191,In_203);
nor U489 (N_489,In_642,In_287);
nor U490 (N_490,In_723,In_477);
nor U491 (N_491,In_855,In_476);
or U492 (N_492,In_376,In_570);
xnor U493 (N_493,In_811,In_416);
nor U494 (N_494,In_681,In_325);
or U495 (N_495,In_716,In_99);
nor U496 (N_496,In_474,In_92);
and U497 (N_497,In_568,In_171);
or U498 (N_498,In_533,In_818);
nor U499 (N_499,In_683,In_569);
and U500 (N_500,In_218,In_235);
nand U501 (N_501,In_423,In_131);
or U502 (N_502,In_809,In_100);
or U503 (N_503,In_102,In_883);
and U504 (N_504,In_113,In_921);
or U505 (N_505,In_812,In_437);
or U506 (N_506,In_512,In_547);
nand U507 (N_507,In_28,In_373);
nor U508 (N_508,In_527,In_359);
nand U509 (N_509,In_420,In_91);
or U510 (N_510,In_626,In_714);
nand U511 (N_511,In_713,In_535);
xnor U512 (N_512,In_697,In_173);
nand U513 (N_513,In_626,In_78);
and U514 (N_514,In_294,In_644);
or U515 (N_515,In_816,In_290);
nand U516 (N_516,In_502,In_640);
or U517 (N_517,In_644,In_104);
nand U518 (N_518,In_488,In_19);
or U519 (N_519,In_344,In_150);
nor U520 (N_520,In_598,In_453);
nand U521 (N_521,In_209,In_971);
and U522 (N_522,In_142,In_849);
and U523 (N_523,In_901,In_783);
nand U524 (N_524,In_616,In_219);
nand U525 (N_525,In_263,In_923);
or U526 (N_526,In_931,In_733);
nand U527 (N_527,In_133,In_66);
nand U528 (N_528,In_867,In_396);
nand U529 (N_529,In_698,In_782);
xor U530 (N_530,In_768,In_726);
nor U531 (N_531,In_622,In_861);
nor U532 (N_532,In_739,In_407);
nor U533 (N_533,In_537,In_844);
nand U534 (N_534,In_653,In_52);
and U535 (N_535,In_14,In_229);
nand U536 (N_536,In_204,In_428);
and U537 (N_537,In_391,In_821);
or U538 (N_538,In_555,In_98);
and U539 (N_539,In_383,In_360);
nor U540 (N_540,In_284,In_700);
and U541 (N_541,In_713,In_403);
nor U542 (N_542,In_115,In_719);
nand U543 (N_543,In_687,In_996);
nand U544 (N_544,In_512,In_466);
nand U545 (N_545,In_905,In_494);
xnor U546 (N_546,In_123,In_918);
or U547 (N_547,In_360,In_838);
nand U548 (N_548,In_91,In_921);
and U549 (N_549,In_64,In_481);
nor U550 (N_550,In_883,In_541);
and U551 (N_551,In_255,In_746);
or U552 (N_552,In_589,In_943);
nand U553 (N_553,In_689,In_668);
nor U554 (N_554,In_711,In_531);
xnor U555 (N_555,In_575,In_876);
and U556 (N_556,In_78,In_778);
or U557 (N_557,In_153,In_689);
xnor U558 (N_558,In_165,In_306);
and U559 (N_559,In_651,In_606);
nand U560 (N_560,In_963,In_462);
xnor U561 (N_561,In_126,In_920);
or U562 (N_562,In_203,In_494);
xor U563 (N_563,In_516,In_471);
or U564 (N_564,In_312,In_587);
or U565 (N_565,In_132,In_792);
xor U566 (N_566,In_199,In_273);
xnor U567 (N_567,In_513,In_772);
nor U568 (N_568,In_218,In_869);
nor U569 (N_569,In_797,In_954);
nor U570 (N_570,In_77,In_530);
nand U571 (N_571,In_71,In_911);
or U572 (N_572,In_219,In_138);
nor U573 (N_573,In_319,In_633);
nor U574 (N_574,In_959,In_706);
and U575 (N_575,In_9,In_248);
nand U576 (N_576,In_396,In_497);
or U577 (N_577,In_631,In_647);
nand U578 (N_578,In_872,In_169);
nor U579 (N_579,In_410,In_224);
or U580 (N_580,In_340,In_817);
nand U581 (N_581,In_543,In_510);
or U582 (N_582,In_880,In_396);
and U583 (N_583,In_588,In_428);
nand U584 (N_584,In_561,In_819);
nor U585 (N_585,In_991,In_422);
nor U586 (N_586,In_370,In_90);
and U587 (N_587,In_391,In_21);
nor U588 (N_588,In_841,In_418);
nor U589 (N_589,In_326,In_947);
nand U590 (N_590,In_943,In_244);
or U591 (N_591,In_414,In_667);
or U592 (N_592,In_48,In_100);
nand U593 (N_593,In_630,In_720);
xor U594 (N_594,In_145,In_278);
or U595 (N_595,In_587,In_395);
nor U596 (N_596,In_382,In_637);
nor U597 (N_597,In_297,In_701);
nand U598 (N_598,In_87,In_657);
nand U599 (N_599,In_137,In_596);
and U600 (N_600,In_829,In_514);
xnor U601 (N_601,In_652,In_19);
or U602 (N_602,In_773,In_920);
nor U603 (N_603,In_955,In_796);
nand U604 (N_604,In_117,In_483);
nor U605 (N_605,In_479,In_672);
nand U606 (N_606,In_818,In_40);
or U607 (N_607,In_654,In_915);
nand U608 (N_608,In_847,In_710);
xor U609 (N_609,In_997,In_690);
nand U610 (N_610,In_377,In_544);
nand U611 (N_611,In_955,In_440);
nor U612 (N_612,In_447,In_737);
nor U613 (N_613,In_737,In_252);
xnor U614 (N_614,In_441,In_599);
or U615 (N_615,In_995,In_672);
and U616 (N_616,In_606,In_6);
or U617 (N_617,In_209,In_801);
and U618 (N_618,In_735,In_676);
nor U619 (N_619,In_233,In_732);
and U620 (N_620,In_233,In_154);
or U621 (N_621,In_10,In_425);
nor U622 (N_622,In_420,In_990);
nor U623 (N_623,In_286,In_813);
nand U624 (N_624,In_595,In_966);
and U625 (N_625,In_432,In_607);
and U626 (N_626,In_158,In_23);
xnor U627 (N_627,In_717,In_386);
nand U628 (N_628,In_939,In_280);
nand U629 (N_629,In_416,In_359);
and U630 (N_630,In_732,In_889);
nor U631 (N_631,In_767,In_805);
nor U632 (N_632,In_138,In_458);
or U633 (N_633,In_682,In_641);
and U634 (N_634,In_139,In_663);
nand U635 (N_635,In_982,In_188);
nor U636 (N_636,In_632,In_344);
or U637 (N_637,In_352,In_219);
nand U638 (N_638,In_364,In_918);
nand U639 (N_639,In_964,In_411);
or U640 (N_640,In_853,In_942);
nand U641 (N_641,In_934,In_847);
nand U642 (N_642,In_730,In_416);
and U643 (N_643,In_183,In_493);
nand U644 (N_644,In_987,In_551);
nand U645 (N_645,In_403,In_295);
nor U646 (N_646,In_200,In_353);
nand U647 (N_647,In_221,In_156);
and U648 (N_648,In_231,In_28);
and U649 (N_649,In_535,In_187);
nor U650 (N_650,In_440,In_177);
xor U651 (N_651,In_290,In_417);
and U652 (N_652,In_692,In_303);
and U653 (N_653,In_3,In_15);
or U654 (N_654,In_116,In_403);
and U655 (N_655,In_319,In_577);
or U656 (N_656,In_438,In_819);
nand U657 (N_657,In_166,In_508);
or U658 (N_658,In_292,In_999);
nor U659 (N_659,In_677,In_174);
nand U660 (N_660,In_672,In_361);
and U661 (N_661,In_250,In_432);
and U662 (N_662,In_398,In_959);
or U663 (N_663,In_201,In_274);
xor U664 (N_664,In_333,In_276);
nor U665 (N_665,In_941,In_622);
or U666 (N_666,In_459,In_24);
nand U667 (N_667,In_496,In_7);
and U668 (N_668,In_893,In_188);
nand U669 (N_669,In_17,In_64);
and U670 (N_670,In_44,In_490);
nor U671 (N_671,In_250,In_444);
or U672 (N_672,In_535,In_134);
or U673 (N_673,In_723,In_217);
nand U674 (N_674,In_938,In_269);
and U675 (N_675,In_220,In_1);
or U676 (N_676,In_881,In_788);
or U677 (N_677,In_885,In_682);
nand U678 (N_678,In_377,In_463);
xnor U679 (N_679,In_646,In_692);
and U680 (N_680,In_258,In_36);
and U681 (N_681,In_694,In_996);
xor U682 (N_682,In_709,In_293);
or U683 (N_683,In_927,In_453);
nand U684 (N_684,In_667,In_15);
and U685 (N_685,In_172,In_794);
nand U686 (N_686,In_973,In_709);
and U687 (N_687,In_489,In_531);
and U688 (N_688,In_887,In_292);
nor U689 (N_689,In_137,In_664);
or U690 (N_690,In_778,In_968);
or U691 (N_691,In_640,In_932);
and U692 (N_692,In_730,In_798);
nor U693 (N_693,In_155,In_73);
and U694 (N_694,In_38,In_84);
nor U695 (N_695,In_975,In_880);
nor U696 (N_696,In_63,In_749);
or U697 (N_697,In_142,In_713);
nand U698 (N_698,In_458,In_210);
nand U699 (N_699,In_306,In_913);
and U700 (N_700,In_661,In_10);
or U701 (N_701,In_828,In_117);
nand U702 (N_702,In_617,In_411);
xnor U703 (N_703,In_461,In_522);
xnor U704 (N_704,In_599,In_264);
or U705 (N_705,In_957,In_312);
and U706 (N_706,In_215,In_289);
and U707 (N_707,In_741,In_819);
and U708 (N_708,In_518,In_387);
nor U709 (N_709,In_540,In_9);
xor U710 (N_710,In_246,In_132);
or U711 (N_711,In_815,In_746);
nor U712 (N_712,In_175,In_246);
xnor U713 (N_713,In_316,In_448);
xor U714 (N_714,In_908,In_169);
nor U715 (N_715,In_780,In_855);
xnor U716 (N_716,In_828,In_316);
xor U717 (N_717,In_160,In_806);
nor U718 (N_718,In_230,In_796);
nand U719 (N_719,In_88,In_481);
xor U720 (N_720,In_85,In_772);
nor U721 (N_721,In_578,In_752);
and U722 (N_722,In_135,In_671);
nand U723 (N_723,In_472,In_942);
and U724 (N_724,In_712,In_277);
or U725 (N_725,In_34,In_894);
nand U726 (N_726,In_105,In_985);
and U727 (N_727,In_432,In_504);
and U728 (N_728,In_285,In_306);
nand U729 (N_729,In_414,In_459);
or U730 (N_730,In_94,In_780);
nand U731 (N_731,In_785,In_989);
or U732 (N_732,In_45,In_438);
or U733 (N_733,In_885,In_67);
and U734 (N_734,In_846,In_407);
nor U735 (N_735,In_553,In_220);
and U736 (N_736,In_857,In_459);
nand U737 (N_737,In_671,In_630);
nor U738 (N_738,In_900,In_738);
or U739 (N_739,In_90,In_448);
and U740 (N_740,In_204,In_270);
nor U741 (N_741,In_718,In_368);
or U742 (N_742,In_418,In_733);
nand U743 (N_743,In_975,In_455);
xor U744 (N_744,In_257,In_857);
and U745 (N_745,In_634,In_627);
nand U746 (N_746,In_117,In_908);
or U747 (N_747,In_330,In_386);
nor U748 (N_748,In_803,In_835);
nor U749 (N_749,In_535,In_137);
and U750 (N_750,In_50,In_351);
xor U751 (N_751,In_574,In_473);
and U752 (N_752,In_565,In_809);
or U753 (N_753,In_185,In_603);
or U754 (N_754,In_81,In_600);
and U755 (N_755,In_651,In_275);
nor U756 (N_756,In_817,In_579);
nand U757 (N_757,In_469,In_699);
xor U758 (N_758,In_196,In_640);
and U759 (N_759,In_82,In_187);
nor U760 (N_760,In_429,In_647);
xnor U761 (N_761,In_300,In_699);
nor U762 (N_762,In_96,In_583);
xnor U763 (N_763,In_957,In_633);
or U764 (N_764,In_565,In_297);
nand U765 (N_765,In_757,In_135);
nand U766 (N_766,In_9,In_913);
or U767 (N_767,In_277,In_38);
and U768 (N_768,In_886,In_753);
or U769 (N_769,In_465,In_271);
nor U770 (N_770,In_966,In_437);
nand U771 (N_771,In_883,In_752);
and U772 (N_772,In_727,In_741);
nand U773 (N_773,In_6,In_210);
nor U774 (N_774,In_469,In_114);
xor U775 (N_775,In_395,In_210);
nand U776 (N_776,In_791,In_112);
nand U777 (N_777,In_539,In_340);
nand U778 (N_778,In_451,In_257);
nor U779 (N_779,In_146,In_828);
and U780 (N_780,In_336,In_354);
or U781 (N_781,In_955,In_893);
nor U782 (N_782,In_854,In_673);
or U783 (N_783,In_968,In_652);
and U784 (N_784,In_813,In_803);
xor U785 (N_785,In_960,In_91);
and U786 (N_786,In_331,In_120);
or U787 (N_787,In_842,In_47);
nand U788 (N_788,In_147,In_970);
nand U789 (N_789,In_687,In_764);
xnor U790 (N_790,In_498,In_452);
xnor U791 (N_791,In_883,In_834);
xnor U792 (N_792,In_785,In_46);
nor U793 (N_793,In_120,In_985);
and U794 (N_794,In_626,In_654);
and U795 (N_795,In_355,In_796);
nand U796 (N_796,In_124,In_218);
nor U797 (N_797,In_635,In_680);
nor U798 (N_798,In_11,In_609);
and U799 (N_799,In_68,In_563);
xnor U800 (N_800,In_419,In_721);
and U801 (N_801,In_168,In_837);
nor U802 (N_802,In_566,In_259);
or U803 (N_803,In_498,In_858);
and U804 (N_804,In_844,In_153);
or U805 (N_805,In_120,In_979);
nor U806 (N_806,In_344,In_349);
nand U807 (N_807,In_305,In_37);
nor U808 (N_808,In_509,In_218);
nand U809 (N_809,In_659,In_241);
and U810 (N_810,In_783,In_937);
nand U811 (N_811,In_899,In_895);
nand U812 (N_812,In_555,In_203);
nand U813 (N_813,In_640,In_191);
nor U814 (N_814,In_267,In_53);
nor U815 (N_815,In_747,In_695);
nor U816 (N_816,In_943,In_694);
and U817 (N_817,In_858,In_290);
nand U818 (N_818,In_744,In_980);
or U819 (N_819,In_528,In_430);
nand U820 (N_820,In_749,In_977);
or U821 (N_821,In_490,In_573);
nor U822 (N_822,In_168,In_294);
nor U823 (N_823,In_710,In_480);
xor U824 (N_824,In_765,In_761);
xnor U825 (N_825,In_83,In_974);
nor U826 (N_826,In_650,In_889);
and U827 (N_827,In_894,In_671);
nor U828 (N_828,In_578,In_57);
and U829 (N_829,In_587,In_358);
xnor U830 (N_830,In_884,In_982);
and U831 (N_831,In_677,In_423);
xnor U832 (N_832,In_931,In_253);
nand U833 (N_833,In_268,In_850);
xor U834 (N_834,In_494,In_288);
and U835 (N_835,In_568,In_775);
nand U836 (N_836,In_152,In_78);
or U837 (N_837,In_195,In_933);
nor U838 (N_838,In_612,In_479);
or U839 (N_839,In_6,In_98);
nand U840 (N_840,In_625,In_668);
xnor U841 (N_841,In_337,In_99);
or U842 (N_842,In_135,In_901);
nand U843 (N_843,In_141,In_335);
or U844 (N_844,In_107,In_372);
nor U845 (N_845,In_668,In_561);
nor U846 (N_846,In_76,In_96);
nand U847 (N_847,In_698,In_891);
or U848 (N_848,In_869,In_314);
nor U849 (N_849,In_763,In_427);
or U850 (N_850,In_806,In_62);
or U851 (N_851,In_532,In_37);
and U852 (N_852,In_883,In_99);
or U853 (N_853,In_503,In_111);
and U854 (N_854,In_998,In_920);
nand U855 (N_855,In_949,In_138);
and U856 (N_856,In_990,In_188);
or U857 (N_857,In_542,In_252);
nor U858 (N_858,In_17,In_216);
nor U859 (N_859,In_611,In_312);
or U860 (N_860,In_3,In_761);
and U861 (N_861,In_849,In_390);
or U862 (N_862,In_284,In_187);
or U863 (N_863,In_715,In_203);
and U864 (N_864,In_946,In_963);
or U865 (N_865,In_793,In_60);
nand U866 (N_866,In_919,In_507);
nor U867 (N_867,In_243,In_359);
or U868 (N_868,In_835,In_25);
nand U869 (N_869,In_729,In_932);
nand U870 (N_870,In_291,In_944);
or U871 (N_871,In_885,In_41);
or U872 (N_872,In_311,In_271);
or U873 (N_873,In_678,In_382);
and U874 (N_874,In_658,In_485);
nand U875 (N_875,In_574,In_6);
xnor U876 (N_876,In_740,In_317);
nor U877 (N_877,In_455,In_839);
nor U878 (N_878,In_214,In_557);
nand U879 (N_879,In_860,In_20);
nor U880 (N_880,In_845,In_924);
nor U881 (N_881,In_256,In_736);
nand U882 (N_882,In_326,In_778);
or U883 (N_883,In_439,In_572);
and U884 (N_884,In_437,In_205);
nand U885 (N_885,In_391,In_748);
nand U886 (N_886,In_768,In_625);
and U887 (N_887,In_948,In_458);
xnor U888 (N_888,In_974,In_243);
or U889 (N_889,In_730,In_92);
and U890 (N_890,In_881,In_860);
nand U891 (N_891,In_251,In_332);
or U892 (N_892,In_52,In_687);
and U893 (N_893,In_622,In_620);
and U894 (N_894,In_137,In_473);
or U895 (N_895,In_490,In_93);
nor U896 (N_896,In_740,In_329);
nand U897 (N_897,In_552,In_82);
nand U898 (N_898,In_205,In_456);
and U899 (N_899,In_443,In_894);
nand U900 (N_900,In_612,In_437);
nand U901 (N_901,In_147,In_154);
nand U902 (N_902,In_993,In_794);
and U903 (N_903,In_160,In_786);
xor U904 (N_904,In_238,In_501);
nand U905 (N_905,In_763,In_447);
and U906 (N_906,In_846,In_516);
nand U907 (N_907,In_692,In_716);
nor U908 (N_908,In_106,In_175);
nor U909 (N_909,In_148,In_548);
and U910 (N_910,In_749,In_272);
nand U911 (N_911,In_9,In_985);
nand U912 (N_912,In_656,In_659);
nand U913 (N_913,In_514,In_353);
and U914 (N_914,In_857,In_152);
nand U915 (N_915,In_976,In_502);
and U916 (N_916,In_736,In_891);
nor U917 (N_917,In_618,In_707);
nand U918 (N_918,In_448,In_935);
nand U919 (N_919,In_786,In_228);
and U920 (N_920,In_293,In_201);
xnor U921 (N_921,In_913,In_365);
nand U922 (N_922,In_47,In_701);
or U923 (N_923,In_486,In_848);
nand U924 (N_924,In_626,In_348);
nor U925 (N_925,In_976,In_32);
xnor U926 (N_926,In_634,In_648);
nand U927 (N_927,In_962,In_243);
nor U928 (N_928,In_661,In_218);
nor U929 (N_929,In_599,In_170);
nand U930 (N_930,In_509,In_768);
and U931 (N_931,In_98,In_836);
and U932 (N_932,In_56,In_787);
xnor U933 (N_933,In_850,In_489);
nor U934 (N_934,In_204,In_551);
nor U935 (N_935,In_891,In_745);
xor U936 (N_936,In_578,In_27);
nor U937 (N_937,In_63,In_39);
nor U938 (N_938,In_365,In_984);
nand U939 (N_939,In_613,In_830);
nor U940 (N_940,In_247,In_642);
or U941 (N_941,In_776,In_202);
nor U942 (N_942,In_501,In_842);
and U943 (N_943,In_861,In_459);
nand U944 (N_944,In_806,In_277);
nor U945 (N_945,In_387,In_467);
and U946 (N_946,In_993,In_817);
nand U947 (N_947,In_5,In_165);
xnor U948 (N_948,In_132,In_27);
or U949 (N_949,In_123,In_444);
nor U950 (N_950,In_495,In_326);
and U951 (N_951,In_88,In_251);
or U952 (N_952,In_688,In_22);
or U953 (N_953,In_654,In_31);
or U954 (N_954,In_460,In_207);
or U955 (N_955,In_745,In_322);
or U956 (N_956,In_730,In_649);
or U957 (N_957,In_879,In_842);
xnor U958 (N_958,In_612,In_908);
nand U959 (N_959,In_127,In_453);
and U960 (N_960,In_729,In_265);
xor U961 (N_961,In_222,In_303);
and U962 (N_962,In_927,In_867);
nor U963 (N_963,In_496,In_285);
or U964 (N_964,In_286,In_585);
nor U965 (N_965,In_44,In_118);
nand U966 (N_966,In_436,In_838);
xnor U967 (N_967,In_615,In_52);
or U968 (N_968,In_139,In_500);
nor U969 (N_969,In_442,In_49);
and U970 (N_970,In_621,In_604);
nor U971 (N_971,In_154,In_459);
xor U972 (N_972,In_785,In_648);
xnor U973 (N_973,In_715,In_889);
and U974 (N_974,In_728,In_318);
and U975 (N_975,In_949,In_866);
or U976 (N_976,In_543,In_725);
nor U977 (N_977,In_493,In_706);
nand U978 (N_978,In_294,In_999);
and U979 (N_979,In_146,In_503);
or U980 (N_980,In_562,In_953);
or U981 (N_981,In_389,In_966);
nor U982 (N_982,In_495,In_372);
nand U983 (N_983,In_40,In_78);
or U984 (N_984,In_735,In_26);
nand U985 (N_985,In_522,In_170);
or U986 (N_986,In_2,In_382);
nand U987 (N_987,In_476,In_961);
and U988 (N_988,In_53,In_207);
nor U989 (N_989,In_581,In_746);
nand U990 (N_990,In_65,In_708);
and U991 (N_991,In_375,In_532);
or U992 (N_992,In_774,In_726);
nand U993 (N_993,In_571,In_247);
nand U994 (N_994,In_518,In_96);
or U995 (N_995,In_606,In_403);
and U996 (N_996,In_714,In_223);
xor U997 (N_997,In_181,In_889);
nand U998 (N_998,In_74,In_326);
xnor U999 (N_999,In_572,In_514);
nor U1000 (N_1000,N_424,N_798);
and U1001 (N_1001,N_894,N_836);
or U1002 (N_1002,N_282,N_514);
nor U1003 (N_1003,N_785,N_824);
nor U1004 (N_1004,N_461,N_857);
nand U1005 (N_1005,N_649,N_290);
and U1006 (N_1006,N_618,N_680);
nand U1007 (N_1007,N_408,N_473);
nor U1008 (N_1008,N_488,N_376);
or U1009 (N_1009,N_257,N_985);
and U1010 (N_1010,N_31,N_792);
nor U1011 (N_1011,N_579,N_839);
or U1012 (N_1012,N_727,N_450);
nand U1013 (N_1013,N_948,N_941);
nor U1014 (N_1014,N_577,N_572);
nor U1015 (N_1015,N_414,N_558);
or U1016 (N_1016,N_858,N_674);
nand U1017 (N_1017,N_964,N_32);
or U1018 (N_1018,N_500,N_402);
nor U1019 (N_1019,N_602,N_411);
xor U1020 (N_1020,N_502,N_813);
nor U1021 (N_1021,N_662,N_404);
and U1022 (N_1022,N_581,N_604);
or U1023 (N_1023,N_217,N_817);
nor U1024 (N_1024,N_534,N_483);
xor U1025 (N_1025,N_56,N_441);
and U1026 (N_1026,N_811,N_999);
nor U1027 (N_1027,N_864,N_417);
and U1028 (N_1028,N_762,N_564);
or U1029 (N_1029,N_748,N_945);
xnor U1030 (N_1030,N_278,N_54);
nand U1031 (N_1031,N_459,N_511);
nand U1032 (N_1032,N_825,N_679);
nand U1033 (N_1033,N_851,N_144);
and U1034 (N_1034,N_816,N_910);
or U1035 (N_1035,N_318,N_261);
or U1036 (N_1036,N_196,N_706);
or U1037 (N_1037,N_177,N_694);
nand U1038 (N_1038,N_353,N_667);
xnor U1039 (N_1039,N_982,N_549);
or U1040 (N_1040,N_430,N_949);
nor U1041 (N_1041,N_886,N_270);
nor U1042 (N_1042,N_340,N_292);
or U1043 (N_1043,N_908,N_291);
nand U1044 (N_1044,N_116,N_763);
or U1045 (N_1045,N_744,N_302);
and U1046 (N_1046,N_573,N_717);
xnor U1047 (N_1047,N_133,N_78);
nand U1048 (N_1048,N_884,N_220);
nor U1049 (N_1049,N_157,N_466);
and U1050 (N_1050,N_223,N_683);
and U1051 (N_1051,N_236,N_963);
nor U1052 (N_1052,N_233,N_974);
nor U1053 (N_1053,N_207,N_400);
xnor U1054 (N_1054,N_969,N_922);
and U1055 (N_1055,N_678,N_94);
and U1056 (N_1056,N_237,N_85);
nand U1057 (N_1057,N_395,N_988);
nand U1058 (N_1058,N_814,N_743);
or U1059 (N_1059,N_383,N_780);
or U1060 (N_1060,N_841,N_164);
and U1061 (N_1061,N_289,N_701);
xor U1062 (N_1062,N_19,N_18);
xor U1063 (N_1063,N_137,N_193);
or U1064 (N_1064,N_854,N_728);
nor U1065 (N_1065,N_457,N_741);
nand U1066 (N_1066,N_893,N_720);
xor U1067 (N_1067,N_877,N_775);
and U1068 (N_1068,N_265,N_664);
and U1069 (N_1069,N_153,N_958);
nor U1070 (N_1070,N_528,N_658);
nor U1071 (N_1071,N_454,N_362);
or U1072 (N_1072,N_175,N_123);
nand U1073 (N_1073,N_156,N_273);
and U1074 (N_1074,N_531,N_169);
nand U1075 (N_1075,N_77,N_6);
nand U1076 (N_1076,N_600,N_889);
and U1077 (N_1077,N_592,N_229);
xnor U1078 (N_1078,N_828,N_248);
nand U1079 (N_1079,N_366,N_612);
nor U1080 (N_1080,N_168,N_632);
nand U1081 (N_1081,N_872,N_891);
or U1082 (N_1082,N_371,N_227);
xnor U1083 (N_1083,N_416,N_176);
or U1084 (N_1084,N_368,N_66);
nand U1085 (N_1085,N_40,N_332);
nor U1086 (N_1086,N_88,N_903);
or U1087 (N_1087,N_840,N_337);
nand U1088 (N_1088,N_946,N_319);
nor U1089 (N_1089,N_101,N_560);
nand U1090 (N_1090,N_323,N_349);
xor U1091 (N_1091,N_293,N_718);
and U1092 (N_1092,N_786,N_228);
nor U1093 (N_1093,N_46,N_996);
or U1094 (N_1094,N_675,N_799);
and U1095 (N_1095,N_342,N_753);
nor U1096 (N_1096,N_730,N_198);
nand U1097 (N_1097,N_484,N_955);
or U1098 (N_1098,N_225,N_757);
and U1099 (N_1099,N_688,N_556);
xor U1100 (N_1100,N_458,N_778);
xnor U1101 (N_1101,N_213,N_513);
and U1102 (N_1102,N_173,N_33);
nand U1103 (N_1103,N_69,N_617);
or U1104 (N_1104,N_83,N_405);
nand U1105 (N_1105,N_686,N_219);
nor U1106 (N_1106,N_682,N_550);
nand U1107 (N_1107,N_385,N_258);
or U1108 (N_1108,N_240,N_28);
or U1109 (N_1109,N_770,N_47);
or U1110 (N_1110,N_609,N_271);
nand U1111 (N_1111,N_546,N_247);
nor U1112 (N_1112,N_719,N_691);
and U1113 (N_1113,N_952,N_482);
and U1114 (N_1114,N_341,N_21);
and U1115 (N_1115,N_24,N_976);
nor U1116 (N_1116,N_328,N_915);
and U1117 (N_1117,N_926,N_774);
and U1118 (N_1118,N_914,N_305);
nor U1119 (N_1119,N_284,N_870);
nand U1120 (N_1120,N_335,N_127);
nor U1121 (N_1121,N_871,N_485);
nand U1122 (N_1122,N_504,N_802);
xnor U1123 (N_1123,N_875,N_852);
or U1124 (N_1124,N_433,N_487);
nor U1125 (N_1125,N_367,N_966);
nor U1126 (N_1126,N_880,N_890);
nand U1127 (N_1127,N_950,N_204);
and U1128 (N_1128,N_160,N_251);
nor U1129 (N_1129,N_876,N_673);
and U1130 (N_1130,N_421,N_288);
and U1131 (N_1131,N_885,N_155);
xnor U1132 (N_1132,N_768,N_707);
or U1133 (N_1133,N_187,N_99);
nand U1134 (N_1134,N_325,N_361);
and U1135 (N_1135,N_529,N_703);
xor U1136 (N_1136,N_315,N_826);
or U1137 (N_1137,N_920,N_252);
nor U1138 (N_1138,N_733,N_943);
nor U1139 (N_1139,N_708,N_312);
nor U1140 (N_1140,N_45,N_320);
nand U1141 (N_1141,N_769,N_585);
and U1142 (N_1142,N_343,N_742);
or U1143 (N_1143,N_723,N_436);
and U1144 (N_1144,N_476,N_820);
and U1145 (N_1145,N_684,N_731);
nor U1146 (N_1146,N_773,N_186);
and U1147 (N_1147,N_166,N_359);
nand U1148 (N_1148,N_189,N_179);
nand U1149 (N_1149,N_784,N_525);
and U1150 (N_1150,N_503,N_566);
and U1151 (N_1151,N_264,N_306);
nand U1152 (N_1152,N_721,N_308);
and U1153 (N_1153,N_406,N_986);
or U1154 (N_1154,N_126,N_953);
and U1155 (N_1155,N_110,N_594);
nor U1156 (N_1156,N_805,N_711);
and U1157 (N_1157,N_388,N_64);
nand U1158 (N_1158,N_418,N_591);
and U1159 (N_1159,N_188,N_972);
and U1160 (N_1160,N_896,N_102);
and U1161 (N_1161,N_118,N_779);
or U1162 (N_1162,N_364,N_317);
or U1163 (N_1163,N_641,N_230);
and U1164 (N_1164,N_981,N_593);
nor U1165 (N_1165,N_146,N_279);
and U1166 (N_1166,N_409,N_389);
nand U1167 (N_1167,N_130,N_382);
nand U1168 (N_1168,N_62,N_739);
nand U1169 (N_1169,N_158,N_689);
nor U1170 (N_1170,N_859,N_475);
and U1171 (N_1171,N_700,N_631);
nor U1172 (N_1172,N_855,N_242);
xnor U1173 (N_1173,N_849,N_4);
nor U1174 (N_1174,N_509,N_378);
nand U1175 (N_1175,N_547,N_401);
nor U1176 (N_1176,N_7,N_899);
nand U1177 (N_1177,N_91,N_874);
and U1178 (N_1178,N_373,N_755);
and U1179 (N_1179,N_676,N_43);
nor U1180 (N_1180,N_627,N_333);
or U1181 (N_1181,N_355,N_125);
and U1182 (N_1182,N_745,N_172);
or U1183 (N_1183,N_449,N_104);
nor U1184 (N_1184,N_109,N_789);
nor U1185 (N_1185,N_912,N_23);
nor U1186 (N_1186,N_842,N_656);
nor U1187 (N_1187,N_70,N_595);
or U1188 (N_1188,N_68,N_788);
nand U1189 (N_1189,N_465,N_202);
nand U1190 (N_1190,N_250,N_660);
and U1191 (N_1191,N_390,N_426);
or U1192 (N_1192,N_865,N_846);
nand U1193 (N_1193,N_951,N_14);
and U1194 (N_1194,N_663,N_338);
and U1195 (N_1195,N_259,N_148);
and U1196 (N_1196,N_931,N_938);
or U1197 (N_1197,N_897,N_506);
nand U1198 (N_1198,N_444,N_224);
or U1199 (N_1199,N_997,N_954);
and U1200 (N_1200,N_422,N_647);
or U1201 (N_1201,N_968,N_274);
or U1202 (N_1202,N_984,N_821);
nand U1203 (N_1203,N_751,N_25);
or U1204 (N_1204,N_470,N_324);
nor U1205 (N_1205,N_336,N_806);
nand U1206 (N_1206,N_736,N_443);
nor U1207 (N_1207,N_214,N_944);
or U1208 (N_1208,N_508,N_149);
or U1209 (N_1209,N_44,N_906);
and U1210 (N_1210,N_603,N_212);
and U1211 (N_1211,N_354,N_911);
and U1212 (N_1212,N_134,N_398);
or U1213 (N_1213,N_128,N_63);
and U1214 (N_1214,N_695,N_266);
xor U1215 (N_1215,N_297,N_630);
nor U1216 (N_1216,N_394,N_86);
nor U1217 (N_1217,N_861,N_568);
nor U1218 (N_1218,N_758,N_139);
and U1219 (N_1219,N_183,N_512);
nor U1220 (N_1220,N_50,N_777);
nand U1221 (N_1221,N_832,N_613);
nand U1222 (N_1222,N_481,N_446);
and U1223 (N_1223,N_881,N_434);
nor U1224 (N_1224,N_119,N_479);
nor U1225 (N_1225,N_921,N_165);
nand U1226 (N_1226,N_793,N_296);
nand U1227 (N_1227,N_794,N_625);
and U1228 (N_1228,N_243,N_704);
or U1229 (N_1229,N_108,N_716);
nand U1230 (N_1230,N_554,N_321);
and U1231 (N_1231,N_440,N_544);
nor U1232 (N_1232,N_956,N_725);
xnor U1233 (N_1233,N_606,N_729);
nor U1234 (N_1234,N_249,N_959);
nand U1235 (N_1235,N_732,N_215);
xnor U1236 (N_1236,N_830,N_524);
nor U1237 (N_1237,N_575,N_211);
nand U1238 (N_1238,N_636,N_490);
xor U1239 (N_1239,N_532,N_451);
xnor U1240 (N_1240,N_559,N_671);
and U1241 (N_1241,N_239,N_231);
xor U1242 (N_1242,N_935,N_590);
nand U1243 (N_1243,N_163,N_919);
and U1244 (N_1244,N_898,N_930);
nor U1245 (N_1245,N_942,N_304);
nor U1246 (N_1246,N_635,N_626);
and U1247 (N_1247,N_665,N_38);
nor U1248 (N_1248,N_882,N_587);
nand U1249 (N_1249,N_49,N_601);
or U1250 (N_1250,N_650,N_979);
or U1251 (N_1251,N_20,N_245);
and U1252 (N_1252,N_790,N_218);
and U1253 (N_1253,N_42,N_838);
nor U1254 (N_1254,N_420,N_697);
nor U1255 (N_1255,N_391,N_275);
and U1256 (N_1256,N_761,N_494);
xor U1257 (N_1257,N_510,N_17);
nor U1258 (N_1258,N_637,N_493);
and U1259 (N_1259,N_92,N_403);
or U1260 (N_1260,N_619,N_991);
or U1261 (N_1261,N_940,N_498);
and U1262 (N_1262,N_344,N_100);
nand U1263 (N_1263,N_55,N_463);
nand U1264 (N_1264,N_58,N_184);
xnor U1265 (N_1265,N_588,N_140);
and U1266 (N_1266,N_151,N_696);
nand U1267 (N_1267,N_299,N_542);
nor U1268 (N_1268,N_582,N_621);
and U1269 (N_1269,N_693,N_11);
and U1270 (N_1270,N_357,N_379);
nand U1271 (N_1271,N_978,N_563);
or U1272 (N_1272,N_37,N_61);
or U1273 (N_1273,N_869,N_862);
xnor U1274 (N_1274,N_765,N_386);
or U1275 (N_1275,N_53,N_276);
nor U1276 (N_1276,N_447,N_272);
nand U1277 (N_1277,N_347,N_90);
xnor U1278 (N_1278,N_659,N_428);
or U1279 (N_1279,N_372,N_644);
and U1280 (N_1280,N_103,N_331);
or U1281 (N_1281,N_486,N_238);
xor U1282 (N_1282,N_269,N_84);
and U1283 (N_1283,N_268,N_87);
xnor U1284 (N_1284,N_505,N_145);
and U1285 (N_1285,N_904,N_285);
and U1286 (N_1286,N_462,N_760);
nand U1287 (N_1287,N_990,N_234);
and U1288 (N_1288,N_34,N_201);
nand U1289 (N_1289,N_819,N_737);
nand U1290 (N_1290,N_822,N_280);
nand U1291 (N_1291,N_75,N_190);
xnor U1292 (N_1292,N_501,N_286);
or U1293 (N_1293,N_622,N_907);
xor U1294 (N_1294,N_967,N_474);
nor U1295 (N_1295,N_995,N_517);
xnor U1296 (N_1296,N_642,N_724);
or U1297 (N_1297,N_262,N_666);
xnor U1298 (N_1298,N_750,N_132);
nand U1299 (N_1299,N_80,N_199);
nand U1300 (N_1300,N_801,N_518);
nand U1301 (N_1301,N_460,N_316);
nor U1302 (N_1302,N_977,N_713);
or U1303 (N_1303,N_455,N_973);
and U1304 (N_1304,N_878,N_516);
and U1305 (N_1305,N_633,N_301);
nor U1306 (N_1306,N_150,N_298);
nand U1307 (N_1307,N_496,N_569);
nand U1308 (N_1308,N_407,N_112);
nor U1309 (N_1309,N_363,N_314);
and U1310 (N_1310,N_927,N_0);
nand U1311 (N_1311,N_471,N_795);
and U1312 (N_1312,N_491,N_530);
xor U1313 (N_1313,N_12,N_384);
nor U1314 (N_1314,N_60,N_749);
or U1315 (N_1315,N_624,N_669);
nor U1316 (N_1316,N_685,N_310);
xnor U1317 (N_1317,N_937,N_432);
nor U1318 (N_1318,N_771,N_690);
and U1319 (N_1319,N_397,N_856);
nand U1320 (N_1320,N_415,N_759);
nand U1321 (N_1321,N_847,N_929);
or U1322 (N_1322,N_216,N_255);
nand U1323 (N_1323,N_161,N_346);
nand U1324 (N_1324,N_431,N_205);
and U1325 (N_1325,N_653,N_71);
xor U1326 (N_1326,N_277,N_81);
and U1327 (N_1327,N_152,N_515);
xor U1328 (N_1328,N_791,N_507);
xor U1329 (N_1329,N_345,N_597);
nand U1330 (N_1330,N_616,N_610);
nand U1331 (N_1331,N_971,N_226);
and U1332 (N_1332,N_987,N_191);
nor U1333 (N_1333,N_135,N_452);
nor U1334 (N_1334,N_468,N_947);
or U1335 (N_1335,N_598,N_369);
nand U1336 (N_1336,N_300,N_72);
nand U1337 (N_1337,N_834,N_185);
or U1338 (N_1338,N_640,N_143);
or U1339 (N_1339,N_360,N_477);
and U1340 (N_1340,N_65,N_787);
nor U1341 (N_1341,N_776,N_52);
nor U1342 (N_1342,N_808,N_925);
nand U1343 (N_1343,N_888,N_93);
nand U1344 (N_1344,N_519,N_147);
or U1345 (N_1345,N_829,N_677);
or U1346 (N_1346,N_467,N_537);
xor U1347 (N_1347,N_327,N_543);
nor U1348 (N_1348,N_283,N_845);
or U1349 (N_1349,N_705,N_197);
nand U1350 (N_1350,N_10,N_767);
and U1351 (N_1351,N_772,N_895);
nor U1352 (N_1352,N_553,N_76);
nand U1353 (N_1353,N_961,N_608);
xor U1354 (N_1354,N_540,N_117);
xor U1355 (N_1355,N_983,N_699);
or U1356 (N_1356,N_3,N_918);
or U1357 (N_1357,N_445,N_709);
or U1358 (N_1358,N_27,N_651);
nand U1359 (N_1359,N_162,N_901);
and U1360 (N_1360,N_2,N_375);
and U1361 (N_1361,N_994,N_628);
nand U1362 (N_1362,N_561,N_965);
nor U1363 (N_1363,N_567,N_263);
or U1364 (N_1364,N_115,N_419);
and U1365 (N_1365,N_48,N_221);
or U1366 (N_1366,N_863,N_339);
nand U1367 (N_1367,N_923,N_648);
or U1368 (N_1368,N_311,N_495);
nor U1369 (N_1369,N_256,N_195);
nand U1370 (N_1370,N_67,N_79);
nor U1371 (N_1371,N_583,N_545);
nor U1372 (N_1372,N_464,N_356);
xor U1373 (N_1373,N_909,N_535);
nor U1374 (N_1374,N_111,N_121);
and U1375 (N_1375,N_710,N_917);
or U1376 (N_1376,N_287,N_370);
or U1377 (N_1377,N_222,N_844);
or U1378 (N_1378,N_330,N_141);
nand U1379 (N_1379,N_348,N_313);
nor U1380 (N_1380,N_351,N_174);
or U1381 (N_1381,N_82,N_818);
nand U1382 (N_1382,N_469,N_281);
nand U1383 (N_1383,N_380,N_107);
and U1384 (N_1384,N_781,N_1);
and U1385 (N_1385,N_634,N_657);
and U1386 (N_1386,N_365,N_393);
and U1387 (N_1387,N_998,N_435);
nand U1388 (N_1388,N_873,N_377);
nand U1389 (N_1389,N_497,N_96);
nand U1390 (N_1390,N_13,N_715);
xor U1391 (N_1391,N_499,N_387);
and U1392 (N_1392,N_933,N_548);
or U1393 (N_1393,N_576,N_902);
and U1394 (N_1394,N_734,N_294);
or U1395 (N_1395,N_578,N_244);
or U1396 (N_1396,N_209,N_924);
nor U1397 (N_1397,N_980,N_934);
or U1398 (N_1398,N_738,N_629);
nor U1399 (N_1399,N_74,N_15);
nand U1400 (N_1400,N_536,N_605);
nand U1401 (N_1401,N_827,N_410);
and U1402 (N_1402,N_480,N_520);
xor U1403 (N_1403,N_900,N_687);
nand U1404 (N_1404,N_932,N_551);
or U1405 (N_1405,N_810,N_260);
nand U1406 (N_1406,N_989,N_136);
or U1407 (N_1407,N_584,N_522);
nand U1408 (N_1408,N_124,N_607);
nand U1409 (N_1409,N_831,N_853);
nor U1410 (N_1410,N_399,N_208);
nand U1411 (N_1411,N_241,N_645);
nand U1412 (N_1412,N_22,N_803);
nor U1413 (N_1413,N_670,N_735);
or U1414 (N_1414,N_565,N_623);
and U1415 (N_1415,N_97,N_620);
and U1416 (N_1416,N_427,N_960);
and U1417 (N_1417,N_639,N_541);
nor U1418 (N_1418,N_246,N_860);
or U1419 (N_1419,N_171,N_714);
nand U1420 (N_1420,N_596,N_200);
nand U1421 (N_1421,N_105,N_823);
nor U1422 (N_1422,N_180,N_866);
nand U1423 (N_1423,N_746,N_804);
and U1424 (N_1424,N_580,N_975);
nand U1425 (N_1425,N_192,N_120);
or U1426 (N_1426,N_586,N_51);
nand U1427 (N_1427,N_492,N_783);
nor U1428 (N_1428,N_712,N_129);
nand U1429 (N_1429,N_41,N_295);
and U1430 (N_1430,N_589,N_523);
and U1431 (N_1431,N_456,N_131);
nor U1432 (N_1432,N_615,N_178);
nand U1433 (N_1433,N_114,N_754);
nand U1434 (N_1434,N_29,N_309);
and U1435 (N_1435,N_599,N_552);
nor U1436 (N_1436,N_235,N_329);
or U1437 (N_1437,N_570,N_425);
nor U1438 (N_1438,N_868,N_437);
nand U1439 (N_1439,N_638,N_59);
nand U1440 (N_1440,N_448,N_89);
nor U1441 (N_1441,N_800,N_835);
nor U1442 (N_1442,N_253,N_655);
and U1443 (N_1443,N_413,N_646);
xnor U1444 (N_1444,N_98,N_307);
nor U1445 (N_1445,N_812,N_957);
nor U1446 (N_1446,N_526,N_892);
nor U1447 (N_1447,N_747,N_833);
or U1448 (N_1448,N_913,N_702);
nand U1449 (N_1449,N_539,N_809);
and U1450 (N_1450,N_992,N_555);
and U1451 (N_1451,N_916,N_322);
or U1452 (N_1452,N_905,N_722);
or U1453 (N_1453,N_611,N_381);
nor U1454 (N_1454,N_843,N_16);
nand U1455 (N_1455,N_181,N_194);
nand U1456 (N_1456,N_170,N_740);
nor U1457 (N_1457,N_392,N_429);
and U1458 (N_1458,N_122,N_962);
nor U1459 (N_1459,N_439,N_681);
nand U1460 (N_1460,N_837,N_159);
or U1461 (N_1461,N_5,N_203);
nor U1462 (N_1462,N_883,N_39);
nand U1463 (N_1463,N_668,N_267);
xor U1464 (N_1464,N_303,N_807);
or U1465 (N_1465,N_887,N_726);
nor U1466 (N_1466,N_106,N_167);
or U1467 (N_1467,N_936,N_928);
xnor U1468 (N_1468,N_182,N_352);
nand U1469 (N_1469,N_797,N_113);
nand U1470 (N_1470,N_527,N_574);
nor U1471 (N_1471,N_661,N_9);
nor U1472 (N_1472,N_654,N_867);
nor U1473 (N_1473,N_326,N_533);
and U1474 (N_1474,N_815,N_138);
xnor U1475 (N_1475,N_232,N_652);
or U1476 (N_1476,N_412,N_154);
nor U1477 (N_1477,N_254,N_692);
nand U1478 (N_1478,N_423,N_8);
and U1479 (N_1479,N_766,N_334);
nor U1480 (N_1480,N_35,N_453);
nor U1481 (N_1481,N_36,N_350);
or U1482 (N_1482,N_142,N_396);
nor U1483 (N_1483,N_26,N_848);
nand U1484 (N_1484,N_30,N_206);
or U1485 (N_1485,N_478,N_358);
and U1486 (N_1486,N_764,N_939);
xnor U1487 (N_1487,N_521,N_210);
nand U1488 (N_1488,N_57,N_850);
and U1489 (N_1489,N_782,N_489);
or U1490 (N_1490,N_698,N_993);
nand U1491 (N_1491,N_672,N_756);
and U1492 (N_1492,N_73,N_752);
or U1493 (N_1493,N_970,N_643);
nor U1494 (N_1494,N_614,N_95);
nand U1495 (N_1495,N_472,N_879);
nand U1496 (N_1496,N_442,N_571);
and U1497 (N_1497,N_796,N_374);
and U1498 (N_1498,N_538,N_438);
nor U1499 (N_1499,N_557,N_562);
and U1500 (N_1500,N_101,N_895);
nor U1501 (N_1501,N_57,N_375);
nor U1502 (N_1502,N_918,N_393);
nand U1503 (N_1503,N_487,N_903);
nor U1504 (N_1504,N_29,N_903);
and U1505 (N_1505,N_95,N_534);
or U1506 (N_1506,N_446,N_695);
and U1507 (N_1507,N_721,N_948);
nor U1508 (N_1508,N_916,N_832);
nor U1509 (N_1509,N_896,N_166);
nor U1510 (N_1510,N_418,N_871);
or U1511 (N_1511,N_381,N_345);
nand U1512 (N_1512,N_541,N_185);
and U1513 (N_1513,N_699,N_769);
or U1514 (N_1514,N_710,N_952);
and U1515 (N_1515,N_655,N_897);
nand U1516 (N_1516,N_183,N_549);
nand U1517 (N_1517,N_227,N_749);
nand U1518 (N_1518,N_70,N_787);
or U1519 (N_1519,N_614,N_339);
nand U1520 (N_1520,N_620,N_887);
nand U1521 (N_1521,N_10,N_677);
and U1522 (N_1522,N_618,N_35);
or U1523 (N_1523,N_111,N_910);
xor U1524 (N_1524,N_831,N_528);
nor U1525 (N_1525,N_966,N_80);
nor U1526 (N_1526,N_261,N_867);
or U1527 (N_1527,N_102,N_987);
or U1528 (N_1528,N_77,N_878);
nand U1529 (N_1529,N_254,N_593);
nor U1530 (N_1530,N_511,N_505);
nor U1531 (N_1531,N_722,N_541);
nand U1532 (N_1532,N_821,N_369);
or U1533 (N_1533,N_40,N_190);
nand U1534 (N_1534,N_457,N_814);
or U1535 (N_1535,N_659,N_909);
or U1536 (N_1536,N_69,N_311);
and U1537 (N_1537,N_427,N_159);
and U1538 (N_1538,N_239,N_286);
nor U1539 (N_1539,N_186,N_339);
xnor U1540 (N_1540,N_197,N_912);
or U1541 (N_1541,N_163,N_36);
nand U1542 (N_1542,N_176,N_982);
and U1543 (N_1543,N_201,N_604);
and U1544 (N_1544,N_435,N_470);
and U1545 (N_1545,N_229,N_962);
and U1546 (N_1546,N_569,N_532);
or U1547 (N_1547,N_392,N_782);
and U1548 (N_1548,N_36,N_818);
and U1549 (N_1549,N_403,N_779);
or U1550 (N_1550,N_904,N_333);
nand U1551 (N_1551,N_904,N_813);
or U1552 (N_1552,N_583,N_521);
nand U1553 (N_1553,N_149,N_272);
and U1554 (N_1554,N_125,N_170);
nor U1555 (N_1555,N_202,N_408);
or U1556 (N_1556,N_218,N_639);
and U1557 (N_1557,N_554,N_46);
or U1558 (N_1558,N_390,N_225);
or U1559 (N_1559,N_736,N_412);
nand U1560 (N_1560,N_41,N_731);
xor U1561 (N_1561,N_745,N_729);
nor U1562 (N_1562,N_111,N_582);
nand U1563 (N_1563,N_198,N_775);
and U1564 (N_1564,N_703,N_945);
nand U1565 (N_1565,N_539,N_287);
and U1566 (N_1566,N_17,N_37);
xnor U1567 (N_1567,N_866,N_956);
nand U1568 (N_1568,N_17,N_699);
nor U1569 (N_1569,N_0,N_366);
and U1570 (N_1570,N_827,N_810);
xor U1571 (N_1571,N_626,N_43);
or U1572 (N_1572,N_720,N_269);
and U1573 (N_1573,N_938,N_562);
nor U1574 (N_1574,N_18,N_180);
or U1575 (N_1575,N_495,N_220);
nand U1576 (N_1576,N_530,N_600);
nand U1577 (N_1577,N_496,N_377);
nand U1578 (N_1578,N_42,N_837);
nor U1579 (N_1579,N_526,N_116);
nor U1580 (N_1580,N_25,N_655);
nand U1581 (N_1581,N_380,N_619);
or U1582 (N_1582,N_800,N_528);
or U1583 (N_1583,N_23,N_397);
xnor U1584 (N_1584,N_294,N_259);
or U1585 (N_1585,N_485,N_197);
nand U1586 (N_1586,N_300,N_874);
nor U1587 (N_1587,N_360,N_550);
or U1588 (N_1588,N_636,N_500);
nor U1589 (N_1589,N_423,N_95);
nor U1590 (N_1590,N_163,N_798);
or U1591 (N_1591,N_261,N_912);
and U1592 (N_1592,N_260,N_11);
and U1593 (N_1593,N_801,N_13);
xor U1594 (N_1594,N_923,N_798);
xnor U1595 (N_1595,N_765,N_183);
and U1596 (N_1596,N_843,N_45);
and U1597 (N_1597,N_426,N_396);
and U1598 (N_1598,N_364,N_524);
nor U1599 (N_1599,N_716,N_34);
nand U1600 (N_1600,N_66,N_63);
nor U1601 (N_1601,N_519,N_126);
nand U1602 (N_1602,N_564,N_731);
nand U1603 (N_1603,N_134,N_976);
nor U1604 (N_1604,N_134,N_961);
or U1605 (N_1605,N_274,N_803);
and U1606 (N_1606,N_875,N_211);
or U1607 (N_1607,N_523,N_119);
and U1608 (N_1608,N_240,N_845);
xor U1609 (N_1609,N_825,N_454);
nor U1610 (N_1610,N_334,N_151);
nor U1611 (N_1611,N_428,N_142);
or U1612 (N_1612,N_484,N_467);
and U1613 (N_1613,N_963,N_13);
xnor U1614 (N_1614,N_775,N_127);
nand U1615 (N_1615,N_220,N_355);
and U1616 (N_1616,N_295,N_216);
or U1617 (N_1617,N_939,N_85);
and U1618 (N_1618,N_577,N_907);
nand U1619 (N_1619,N_283,N_823);
and U1620 (N_1620,N_448,N_772);
and U1621 (N_1621,N_104,N_688);
nand U1622 (N_1622,N_294,N_64);
nor U1623 (N_1623,N_476,N_487);
nor U1624 (N_1624,N_193,N_276);
nand U1625 (N_1625,N_297,N_471);
and U1626 (N_1626,N_351,N_418);
or U1627 (N_1627,N_46,N_89);
nand U1628 (N_1628,N_231,N_909);
and U1629 (N_1629,N_763,N_654);
or U1630 (N_1630,N_794,N_45);
nor U1631 (N_1631,N_839,N_468);
and U1632 (N_1632,N_838,N_771);
nand U1633 (N_1633,N_576,N_676);
nand U1634 (N_1634,N_459,N_546);
or U1635 (N_1635,N_974,N_242);
xnor U1636 (N_1636,N_780,N_219);
or U1637 (N_1637,N_734,N_142);
nand U1638 (N_1638,N_425,N_166);
and U1639 (N_1639,N_111,N_215);
or U1640 (N_1640,N_474,N_104);
nor U1641 (N_1641,N_743,N_910);
or U1642 (N_1642,N_138,N_698);
or U1643 (N_1643,N_696,N_431);
or U1644 (N_1644,N_919,N_683);
nand U1645 (N_1645,N_358,N_486);
or U1646 (N_1646,N_589,N_38);
nor U1647 (N_1647,N_149,N_866);
nand U1648 (N_1648,N_998,N_454);
or U1649 (N_1649,N_769,N_971);
xnor U1650 (N_1650,N_850,N_638);
or U1651 (N_1651,N_280,N_41);
xor U1652 (N_1652,N_769,N_624);
and U1653 (N_1653,N_564,N_808);
and U1654 (N_1654,N_989,N_898);
nand U1655 (N_1655,N_234,N_231);
and U1656 (N_1656,N_474,N_106);
nor U1657 (N_1657,N_462,N_794);
and U1658 (N_1658,N_744,N_400);
or U1659 (N_1659,N_807,N_313);
or U1660 (N_1660,N_218,N_870);
xnor U1661 (N_1661,N_365,N_498);
and U1662 (N_1662,N_155,N_402);
nor U1663 (N_1663,N_11,N_854);
nor U1664 (N_1664,N_587,N_415);
or U1665 (N_1665,N_86,N_160);
nor U1666 (N_1666,N_137,N_135);
xnor U1667 (N_1667,N_947,N_741);
and U1668 (N_1668,N_854,N_686);
xor U1669 (N_1669,N_666,N_128);
or U1670 (N_1670,N_182,N_952);
nand U1671 (N_1671,N_502,N_89);
and U1672 (N_1672,N_839,N_699);
and U1673 (N_1673,N_642,N_407);
nor U1674 (N_1674,N_325,N_247);
nor U1675 (N_1675,N_96,N_332);
and U1676 (N_1676,N_747,N_226);
and U1677 (N_1677,N_173,N_693);
or U1678 (N_1678,N_292,N_874);
and U1679 (N_1679,N_46,N_737);
and U1680 (N_1680,N_310,N_574);
nand U1681 (N_1681,N_673,N_433);
nor U1682 (N_1682,N_519,N_461);
nand U1683 (N_1683,N_768,N_620);
nand U1684 (N_1684,N_434,N_759);
or U1685 (N_1685,N_687,N_912);
and U1686 (N_1686,N_682,N_383);
or U1687 (N_1687,N_624,N_402);
or U1688 (N_1688,N_572,N_664);
or U1689 (N_1689,N_561,N_859);
xnor U1690 (N_1690,N_212,N_732);
and U1691 (N_1691,N_657,N_86);
xnor U1692 (N_1692,N_365,N_123);
xor U1693 (N_1693,N_137,N_229);
xor U1694 (N_1694,N_605,N_402);
xor U1695 (N_1695,N_94,N_948);
and U1696 (N_1696,N_574,N_965);
nand U1697 (N_1697,N_630,N_38);
and U1698 (N_1698,N_926,N_499);
and U1699 (N_1699,N_843,N_354);
or U1700 (N_1700,N_196,N_566);
or U1701 (N_1701,N_892,N_360);
and U1702 (N_1702,N_319,N_535);
or U1703 (N_1703,N_718,N_128);
and U1704 (N_1704,N_748,N_812);
xor U1705 (N_1705,N_756,N_910);
nand U1706 (N_1706,N_523,N_629);
nor U1707 (N_1707,N_510,N_315);
nor U1708 (N_1708,N_762,N_257);
xnor U1709 (N_1709,N_714,N_856);
nand U1710 (N_1710,N_290,N_318);
nand U1711 (N_1711,N_17,N_766);
and U1712 (N_1712,N_45,N_704);
or U1713 (N_1713,N_464,N_938);
or U1714 (N_1714,N_144,N_260);
and U1715 (N_1715,N_424,N_834);
nor U1716 (N_1716,N_155,N_35);
and U1717 (N_1717,N_897,N_266);
nand U1718 (N_1718,N_75,N_548);
and U1719 (N_1719,N_32,N_578);
nor U1720 (N_1720,N_295,N_982);
or U1721 (N_1721,N_721,N_243);
xnor U1722 (N_1722,N_226,N_593);
nand U1723 (N_1723,N_839,N_550);
and U1724 (N_1724,N_445,N_400);
or U1725 (N_1725,N_299,N_763);
nor U1726 (N_1726,N_767,N_989);
nor U1727 (N_1727,N_646,N_895);
nand U1728 (N_1728,N_465,N_191);
or U1729 (N_1729,N_248,N_687);
or U1730 (N_1730,N_396,N_943);
and U1731 (N_1731,N_624,N_352);
nand U1732 (N_1732,N_1,N_579);
nor U1733 (N_1733,N_213,N_607);
or U1734 (N_1734,N_852,N_148);
and U1735 (N_1735,N_65,N_503);
nand U1736 (N_1736,N_358,N_936);
nand U1737 (N_1737,N_216,N_701);
nor U1738 (N_1738,N_955,N_17);
nor U1739 (N_1739,N_417,N_956);
or U1740 (N_1740,N_936,N_988);
xnor U1741 (N_1741,N_475,N_162);
and U1742 (N_1742,N_168,N_339);
nand U1743 (N_1743,N_210,N_433);
nand U1744 (N_1744,N_191,N_98);
and U1745 (N_1745,N_807,N_281);
and U1746 (N_1746,N_332,N_428);
and U1747 (N_1747,N_486,N_986);
xnor U1748 (N_1748,N_220,N_405);
nand U1749 (N_1749,N_391,N_576);
nor U1750 (N_1750,N_217,N_221);
nor U1751 (N_1751,N_688,N_694);
nor U1752 (N_1752,N_975,N_928);
xor U1753 (N_1753,N_103,N_371);
xnor U1754 (N_1754,N_87,N_107);
and U1755 (N_1755,N_664,N_331);
xnor U1756 (N_1756,N_731,N_674);
nor U1757 (N_1757,N_494,N_830);
nor U1758 (N_1758,N_323,N_511);
nor U1759 (N_1759,N_659,N_10);
nand U1760 (N_1760,N_654,N_287);
xor U1761 (N_1761,N_978,N_575);
xor U1762 (N_1762,N_888,N_649);
nand U1763 (N_1763,N_121,N_291);
nand U1764 (N_1764,N_961,N_287);
and U1765 (N_1765,N_966,N_694);
and U1766 (N_1766,N_246,N_269);
xor U1767 (N_1767,N_554,N_89);
nand U1768 (N_1768,N_62,N_378);
or U1769 (N_1769,N_413,N_94);
and U1770 (N_1770,N_716,N_797);
or U1771 (N_1771,N_764,N_712);
xnor U1772 (N_1772,N_333,N_704);
nand U1773 (N_1773,N_395,N_10);
and U1774 (N_1774,N_143,N_249);
nand U1775 (N_1775,N_870,N_181);
xor U1776 (N_1776,N_531,N_731);
and U1777 (N_1777,N_660,N_847);
xor U1778 (N_1778,N_261,N_673);
or U1779 (N_1779,N_942,N_732);
and U1780 (N_1780,N_195,N_270);
nor U1781 (N_1781,N_13,N_923);
nor U1782 (N_1782,N_728,N_698);
nor U1783 (N_1783,N_306,N_370);
or U1784 (N_1784,N_866,N_110);
nand U1785 (N_1785,N_427,N_186);
and U1786 (N_1786,N_924,N_351);
or U1787 (N_1787,N_491,N_926);
nor U1788 (N_1788,N_817,N_639);
xnor U1789 (N_1789,N_966,N_645);
xnor U1790 (N_1790,N_781,N_249);
or U1791 (N_1791,N_426,N_981);
nor U1792 (N_1792,N_590,N_473);
nor U1793 (N_1793,N_163,N_803);
nand U1794 (N_1794,N_819,N_194);
and U1795 (N_1795,N_607,N_646);
or U1796 (N_1796,N_871,N_393);
and U1797 (N_1797,N_634,N_190);
or U1798 (N_1798,N_294,N_828);
or U1799 (N_1799,N_357,N_951);
or U1800 (N_1800,N_835,N_153);
nand U1801 (N_1801,N_176,N_303);
and U1802 (N_1802,N_840,N_488);
nor U1803 (N_1803,N_753,N_295);
xnor U1804 (N_1804,N_236,N_265);
nor U1805 (N_1805,N_662,N_863);
and U1806 (N_1806,N_563,N_949);
xor U1807 (N_1807,N_562,N_387);
nor U1808 (N_1808,N_420,N_458);
or U1809 (N_1809,N_520,N_529);
xnor U1810 (N_1810,N_419,N_634);
nor U1811 (N_1811,N_216,N_624);
and U1812 (N_1812,N_450,N_690);
nor U1813 (N_1813,N_624,N_215);
or U1814 (N_1814,N_451,N_77);
and U1815 (N_1815,N_880,N_621);
or U1816 (N_1816,N_459,N_150);
nand U1817 (N_1817,N_169,N_339);
nand U1818 (N_1818,N_61,N_730);
nand U1819 (N_1819,N_790,N_906);
and U1820 (N_1820,N_75,N_608);
nand U1821 (N_1821,N_545,N_566);
nor U1822 (N_1822,N_633,N_915);
nand U1823 (N_1823,N_416,N_952);
or U1824 (N_1824,N_131,N_861);
nor U1825 (N_1825,N_739,N_896);
or U1826 (N_1826,N_883,N_73);
or U1827 (N_1827,N_270,N_887);
nand U1828 (N_1828,N_628,N_273);
nor U1829 (N_1829,N_484,N_13);
nand U1830 (N_1830,N_50,N_861);
or U1831 (N_1831,N_969,N_123);
and U1832 (N_1832,N_383,N_45);
xnor U1833 (N_1833,N_406,N_962);
nand U1834 (N_1834,N_654,N_48);
nor U1835 (N_1835,N_524,N_995);
nand U1836 (N_1836,N_291,N_360);
and U1837 (N_1837,N_456,N_212);
and U1838 (N_1838,N_499,N_424);
nor U1839 (N_1839,N_507,N_648);
and U1840 (N_1840,N_353,N_880);
xor U1841 (N_1841,N_241,N_269);
and U1842 (N_1842,N_756,N_860);
nor U1843 (N_1843,N_665,N_286);
nor U1844 (N_1844,N_763,N_933);
and U1845 (N_1845,N_308,N_347);
nand U1846 (N_1846,N_973,N_407);
or U1847 (N_1847,N_570,N_513);
nand U1848 (N_1848,N_921,N_60);
or U1849 (N_1849,N_100,N_860);
and U1850 (N_1850,N_454,N_732);
nor U1851 (N_1851,N_538,N_976);
nor U1852 (N_1852,N_267,N_285);
nand U1853 (N_1853,N_142,N_936);
nand U1854 (N_1854,N_873,N_376);
nor U1855 (N_1855,N_43,N_193);
nand U1856 (N_1856,N_495,N_769);
nor U1857 (N_1857,N_35,N_801);
nand U1858 (N_1858,N_243,N_611);
and U1859 (N_1859,N_528,N_984);
and U1860 (N_1860,N_84,N_81);
xnor U1861 (N_1861,N_173,N_780);
nor U1862 (N_1862,N_110,N_234);
and U1863 (N_1863,N_568,N_406);
nor U1864 (N_1864,N_797,N_899);
nor U1865 (N_1865,N_647,N_578);
nand U1866 (N_1866,N_786,N_0);
nor U1867 (N_1867,N_235,N_469);
nand U1868 (N_1868,N_541,N_803);
xor U1869 (N_1869,N_256,N_289);
or U1870 (N_1870,N_263,N_167);
or U1871 (N_1871,N_276,N_755);
or U1872 (N_1872,N_375,N_419);
and U1873 (N_1873,N_960,N_51);
nor U1874 (N_1874,N_647,N_413);
xnor U1875 (N_1875,N_872,N_89);
xor U1876 (N_1876,N_601,N_4);
nand U1877 (N_1877,N_903,N_439);
nand U1878 (N_1878,N_455,N_760);
or U1879 (N_1879,N_339,N_814);
or U1880 (N_1880,N_230,N_414);
nand U1881 (N_1881,N_655,N_987);
and U1882 (N_1882,N_286,N_168);
and U1883 (N_1883,N_344,N_429);
nand U1884 (N_1884,N_158,N_780);
and U1885 (N_1885,N_625,N_887);
nor U1886 (N_1886,N_884,N_705);
nor U1887 (N_1887,N_82,N_134);
nor U1888 (N_1888,N_33,N_287);
and U1889 (N_1889,N_910,N_696);
nor U1890 (N_1890,N_256,N_929);
nand U1891 (N_1891,N_121,N_954);
nand U1892 (N_1892,N_403,N_446);
and U1893 (N_1893,N_950,N_373);
nor U1894 (N_1894,N_622,N_169);
or U1895 (N_1895,N_917,N_729);
and U1896 (N_1896,N_802,N_567);
or U1897 (N_1897,N_622,N_264);
or U1898 (N_1898,N_921,N_923);
nor U1899 (N_1899,N_91,N_949);
or U1900 (N_1900,N_271,N_116);
or U1901 (N_1901,N_186,N_374);
and U1902 (N_1902,N_458,N_341);
nand U1903 (N_1903,N_366,N_118);
and U1904 (N_1904,N_283,N_188);
nand U1905 (N_1905,N_106,N_3);
and U1906 (N_1906,N_66,N_822);
or U1907 (N_1907,N_940,N_461);
and U1908 (N_1908,N_828,N_767);
or U1909 (N_1909,N_870,N_388);
nand U1910 (N_1910,N_940,N_257);
or U1911 (N_1911,N_201,N_790);
nor U1912 (N_1912,N_30,N_267);
and U1913 (N_1913,N_628,N_841);
nor U1914 (N_1914,N_567,N_425);
nand U1915 (N_1915,N_335,N_526);
and U1916 (N_1916,N_545,N_735);
nand U1917 (N_1917,N_796,N_851);
xor U1918 (N_1918,N_557,N_944);
nor U1919 (N_1919,N_126,N_949);
nand U1920 (N_1920,N_717,N_845);
or U1921 (N_1921,N_581,N_441);
nor U1922 (N_1922,N_571,N_39);
nand U1923 (N_1923,N_79,N_634);
nor U1924 (N_1924,N_793,N_659);
nor U1925 (N_1925,N_419,N_759);
nor U1926 (N_1926,N_953,N_11);
and U1927 (N_1927,N_899,N_572);
nand U1928 (N_1928,N_437,N_73);
nand U1929 (N_1929,N_17,N_737);
or U1930 (N_1930,N_859,N_332);
or U1931 (N_1931,N_198,N_590);
nor U1932 (N_1932,N_202,N_39);
nor U1933 (N_1933,N_774,N_771);
or U1934 (N_1934,N_544,N_868);
or U1935 (N_1935,N_910,N_704);
nand U1936 (N_1936,N_822,N_924);
and U1937 (N_1937,N_38,N_323);
nor U1938 (N_1938,N_938,N_206);
and U1939 (N_1939,N_252,N_309);
or U1940 (N_1940,N_744,N_528);
nand U1941 (N_1941,N_279,N_907);
or U1942 (N_1942,N_808,N_422);
or U1943 (N_1943,N_205,N_290);
or U1944 (N_1944,N_195,N_666);
nand U1945 (N_1945,N_159,N_318);
nand U1946 (N_1946,N_146,N_210);
nor U1947 (N_1947,N_721,N_208);
nor U1948 (N_1948,N_429,N_920);
nor U1949 (N_1949,N_399,N_887);
and U1950 (N_1950,N_801,N_685);
or U1951 (N_1951,N_759,N_400);
or U1952 (N_1952,N_894,N_608);
or U1953 (N_1953,N_100,N_486);
or U1954 (N_1954,N_74,N_715);
nand U1955 (N_1955,N_670,N_690);
and U1956 (N_1956,N_540,N_681);
nor U1957 (N_1957,N_339,N_639);
or U1958 (N_1958,N_812,N_366);
or U1959 (N_1959,N_108,N_460);
xor U1960 (N_1960,N_66,N_989);
nor U1961 (N_1961,N_566,N_422);
or U1962 (N_1962,N_238,N_633);
and U1963 (N_1963,N_134,N_670);
nand U1964 (N_1964,N_727,N_188);
or U1965 (N_1965,N_66,N_489);
and U1966 (N_1966,N_235,N_410);
nand U1967 (N_1967,N_984,N_520);
xnor U1968 (N_1968,N_794,N_106);
and U1969 (N_1969,N_354,N_699);
nand U1970 (N_1970,N_926,N_603);
nor U1971 (N_1971,N_98,N_208);
nand U1972 (N_1972,N_243,N_182);
nand U1973 (N_1973,N_111,N_684);
nand U1974 (N_1974,N_721,N_371);
xor U1975 (N_1975,N_963,N_520);
or U1976 (N_1976,N_933,N_810);
or U1977 (N_1977,N_190,N_2);
nand U1978 (N_1978,N_256,N_54);
or U1979 (N_1979,N_143,N_595);
nor U1980 (N_1980,N_620,N_246);
nand U1981 (N_1981,N_28,N_113);
nor U1982 (N_1982,N_293,N_487);
or U1983 (N_1983,N_869,N_386);
xor U1984 (N_1984,N_64,N_722);
and U1985 (N_1985,N_894,N_242);
nand U1986 (N_1986,N_853,N_237);
and U1987 (N_1987,N_294,N_988);
or U1988 (N_1988,N_497,N_209);
nor U1989 (N_1989,N_584,N_992);
nor U1990 (N_1990,N_688,N_309);
and U1991 (N_1991,N_45,N_5);
nor U1992 (N_1992,N_886,N_739);
nand U1993 (N_1993,N_344,N_975);
and U1994 (N_1994,N_8,N_58);
and U1995 (N_1995,N_644,N_221);
nor U1996 (N_1996,N_485,N_66);
or U1997 (N_1997,N_251,N_401);
nor U1998 (N_1998,N_462,N_418);
nor U1999 (N_1999,N_870,N_906);
nand U2000 (N_2000,N_1191,N_1089);
or U2001 (N_2001,N_1661,N_1496);
nand U2002 (N_2002,N_1177,N_1378);
nand U2003 (N_2003,N_1522,N_1779);
and U2004 (N_2004,N_1977,N_1428);
and U2005 (N_2005,N_1229,N_1876);
and U2006 (N_2006,N_1572,N_1722);
nor U2007 (N_2007,N_1628,N_1888);
xor U2008 (N_2008,N_1725,N_1968);
and U2009 (N_2009,N_1846,N_1823);
and U2010 (N_2010,N_1466,N_1623);
and U2011 (N_2011,N_1656,N_1692);
nand U2012 (N_2012,N_1763,N_1591);
or U2013 (N_2013,N_1135,N_1875);
and U2014 (N_2014,N_1465,N_1903);
xor U2015 (N_2015,N_1881,N_1862);
nor U2016 (N_2016,N_1784,N_1321);
nand U2017 (N_2017,N_1417,N_1695);
nor U2018 (N_2018,N_1140,N_1458);
or U2019 (N_2019,N_1964,N_1296);
or U2020 (N_2020,N_1363,N_1821);
nand U2021 (N_2021,N_1454,N_1643);
nand U2022 (N_2022,N_1293,N_1445);
and U2023 (N_2023,N_1058,N_1648);
and U2024 (N_2024,N_1502,N_1832);
or U2025 (N_2025,N_1124,N_1556);
or U2026 (N_2026,N_1141,N_1901);
and U2027 (N_2027,N_1283,N_1434);
or U2028 (N_2028,N_1227,N_1604);
or U2029 (N_2029,N_1536,N_1091);
nor U2030 (N_2030,N_1994,N_1511);
or U2031 (N_2031,N_1517,N_1199);
nor U2032 (N_2032,N_1398,N_1214);
and U2033 (N_2033,N_1811,N_1059);
nor U2034 (N_2034,N_1577,N_1733);
xor U2035 (N_2035,N_1279,N_1807);
nand U2036 (N_2036,N_1772,N_1006);
nand U2037 (N_2037,N_1097,N_1701);
or U2038 (N_2038,N_1554,N_1965);
or U2039 (N_2039,N_1009,N_1143);
nand U2040 (N_2040,N_1337,N_1838);
or U2041 (N_2041,N_1081,N_1034);
nand U2042 (N_2042,N_1063,N_1858);
or U2043 (N_2043,N_1826,N_1737);
nand U2044 (N_2044,N_1674,N_1381);
nor U2045 (N_2045,N_1017,N_1074);
or U2046 (N_2046,N_1213,N_1793);
nor U2047 (N_2047,N_1208,N_1548);
nor U2048 (N_2048,N_1840,N_1112);
nand U2049 (N_2049,N_1192,N_1524);
nor U2050 (N_2050,N_1746,N_1877);
nor U2051 (N_2051,N_1892,N_1275);
and U2052 (N_2052,N_1658,N_1889);
and U2053 (N_2053,N_1675,N_1553);
or U2054 (N_2054,N_1188,N_1549);
xnor U2055 (N_2055,N_1365,N_1108);
and U2056 (N_2056,N_1935,N_1709);
and U2057 (N_2057,N_1714,N_1393);
nand U2058 (N_2058,N_1236,N_1072);
nor U2059 (N_2059,N_1167,N_1665);
nor U2060 (N_2060,N_1024,N_1110);
or U2061 (N_2061,N_1054,N_1232);
nand U2062 (N_2062,N_1376,N_1016);
nor U2063 (N_2063,N_1891,N_1197);
or U2064 (N_2064,N_1806,N_1996);
and U2065 (N_2065,N_1479,N_1298);
xnor U2066 (N_2066,N_1587,N_1045);
and U2067 (N_2067,N_1314,N_1448);
or U2068 (N_2068,N_1038,N_1865);
nor U2069 (N_2069,N_1134,N_1543);
nand U2070 (N_2070,N_1264,N_1348);
or U2071 (N_2071,N_1914,N_1230);
and U2072 (N_2072,N_1401,N_1406);
or U2073 (N_2073,N_1861,N_1367);
or U2074 (N_2074,N_1211,N_1362);
or U2075 (N_2075,N_1286,N_1446);
nand U2076 (N_2076,N_1924,N_1592);
or U2077 (N_2077,N_1262,N_1802);
and U2078 (N_2078,N_1392,N_1305);
and U2079 (N_2079,N_1269,N_1715);
or U2080 (N_2080,N_1079,N_1583);
or U2081 (N_2081,N_1099,N_1154);
nor U2082 (N_2082,N_1571,N_1245);
nor U2083 (N_2083,N_1650,N_1796);
or U2084 (N_2084,N_1787,N_1541);
and U2085 (N_2085,N_1451,N_1330);
nor U2086 (N_2086,N_1165,N_1655);
or U2087 (N_2087,N_1982,N_1537);
nor U2088 (N_2088,N_1387,N_1927);
or U2089 (N_2089,N_1345,N_1101);
nand U2090 (N_2090,N_1760,N_1723);
and U2091 (N_2091,N_1841,N_1683);
xor U2092 (N_2092,N_1341,N_1313);
nand U2093 (N_2093,N_1855,N_1637);
nand U2094 (N_2094,N_1237,N_1620);
nand U2095 (N_2095,N_1594,N_1023);
nor U2096 (N_2096,N_1538,N_1453);
and U2097 (N_2097,N_1086,N_1781);
or U2098 (N_2098,N_1829,N_1506);
nor U2099 (N_2099,N_1552,N_1622);
xnor U2100 (N_2100,N_1630,N_1680);
and U2101 (N_2101,N_1120,N_1696);
or U2102 (N_2102,N_1767,N_1164);
or U2103 (N_2103,N_1886,N_1126);
nor U2104 (N_2104,N_1920,N_1021);
nor U2105 (N_2105,N_1952,N_1973);
and U2106 (N_2106,N_1360,N_1752);
or U2107 (N_2107,N_1997,N_1989);
or U2108 (N_2108,N_1272,N_1399);
or U2109 (N_2109,N_1910,N_1971);
nand U2110 (N_2110,N_1719,N_1057);
and U2111 (N_2111,N_1642,N_1336);
nand U2112 (N_2112,N_1672,N_1581);
nor U2113 (N_2113,N_1419,N_1922);
or U2114 (N_2114,N_1640,N_1307);
nand U2115 (N_2115,N_1944,N_1000);
nand U2116 (N_2116,N_1349,N_1870);
or U2117 (N_2117,N_1457,N_1487);
xor U2118 (N_2118,N_1596,N_1555);
nor U2119 (N_2119,N_1686,N_1347);
nor U2120 (N_2120,N_1344,N_1312);
and U2121 (N_2121,N_1357,N_1991);
xor U2122 (N_2122,N_1516,N_1193);
or U2123 (N_2123,N_1615,N_1815);
nand U2124 (N_2124,N_1817,N_1663);
and U2125 (N_2125,N_1909,N_1681);
xor U2126 (N_2126,N_1106,N_1383);
nor U2127 (N_2127,N_1477,N_1289);
nand U2128 (N_2128,N_1624,N_1184);
nand U2129 (N_2129,N_1573,N_1762);
and U2130 (N_2130,N_1856,N_1201);
xor U2131 (N_2131,N_1593,N_1353);
nand U2132 (N_2132,N_1327,N_1791);
or U2133 (N_2133,N_1439,N_1157);
nand U2134 (N_2134,N_1693,N_1519);
xor U2135 (N_2135,N_1810,N_1566);
and U2136 (N_2136,N_1361,N_1651);
nor U2137 (N_2137,N_1716,N_1690);
and U2138 (N_2138,N_1073,N_1843);
or U2139 (N_2139,N_1472,N_1700);
nor U2140 (N_2140,N_1761,N_1462);
or U2141 (N_2141,N_1249,N_1318);
or U2142 (N_2142,N_1179,N_1122);
nand U2143 (N_2143,N_1409,N_1638);
xor U2144 (N_2144,N_1437,N_1268);
nand U2145 (N_2145,N_1530,N_1489);
and U2146 (N_2146,N_1037,N_1426);
nor U2147 (N_2147,N_1026,N_1464);
and U2148 (N_2148,N_1917,N_1092);
or U2149 (N_2149,N_1677,N_1299);
or U2150 (N_2150,N_1742,N_1241);
nor U2151 (N_2151,N_1359,N_1443);
and U2152 (N_2152,N_1325,N_1463);
and U2153 (N_2153,N_1768,N_1985);
and U2154 (N_2154,N_1030,N_1206);
or U2155 (N_2155,N_1839,N_1253);
nand U2156 (N_2156,N_1107,N_1565);
and U2157 (N_2157,N_1906,N_1231);
or U2158 (N_2158,N_1266,N_1720);
nand U2159 (N_2159,N_1388,N_1939);
xor U2160 (N_2160,N_1609,N_1644);
xor U2161 (N_2161,N_1830,N_1647);
or U2162 (N_2162,N_1532,N_1560);
nor U2163 (N_2163,N_1137,N_1261);
nor U2164 (N_2164,N_1744,N_1412);
nor U2165 (N_2165,N_1402,N_1127);
nand U2166 (N_2166,N_1780,N_1494);
and U2167 (N_2167,N_1189,N_1055);
xnor U2168 (N_2168,N_1669,N_1645);
nor U2169 (N_2169,N_1308,N_1271);
nor U2170 (N_2170,N_1745,N_1297);
and U2171 (N_2171,N_1528,N_1602);
xnor U2172 (N_2172,N_1194,N_1350);
nor U2173 (N_2173,N_1667,N_1795);
xor U2174 (N_2174,N_1851,N_1697);
nor U2175 (N_2175,N_1246,N_1435);
nand U2176 (N_2176,N_1385,N_1694);
nor U2177 (N_2177,N_1514,N_1042);
and U2178 (N_2178,N_1270,N_1688);
or U2179 (N_2179,N_1684,N_1216);
nand U2180 (N_2180,N_1473,N_1371);
or U2181 (N_2181,N_1918,N_1203);
nand U2182 (N_2182,N_1222,N_1377);
and U2183 (N_2183,N_1526,N_1163);
and U2184 (N_2184,N_1751,N_1614);
nand U2185 (N_2185,N_1803,N_1929);
xor U2186 (N_2186,N_1984,N_1934);
or U2187 (N_2187,N_1508,N_1764);
nand U2188 (N_2188,N_1049,N_1225);
or U2189 (N_2189,N_1953,N_1332);
and U2190 (N_2190,N_1682,N_1204);
nand U2191 (N_2191,N_1404,N_1905);
and U2192 (N_2192,N_1427,N_1324);
xnor U2193 (N_2193,N_1588,N_1224);
nand U2194 (N_2194,N_1162,N_1090);
nor U2195 (N_2195,N_1217,N_1729);
or U2196 (N_2196,N_1257,N_1657);
and U2197 (N_2197,N_1626,N_1575);
nand U2198 (N_2198,N_1255,N_1662);
nand U2199 (N_2199,N_1469,N_1703);
nor U2200 (N_2200,N_1827,N_1652);
xor U2201 (N_2201,N_1080,N_1105);
nor U2202 (N_2202,N_1062,N_1600);
xor U2203 (N_2203,N_1860,N_1713);
nor U2204 (N_2204,N_1818,N_1961);
nor U2205 (N_2205,N_1083,N_1295);
nand U2206 (N_2206,N_1864,N_1056);
nand U2207 (N_2207,N_1040,N_1979);
nand U2208 (N_2208,N_1012,N_1576);
nor U2209 (N_2209,N_1708,N_1902);
nand U2210 (N_2210,N_1178,N_1774);
and U2211 (N_2211,N_1287,N_1853);
and U2212 (N_2212,N_1616,N_1405);
nor U2213 (N_2213,N_1254,N_1195);
nand U2214 (N_2214,N_1625,N_1075);
and U2215 (N_2215,N_1753,N_1945);
xor U2216 (N_2216,N_1574,N_1407);
and U2217 (N_2217,N_1433,N_1460);
nor U2218 (N_2218,N_1171,N_1689);
nand U2219 (N_2219,N_1260,N_1323);
or U2220 (N_2220,N_1242,N_1601);
xnor U2221 (N_2221,N_1666,N_1095);
and U2222 (N_2222,N_1699,N_1797);
or U2223 (N_2223,N_1520,N_1098);
nand U2224 (N_2224,N_1276,N_1033);
nand U2225 (N_2225,N_1887,N_1147);
nand U2226 (N_2226,N_1316,N_1133);
nor U2227 (N_2227,N_1585,N_1990);
nor U2228 (N_2228,N_1161,N_1183);
or U2229 (N_2229,N_1738,N_1702);
nand U2230 (N_2230,N_1495,N_1317);
and U2231 (N_2231,N_1710,N_1442);
and U2232 (N_2232,N_1863,N_1370);
xor U2233 (N_2233,N_1440,N_1082);
or U2234 (N_2234,N_1529,N_1410);
or U2235 (N_2235,N_1156,N_1597);
nor U2236 (N_2236,N_1919,N_1676);
nor U2237 (N_2237,N_1704,N_1957);
nand U2238 (N_2238,N_1390,N_1885);
nand U2239 (N_2239,N_1724,N_1088);
nor U2240 (N_2240,N_1804,N_1436);
nand U2241 (N_2241,N_1455,N_1819);
or U2242 (N_2242,N_1010,N_1938);
and U2243 (N_2243,N_1564,N_1247);
or U2244 (N_2244,N_1131,N_1825);
nand U2245 (N_2245,N_1338,N_1567);
xor U2246 (N_2246,N_1734,N_1234);
or U2247 (N_2247,N_1485,N_1265);
or U2248 (N_2248,N_1782,N_1568);
and U2249 (N_2249,N_1498,N_1955);
nor U2250 (N_2250,N_1562,N_1756);
nand U2251 (N_2251,N_1300,N_1022);
and U2252 (N_2252,N_1940,N_1066);
or U2253 (N_2253,N_1490,N_1612);
xnor U2254 (N_2254,N_1326,N_1857);
nand U2255 (N_2255,N_1976,N_1218);
and U2256 (N_2256,N_1028,N_1874);
nand U2257 (N_2257,N_1850,N_1783);
nor U2258 (N_2258,N_1333,N_1907);
xnor U2259 (N_2259,N_1431,N_1963);
nand U2260 (N_2260,N_1303,N_1306);
nor U2261 (N_2261,N_1027,N_1175);
nor U2262 (N_2262,N_1911,N_1174);
nand U2263 (N_2263,N_1480,N_1966);
nor U2264 (N_2264,N_1356,N_1117);
nor U2265 (N_2265,N_1041,N_1138);
or U2266 (N_2266,N_1032,N_1233);
nor U2267 (N_2267,N_1925,N_1284);
nor U2268 (N_2268,N_1928,N_1605);
xnor U2269 (N_2269,N_1967,N_1239);
or U2270 (N_2270,N_1153,N_1915);
nand U2271 (N_2271,N_1382,N_1053);
and U2272 (N_2272,N_1280,N_1582);
xor U2273 (N_2273,N_1736,N_1396);
or U2274 (N_2274,N_1546,N_1606);
nand U2275 (N_2275,N_1301,N_1430);
nor U2276 (N_2276,N_1450,N_1292);
nor U2277 (N_2277,N_1949,N_1842);
xnor U2278 (N_2278,N_1834,N_1411);
nand U2279 (N_2279,N_1951,N_1687);
nor U2280 (N_2280,N_1486,N_1150);
or U2281 (N_2281,N_1854,N_1882);
nor U2282 (N_2282,N_1794,N_1429);
nand U2283 (N_2283,N_1664,N_1148);
nor U2284 (N_2284,N_1007,N_1956);
or U2285 (N_2285,N_1867,N_1334);
or U2286 (N_2286,N_1400,N_1375);
nand U2287 (N_2287,N_1019,N_1173);
or U2288 (N_2288,N_1987,N_1152);
nand U2289 (N_2289,N_1717,N_1413);
nor U2290 (N_2290,N_1619,N_1879);
or U2291 (N_2291,N_1483,N_1908);
nand U2292 (N_2292,N_1001,N_1223);
nor U2293 (N_2293,N_1482,N_1481);
and U2294 (N_2294,N_1848,N_1921);
nor U2295 (N_2295,N_1077,N_1880);
and U2296 (N_2296,N_1579,N_1765);
nor U2297 (N_2297,N_1043,N_1852);
nand U2298 (N_2298,N_1789,N_1273);
nor U2299 (N_2299,N_1476,N_1711);
or U2300 (N_2300,N_1277,N_1492);
or U2301 (N_2301,N_1364,N_1207);
or U2302 (N_2302,N_1475,N_1603);
and U2303 (N_2303,N_1691,N_1598);
and U2304 (N_2304,N_1172,N_1386);
nor U2305 (N_2305,N_1618,N_1859);
or U2306 (N_2306,N_1978,N_1160);
or U2307 (N_2307,N_1397,N_1766);
and U2308 (N_2308,N_1732,N_1534);
and U2309 (N_2309,N_1707,N_1563);
and U2310 (N_2310,N_1226,N_1116);
nand U2311 (N_2311,N_1893,N_1251);
and U2312 (N_2312,N_1493,N_1315);
or U2313 (N_2313,N_1969,N_1258);
and U2314 (N_2314,N_1182,N_1035);
nand U2315 (N_2315,N_1039,N_1649);
nand U2316 (N_2316,N_1470,N_1243);
and U2317 (N_2317,N_1739,N_1671);
or U2318 (N_2318,N_1025,N_1747);
nor U2319 (N_2319,N_1240,N_1219);
or U2320 (N_2320,N_1942,N_1559);
nor U2321 (N_2321,N_1916,N_1561);
nand U2322 (N_2322,N_1912,N_1136);
nand U2323 (N_2323,N_1020,N_1181);
or U2324 (N_2324,N_1960,N_1139);
nor U2325 (N_2325,N_1111,N_1515);
nor U2326 (N_2326,N_1633,N_1721);
nor U2327 (N_2327,N_1584,N_1629);
nand U2328 (N_2328,N_1970,N_1061);
or U2329 (N_2329,N_1558,N_1046);
nand U2330 (N_2330,N_1256,N_1557);
nor U2331 (N_2331,N_1510,N_1048);
nand U2332 (N_2332,N_1569,N_1551);
or U2333 (N_2333,N_1718,N_1076);
nor U2334 (N_2334,N_1169,N_1894);
nand U2335 (N_2335,N_1769,N_1113);
nor U2336 (N_2336,N_1340,N_1813);
and U2337 (N_2337,N_1754,N_1706);
and U2338 (N_2338,N_1883,N_1958);
and U2339 (N_2339,N_1513,N_1444);
nor U2340 (N_2340,N_1159,N_1221);
xor U2341 (N_2341,N_1414,N_1125);
nor U2342 (N_2342,N_1259,N_1758);
nor U2343 (N_2343,N_1743,N_1844);
or U2344 (N_2344,N_1084,N_1339);
or U2345 (N_2345,N_1008,N_1394);
or U2346 (N_2346,N_1202,N_1471);
xor U2347 (N_2347,N_1452,N_1186);
nand U2348 (N_2348,N_1896,N_1085);
xnor U2349 (N_2349,N_1087,N_1635);
or U2350 (N_2350,N_1613,N_1974);
and U2351 (N_2351,N_1004,N_1750);
nand U2352 (N_2352,N_1212,N_1959);
or U2353 (N_2353,N_1748,N_1389);
xor U2354 (N_2354,N_1812,N_1930);
and U2355 (N_2355,N_1267,N_1932);
nor U2356 (N_2356,N_1941,N_1828);
nand U2357 (N_2357,N_1068,N_1238);
and U2358 (N_2358,N_1878,N_1119);
or U2359 (N_2359,N_1384,N_1015);
nand U2360 (N_2360,N_1972,N_1070);
and U2361 (N_2361,N_1118,N_1726);
or U2362 (N_2362,N_1302,N_1474);
nor U2363 (N_2363,N_1948,N_1636);
or U2364 (N_2364,N_1755,N_1031);
or U2365 (N_2365,N_1155,N_1003);
or U2366 (N_2366,N_1809,N_1209);
nand U2367 (N_2367,N_1790,N_1491);
nand U2368 (N_2368,N_1539,N_1503);
nand U2369 (N_2369,N_1607,N_1190);
nand U2370 (N_2370,N_1067,N_1728);
or U2371 (N_2371,N_1531,N_1586);
and U2372 (N_2372,N_1425,N_1540);
and U2373 (N_2373,N_1309,N_1759);
nand U2374 (N_2374,N_1547,N_1773);
or U2375 (N_2375,N_1252,N_1343);
or U2376 (N_2376,N_1320,N_1798);
nand U2377 (N_2377,N_1328,N_1980);
nand U2378 (N_2378,N_1497,N_1873);
nand U2379 (N_2379,N_1776,N_1044);
nor U2380 (N_2380,N_1158,N_1422);
nor U2381 (N_2381,N_1771,N_1527);
nor U2382 (N_2382,N_1947,N_1198);
and U2383 (N_2383,N_1653,N_1580);
nor U2384 (N_2384,N_1712,N_1005);
xor U2385 (N_2385,N_1632,N_1282);
and U2386 (N_2386,N_1500,N_1176);
nor U2387 (N_2387,N_1578,N_1975);
and U2388 (N_2388,N_1535,N_1962);
or U2389 (N_2389,N_1641,N_1052);
and U2390 (N_2390,N_1215,N_1329);
and U2391 (N_2391,N_1488,N_1395);
xor U2392 (N_2392,N_1673,N_1166);
nand U2393 (N_2393,N_1368,N_1121);
and U2394 (N_2394,N_1310,N_1542);
nand U2395 (N_2395,N_1011,N_1931);
or U2396 (N_2396,N_1069,N_1335);
xor U2397 (N_2397,N_1461,N_1685);
nor U2398 (N_2398,N_1824,N_1484);
and U2399 (N_2399,N_1468,N_1646);
or U2400 (N_2400,N_1668,N_1499);
and U2401 (N_2401,N_1346,N_1847);
nand U2402 (N_2402,N_1518,N_1456);
xnor U2403 (N_2403,N_1094,N_1109);
or U2404 (N_2404,N_1200,N_1936);
and U2405 (N_2405,N_1801,N_1051);
nor U2406 (N_2406,N_1814,N_1570);
and U2407 (N_2407,N_1248,N_1129);
and U2408 (N_2408,N_1670,N_1884);
nor U2409 (N_2409,N_1278,N_1988);
nor U2410 (N_2410,N_1868,N_1244);
nor U2411 (N_2411,N_1014,N_1142);
nand U2412 (N_2412,N_1123,N_1898);
xor U2413 (N_2413,N_1047,N_1775);
nor U2414 (N_2414,N_1441,N_1130);
nor U2415 (N_2415,N_1342,N_1291);
nor U2416 (N_2416,N_1210,N_1416);
or U2417 (N_2417,N_1180,N_1995);
xnor U2418 (N_2418,N_1599,N_1352);
and U2419 (N_2419,N_1836,N_1808);
nand U2420 (N_2420,N_1816,N_1835);
and U2421 (N_2421,N_1029,N_1504);
nor U2422 (N_2422,N_1369,N_1355);
nor U2423 (N_2423,N_1115,N_1403);
or U2424 (N_2424,N_1679,N_1235);
xor U2425 (N_2425,N_1505,N_1950);
xnor U2426 (N_2426,N_1698,N_1447);
xnor U2427 (N_2427,N_1890,N_1220);
and U2428 (N_2428,N_1170,N_1071);
and U2429 (N_2429,N_1128,N_1380);
nor U2430 (N_2430,N_1866,N_1731);
nand U2431 (N_2431,N_1899,N_1096);
nand U2432 (N_2432,N_1943,N_1590);
nor U2433 (N_2433,N_1923,N_1151);
or U2434 (N_2434,N_1168,N_1322);
nand U2435 (N_2435,N_1250,N_1610);
nand U2436 (N_2436,N_1871,N_1438);
and U2437 (N_2437,N_1478,N_1512);
nor U2438 (N_2438,N_1294,N_1523);
xor U2439 (N_2439,N_1904,N_1981);
or U2440 (N_2440,N_1374,N_1228);
nor U2441 (N_2441,N_1897,N_1833);
xnor U2442 (N_2442,N_1449,N_1872);
or U2443 (N_2443,N_1196,N_1432);
nor U2444 (N_2444,N_1589,N_1705);
and U2445 (N_2445,N_1002,N_1913);
nor U2446 (N_2446,N_1820,N_1986);
and U2447 (N_2447,N_1792,N_1281);
nor U2448 (N_2448,N_1730,N_1946);
nor U2449 (N_2449,N_1509,N_1845);
xnor U2450 (N_2450,N_1786,N_1351);
and U2451 (N_2451,N_1205,N_1926);
nor U2452 (N_2452,N_1185,N_1093);
nor U2453 (N_2453,N_1521,N_1634);
nor U2454 (N_2454,N_1421,N_1102);
and U2455 (N_2455,N_1608,N_1036);
and U2456 (N_2456,N_1741,N_1418);
nand U2457 (N_2457,N_1999,N_1900);
or U2458 (N_2458,N_1785,N_1937);
nor U2459 (N_2459,N_1501,N_1983);
or U2460 (N_2460,N_1100,N_1415);
xnor U2461 (N_2461,N_1533,N_1993);
nand U2462 (N_2462,N_1805,N_1274);
nor U2463 (N_2463,N_1373,N_1103);
nand U2464 (N_2464,N_1895,N_1132);
nand U2465 (N_2465,N_1065,N_1617);
and U2466 (N_2466,N_1263,N_1354);
or U2467 (N_2467,N_1777,N_1379);
or U2468 (N_2468,N_1992,N_1631);
or U2469 (N_2469,N_1060,N_1064);
nor U2470 (N_2470,N_1545,N_1933);
nand U2471 (N_2471,N_1998,N_1459);
or U2472 (N_2472,N_1660,N_1366);
nand U2473 (N_2473,N_1146,N_1869);
or U2474 (N_2474,N_1285,N_1358);
or U2475 (N_2475,N_1757,N_1639);
nor U2476 (N_2476,N_1544,N_1078);
and U2477 (N_2477,N_1423,N_1144);
or U2478 (N_2478,N_1467,N_1408);
xor U2479 (N_2479,N_1659,N_1319);
nand U2480 (N_2480,N_1595,N_1104);
nor U2481 (N_2481,N_1331,N_1954);
nand U2482 (N_2482,N_1391,N_1735);
and U2483 (N_2483,N_1770,N_1013);
and U2484 (N_2484,N_1727,N_1050);
or U2485 (N_2485,N_1778,N_1654);
and U2486 (N_2486,N_1145,N_1424);
or U2487 (N_2487,N_1507,N_1550);
or U2488 (N_2488,N_1018,N_1740);
nand U2489 (N_2489,N_1822,N_1311);
nor U2490 (N_2490,N_1304,N_1837);
or U2491 (N_2491,N_1372,N_1627);
and U2492 (N_2492,N_1149,N_1187);
and U2493 (N_2493,N_1290,N_1621);
nand U2494 (N_2494,N_1749,N_1288);
nor U2495 (N_2495,N_1678,N_1799);
nand U2496 (N_2496,N_1849,N_1525);
xnor U2497 (N_2497,N_1831,N_1114);
nor U2498 (N_2498,N_1788,N_1800);
nand U2499 (N_2499,N_1611,N_1420);
or U2500 (N_2500,N_1865,N_1529);
and U2501 (N_2501,N_1814,N_1265);
or U2502 (N_2502,N_1266,N_1483);
and U2503 (N_2503,N_1326,N_1492);
or U2504 (N_2504,N_1126,N_1561);
and U2505 (N_2505,N_1128,N_1063);
nor U2506 (N_2506,N_1134,N_1030);
or U2507 (N_2507,N_1332,N_1689);
nor U2508 (N_2508,N_1067,N_1394);
xnor U2509 (N_2509,N_1678,N_1166);
and U2510 (N_2510,N_1628,N_1976);
nor U2511 (N_2511,N_1752,N_1204);
or U2512 (N_2512,N_1950,N_1231);
or U2513 (N_2513,N_1015,N_1601);
or U2514 (N_2514,N_1211,N_1798);
or U2515 (N_2515,N_1561,N_1125);
or U2516 (N_2516,N_1863,N_1300);
nor U2517 (N_2517,N_1852,N_1187);
or U2518 (N_2518,N_1413,N_1514);
or U2519 (N_2519,N_1969,N_1334);
or U2520 (N_2520,N_1130,N_1297);
nand U2521 (N_2521,N_1734,N_1533);
and U2522 (N_2522,N_1672,N_1726);
or U2523 (N_2523,N_1316,N_1444);
nand U2524 (N_2524,N_1156,N_1903);
and U2525 (N_2525,N_1610,N_1445);
or U2526 (N_2526,N_1113,N_1561);
nand U2527 (N_2527,N_1712,N_1102);
nand U2528 (N_2528,N_1770,N_1692);
and U2529 (N_2529,N_1810,N_1087);
xor U2530 (N_2530,N_1650,N_1482);
and U2531 (N_2531,N_1599,N_1965);
or U2532 (N_2532,N_1034,N_1449);
or U2533 (N_2533,N_1395,N_1892);
nor U2534 (N_2534,N_1072,N_1553);
nand U2535 (N_2535,N_1386,N_1035);
nand U2536 (N_2536,N_1830,N_1709);
or U2537 (N_2537,N_1804,N_1618);
and U2538 (N_2538,N_1000,N_1834);
nor U2539 (N_2539,N_1022,N_1319);
nor U2540 (N_2540,N_1229,N_1389);
or U2541 (N_2541,N_1285,N_1641);
or U2542 (N_2542,N_1244,N_1363);
and U2543 (N_2543,N_1760,N_1652);
or U2544 (N_2544,N_1630,N_1492);
or U2545 (N_2545,N_1691,N_1139);
nand U2546 (N_2546,N_1911,N_1018);
nand U2547 (N_2547,N_1428,N_1988);
nor U2548 (N_2548,N_1756,N_1553);
nor U2549 (N_2549,N_1137,N_1681);
nor U2550 (N_2550,N_1657,N_1767);
or U2551 (N_2551,N_1974,N_1936);
nand U2552 (N_2552,N_1118,N_1314);
nand U2553 (N_2553,N_1873,N_1427);
nand U2554 (N_2554,N_1189,N_1938);
or U2555 (N_2555,N_1429,N_1170);
or U2556 (N_2556,N_1378,N_1613);
and U2557 (N_2557,N_1970,N_1456);
xnor U2558 (N_2558,N_1917,N_1644);
or U2559 (N_2559,N_1767,N_1374);
nor U2560 (N_2560,N_1453,N_1090);
and U2561 (N_2561,N_1113,N_1504);
nand U2562 (N_2562,N_1107,N_1236);
nor U2563 (N_2563,N_1581,N_1811);
nor U2564 (N_2564,N_1077,N_1167);
and U2565 (N_2565,N_1010,N_1718);
and U2566 (N_2566,N_1627,N_1485);
nand U2567 (N_2567,N_1119,N_1291);
and U2568 (N_2568,N_1646,N_1016);
nor U2569 (N_2569,N_1749,N_1745);
or U2570 (N_2570,N_1620,N_1835);
or U2571 (N_2571,N_1332,N_1338);
and U2572 (N_2572,N_1781,N_1980);
and U2573 (N_2573,N_1267,N_1821);
or U2574 (N_2574,N_1937,N_1000);
or U2575 (N_2575,N_1547,N_1694);
xor U2576 (N_2576,N_1495,N_1120);
or U2577 (N_2577,N_1548,N_1478);
nor U2578 (N_2578,N_1282,N_1898);
or U2579 (N_2579,N_1307,N_1729);
nand U2580 (N_2580,N_1220,N_1960);
nor U2581 (N_2581,N_1849,N_1239);
and U2582 (N_2582,N_1098,N_1340);
nor U2583 (N_2583,N_1797,N_1197);
nor U2584 (N_2584,N_1170,N_1505);
nand U2585 (N_2585,N_1190,N_1368);
xnor U2586 (N_2586,N_1521,N_1397);
or U2587 (N_2587,N_1285,N_1628);
nand U2588 (N_2588,N_1983,N_1436);
xnor U2589 (N_2589,N_1496,N_1751);
nor U2590 (N_2590,N_1050,N_1982);
xor U2591 (N_2591,N_1020,N_1420);
and U2592 (N_2592,N_1003,N_1906);
or U2593 (N_2593,N_1480,N_1291);
nor U2594 (N_2594,N_1881,N_1641);
nand U2595 (N_2595,N_1156,N_1387);
nand U2596 (N_2596,N_1741,N_1760);
or U2597 (N_2597,N_1277,N_1010);
or U2598 (N_2598,N_1716,N_1805);
or U2599 (N_2599,N_1180,N_1030);
or U2600 (N_2600,N_1081,N_1541);
or U2601 (N_2601,N_1881,N_1796);
and U2602 (N_2602,N_1583,N_1631);
or U2603 (N_2603,N_1404,N_1166);
nand U2604 (N_2604,N_1244,N_1713);
or U2605 (N_2605,N_1239,N_1325);
and U2606 (N_2606,N_1833,N_1629);
and U2607 (N_2607,N_1806,N_1144);
and U2608 (N_2608,N_1292,N_1279);
and U2609 (N_2609,N_1263,N_1555);
nand U2610 (N_2610,N_1597,N_1623);
nor U2611 (N_2611,N_1030,N_1583);
xor U2612 (N_2612,N_1625,N_1751);
xnor U2613 (N_2613,N_1898,N_1939);
nand U2614 (N_2614,N_1307,N_1933);
or U2615 (N_2615,N_1885,N_1193);
nor U2616 (N_2616,N_1264,N_1399);
xnor U2617 (N_2617,N_1969,N_1593);
nor U2618 (N_2618,N_1305,N_1057);
nor U2619 (N_2619,N_1175,N_1334);
nand U2620 (N_2620,N_1220,N_1955);
nand U2621 (N_2621,N_1768,N_1615);
nand U2622 (N_2622,N_1089,N_1227);
and U2623 (N_2623,N_1948,N_1504);
nor U2624 (N_2624,N_1083,N_1968);
and U2625 (N_2625,N_1316,N_1403);
nand U2626 (N_2626,N_1201,N_1709);
or U2627 (N_2627,N_1682,N_1519);
and U2628 (N_2628,N_1374,N_1525);
nor U2629 (N_2629,N_1718,N_1211);
nand U2630 (N_2630,N_1434,N_1245);
nor U2631 (N_2631,N_1898,N_1183);
or U2632 (N_2632,N_1841,N_1936);
and U2633 (N_2633,N_1394,N_1727);
nand U2634 (N_2634,N_1869,N_1820);
nand U2635 (N_2635,N_1294,N_1386);
and U2636 (N_2636,N_1590,N_1592);
xor U2637 (N_2637,N_1487,N_1995);
or U2638 (N_2638,N_1316,N_1872);
nor U2639 (N_2639,N_1315,N_1807);
nand U2640 (N_2640,N_1540,N_1975);
nor U2641 (N_2641,N_1996,N_1465);
nor U2642 (N_2642,N_1537,N_1114);
xnor U2643 (N_2643,N_1237,N_1143);
nand U2644 (N_2644,N_1021,N_1020);
nor U2645 (N_2645,N_1576,N_1261);
and U2646 (N_2646,N_1452,N_1364);
nor U2647 (N_2647,N_1591,N_1751);
xor U2648 (N_2648,N_1506,N_1230);
nand U2649 (N_2649,N_1792,N_1483);
xor U2650 (N_2650,N_1961,N_1215);
or U2651 (N_2651,N_1170,N_1259);
and U2652 (N_2652,N_1396,N_1371);
or U2653 (N_2653,N_1931,N_1095);
and U2654 (N_2654,N_1191,N_1305);
and U2655 (N_2655,N_1230,N_1980);
and U2656 (N_2656,N_1821,N_1076);
nand U2657 (N_2657,N_1837,N_1713);
xor U2658 (N_2658,N_1846,N_1150);
and U2659 (N_2659,N_1171,N_1901);
and U2660 (N_2660,N_1567,N_1156);
nor U2661 (N_2661,N_1998,N_1076);
and U2662 (N_2662,N_1256,N_1764);
and U2663 (N_2663,N_1907,N_1390);
nor U2664 (N_2664,N_1284,N_1896);
or U2665 (N_2665,N_1254,N_1620);
nor U2666 (N_2666,N_1316,N_1926);
and U2667 (N_2667,N_1712,N_1615);
or U2668 (N_2668,N_1790,N_1819);
nor U2669 (N_2669,N_1827,N_1759);
or U2670 (N_2670,N_1047,N_1137);
nor U2671 (N_2671,N_1376,N_1157);
nor U2672 (N_2672,N_1154,N_1043);
and U2673 (N_2673,N_1350,N_1694);
and U2674 (N_2674,N_1807,N_1992);
and U2675 (N_2675,N_1035,N_1864);
nand U2676 (N_2676,N_1594,N_1152);
nand U2677 (N_2677,N_1202,N_1284);
nand U2678 (N_2678,N_1425,N_1088);
nand U2679 (N_2679,N_1608,N_1592);
nor U2680 (N_2680,N_1381,N_1248);
xor U2681 (N_2681,N_1846,N_1705);
nor U2682 (N_2682,N_1788,N_1361);
or U2683 (N_2683,N_1584,N_1645);
and U2684 (N_2684,N_1010,N_1157);
or U2685 (N_2685,N_1611,N_1538);
nand U2686 (N_2686,N_1766,N_1833);
or U2687 (N_2687,N_1393,N_1476);
nand U2688 (N_2688,N_1348,N_1460);
nand U2689 (N_2689,N_1710,N_1822);
or U2690 (N_2690,N_1998,N_1357);
and U2691 (N_2691,N_1215,N_1861);
nand U2692 (N_2692,N_1851,N_1121);
and U2693 (N_2693,N_1957,N_1074);
nor U2694 (N_2694,N_1031,N_1949);
nand U2695 (N_2695,N_1266,N_1531);
and U2696 (N_2696,N_1162,N_1945);
xnor U2697 (N_2697,N_1280,N_1304);
and U2698 (N_2698,N_1645,N_1028);
and U2699 (N_2699,N_1262,N_1142);
nand U2700 (N_2700,N_1261,N_1930);
or U2701 (N_2701,N_1861,N_1175);
nor U2702 (N_2702,N_1532,N_1357);
and U2703 (N_2703,N_1214,N_1712);
xnor U2704 (N_2704,N_1059,N_1506);
nor U2705 (N_2705,N_1384,N_1895);
nor U2706 (N_2706,N_1270,N_1405);
and U2707 (N_2707,N_1149,N_1688);
nor U2708 (N_2708,N_1492,N_1664);
nor U2709 (N_2709,N_1011,N_1897);
nand U2710 (N_2710,N_1894,N_1588);
and U2711 (N_2711,N_1236,N_1115);
nand U2712 (N_2712,N_1747,N_1453);
or U2713 (N_2713,N_1945,N_1375);
nor U2714 (N_2714,N_1649,N_1162);
nor U2715 (N_2715,N_1685,N_1153);
or U2716 (N_2716,N_1252,N_1013);
and U2717 (N_2717,N_1699,N_1930);
xnor U2718 (N_2718,N_1438,N_1260);
or U2719 (N_2719,N_1490,N_1891);
nor U2720 (N_2720,N_1645,N_1994);
or U2721 (N_2721,N_1116,N_1033);
or U2722 (N_2722,N_1477,N_1914);
nand U2723 (N_2723,N_1831,N_1692);
nand U2724 (N_2724,N_1727,N_1796);
nor U2725 (N_2725,N_1592,N_1366);
or U2726 (N_2726,N_1951,N_1795);
nand U2727 (N_2727,N_1493,N_1517);
nand U2728 (N_2728,N_1176,N_1730);
and U2729 (N_2729,N_1491,N_1735);
xor U2730 (N_2730,N_1421,N_1240);
and U2731 (N_2731,N_1677,N_1313);
nand U2732 (N_2732,N_1528,N_1200);
and U2733 (N_2733,N_1557,N_1546);
nand U2734 (N_2734,N_1898,N_1284);
or U2735 (N_2735,N_1608,N_1681);
or U2736 (N_2736,N_1787,N_1566);
nor U2737 (N_2737,N_1068,N_1800);
and U2738 (N_2738,N_1590,N_1946);
or U2739 (N_2739,N_1798,N_1451);
or U2740 (N_2740,N_1373,N_1110);
nor U2741 (N_2741,N_1313,N_1202);
nor U2742 (N_2742,N_1359,N_1769);
nand U2743 (N_2743,N_1886,N_1757);
nor U2744 (N_2744,N_1572,N_1339);
and U2745 (N_2745,N_1611,N_1771);
nand U2746 (N_2746,N_1382,N_1890);
nor U2747 (N_2747,N_1620,N_1569);
nand U2748 (N_2748,N_1352,N_1149);
nor U2749 (N_2749,N_1322,N_1599);
and U2750 (N_2750,N_1872,N_1791);
and U2751 (N_2751,N_1638,N_1278);
or U2752 (N_2752,N_1392,N_1573);
xnor U2753 (N_2753,N_1770,N_1707);
and U2754 (N_2754,N_1877,N_1854);
nor U2755 (N_2755,N_1254,N_1982);
nand U2756 (N_2756,N_1316,N_1922);
or U2757 (N_2757,N_1920,N_1275);
nor U2758 (N_2758,N_1199,N_1798);
nand U2759 (N_2759,N_1540,N_1072);
nor U2760 (N_2760,N_1286,N_1769);
nor U2761 (N_2761,N_1092,N_1076);
and U2762 (N_2762,N_1058,N_1775);
or U2763 (N_2763,N_1586,N_1267);
or U2764 (N_2764,N_1363,N_1055);
or U2765 (N_2765,N_1329,N_1788);
nor U2766 (N_2766,N_1476,N_1207);
nor U2767 (N_2767,N_1704,N_1094);
nand U2768 (N_2768,N_1160,N_1113);
xor U2769 (N_2769,N_1004,N_1310);
and U2770 (N_2770,N_1509,N_1887);
and U2771 (N_2771,N_1649,N_1294);
and U2772 (N_2772,N_1700,N_1103);
nor U2773 (N_2773,N_1336,N_1745);
nor U2774 (N_2774,N_1944,N_1685);
nand U2775 (N_2775,N_1963,N_1695);
nand U2776 (N_2776,N_1771,N_1080);
nor U2777 (N_2777,N_1729,N_1559);
and U2778 (N_2778,N_1759,N_1706);
xnor U2779 (N_2779,N_1971,N_1612);
nand U2780 (N_2780,N_1436,N_1428);
nand U2781 (N_2781,N_1966,N_1958);
and U2782 (N_2782,N_1099,N_1494);
nand U2783 (N_2783,N_1398,N_1490);
and U2784 (N_2784,N_1142,N_1201);
and U2785 (N_2785,N_1659,N_1524);
or U2786 (N_2786,N_1133,N_1751);
nor U2787 (N_2787,N_1987,N_1934);
nor U2788 (N_2788,N_1037,N_1592);
or U2789 (N_2789,N_1983,N_1060);
nand U2790 (N_2790,N_1549,N_1012);
nand U2791 (N_2791,N_1487,N_1718);
nor U2792 (N_2792,N_1188,N_1387);
nand U2793 (N_2793,N_1645,N_1944);
nand U2794 (N_2794,N_1756,N_1994);
nand U2795 (N_2795,N_1481,N_1426);
and U2796 (N_2796,N_1003,N_1207);
and U2797 (N_2797,N_1201,N_1813);
nor U2798 (N_2798,N_1966,N_1235);
nor U2799 (N_2799,N_1817,N_1727);
nand U2800 (N_2800,N_1965,N_1389);
nor U2801 (N_2801,N_1832,N_1144);
nor U2802 (N_2802,N_1555,N_1521);
nor U2803 (N_2803,N_1654,N_1416);
and U2804 (N_2804,N_1632,N_1073);
nand U2805 (N_2805,N_1994,N_1376);
nand U2806 (N_2806,N_1684,N_1962);
and U2807 (N_2807,N_1206,N_1059);
xor U2808 (N_2808,N_1092,N_1008);
or U2809 (N_2809,N_1086,N_1378);
or U2810 (N_2810,N_1578,N_1519);
nor U2811 (N_2811,N_1898,N_1924);
xnor U2812 (N_2812,N_1187,N_1107);
and U2813 (N_2813,N_1652,N_1861);
and U2814 (N_2814,N_1949,N_1684);
nand U2815 (N_2815,N_1757,N_1916);
and U2816 (N_2816,N_1004,N_1147);
nor U2817 (N_2817,N_1112,N_1536);
nor U2818 (N_2818,N_1095,N_1285);
nand U2819 (N_2819,N_1957,N_1938);
nand U2820 (N_2820,N_1484,N_1364);
or U2821 (N_2821,N_1904,N_1151);
nor U2822 (N_2822,N_1560,N_1182);
nor U2823 (N_2823,N_1014,N_1983);
nor U2824 (N_2824,N_1852,N_1448);
or U2825 (N_2825,N_1505,N_1032);
nor U2826 (N_2826,N_1476,N_1349);
nand U2827 (N_2827,N_1770,N_1724);
and U2828 (N_2828,N_1202,N_1177);
nor U2829 (N_2829,N_1914,N_1454);
or U2830 (N_2830,N_1585,N_1161);
and U2831 (N_2831,N_1842,N_1665);
xnor U2832 (N_2832,N_1499,N_1802);
and U2833 (N_2833,N_1058,N_1778);
nor U2834 (N_2834,N_1557,N_1835);
nand U2835 (N_2835,N_1407,N_1488);
or U2836 (N_2836,N_1196,N_1272);
nor U2837 (N_2837,N_1459,N_1295);
and U2838 (N_2838,N_1177,N_1537);
nor U2839 (N_2839,N_1060,N_1357);
nand U2840 (N_2840,N_1976,N_1811);
xnor U2841 (N_2841,N_1039,N_1175);
or U2842 (N_2842,N_1645,N_1711);
and U2843 (N_2843,N_1201,N_1170);
nor U2844 (N_2844,N_1892,N_1195);
and U2845 (N_2845,N_1469,N_1035);
or U2846 (N_2846,N_1230,N_1205);
or U2847 (N_2847,N_1068,N_1281);
or U2848 (N_2848,N_1722,N_1550);
nor U2849 (N_2849,N_1242,N_1836);
nor U2850 (N_2850,N_1123,N_1313);
nand U2851 (N_2851,N_1866,N_1815);
nor U2852 (N_2852,N_1022,N_1366);
nand U2853 (N_2853,N_1111,N_1486);
nand U2854 (N_2854,N_1412,N_1236);
or U2855 (N_2855,N_1595,N_1777);
and U2856 (N_2856,N_1521,N_1440);
and U2857 (N_2857,N_1074,N_1534);
nor U2858 (N_2858,N_1642,N_1948);
nor U2859 (N_2859,N_1394,N_1973);
nor U2860 (N_2860,N_1796,N_1808);
or U2861 (N_2861,N_1426,N_1914);
nor U2862 (N_2862,N_1649,N_1851);
xor U2863 (N_2863,N_1636,N_1856);
nand U2864 (N_2864,N_1189,N_1393);
or U2865 (N_2865,N_1582,N_1378);
nor U2866 (N_2866,N_1417,N_1175);
xor U2867 (N_2867,N_1714,N_1902);
and U2868 (N_2868,N_1546,N_1478);
nand U2869 (N_2869,N_1439,N_1132);
nand U2870 (N_2870,N_1192,N_1526);
nor U2871 (N_2871,N_1205,N_1904);
nand U2872 (N_2872,N_1858,N_1905);
nand U2873 (N_2873,N_1553,N_1045);
nand U2874 (N_2874,N_1348,N_1618);
nor U2875 (N_2875,N_1122,N_1660);
nor U2876 (N_2876,N_1642,N_1249);
and U2877 (N_2877,N_1403,N_1516);
or U2878 (N_2878,N_1622,N_1058);
nand U2879 (N_2879,N_1331,N_1102);
xor U2880 (N_2880,N_1270,N_1776);
nand U2881 (N_2881,N_1765,N_1082);
nand U2882 (N_2882,N_1944,N_1307);
nand U2883 (N_2883,N_1353,N_1559);
and U2884 (N_2884,N_1482,N_1722);
nor U2885 (N_2885,N_1806,N_1598);
and U2886 (N_2886,N_1189,N_1018);
nand U2887 (N_2887,N_1215,N_1224);
nor U2888 (N_2888,N_1593,N_1058);
or U2889 (N_2889,N_1020,N_1648);
nor U2890 (N_2890,N_1162,N_1782);
and U2891 (N_2891,N_1780,N_1147);
nor U2892 (N_2892,N_1251,N_1998);
nand U2893 (N_2893,N_1282,N_1547);
and U2894 (N_2894,N_1402,N_1123);
or U2895 (N_2895,N_1229,N_1013);
nor U2896 (N_2896,N_1606,N_1151);
nor U2897 (N_2897,N_1072,N_1063);
and U2898 (N_2898,N_1641,N_1369);
or U2899 (N_2899,N_1956,N_1330);
or U2900 (N_2900,N_1152,N_1250);
or U2901 (N_2901,N_1662,N_1183);
nand U2902 (N_2902,N_1763,N_1972);
and U2903 (N_2903,N_1369,N_1112);
nor U2904 (N_2904,N_1104,N_1968);
or U2905 (N_2905,N_1679,N_1613);
nor U2906 (N_2906,N_1924,N_1587);
nand U2907 (N_2907,N_1036,N_1768);
or U2908 (N_2908,N_1118,N_1321);
or U2909 (N_2909,N_1684,N_1495);
nor U2910 (N_2910,N_1414,N_1497);
or U2911 (N_2911,N_1420,N_1392);
or U2912 (N_2912,N_1988,N_1807);
or U2913 (N_2913,N_1767,N_1661);
nor U2914 (N_2914,N_1861,N_1903);
nor U2915 (N_2915,N_1965,N_1900);
nand U2916 (N_2916,N_1045,N_1939);
or U2917 (N_2917,N_1639,N_1073);
nor U2918 (N_2918,N_1514,N_1646);
or U2919 (N_2919,N_1441,N_1922);
xnor U2920 (N_2920,N_1121,N_1077);
nand U2921 (N_2921,N_1706,N_1277);
nand U2922 (N_2922,N_1365,N_1468);
or U2923 (N_2923,N_1123,N_1088);
nand U2924 (N_2924,N_1385,N_1692);
nor U2925 (N_2925,N_1591,N_1856);
or U2926 (N_2926,N_1595,N_1975);
and U2927 (N_2927,N_1102,N_1868);
and U2928 (N_2928,N_1016,N_1710);
and U2929 (N_2929,N_1917,N_1495);
and U2930 (N_2930,N_1648,N_1988);
nand U2931 (N_2931,N_1822,N_1065);
or U2932 (N_2932,N_1371,N_1334);
and U2933 (N_2933,N_1409,N_1495);
nand U2934 (N_2934,N_1411,N_1677);
nand U2935 (N_2935,N_1523,N_1706);
nor U2936 (N_2936,N_1555,N_1222);
nand U2937 (N_2937,N_1958,N_1663);
nand U2938 (N_2938,N_1395,N_1732);
and U2939 (N_2939,N_1480,N_1721);
or U2940 (N_2940,N_1900,N_1082);
and U2941 (N_2941,N_1111,N_1454);
and U2942 (N_2942,N_1017,N_1103);
nor U2943 (N_2943,N_1841,N_1833);
and U2944 (N_2944,N_1028,N_1048);
and U2945 (N_2945,N_1600,N_1903);
nand U2946 (N_2946,N_1151,N_1306);
nand U2947 (N_2947,N_1664,N_1470);
and U2948 (N_2948,N_1003,N_1295);
and U2949 (N_2949,N_1332,N_1576);
or U2950 (N_2950,N_1907,N_1668);
xnor U2951 (N_2951,N_1222,N_1183);
nand U2952 (N_2952,N_1813,N_1887);
and U2953 (N_2953,N_1018,N_1299);
nand U2954 (N_2954,N_1211,N_1328);
nand U2955 (N_2955,N_1972,N_1078);
and U2956 (N_2956,N_1136,N_1697);
nor U2957 (N_2957,N_1183,N_1512);
or U2958 (N_2958,N_1787,N_1162);
and U2959 (N_2959,N_1746,N_1738);
and U2960 (N_2960,N_1057,N_1560);
and U2961 (N_2961,N_1140,N_1363);
and U2962 (N_2962,N_1131,N_1817);
or U2963 (N_2963,N_1996,N_1423);
or U2964 (N_2964,N_1146,N_1519);
nand U2965 (N_2965,N_1834,N_1988);
or U2966 (N_2966,N_1473,N_1495);
nand U2967 (N_2967,N_1585,N_1149);
nand U2968 (N_2968,N_1636,N_1296);
nor U2969 (N_2969,N_1264,N_1052);
or U2970 (N_2970,N_1402,N_1485);
or U2971 (N_2971,N_1479,N_1864);
nor U2972 (N_2972,N_1858,N_1675);
nor U2973 (N_2973,N_1804,N_1192);
nand U2974 (N_2974,N_1530,N_1119);
or U2975 (N_2975,N_1366,N_1051);
or U2976 (N_2976,N_1865,N_1191);
and U2977 (N_2977,N_1603,N_1039);
nor U2978 (N_2978,N_1320,N_1978);
nand U2979 (N_2979,N_1384,N_1191);
or U2980 (N_2980,N_1412,N_1771);
nor U2981 (N_2981,N_1563,N_1219);
or U2982 (N_2982,N_1248,N_1340);
nand U2983 (N_2983,N_1350,N_1660);
nand U2984 (N_2984,N_1341,N_1448);
or U2985 (N_2985,N_1434,N_1585);
or U2986 (N_2986,N_1073,N_1811);
nand U2987 (N_2987,N_1010,N_1874);
and U2988 (N_2988,N_1254,N_1926);
nor U2989 (N_2989,N_1474,N_1120);
and U2990 (N_2990,N_1935,N_1804);
nand U2991 (N_2991,N_1527,N_1755);
nand U2992 (N_2992,N_1795,N_1367);
or U2993 (N_2993,N_1037,N_1564);
nand U2994 (N_2994,N_1793,N_1686);
xor U2995 (N_2995,N_1636,N_1799);
xor U2996 (N_2996,N_1891,N_1202);
xor U2997 (N_2997,N_1372,N_1990);
and U2998 (N_2998,N_1829,N_1663);
nor U2999 (N_2999,N_1484,N_1581);
or U3000 (N_3000,N_2068,N_2372);
nand U3001 (N_3001,N_2889,N_2774);
nor U3002 (N_3002,N_2916,N_2004);
or U3003 (N_3003,N_2063,N_2223);
nor U3004 (N_3004,N_2328,N_2734);
and U3005 (N_3005,N_2576,N_2362);
or U3006 (N_3006,N_2943,N_2902);
nand U3007 (N_3007,N_2151,N_2994);
or U3008 (N_3008,N_2516,N_2565);
nor U3009 (N_3009,N_2700,N_2908);
or U3010 (N_3010,N_2810,N_2121);
and U3011 (N_3011,N_2976,N_2593);
or U3012 (N_3012,N_2521,N_2118);
or U3013 (N_3013,N_2541,N_2905);
and U3014 (N_3014,N_2125,N_2083);
nand U3015 (N_3015,N_2801,N_2071);
xnor U3016 (N_3016,N_2381,N_2386);
or U3017 (N_3017,N_2210,N_2193);
or U3018 (N_3018,N_2424,N_2980);
or U3019 (N_3019,N_2329,N_2335);
xor U3020 (N_3020,N_2675,N_2251);
and U3021 (N_3021,N_2697,N_2970);
and U3022 (N_3022,N_2244,N_2715);
and U3023 (N_3023,N_2499,N_2863);
xnor U3024 (N_3024,N_2594,N_2556);
nand U3025 (N_3025,N_2950,N_2147);
nor U3026 (N_3026,N_2764,N_2685);
xor U3027 (N_3027,N_2481,N_2699);
or U3028 (N_3028,N_2129,N_2038);
or U3029 (N_3029,N_2958,N_2641);
nand U3030 (N_3030,N_2072,N_2377);
or U3031 (N_3031,N_2874,N_2318);
nand U3032 (N_3032,N_2037,N_2572);
nand U3033 (N_3033,N_2538,N_2163);
or U3034 (N_3034,N_2804,N_2830);
xor U3035 (N_3035,N_2107,N_2834);
and U3036 (N_3036,N_2089,N_2585);
xnor U3037 (N_3037,N_2342,N_2455);
and U3038 (N_3038,N_2837,N_2380);
nand U3039 (N_3039,N_2947,N_2102);
and U3040 (N_3040,N_2618,N_2885);
xor U3041 (N_3041,N_2190,N_2751);
nor U3042 (N_3042,N_2939,N_2621);
nand U3043 (N_3043,N_2928,N_2997);
or U3044 (N_3044,N_2561,N_2531);
nand U3045 (N_3045,N_2303,N_2130);
and U3046 (N_3046,N_2974,N_2838);
xnor U3047 (N_3047,N_2881,N_2247);
nor U3048 (N_3048,N_2176,N_2602);
nor U3049 (N_3049,N_2274,N_2201);
or U3050 (N_3050,N_2097,N_2255);
nand U3051 (N_3051,N_2018,N_2315);
nand U3052 (N_3052,N_2194,N_2983);
xor U3053 (N_3053,N_2705,N_2748);
or U3054 (N_3054,N_2217,N_2023);
and U3055 (N_3055,N_2442,N_2695);
nor U3056 (N_3056,N_2478,N_2722);
and U3057 (N_3057,N_2321,N_2373);
or U3058 (N_3058,N_2806,N_2235);
nand U3059 (N_3059,N_2485,N_2884);
and U3060 (N_3060,N_2589,N_2419);
or U3061 (N_3061,N_2461,N_2297);
nor U3062 (N_3062,N_2486,N_2866);
xor U3063 (N_3063,N_2827,N_2009);
and U3064 (N_3064,N_2729,N_2920);
nor U3065 (N_3065,N_2987,N_2719);
or U3066 (N_3066,N_2530,N_2300);
nor U3067 (N_3067,N_2773,N_2532);
nand U3068 (N_3068,N_2620,N_2649);
nor U3069 (N_3069,N_2935,N_2665);
xnor U3070 (N_3070,N_2723,N_2820);
and U3071 (N_3071,N_2271,N_2917);
and U3072 (N_3072,N_2322,N_2805);
xnor U3073 (N_3073,N_2747,N_2379);
nand U3074 (N_3074,N_2757,N_2095);
or U3075 (N_3075,N_2267,N_2567);
nor U3076 (N_3076,N_2367,N_2616);
nor U3077 (N_3077,N_2829,N_2628);
or U3078 (N_3078,N_2140,N_2412);
or U3079 (N_3079,N_2003,N_2092);
nor U3080 (N_3080,N_2173,N_2915);
or U3081 (N_3081,N_2413,N_2488);
or U3082 (N_3082,N_2370,N_2306);
nor U3083 (N_3083,N_2555,N_2430);
or U3084 (N_3084,N_2350,N_2647);
nor U3085 (N_3085,N_2220,N_2636);
nor U3086 (N_3086,N_2355,N_2765);
nor U3087 (N_3087,N_2264,N_2382);
or U3088 (N_3088,N_2635,N_2361);
xnor U3089 (N_3089,N_2959,N_2960);
or U3090 (N_3090,N_2100,N_2547);
and U3091 (N_3091,N_2758,N_2421);
nand U3092 (N_3092,N_2661,N_2208);
and U3093 (N_3093,N_2592,N_2347);
or U3094 (N_3094,N_2629,N_2060);
or U3095 (N_3095,N_2019,N_2473);
nor U3096 (N_3096,N_2262,N_2079);
nand U3097 (N_3097,N_2826,N_2243);
xor U3098 (N_3098,N_2433,N_2680);
nand U3099 (N_3099,N_2964,N_2448);
nand U3100 (N_3100,N_2750,N_2093);
or U3101 (N_3101,N_2090,N_2245);
nand U3102 (N_3102,N_2405,N_2269);
and U3103 (N_3103,N_2371,N_2042);
and U3104 (N_3104,N_2515,N_2214);
and U3105 (N_3105,N_2776,N_2518);
nor U3106 (N_3106,N_2792,N_2154);
nor U3107 (N_3107,N_2293,N_2780);
or U3108 (N_3108,N_2465,N_2510);
or U3109 (N_3109,N_2180,N_2967);
nor U3110 (N_3110,N_2497,N_2080);
and U3111 (N_3111,N_2384,N_2698);
nand U3112 (N_3112,N_2183,N_2795);
or U3113 (N_3113,N_2257,N_2623);
or U3114 (N_3114,N_2877,N_2085);
or U3115 (N_3115,N_2663,N_2517);
and U3116 (N_3116,N_2520,N_2209);
nand U3117 (N_3117,N_2798,N_2016);
and U3118 (N_3118,N_2617,N_2053);
nand U3119 (N_3119,N_2763,N_2423);
nor U3120 (N_3120,N_2584,N_2638);
nand U3121 (N_3121,N_2164,N_2477);
and U3122 (N_3122,N_2039,N_2912);
xnor U3123 (N_3123,N_2484,N_2756);
nor U3124 (N_3124,N_2134,N_2445);
or U3125 (N_3125,N_2200,N_2848);
nor U3126 (N_3126,N_2112,N_2853);
nor U3127 (N_3127,N_2203,N_2311);
or U3128 (N_3128,N_2177,N_2010);
xor U3129 (N_3129,N_2032,N_2082);
xnor U3130 (N_3130,N_2470,N_2137);
nor U3131 (N_3131,N_2767,N_2150);
or U3132 (N_3132,N_2880,N_2811);
or U3133 (N_3133,N_2279,N_2106);
and U3134 (N_3134,N_2206,N_2110);
or U3135 (N_3135,N_2027,N_2446);
or U3136 (N_3136,N_2721,N_2356);
xor U3137 (N_3137,N_2172,N_2703);
xor U3138 (N_3138,N_2779,N_2736);
nor U3139 (N_3139,N_2332,N_2644);
or U3140 (N_3140,N_2344,N_2054);
xnor U3141 (N_3141,N_2526,N_2535);
nor U3142 (N_3142,N_2813,N_2545);
nor U3143 (N_3143,N_2396,N_2727);
and U3144 (N_3144,N_2021,N_2364);
nor U3145 (N_3145,N_2058,N_2873);
or U3146 (N_3146,N_2077,N_2993);
nor U3147 (N_3147,N_2938,N_2115);
and U3148 (N_3148,N_2733,N_2232);
and U3149 (N_3149,N_2226,N_2393);
nor U3150 (N_3150,N_2427,N_2968);
xnor U3151 (N_3151,N_2444,N_2047);
nand U3152 (N_3152,N_2849,N_2288);
and U3153 (N_3153,N_2654,N_2353);
or U3154 (N_3154,N_2932,N_2913);
or U3155 (N_3155,N_2296,N_2261);
or U3156 (N_3156,N_2476,N_2045);
nor U3157 (N_3157,N_2791,N_2982);
or U3158 (N_3158,N_2743,N_2013);
nor U3159 (N_3159,N_2453,N_2240);
and U3160 (N_3160,N_2450,N_2138);
or U3161 (N_3161,N_2854,N_2590);
nor U3162 (N_3162,N_2025,N_2120);
or U3163 (N_3163,N_2146,N_2454);
or U3164 (N_3164,N_2229,N_2923);
or U3165 (N_3165,N_2651,N_2495);
nand U3166 (N_3166,N_2363,N_2113);
nor U3167 (N_3167,N_2052,N_2298);
nand U3168 (N_3168,N_2921,N_2918);
or U3169 (N_3169,N_2957,N_2343);
nand U3170 (N_3170,N_2055,N_2438);
nor U3171 (N_3171,N_2728,N_2466);
nor U3172 (N_3172,N_2892,N_2761);
nand U3173 (N_3173,N_2281,N_2711);
or U3174 (N_3174,N_2028,N_2979);
nor U3175 (N_3175,N_2278,N_2606);
nor U3176 (N_3176,N_2614,N_2570);
or U3177 (N_3177,N_2034,N_2653);
nor U3178 (N_3178,N_2337,N_2316);
xor U3179 (N_3179,N_2607,N_2667);
and U3180 (N_3180,N_2844,N_2511);
and U3181 (N_3181,N_2542,N_2469);
or U3182 (N_3182,N_2833,N_2999);
or U3183 (N_3183,N_2946,N_2338);
and U3184 (N_3184,N_2124,N_2272);
xnor U3185 (N_3185,N_2707,N_2809);
or U3186 (N_3186,N_2642,N_2586);
or U3187 (N_3187,N_2744,N_2677);
nand U3188 (N_3188,N_2903,N_2775);
or U3189 (N_3189,N_2304,N_2241);
nand U3190 (N_3190,N_2289,N_2883);
and U3191 (N_3191,N_2493,N_2899);
or U3192 (N_3192,N_2070,N_2718);
nor U3193 (N_3193,N_2452,N_2182);
or U3194 (N_3194,N_2753,N_2144);
nand U3195 (N_3195,N_2560,N_2165);
nand U3196 (N_3196,N_2929,N_2961);
or U3197 (N_3197,N_2418,N_2689);
nor U3198 (N_3198,N_2683,N_2745);
nor U3199 (N_3199,N_2988,N_2568);
nor U3200 (N_3200,N_2299,N_2152);
nand U3201 (N_3201,N_2738,N_2199);
nand U3202 (N_3202,N_2778,N_2600);
or U3203 (N_3203,N_2333,N_2949);
nor U3204 (N_3204,N_2553,N_2391);
xor U3205 (N_3205,N_2400,N_2836);
xor U3206 (N_3206,N_2330,N_2451);
or U3207 (N_3207,N_2479,N_2816);
or U3208 (N_3208,N_2907,N_2981);
xor U3209 (N_3209,N_2313,N_2640);
and U3210 (N_3210,N_2491,N_2784);
or U3211 (N_3211,N_2832,N_2867);
xnor U3212 (N_3212,N_2524,N_2672);
and U3213 (N_3213,N_2178,N_2062);
xor U3214 (N_3214,N_2684,N_2771);
or U3215 (N_3215,N_2392,N_2117);
and U3216 (N_3216,N_2160,N_2682);
and U3217 (N_3217,N_2580,N_2523);
and U3218 (N_3218,N_2670,N_2195);
and U3219 (N_3219,N_2108,N_2031);
nand U3220 (N_3220,N_2704,N_2189);
xor U3221 (N_3221,N_2105,N_2390);
nor U3222 (N_3222,N_2507,N_2197);
nand U3223 (N_3223,N_2148,N_2582);
nor U3224 (N_3224,N_2415,N_2216);
nand U3225 (N_3225,N_2875,N_2383);
and U3226 (N_3226,N_2543,N_2503);
nand U3227 (N_3227,N_2360,N_2861);
and U3228 (N_3228,N_2369,N_2078);
nand U3229 (N_3229,N_2835,N_2702);
nand U3230 (N_3230,N_2955,N_2862);
nand U3231 (N_3231,N_2327,N_2619);
or U3232 (N_3232,N_2001,N_2894);
or U3233 (N_3233,N_2266,N_2528);
and U3234 (N_3234,N_2073,N_2740);
nor U3235 (N_3235,N_2227,N_2726);
and U3236 (N_3236,N_2191,N_2301);
or U3237 (N_3237,N_2345,N_2401);
and U3238 (N_3238,N_2659,N_2566);
nand U3239 (N_3239,N_2822,N_2171);
or U3240 (N_3240,N_2712,N_2852);
and U3241 (N_3241,N_2346,N_2910);
nand U3242 (N_3242,N_2119,N_2033);
nand U3243 (N_3243,N_2911,N_2219);
or U3244 (N_3244,N_2046,N_2870);
nand U3245 (N_3245,N_2887,N_2467);
nand U3246 (N_3246,N_2035,N_2049);
nand U3247 (N_3247,N_2886,N_2480);
and U3248 (N_3248,N_2643,N_2006);
nor U3249 (N_3249,N_2284,N_2314);
nor U3250 (N_3250,N_2890,N_2637);
nand U3251 (N_3251,N_2856,N_2462);
or U3252 (N_3252,N_2447,N_2259);
or U3253 (N_3253,N_2857,N_2845);
and U3254 (N_3254,N_2387,N_2839);
nor U3255 (N_3255,N_2326,N_2127);
or U3256 (N_3256,N_2253,N_2029);
xor U3257 (N_3257,N_2443,N_2591);
or U3258 (N_3258,N_2996,N_2739);
nand U3259 (N_3259,N_2896,N_2002);
nand U3260 (N_3260,N_2897,N_2351);
nor U3261 (N_3261,N_2136,N_2552);
and U3262 (N_3262,N_2558,N_2666);
nand U3263 (N_3263,N_2842,N_2630);
or U3264 (N_3264,N_2325,N_2131);
and U3265 (N_3265,N_2048,N_2671);
nand U3266 (N_3266,N_2114,N_2490);
xnor U3267 (N_3267,N_2472,N_2086);
nor U3268 (N_3268,N_2143,N_2563);
nand U3269 (N_3269,N_2188,N_2500);
nand U3270 (N_3270,N_2888,N_2688);
or U3271 (N_3271,N_2709,N_2205);
nor U3272 (N_3272,N_2043,N_2597);
and U3273 (N_3273,N_2224,N_2971);
nor U3274 (N_3274,N_2291,N_2239);
and U3275 (N_3275,N_2871,N_2797);
nor U3276 (N_3276,N_2762,N_2057);
or U3277 (N_3277,N_2290,N_2948);
or U3278 (N_3278,N_2922,N_2170);
nor U3279 (N_3279,N_2181,N_2411);
or U3280 (N_3280,N_2404,N_2075);
nor U3281 (N_3281,N_2422,N_2265);
nand U3282 (N_3282,N_2233,N_2679);
and U3283 (N_3283,N_2799,N_2319);
or U3284 (N_3284,N_2514,N_2676);
and U3285 (N_3285,N_2513,N_2126);
nor U3286 (N_3286,N_2550,N_2752);
and U3287 (N_3287,N_2192,N_2036);
nor U3288 (N_3288,N_2904,N_2690);
nand U3289 (N_3289,N_2385,N_2277);
nand U3290 (N_3290,N_2302,N_2693);
nand U3291 (N_3291,N_2416,N_2204);
and U3292 (N_3292,N_2094,N_2436);
xor U3293 (N_3293,N_2218,N_2645);
nand U3294 (N_3294,N_2365,N_2882);
and U3295 (N_3295,N_2575,N_2794);
nand U3296 (N_3296,N_2796,N_2354);
nor U3297 (N_3297,N_2331,N_2283);
nor U3298 (N_3298,N_2434,N_2287);
and U3299 (N_3299,N_2024,N_2336);
nor U3300 (N_3300,N_2901,N_2258);
or U3301 (N_3301,N_2787,N_2020);
and U3302 (N_3302,N_2366,N_2389);
and U3303 (N_3303,N_2931,N_2158);
and U3304 (N_3304,N_2846,N_2498);
and U3305 (N_3305,N_2044,N_2458);
and U3306 (N_3306,N_2782,N_2168);
and U3307 (N_3307,N_2612,N_2579);
and U3308 (N_3308,N_2710,N_2864);
nor U3309 (N_3309,N_2339,N_2305);
nand U3310 (N_3310,N_2940,N_2487);
or U3311 (N_3311,N_2139,N_2464);
and U3312 (N_3312,N_2292,N_2323);
nand U3313 (N_3313,N_2273,N_2803);
nor U3314 (N_3314,N_2309,N_2425);
nand U3315 (N_3315,N_2622,N_2238);
and U3316 (N_3316,N_2228,N_2174);
or U3317 (N_3317,N_2615,N_2924);
nand U3318 (N_3318,N_2128,N_2588);
nor U3319 (N_3319,N_2587,N_2732);
and U3320 (N_3320,N_2410,N_2657);
nor U3321 (N_3321,N_2668,N_2375);
nor U3322 (N_3322,N_2562,N_2914);
nor U3323 (N_3323,N_2417,N_2706);
nand U3324 (N_3324,N_2236,N_2474);
or U3325 (N_3325,N_2508,N_2403);
and U3326 (N_3326,N_2022,N_2985);
nand U3327 (N_3327,N_2781,N_2007);
or U3328 (N_3328,N_2186,N_2992);
nand U3329 (N_3329,N_2951,N_2944);
nor U3330 (N_3330,N_2059,N_2076);
or U3331 (N_3331,N_2051,N_2598);
nor U3332 (N_3332,N_2398,N_2101);
nor U3333 (N_3333,N_2754,N_2142);
nand U3334 (N_3334,N_2658,N_2463);
or U3335 (N_3335,N_2694,N_2155);
xnor U3336 (N_3336,N_2483,N_2394);
or U3337 (N_3337,N_2496,N_2962);
nor U3338 (N_3338,N_2840,N_2656);
xor U3339 (N_3339,N_2601,N_2956);
nor U3340 (N_3340,N_2858,N_2359);
nor U3341 (N_3341,N_2821,N_2167);
and U3342 (N_3342,N_2527,N_2673);
nand U3343 (N_3343,N_2793,N_2502);
nand U3344 (N_3344,N_2334,N_2998);
nor U3345 (N_3345,N_2091,N_2407);
nor U3346 (N_3346,N_2969,N_2536);
nor U3347 (N_3347,N_2571,N_2285);
and U3348 (N_3348,N_2270,N_2159);
nor U3349 (N_3349,N_2432,N_2634);
and U3350 (N_3350,N_2687,N_2166);
or U3351 (N_3351,N_2109,N_2574);
nand U3352 (N_3352,N_2397,N_2246);
nor U3353 (N_3353,N_2509,N_2494);
nor U3354 (N_3354,N_2724,N_2868);
nor U3355 (N_3355,N_2934,N_2196);
nand U3356 (N_3356,N_2312,N_2851);
and U3357 (N_3357,N_2198,N_2633);
xor U3358 (N_3358,N_2990,N_2989);
nand U3359 (N_3359,N_2308,N_2737);
nor U3360 (N_3360,N_2730,N_2428);
and U3361 (N_3361,N_2122,N_2014);
nand U3362 (N_3362,N_2185,N_2435);
nor U3363 (N_3363,N_2030,N_2789);
nand U3364 (N_3364,N_2161,N_2276);
or U3365 (N_3365,N_2263,N_2879);
and U3366 (N_3366,N_2522,N_2919);
and U3367 (N_3367,N_2686,N_2841);
or U3368 (N_3368,N_2759,N_2603);
nand U3369 (N_3369,N_2000,N_2040);
and U3370 (N_3370,N_2624,N_2162);
nand U3371 (N_3371,N_2157,N_2111);
and U3372 (N_3372,N_2605,N_2626);
or U3373 (N_3373,N_2708,N_2770);
and U3374 (N_3374,N_2828,N_2320);
nand U3375 (N_3375,N_2909,N_2549);
or U3376 (N_3376,N_2613,N_2604);
nand U3377 (N_3377,N_2650,N_2741);
and U3378 (N_3378,N_2749,N_2772);
and U3379 (N_3379,N_2578,N_2696);
nor U3380 (N_3380,N_2984,N_2475);
and U3381 (N_3381,N_2986,N_2608);
nor U3382 (N_3382,N_2945,N_2225);
nor U3383 (N_3383,N_2891,N_2977);
nor U3384 (N_3384,N_2050,N_2268);
nor U3385 (N_3385,N_2893,N_2627);
or U3386 (N_3386,N_2878,N_2457);
or U3387 (N_3387,N_2153,N_2610);
nand U3388 (N_3388,N_2954,N_2800);
nor U3389 (N_3389,N_2250,N_2256);
and U3390 (N_3390,N_2099,N_2234);
nand U3391 (N_3391,N_2123,N_2933);
xnor U3392 (N_3392,N_2664,N_2088);
and U3393 (N_3393,N_2554,N_2652);
nand U3394 (N_3394,N_2978,N_2639);
nand U3395 (N_3395,N_2248,N_2860);
or U3396 (N_3396,N_2011,N_2212);
nor U3397 (N_3397,N_2376,N_2669);
or U3398 (N_3398,N_2074,N_2595);
and U3399 (N_3399,N_2625,N_2017);
nand U3400 (N_3400,N_2768,N_2441);
nand U3401 (N_3401,N_2831,N_2395);
nand U3402 (N_3402,N_2559,N_2540);
xnor U3403 (N_3403,N_2439,N_2539);
nor U3404 (N_3404,N_2202,N_2952);
nor U3405 (N_3405,N_2785,N_2850);
or U3406 (N_3406,N_2286,N_2408);
and U3407 (N_3407,N_2648,N_2349);
xnor U3408 (N_3408,N_2098,N_2015);
nand U3409 (N_3409,N_2374,N_2294);
nor U3410 (N_3410,N_2087,N_2179);
nand U3411 (N_3411,N_2975,N_2537);
nor U3412 (N_3412,N_2812,N_2818);
or U3413 (N_3413,N_2460,N_2662);
nor U3414 (N_3414,N_2175,N_2081);
and U3415 (N_3415,N_2925,N_2280);
nand U3416 (N_3416,N_2169,N_2786);
nand U3417 (N_3417,N_2116,N_2207);
nand U3418 (N_3418,N_2581,N_2402);
or U3419 (N_3419,N_2865,N_2409);
xor U3420 (N_3420,N_2872,N_2611);
nor U3421 (N_3421,N_2599,N_2746);
and U3422 (N_3422,N_2066,N_2008);
or U3423 (N_3423,N_2714,N_2973);
or U3424 (N_3424,N_2471,N_2440);
xnor U3425 (N_3425,N_2104,N_2388);
or U3426 (N_3426,N_2064,N_2674);
xor U3427 (N_3427,N_2717,N_2817);
nand U3428 (N_3428,N_2211,N_2295);
nor U3429 (N_3429,N_2340,N_2815);
nand U3430 (N_3430,N_2678,N_2548);
and U3431 (N_3431,N_2681,N_2230);
xor U3432 (N_3432,N_2252,N_2655);
or U3433 (N_3433,N_2725,N_2544);
nand U3434 (N_3434,N_2583,N_2005);
or U3435 (N_3435,N_2317,N_2546);
or U3436 (N_3436,N_2847,N_2631);
or U3437 (N_3437,N_2489,N_2855);
nor U3438 (N_3438,N_2557,N_2482);
nand U3439 (N_3439,N_2742,N_2282);
nand U3440 (N_3440,N_2242,N_2808);
nand U3441 (N_3441,N_2096,N_2596);
xor U3442 (N_3442,N_2310,N_2927);
nand U3443 (N_3443,N_2187,N_2067);
and U3444 (N_3444,N_2069,N_2632);
and U3445 (N_3445,N_2609,N_2149);
xor U3446 (N_3446,N_2135,N_2231);
or U3447 (N_3447,N_2783,N_2691);
and U3448 (N_3448,N_2941,N_2819);
or U3449 (N_3449,N_2814,N_2254);
nor U3450 (N_3450,N_2506,N_2429);
or U3451 (N_3451,N_2237,N_2533);
or U3452 (N_3452,N_2790,N_2824);
nor U3453 (N_3453,N_2156,N_2991);
and U3454 (N_3454,N_2731,N_2660);
and U3455 (N_3455,N_2577,N_2926);
and U3456 (N_3456,N_2378,N_2766);
nor U3457 (N_3457,N_2720,N_2716);
and U3458 (N_3458,N_2963,N_2501);
nand U3459 (N_3459,N_2012,N_2760);
nand U3460 (N_3460,N_2869,N_2406);
nor U3461 (N_3461,N_2930,N_2802);
xor U3462 (N_3462,N_2505,N_2468);
or U3463 (N_3463,N_2755,N_2825);
and U3464 (N_3464,N_2026,N_2942);
xnor U3465 (N_3465,N_2525,N_2492);
xor U3466 (N_3466,N_2701,N_2065);
nand U3467 (N_3467,N_2084,N_2449);
nor U3468 (N_3468,N_2573,N_2788);
nor U3469 (N_3469,N_2221,N_2512);
or U3470 (N_3470,N_2132,N_2459);
nor U3471 (N_3471,N_2368,N_2357);
nand U3472 (N_3472,N_2260,N_2972);
or U3473 (N_3473,N_2275,N_2456);
or U3474 (N_3474,N_2551,N_2906);
and U3475 (N_3475,N_2213,N_2900);
xnor U3476 (N_3476,N_2735,N_2324);
nand U3477 (N_3477,N_2713,N_2145);
and U3478 (N_3478,N_2898,N_2966);
nand U3479 (N_3479,N_2936,N_2041);
xnor U3480 (N_3480,N_2859,N_2215);
nor U3481 (N_3481,N_2352,N_2965);
nand U3482 (N_3482,N_2823,N_2341);
and U3483 (N_3483,N_2569,N_2769);
and U3484 (N_3484,N_2056,N_2133);
or U3485 (N_3485,N_2529,N_2307);
or U3486 (N_3486,N_2895,N_2692);
nand U3487 (N_3487,N_2141,N_2358);
or U3488 (N_3488,N_2995,N_2504);
nor U3489 (N_3489,N_2061,N_2399);
and U3490 (N_3490,N_2420,N_2222);
and U3491 (N_3491,N_2249,N_2414);
or U3492 (N_3492,N_2876,N_2937);
nand U3493 (N_3493,N_2843,N_2646);
nor U3494 (N_3494,N_2564,N_2348);
and U3495 (N_3495,N_2184,N_2431);
xor U3496 (N_3496,N_2519,N_2103);
nand U3497 (N_3497,N_2534,N_2807);
or U3498 (N_3498,N_2437,N_2953);
and U3499 (N_3499,N_2777,N_2426);
or U3500 (N_3500,N_2148,N_2089);
or U3501 (N_3501,N_2664,N_2430);
or U3502 (N_3502,N_2672,N_2522);
and U3503 (N_3503,N_2624,N_2464);
and U3504 (N_3504,N_2634,N_2485);
or U3505 (N_3505,N_2060,N_2235);
and U3506 (N_3506,N_2814,N_2182);
and U3507 (N_3507,N_2812,N_2929);
or U3508 (N_3508,N_2310,N_2567);
or U3509 (N_3509,N_2497,N_2965);
nand U3510 (N_3510,N_2203,N_2932);
nor U3511 (N_3511,N_2237,N_2993);
nand U3512 (N_3512,N_2909,N_2346);
nand U3513 (N_3513,N_2884,N_2755);
nor U3514 (N_3514,N_2839,N_2200);
nor U3515 (N_3515,N_2930,N_2739);
nor U3516 (N_3516,N_2840,N_2812);
and U3517 (N_3517,N_2514,N_2286);
nand U3518 (N_3518,N_2378,N_2352);
nand U3519 (N_3519,N_2397,N_2464);
xor U3520 (N_3520,N_2827,N_2665);
nand U3521 (N_3521,N_2731,N_2334);
nand U3522 (N_3522,N_2085,N_2420);
or U3523 (N_3523,N_2991,N_2385);
nor U3524 (N_3524,N_2691,N_2672);
or U3525 (N_3525,N_2170,N_2694);
and U3526 (N_3526,N_2652,N_2344);
and U3527 (N_3527,N_2633,N_2620);
and U3528 (N_3528,N_2717,N_2008);
nand U3529 (N_3529,N_2961,N_2932);
and U3530 (N_3530,N_2536,N_2646);
or U3531 (N_3531,N_2353,N_2210);
nor U3532 (N_3532,N_2701,N_2041);
nor U3533 (N_3533,N_2795,N_2572);
nand U3534 (N_3534,N_2171,N_2663);
nor U3535 (N_3535,N_2679,N_2598);
nand U3536 (N_3536,N_2006,N_2082);
or U3537 (N_3537,N_2111,N_2680);
nor U3538 (N_3538,N_2840,N_2549);
xnor U3539 (N_3539,N_2331,N_2135);
or U3540 (N_3540,N_2234,N_2053);
nand U3541 (N_3541,N_2622,N_2087);
or U3542 (N_3542,N_2642,N_2561);
or U3543 (N_3543,N_2809,N_2408);
nor U3544 (N_3544,N_2322,N_2920);
nor U3545 (N_3545,N_2444,N_2470);
or U3546 (N_3546,N_2694,N_2237);
nand U3547 (N_3547,N_2316,N_2533);
or U3548 (N_3548,N_2774,N_2304);
or U3549 (N_3549,N_2626,N_2155);
nand U3550 (N_3550,N_2812,N_2693);
or U3551 (N_3551,N_2365,N_2101);
nor U3552 (N_3552,N_2889,N_2993);
nand U3553 (N_3553,N_2155,N_2530);
or U3554 (N_3554,N_2789,N_2266);
and U3555 (N_3555,N_2715,N_2616);
or U3556 (N_3556,N_2126,N_2082);
xnor U3557 (N_3557,N_2004,N_2226);
nand U3558 (N_3558,N_2086,N_2485);
nand U3559 (N_3559,N_2564,N_2630);
nand U3560 (N_3560,N_2687,N_2024);
and U3561 (N_3561,N_2222,N_2436);
or U3562 (N_3562,N_2647,N_2872);
nand U3563 (N_3563,N_2880,N_2612);
nand U3564 (N_3564,N_2294,N_2427);
nor U3565 (N_3565,N_2676,N_2853);
or U3566 (N_3566,N_2617,N_2552);
or U3567 (N_3567,N_2840,N_2613);
and U3568 (N_3568,N_2832,N_2459);
and U3569 (N_3569,N_2949,N_2204);
nor U3570 (N_3570,N_2253,N_2216);
nor U3571 (N_3571,N_2238,N_2936);
or U3572 (N_3572,N_2488,N_2435);
nor U3573 (N_3573,N_2336,N_2541);
xor U3574 (N_3574,N_2918,N_2654);
and U3575 (N_3575,N_2623,N_2180);
nor U3576 (N_3576,N_2223,N_2989);
or U3577 (N_3577,N_2124,N_2949);
nor U3578 (N_3578,N_2273,N_2413);
nand U3579 (N_3579,N_2309,N_2986);
or U3580 (N_3580,N_2400,N_2462);
nand U3581 (N_3581,N_2049,N_2900);
and U3582 (N_3582,N_2501,N_2883);
or U3583 (N_3583,N_2165,N_2118);
or U3584 (N_3584,N_2346,N_2948);
nand U3585 (N_3585,N_2676,N_2936);
nor U3586 (N_3586,N_2713,N_2136);
nor U3587 (N_3587,N_2588,N_2948);
and U3588 (N_3588,N_2128,N_2333);
and U3589 (N_3589,N_2607,N_2605);
nor U3590 (N_3590,N_2897,N_2102);
or U3591 (N_3591,N_2054,N_2294);
nor U3592 (N_3592,N_2142,N_2479);
nor U3593 (N_3593,N_2243,N_2783);
xnor U3594 (N_3594,N_2852,N_2771);
or U3595 (N_3595,N_2530,N_2949);
or U3596 (N_3596,N_2247,N_2376);
nand U3597 (N_3597,N_2147,N_2464);
nor U3598 (N_3598,N_2080,N_2525);
and U3599 (N_3599,N_2254,N_2282);
nand U3600 (N_3600,N_2824,N_2732);
or U3601 (N_3601,N_2446,N_2151);
nand U3602 (N_3602,N_2213,N_2991);
xnor U3603 (N_3603,N_2283,N_2423);
nand U3604 (N_3604,N_2346,N_2772);
and U3605 (N_3605,N_2789,N_2118);
or U3606 (N_3606,N_2858,N_2099);
nor U3607 (N_3607,N_2260,N_2988);
and U3608 (N_3608,N_2097,N_2198);
nor U3609 (N_3609,N_2699,N_2117);
nor U3610 (N_3610,N_2259,N_2423);
nor U3611 (N_3611,N_2366,N_2355);
nand U3612 (N_3612,N_2631,N_2244);
or U3613 (N_3613,N_2435,N_2098);
xor U3614 (N_3614,N_2757,N_2548);
xnor U3615 (N_3615,N_2162,N_2399);
nor U3616 (N_3616,N_2686,N_2422);
nor U3617 (N_3617,N_2582,N_2534);
xor U3618 (N_3618,N_2855,N_2107);
or U3619 (N_3619,N_2596,N_2433);
nor U3620 (N_3620,N_2028,N_2296);
nand U3621 (N_3621,N_2006,N_2785);
nor U3622 (N_3622,N_2802,N_2607);
nand U3623 (N_3623,N_2695,N_2260);
and U3624 (N_3624,N_2705,N_2292);
nand U3625 (N_3625,N_2118,N_2858);
xor U3626 (N_3626,N_2480,N_2426);
nor U3627 (N_3627,N_2323,N_2055);
and U3628 (N_3628,N_2349,N_2632);
nand U3629 (N_3629,N_2918,N_2583);
and U3630 (N_3630,N_2168,N_2060);
nor U3631 (N_3631,N_2435,N_2047);
nand U3632 (N_3632,N_2060,N_2595);
xor U3633 (N_3633,N_2680,N_2404);
and U3634 (N_3634,N_2805,N_2552);
nand U3635 (N_3635,N_2660,N_2434);
or U3636 (N_3636,N_2569,N_2670);
nand U3637 (N_3637,N_2063,N_2208);
or U3638 (N_3638,N_2613,N_2228);
nand U3639 (N_3639,N_2210,N_2376);
nor U3640 (N_3640,N_2032,N_2099);
and U3641 (N_3641,N_2454,N_2689);
nor U3642 (N_3642,N_2136,N_2897);
nor U3643 (N_3643,N_2850,N_2934);
xnor U3644 (N_3644,N_2617,N_2105);
xor U3645 (N_3645,N_2589,N_2426);
nand U3646 (N_3646,N_2200,N_2930);
or U3647 (N_3647,N_2521,N_2554);
and U3648 (N_3648,N_2176,N_2391);
nor U3649 (N_3649,N_2824,N_2751);
and U3650 (N_3650,N_2807,N_2145);
and U3651 (N_3651,N_2871,N_2175);
nand U3652 (N_3652,N_2308,N_2635);
nand U3653 (N_3653,N_2621,N_2099);
and U3654 (N_3654,N_2041,N_2619);
nor U3655 (N_3655,N_2437,N_2985);
nand U3656 (N_3656,N_2856,N_2124);
nand U3657 (N_3657,N_2989,N_2051);
xor U3658 (N_3658,N_2824,N_2411);
and U3659 (N_3659,N_2140,N_2992);
or U3660 (N_3660,N_2379,N_2195);
or U3661 (N_3661,N_2943,N_2194);
and U3662 (N_3662,N_2925,N_2292);
nor U3663 (N_3663,N_2115,N_2277);
and U3664 (N_3664,N_2055,N_2860);
and U3665 (N_3665,N_2864,N_2450);
nor U3666 (N_3666,N_2270,N_2476);
xor U3667 (N_3667,N_2160,N_2839);
xnor U3668 (N_3668,N_2176,N_2048);
or U3669 (N_3669,N_2466,N_2656);
and U3670 (N_3670,N_2816,N_2905);
xor U3671 (N_3671,N_2493,N_2705);
nor U3672 (N_3672,N_2211,N_2592);
xnor U3673 (N_3673,N_2768,N_2802);
nand U3674 (N_3674,N_2910,N_2829);
nand U3675 (N_3675,N_2892,N_2742);
nand U3676 (N_3676,N_2440,N_2489);
xor U3677 (N_3677,N_2220,N_2055);
nor U3678 (N_3678,N_2136,N_2135);
nor U3679 (N_3679,N_2402,N_2191);
nor U3680 (N_3680,N_2041,N_2520);
and U3681 (N_3681,N_2696,N_2887);
or U3682 (N_3682,N_2426,N_2174);
nand U3683 (N_3683,N_2889,N_2803);
nand U3684 (N_3684,N_2010,N_2633);
and U3685 (N_3685,N_2592,N_2061);
nand U3686 (N_3686,N_2199,N_2200);
nand U3687 (N_3687,N_2679,N_2989);
nand U3688 (N_3688,N_2407,N_2509);
or U3689 (N_3689,N_2012,N_2068);
nand U3690 (N_3690,N_2920,N_2526);
or U3691 (N_3691,N_2271,N_2687);
nand U3692 (N_3692,N_2728,N_2713);
nand U3693 (N_3693,N_2461,N_2501);
or U3694 (N_3694,N_2269,N_2758);
or U3695 (N_3695,N_2270,N_2338);
xor U3696 (N_3696,N_2288,N_2686);
nor U3697 (N_3697,N_2992,N_2834);
nand U3698 (N_3698,N_2065,N_2141);
or U3699 (N_3699,N_2657,N_2584);
and U3700 (N_3700,N_2805,N_2684);
or U3701 (N_3701,N_2420,N_2892);
or U3702 (N_3702,N_2502,N_2951);
and U3703 (N_3703,N_2885,N_2120);
and U3704 (N_3704,N_2084,N_2514);
nand U3705 (N_3705,N_2979,N_2382);
or U3706 (N_3706,N_2024,N_2293);
or U3707 (N_3707,N_2648,N_2845);
nor U3708 (N_3708,N_2531,N_2509);
and U3709 (N_3709,N_2455,N_2398);
xnor U3710 (N_3710,N_2052,N_2968);
nor U3711 (N_3711,N_2960,N_2277);
nor U3712 (N_3712,N_2928,N_2458);
nor U3713 (N_3713,N_2867,N_2388);
and U3714 (N_3714,N_2261,N_2341);
or U3715 (N_3715,N_2027,N_2872);
nor U3716 (N_3716,N_2032,N_2150);
nand U3717 (N_3717,N_2640,N_2116);
nor U3718 (N_3718,N_2032,N_2989);
nand U3719 (N_3719,N_2214,N_2544);
nand U3720 (N_3720,N_2813,N_2968);
nor U3721 (N_3721,N_2100,N_2407);
nor U3722 (N_3722,N_2514,N_2769);
nand U3723 (N_3723,N_2033,N_2373);
and U3724 (N_3724,N_2790,N_2443);
or U3725 (N_3725,N_2306,N_2625);
nor U3726 (N_3726,N_2440,N_2876);
or U3727 (N_3727,N_2402,N_2352);
nand U3728 (N_3728,N_2923,N_2350);
and U3729 (N_3729,N_2709,N_2577);
or U3730 (N_3730,N_2101,N_2916);
or U3731 (N_3731,N_2034,N_2379);
nor U3732 (N_3732,N_2795,N_2594);
nor U3733 (N_3733,N_2956,N_2834);
and U3734 (N_3734,N_2076,N_2093);
nand U3735 (N_3735,N_2357,N_2401);
xor U3736 (N_3736,N_2911,N_2994);
and U3737 (N_3737,N_2248,N_2108);
or U3738 (N_3738,N_2167,N_2671);
nand U3739 (N_3739,N_2273,N_2951);
or U3740 (N_3740,N_2559,N_2256);
nor U3741 (N_3741,N_2257,N_2379);
nand U3742 (N_3742,N_2963,N_2589);
xnor U3743 (N_3743,N_2372,N_2674);
and U3744 (N_3744,N_2036,N_2936);
nor U3745 (N_3745,N_2031,N_2611);
nand U3746 (N_3746,N_2379,N_2209);
or U3747 (N_3747,N_2204,N_2500);
and U3748 (N_3748,N_2713,N_2284);
or U3749 (N_3749,N_2267,N_2499);
nand U3750 (N_3750,N_2889,N_2567);
or U3751 (N_3751,N_2351,N_2391);
xnor U3752 (N_3752,N_2624,N_2943);
nand U3753 (N_3753,N_2163,N_2348);
or U3754 (N_3754,N_2221,N_2076);
or U3755 (N_3755,N_2947,N_2347);
nor U3756 (N_3756,N_2329,N_2743);
xor U3757 (N_3757,N_2606,N_2099);
or U3758 (N_3758,N_2661,N_2487);
nor U3759 (N_3759,N_2626,N_2956);
and U3760 (N_3760,N_2468,N_2333);
or U3761 (N_3761,N_2345,N_2029);
or U3762 (N_3762,N_2770,N_2397);
and U3763 (N_3763,N_2535,N_2746);
and U3764 (N_3764,N_2667,N_2268);
or U3765 (N_3765,N_2163,N_2657);
nor U3766 (N_3766,N_2824,N_2380);
xnor U3767 (N_3767,N_2267,N_2178);
or U3768 (N_3768,N_2452,N_2150);
or U3769 (N_3769,N_2105,N_2553);
nand U3770 (N_3770,N_2646,N_2455);
and U3771 (N_3771,N_2532,N_2314);
and U3772 (N_3772,N_2009,N_2188);
xor U3773 (N_3773,N_2626,N_2792);
nand U3774 (N_3774,N_2867,N_2725);
nor U3775 (N_3775,N_2970,N_2291);
nor U3776 (N_3776,N_2688,N_2976);
nand U3777 (N_3777,N_2838,N_2957);
xnor U3778 (N_3778,N_2680,N_2145);
or U3779 (N_3779,N_2376,N_2758);
nor U3780 (N_3780,N_2937,N_2921);
xor U3781 (N_3781,N_2710,N_2333);
xor U3782 (N_3782,N_2650,N_2064);
nor U3783 (N_3783,N_2652,N_2500);
and U3784 (N_3784,N_2058,N_2645);
and U3785 (N_3785,N_2289,N_2739);
nor U3786 (N_3786,N_2905,N_2595);
or U3787 (N_3787,N_2099,N_2947);
nand U3788 (N_3788,N_2758,N_2283);
nand U3789 (N_3789,N_2229,N_2566);
xnor U3790 (N_3790,N_2246,N_2721);
and U3791 (N_3791,N_2438,N_2014);
nor U3792 (N_3792,N_2569,N_2641);
or U3793 (N_3793,N_2060,N_2178);
or U3794 (N_3794,N_2816,N_2554);
or U3795 (N_3795,N_2068,N_2015);
and U3796 (N_3796,N_2148,N_2866);
and U3797 (N_3797,N_2071,N_2777);
and U3798 (N_3798,N_2230,N_2143);
and U3799 (N_3799,N_2707,N_2107);
or U3800 (N_3800,N_2034,N_2324);
nor U3801 (N_3801,N_2655,N_2727);
nand U3802 (N_3802,N_2482,N_2003);
nand U3803 (N_3803,N_2790,N_2008);
and U3804 (N_3804,N_2098,N_2183);
and U3805 (N_3805,N_2027,N_2926);
nand U3806 (N_3806,N_2590,N_2023);
or U3807 (N_3807,N_2995,N_2641);
or U3808 (N_3808,N_2650,N_2158);
xor U3809 (N_3809,N_2834,N_2486);
nand U3810 (N_3810,N_2062,N_2803);
or U3811 (N_3811,N_2138,N_2545);
or U3812 (N_3812,N_2319,N_2464);
and U3813 (N_3813,N_2596,N_2616);
nand U3814 (N_3814,N_2507,N_2608);
xor U3815 (N_3815,N_2101,N_2384);
nor U3816 (N_3816,N_2889,N_2895);
or U3817 (N_3817,N_2729,N_2457);
or U3818 (N_3818,N_2018,N_2867);
xor U3819 (N_3819,N_2023,N_2834);
or U3820 (N_3820,N_2908,N_2900);
or U3821 (N_3821,N_2175,N_2141);
nor U3822 (N_3822,N_2402,N_2983);
or U3823 (N_3823,N_2206,N_2464);
and U3824 (N_3824,N_2717,N_2744);
nor U3825 (N_3825,N_2174,N_2239);
or U3826 (N_3826,N_2162,N_2708);
or U3827 (N_3827,N_2426,N_2703);
and U3828 (N_3828,N_2456,N_2496);
nand U3829 (N_3829,N_2475,N_2326);
nand U3830 (N_3830,N_2617,N_2402);
nand U3831 (N_3831,N_2016,N_2160);
and U3832 (N_3832,N_2861,N_2833);
and U3833 (N_3833,N_2710,N_2385);
nor U3834 (N_3834,N_2448,N_2693);
and U3835 (N_3835,N_2790,N_2507);
nor U3836 (N_3836,N_2263,N_2868);
or U3837 (N_3837,N_2477,N_2923);
and U3838 (N_3838,N_2854,N_2084);
nand U3839 (N_3839,N_2457,N_2246);
nand U3840 (N_3840,N_2511,N_2887);
xor U3841 (N_3841,N_2345,N_2463);
or U3842 (N_3842,N_2603,N_2524);
or U3843 (N_3843,N_2263,N_2086);
or U3844 (N_3844,N_2344,N_2288);
and U3845 (N_3845,N_2505,N_2081);
or U3846 (N_3846,N_2434,N_2572);
nor U3847 (N_3847,N_2312,N_2787);
or U3848 (N_3848,N_2923,N_2028);
nor U3849 (N_3849,N_2070,N_2387);
or U3850 (N_3850,N_2782,N_2575);
and U3851 (N_3851,N_2855,N_2720);
or U3852 (N_3852,N_2091,N_2318);
nor U3853 (N_3853,N_2701,N_2216);
xor U3854 (N_3854,N_2598,N_2530);
and U3855 (N_3855,N_2798,N_2749);
nand U3856 (N_3856,N_2778,N_2806);
nand U3857 (N_3857,N_2373,N_2333);
nor U3858 (N_3858,N_2424,N_2518);
nor U3859 (N_3859,N_2538,N_2260);
or U3860 (N_3860,N_2971,N_2544);
nor U3861 (N_3861,N_2742,N_2337);
or U3862 (N_3862,N_2393,N_2390);
nor U3863 (N_3863,N_2648,N_2392);
and U3864 (N_3864,N_2886,N_2789);
or U3865 (N_3865,N_2204,N_2165);
nand U3866 (N_3866,N_2518,N_2709);
nor U3867 (N_3867,N_2011,N_2771);
nor U3868 (N_3868,N_2162,N_2608);
or U3869 (N_3869,N_2273,N_2541);
nand U3870 (N_3870,N_2772,N_2548);
nor U3871 (N_3871,N_2012,N_2629);
and U3872 (N_3872,N_2782,N_2786);
or U3873 (N_3873,N_2361,N_2206);
and U3874 (N_3874,N_2773,N_2913);
and U3875 (N_3875,N_2282,N_2530);
nand U3876 (N_3876,N_2954,N_2711);
nor U3877 (N_3877,N_2330,N_2152);
nor U3878 (N_3878,N_2769,N_2515);
nor U3879 (N_3879,N_2515,N_2445);
and U3880 (N_3880,N_2395,N_2155);
nor U3881 (N_3881,N_2613,N_2099);
and U3882 (N_3882,N_2145,N_2622);
or U3883 (N_3883,N_2895,N_2325);
xor U3884 (N_3884,N_2606,N_2484);
nor U3885 (N_3885,N_2646,N_2308);
nor U3886 (N_3886,N_2347,N_2965);
nand U3887 (N_3887,N_2948,N_2320);
or U3888 (N_3888,N_2540,N_2421);
and U3889 (N_3889,N_2413,N_2838);
and U3890 (N_3890,N_2764,N_2778);
and U3891 (N_3891,N_2009,N_2439);
or U3892 (N_3892,N_2875,N_2211);
or U3893 (N_3893,N_2720,N_2750);
nand U3894 (N_3894,N_2368,N_2003);
or U3895 (N_3895,N_2400,N_2459);
nand U3896 (N_3896,N_2102,N_2700);
or U3897 (N_3897,N_2714,N_2531);
xor U3898 (N_3898,N_2936,N_2980);
nor U3899 (N_3899,N_2310,N_2972);
xor U3900 (N_3900,N_2339,N_2314);
nand U3901 (N_3901,N_2646,N_2902);
nor U3902 (N_3902,N_2427,N_2016);
nor U3903 (N_3903,N_2617,N_2222);
xor U3904 (N_3904,N_2643,N_2287);
or U3905 (N_3905,N_2284,N_2418);
nor U3906 (N_3906,N_2910,N_2307);
and U3907 (N_3907,N_2255,N_2505);
nor U3908 (N_3908,N_2260,N_2576);
and U3909 (N_3909,N_2435,N_2607);
nor U3910 (N_3910,N_2277,N_2974);
xnor U3911 (N_3911,N_2967,N_2931);
nand U3912 (N_3912,N_2423,N_2398);
and U3913 (N_3913,N_2581,N_2847);
and U3914 (N_3914,N_2526,N_2301);
xnor U3915 (N_3915,N_2683,N_2565);
nor U3916 (N_3916,N_2275,N_2728);
or U3917 (N_3917,N_2759,N_2791);
or U3918 (N_3918,N_2804,N_2846);
or U3919 (N_3919,N_2130,N_2150);
nor U3920 (N_3920,N_2803,N_2011);
or U3921 (N_3921,N_2189,N_2418);
or U3922 (N_3922,N_2648,N_2871);
and U3923 (N_3923,N_2328,N_2579);
and U3924 (N_3924,N_2205,N_2518);
and U3925 (N_3925,N_2648,N_2618);
or U3926 (N_3926,N_2144,N_2845);
and U3927 (N_3927,N_2042,N_2890);
xor U3928 (N_3928,N_2672,N_2275);
nor U3929 (N_3929,N_2583,N_2550);
xnor U3930 (N_3930,N_2300,N_2157);
and U3931 (N_3931,N_2763,N_2521);
nor U3932 (N_3932,N_2214,N_2351);
and U3933 (N_3933,N_2654,N_2343);
nor U3934 (N_3934,N_2214,N_2629);
or U3935 (N_3935,N_2089,N_2766);
nand U3936 (N_3936,N_2343,N_2212);
xnor U3937 (N_3937,N_2891,N_2515);
nand U3938 (N_3938,N_2312,N_2333);
nor U3939 (N_3939,N_2634,N_2530);
nand U3940 (N_3940,N_2821,N_2884);
nor U3941 (N_3941,N_2529,N_2055);
nor U3942 (N_3942,N_2090,N_2963);
nand U3943 (N_3943,N_2892,N_2008);
xnor U3944 (N_3944,N_2638,N_2068);
xnor U3945 (N_3945,N_2345,N_2914);
nor U3946 (N_3946,N_2832,N_2078);
or U3947 (N_3947,N_2884,N_2671);
nor U3948 (N_3948,N_2835,N_2766);
nand U3949 (N_3949,N_2591,N_2018);
or U3950 (N_3950,N_2734,N_2155);
or U3951 (N_3951,N_2746,N_2120);
xnor U3952 (N_3952,N_2208,N_2707);
nand U3953 (N_3953,N_2007,N_2068);
nor U3954 (N_3954,N_2508,N_2099);
nand U3955 (N_3955,N_2281,N_2847);
and U3956 (N_3956,N_2231,N_2431);
nor U3957 (N_3957,N_2522,N_2678);
and U3958 (N_3958,N_2052,N_2873);
nor U3959 (N_3959,N_2751,N_2397);
nor U3960 (N_3960,N_2838,N_2380);
nand U3961 (N_3961,N_2378,N_2206);
nand U3962 (N_3962,N_2739,N_2696);
nor U3963 (N_3963,N_2952,N_2041);
and U3964 (N_3964,N_2723,N_2977);
and U3965 (N_3965,N_2201,N_2452);
nor U3966 (N_3966,N_2418,N_2134);
nor U3967 (N_3967,N_2916,N_2165);
or U3968 (N_3968,N_2215,N_2943);
nand U3969 (N_3969,N_2093,N_2146);
or U3970 (N_3970,N_2585,N_2775);
nand U3971 (N_3971,N_2185,N_2008);
or U3972 (N_3972,N_2527,N_2386);
nand U3973 (N_3973,N_2792,N_2564);
nand U3974 (N_3974,N_2037,N_2046);
nor U3975 (N_3975,N_2656,N_2789);
or U3976 (N_3976,N_2101,N_2299);
or U3977 (N_3977,N_2021,N_2403);
nor U3978 (N_3978,N_2685,N_2698);
nor U3979 (N_3979,N_2012,N_2657);
or U3980 (N_3980,N_2640,N_2866);
and U3981 (N_3981,N_2438,N_2661);
nor U3982 (N_3982,N_2191,N_2188);
or U3983 (N_3983,N_2821,N_2798);
nor U3984 (N_3984,N_2339,N_2157);
nand U3985 (N_3985,N_2236,N_2161);
xor U3986 (N_3986,N_2998,N_2053);
nand U3987 (N_3987,N_2139,N_2419);
nor U3988 (N_3988,N_2399,N_2481);
nor U3989 (N_3989,N_2030,N_2673);
nand U3990 (N_3990,N_2475,N_2110);
nand U3991 (N_3991,N_2948,N_2925);
or U3992 (N_3992,N_2597,N_2673);
nor U3993 (N_3993,N_2900,N_2250);
nand U3994 (N_3994,N_2176,N_2273);
or U3995 (N_3995,N_2889,N_2608);
and U3996 (N_3996,N_2136,N_2874);
nand U3997 (N_3997,N_2518,N_2358);
nand U3998 (N_3998,N_2291,N_2809);
and U3999 (N_3999,N_2718,N_2638);
nand U4000 (N_4000,N_3936,N_3660);
nor U4001 (N_4001,N_3545,N_3135);
and U4002 (N_4002,N_3589,N_3709);
and U4003 (N_4003,N_3512,N_3729);
or U4004 (N_4004,N_3262,N_3178);
nand U4005 (N_4005,N_3510,N_3854);
and U4006 (N_4006,N_3043,N_3045);
and U4007 (N_4007,N_3464,N_3669);
or U4008 (N_4008,N_3006,N_3180);
and U4009 (N_4009,N_3557,N_3711);
and U4010 (N_4010,N_3395,N_3671);
nor U4011 (N_4011,N_3419,N_3315);
nor U4012 (N_4012,N_3573,N_3959);
and U4013 (N_4013,N_3962,N_3456);
or U4014 (N_4014,N_3868,N_3275);
and U4015 (N_4015,N_3703,N_3147);
nor U4016 (N_4016,N_3287,N_3273);
nand U4017 (N_4017,N_3359,N_3129);
and U4018 (N_4018,N_3363,N_3821);
nand U4019 (N_4019,N_3564,N_3004);
and U4020 (N_4020,N_3836,N_3839);
and U4021 (N_4021,N_3768,N_3439);
nor U4022 (N_4022,N_3370,N_3113);
nor U4023 (N_4023,N_3747,N_3442);
xor U4024 (N_4024,N_3975,N_3141);
or U4025 (N_4025,N_3591,N_3846);
or U4026 (N_4026,N_3584,N_3354);
or U4027 (N_4027,N_3949,N_3222);
or U4028 (N_4028,N_3960,N_3505);
and U4029 (N_4029,N_3320,N_3683);
nor U4030 (N_4030,N_3025,N_3874);
and U4031 (N_4031,N_3264,N_3828);
nand U4032 (N_4032,N_3724,N_3504);
nor U4033 (N_4033,N_3713,N_3356);
nor U4034 (N_4034,N_3654,N_3843);
and U4035 (N_4035,N_3385,N_3721);
nor U4036 (N_4036,N_3571,N_3106);
or U4037 (N_4037,N_3842,N_3666);
or U4038 (N_4038,N_3070,N_3636);
nor U4039 (N_4039,N_3425,N_3668);
or U4040 (N_4040,N_3769,N_3398);
or U4041 (N_4041,N_3110,N_3487);
or U4042 (N_4042,N_3736,N_3889);
nand U4043 (N_4043,N_3390,N_3224);
nor U4044 (N_4044,N_3463,N_3190);
xor U4045 (N_4045,N_3026,N_3319);
nor U4046 (N_4046,N_3422,N_3833);
nand U4047 (N_4047,N_3614,N_3167);
nor U4048 (N_4048,N_3509,N_3714);
or U4049 (N_4049,N_3230,N_3097);
nor U4050 (N_4050,N_3211,N_3820);
or U4051 (N_4051,N_3470,N_3686);
and U4052 (N_4052,N_3689,N_3341);
nand U4053 (N_4053,N_3128,N_3396);
or U4054 (N_4054,N_3687,N_3444);
nand U4055 (N_4055,N_3594,N_3154);
nor U4056 (N_4056,N_3270,N_3725);
and U4057 (N_4057,N_3677,N_3336);
or U4058 (N_4058,N_3355,N_3892);
nand U4059 (N_4059,N_3126,N_3939);
nor U4060 (N_4060,N_3330,N_3732);
nand U4061 (N_4061,N_3517,N_3041);
and U4062 (N_4062,N_3184,N_3475);
nor U4063 (N_4063,N_3700,N_3968);
or U4064 (N_4064,N_3495,N_3688);
and U4065 (N_4065,N_3832,N_3965);
xnor U4066 (N_4066,N_3650,N_3643);
xor U4067 (N_4067,N_3998,N_3247);
nor U4068 (N_4068,N_3902,N_3292);
nand U4069 (N_4069,N_3883,N_3427);
or U4070 (N_4070,N_3088,N_3234);
nor U4071 (N_4071,N_3790,N_3640);
xor U4072 (N_4072,N_3116,N_3752);
nor U4073 (N_4073,N_3554,N_3611);
or U4074 (N_4074,N_3556,N_3193);
or U4075 (N_4075,N_3170,N_3802);
nand U4076 (N_4076,N_3679,N_3623);
nor U4077 (N_4077,N_3777,N_3108);
and U4078 (N_4078,N_3885,N_3133);
and U4079 (N_4079,N_3192,N_3327);
or U4080 (N_4080,N_3114,N_3226);
nand U4081 (N_4081,N_3277,N_3387);
nand U4082 (N_4082,N_3406,N_3418);
and U4083 (N_4083,N_3888,N_3825);
or U4084 (N_4084,N_3502,N_3699);
and U4085 (N_4085,N_3194,N_3749);
nand U4086 (N_4086,N_3855,N_3302);
nand U4087 (N_4087,N_3488,N_3956);
nor U4088 (N_4088,N_3196,N_3508);
nand U4089 (N_4089,N_3239,N_3117);
and U4090 (N_4090,N_3221,N_3250);
nor U4091 (N_4091,N_3243,N_3325);
xnor U4092 (N_4092,N_3417,N_3134);
or U4093 (N_4093,N_3220,N_3314);
or U4094 (N_4094,N_3143,N_3943);
nor U4095 (N_4095,N_3274,N_3581);
and U4096 (N_4096,N_3291,N_3467);
xnor U4097 (N_4097,N_3626,N_3791);
or U4098 (N_4098,N_3079,N_3754);
xor U4099 (N_4099,N_3829,N_3983);
or U4100 (N_4100,N_3259,N_3600);
or U4101 (N_4101,N_3657,N_3403);
and U4102 (N_4102,N_3461,N_3493);
or U4103 (N_4103,N_3438,N_3358);
nor U4104 (N_4104,N_3596,N_3524);
or U4105 (N_4105,N_3908,N_3718);
nor U4106 (N_4106,N_3503,N_3880);
nor U4107 (N_4107,N_3413,N_3381);
and U4108 (N_4108,N_3945,N_3818);
nand U4109 (N_4109,N_3434,N_3459);
nor U4110 (N_4110,N_3912,N_3536);
xnor U4111 (N_4111,N_3979,N_3534);
nor U4112 (N_4112,N_3012,N_3916);
nor U4113 (N_4113,N_3051,N_3360);
nor U4114 (N_4114,N_3175,N_3044);
nor U4115 (N_4115,N_3954,N_3022);
or U4116 (N_4116,N_3307,N_3269);
nor U4117 (N_4117,N_3995,N_3593);
and U4118 (N_4118,N_3870,N_3506);
xor U4119 (N_4119,N_3760,N_3347);
and U4120 (N_4120,N_3156,N_3538);
or U4121 (N_4121,N_3055,N_3844);
or U4122 (N_4122,N_3095,N_3249);
or U4123 (N_4123,N_3719,N_3858);
nand U4124 (N_4124,N_3994,N_3382);
xor U4125 (N_4125,N_3860,N_3380);
and U4126 (N_4126,N_3225,N_3678);
and U4127 (N_4127,N_3921,N_3674);
nand U4128 (N_4128,N_3089,N_3214);
nand U4129 (N_4129,N_3151,N_3102);
nand U4130 (N_4130,N_3290,N_3195);
and U4131 (N_4131,N_3105,N_3468);
nand U4132 (N_4132,N_3986,N_3693);
and U4133 (N_4133,N_3951,N_3827);
or U4134 (N_4134,N_3241,N_3778);
nand U4135 (N_4135,N_3970,N_3308);
and U4136 (N_4136,N_3383,N_3809);
nand U4137 (N_4137,N_3484,N_3608);
nand U4138 (N_4138,N_3852,N_3811);
nand U4139 (N_4139,N_3553,N_3685);
nand U4140 (N_4140,N_3201,N_3293);
and U4141 (N_4141,N_3755,N_3924);
or U4142 (N_4142,N_3021,N_3751);
or U4143 (N_4143,N_3710,N_3357);
and U4144 (N_4144,N_3915,N_3013);
and U4145 (N_4145,N_3007,N_3499);
or U4146 (N_4146,N_3324,N_3212);
nand U4147 (N_4147,N_3233,N_3256);
nor U4148 (N_4148,N_3672,N_3216);
xnor U4149 (N_4149,N_3447,N_3339);
xnor U4150 (N_4150,N_3078,N_3851);
or U4151 (N_4151,N_3937,N_3601);
nand U4152 (N_4152,N_3345,N_3062);
and U4153 (N_4153,N_3823,N_3947);
nand U4154 (N_4154,N_3440,N_3279);
nor U4155 (N_4155,N_3120,N_3466);
and U4156 (N_4156,N_3263,N_3624);
nand U4157 (N_4157,N_3046,N_3077);
and U4158 (N_4158,N_3801,N_3261);
nor U4159 (N_4159,N_3486,N_3260);
nand U4160 (N_4160,N_3558,N_3452);
and U4161 (N_4161,N_3866,N_3559);
nand U4162 (N_4162,N_3410,N_3798);
nand U4163 (N_4163,N_3472,N_3784);
and U4164 (N_4164,N_3938,N_3348);
and U4165 (N_4165,N_3638,N_3750);
nor U4166 (N_4166,N_3819,N_3146);
nand U4167 (N_4167,N_3779,N_3988);
xnor U4168 (N_4168,N_3774,N_3276);
and U4169 (N_4169,N_3029,N_3030);
nand U4170 (N_4170,N_3739,N_3935);
nand U4171 (N_4171,N_3177,N_3333);
or U4172 (N_4172,N_3618,N_3627);
nor U4173 (N_4173,N_3926,N_3625);
and U4174 (N_4174,N_3014,N_3730);
xor U4175 (N_4175,N_3615,N_3125);
nor U4176 (N_4176,N_3658,N_3609);
or U4177 (N_4177,N_3997,N_3927);
nand U4178 (N_4178,N_3197,N_3881);
and U4179 (N_4179,N_3349,N_3082);
or U4180 (N_4180,N_3155,N_3034);
or U4181 (N_4181,N_3255,N_3490);
or U4182 (N_4182,N_3465,N_3432);
nor U4183 (N_4183,N_3577,N_3240);
or U4184 (N_4184,N_3987,N_3622);
and U4185 (N_4185,N_3568,N_3326);
nor U4186 (N_4186,N_3285,N_3950);
nand U4187 (N_4187,N_3879,N_3610);
or U4188 (N_4188,N_3152,N_3223);
nor U4189 (N_4189,N_3052,N_3098);
and U4190 (N_4190,N_3887,N_3058);
nand U4191 (N_4191,N_3210,N_3074);
nand U4192 (N_4192,N_3335,N_3920);
or U4193 (N_4193,N_3236,N_3587);
or U4194 (N_4194,N_3049,N_3598);
and U4195 (N_4195,N_3597,N_3788);
or U4196 (N_4196,N_3379,N_3780);
nor U4197 (N_4197,N_3961,N_3928);
and U4198 (N_4198,N_3616,N_3080);
and U4199 (N_4199,N_3507,N_3925);
and U4200 (N_4200,N_3585,N_3796);
nand U4201 (N_4201,N_3757,N_3284);
nor U4202 (N_4202,N_3017,N_3183);
nor U4203 (N_4203,N_3914,N_3712);
nand U4204 (N_4204,N_3065,N_3057);
and U4205 (N_4205,N_3163,N_3569);
nand U4206 (N_4206,N_3992,N_3199);
nand U4207 (N_4207,N_3016,N_3451);
or U4208 (N_4208,N_3518,N_3416);
or U4209 (N_4209,N_3815,N_3373);
xnor U4210 (N_4210,N_3421,N_3064);
or U4211 (N_4211,N_3181,N_3482);
nand U4212 (N_4212,N_3480,N_3394);
and U4213 (N_4213,N_3800,N_3771);
nor U4214 (N_4214,N_3955,N_3588);
or U4215 (N_4215,N_3450,N_3966);
nor U4216 (N_4216,N_3140,N_3613);
nor U4217 (N_4217,N_3758,N_3932);
nor U4218 (N_4218,N_3541,N_3745);
or U4219 (N_4219,N_3549,N_3377);
nand U4220 (N_4220,N_3980,N_3822);
and U4221 (N_4221,N_3894,N_3002);
and U4222 (N_4222,N_3940,N_3171);
and U4223 (N_4223,N_3378,N_3306);
or U4224 (N_4224,N_3574,N_3922);
and U4225 (N_4225,N_3008,N_3783);
nor U4226 (N_4226,N_3934,N_3513);
or U4227 (N_4227,N_3492,N_3740);
xor U4228 (N_4228,N_3407,N_3069);
nor U4229 (N_4229,N_3412,N_3728);
and U4230 (N_4230,N_3019,N_3743);
nor U4231 (N_4231,N_3787,N_3096);
or U4232 (N_4232,N_3853,N_3294);
nor U4233 (N_4233,N_3899,N_3834);
nand U4234 (N_4234,N_3115,N_3453);
nand U4235 (N_4235,N_3414,N_3401);
or U4236 (N_4236,N_3411,N_3352);
or U4237 (N_4237,N_3298,N_3350);
nor U4238 (N_4238,N_3435,N_3873);
xnor U4239 (N_4239,N_3696,N_3301);
xnor U4240 (N_4240,N_3578,N_3715);
and U4241 (N_4241,N_3267,N_3476);
nor U4242 (N_4242,N_3648,N_3165);
or U4243 (N_4243,N_3905,N_3628);
xor U4244 (N_4244,N_3191,N_3941);
or U4245 (N_4245,N_3061,N_3797);
or U4246 (N_4246,N_3582,N_3701);
or U4247 (N_4247,N_3691,N_3066);
nor U4248 (N_4248,N_3288,N_3166);
nand U4249 (N_4249,N_3519,N_3551);
nand U4250 (N_4250,N_3405,N_3856);
or U4251 (N_4251,N_3875,N_3977);
and U4252 (N_4252,N_3209,N_3521);
xor U4253 (N_4253,N_3112,N_3281);
nor U4254 (N_4254,N_3984,N_3698);
or U4255 (N_4255,N_3297,N_3520);
nor U4256 (N_4256,N_3911,N_3397);
and U4257 (N_4257,N_3664,N_3299);
nor U4258 (N_4258,N_3500,N_3957);
and U4259 (N_4259,N_3393,N_3682);
nor U4260 (N_4260,N_3121,N_3127);
or U4261 (N_4261,N_3599,N_3633);
nor U4262 (N_4262,N_3042,N_3958);
xor U4263 (N_4263,N_3849,N_3100);
nor U4264 (N_4264,N_3087,N_3772);
or U4265 (N_4265,N_3895,N_3550);
nor U4266 (N_4266,N_3428,N_3562);
and U4267 (N_4267,N_3479,N_3020);
xnor U4268 (N_4268,N_3072,N_3543);
nand U4269 (N_4269,N_3807,N_3471);
or U4270 (N_4270,N_3238,N_3501);
nand U4271 (N_4271,N_3384,N_3090);
nand U4272 (N_4272,N_3056,N_3865);
nor U4273 (N_4273,N_3590,N_3604);
nand U4274 (N_4274,N_3632,N_3010);
nand U4275 (N_4275,N_3532,N_3877);
nor U4276 (N_4276,N_3185,N_3123);
or U4277 (N_4277,N_3789,N_3018);
nand U4278 (N_4278,N_3716,N_3570);
nand U4279 (N_4279,N_3522,N_3148);
nand U4280 (N_4280,N_3910,N_3316);
or U4281 (N_4281,N_3900,N_3734);
xor U4282 (N_4282,N_3252,N_3000);
nand U4283 (N_4283,N_3835,N_3169);
nor U4284 (N_4284,N_3001,N_3283);
nand U4285 (N_4285,N_3477,N_3303);
and U4286 (N_4286,N_3737,N_3544);
or U4287 (N_4287,N_3652,N_3469);
and U4288 (N_4288,N_3481,N_3727);
and U4289 (N_4289,N_3491,N_3153);
nand U4290 (N_4290,N_3909,N_3068);
nor U4291 (N_4291,N_3142,N_3048);
and U4292 (N_4292,N_3770,N_3651);
nand U4293 (N_4293,N_3762,N_3704);
nand U4294 (N_4294,N_3423,N_3202);
or U4295 (N_4295,N_3258,N_3071);
nand U4296 (N_4296,N_3646,N_3974);
nor U4297 (N_4297,N_3906,N_3309);
or U4298 (N_4298,N_3795,N_3645);
nand U4299 (N_4299,N_3478,N_3132);
or U4300 (N_4300,N_3838,N_3918);
xnor U4301 (N_4301,N_3158,N_3841);
nand U4302 (N_4302,N_3160,N_3187);
xnor U4303 (N_4303,N_3665,N_3804);
nor U4304 (N_4304,N_3207,N_3996);
or U4305 (N_4305,N_3620,N_3436);
nor U4306 (N_4306,N_3602,N_3989);
or U4307 (N_4307,N_3205,N_3566);
nor U4308 (N_4308,N_3514,N_3386);
or U4309 (N_4309,N_3540,N_3878);
or U4310 (N_4310,N_3639,N_3203);
or U4311 (N_4311,N_3946,N_3840);
nor U4312 (N_4312,N_3329,N_3555);
xnor U4313 (N_4313,N_3867,N_3122);
and U4314 (N_4314,N_3433,N_3653);
or U4315 (N_4315,N_3015,N_3431);
and U4316 (N_4316,N_3038,N_3913);
or U4317 (N_4317,N_3675,N_3159);
xor U4318 (N_4318,N_3535,N_3978);
nand U4319 (N_4319,N_3150,N_3473);
or U4320 (N_4320,N_3861,N_3104);
nand U4321 (N_4321,N_3157,N_3647);
xor U4322 (N_4322,N_3605,N_3826);
or U4323 (N_4323,N_3705,N_3107);
and U4324 (N_4324,N_3776,N_3092);
nor U4325 (N_4325,N_3923,N_3857);
and U4326 (N_4326,N_3680,N_3863);
nor U4327 (N_4327,N_3035,N_3805);
xor U4328 (N_4328,N_3898,N_3312);
and U4329 (N_4329,N_3245,N_3340);
and U4330 (N_4330,N_3830,N_3869);
nand U4331 (N_4331,N_3408,N_3635);
xor U4332 (N_4332,N_3286,N_3229);
or U4333 (N_4333,N_3321,N_3717);
nor U4334 (N_4334,N_3268,N_3546);
nand U4335 (N_4335,N_3586,N_3351);
nor U4336 (N_4336,N_3457,N_3528);
nand U4337 (N_4337,N_3455,N_3374);
nor U4338 (N_4338,N_3149,N_3039);
or U4339 (N_4339,N_3901,N_3563);
or U4340 (N_4340,N_3931,N_3793);
and U4341 (N_4341,N_3454,N_3215);
xor U4342 (N_4342,N_3368,N_3575);
and U4343 (N_4343,N_3024,N_3673);
nor U4344 (N_4344,N_3031,N_3952);
nor U4345 (N_4345,N_3969,N_3164);
and U4346 (N_4346,N_3257,N_3547);
nand U4347 (N_4347,N_3756,N_3253);
or U4348 (N_4348,N_3806,N_3763);
or U4349 (N_4349,N_3726,N_3168);
nand U4350 (N_4350,N_3649,N_3036);
or U4351 (N_4351,N_3161,N_3060);
or U4352 (N_4352,N_3430,N_3744);
nand U4353 (N_4353,N_3897,N_3985);
nand U4354 (N_4354,N_3073,N_3265);
nand U4355 (N_4355,N_3404,N_3667);
nand U4356 (N_4356,N_3991,N_3848);
nand U4357 (N_4357,N_3812,N_3859);
or U4358 (N_4358,N_3967,N_3526);
or U4359 (N_4359,N_3278,N_3748);
or U4360 (N_4360,N_3742,N_3738);
and U4361 (N_4361,N_3990,N_3655);
nor U4362 (N_4362,N_3733,N_3891);
or U4363 (N_4363,N_3872,N_3172);
nor U4364 (N_4364,N_3248,N_3824);
nor U4365 (N_4365,N_3572,N_3353);
xnor U4366 (N_4366,N_3346,N_3145);
nor U4367 (N_4367,N_3136,N_3235);
nor U4368 (N_4368,N_3702,N_3244);
or U4369 (N_4369,N_3612,N_3871);
or U4370 (N_4370,N_3219,N_3595);
nor U4371 (N_4371,N_3515,N_3903);
xor U4372 (N_4372,N_3059,N_3198);
nor U4373 (N_4373,N_3311,N_3409);
nor U4374 (N_4374,N_3027,N_3695);
nand U4375 (N_4375,N_3206,N_3919);
or U4376 (N_4376,N_3567,N_3003);
or U4377 (N_4377,N_3103,N_3525);
xor U4378 (N_4378,N_3334,N_3489);
nor U4379 (N_4379,N_3282,N_3753);
or U4380 (N_4380,N_3579,N_3964);
nand U4381 (N_4381,N_3429,N_3982);
nand U4382 (N_4382,N_3213,N_3322);
nor U4383 (N_4383,N_3993,N_3295);
nor U4384 (N_4384,N_3933,N_3289);
and U4385 (N_4385,N_3449,N_3228);
and U4386 (N_4386,N_3972,N_3011);
nand U4387 (N_4387,N_3782,N_3005);
and U4388 (N_4388,N_3366,N_3317);
nand U4389 (N_4389,N_3342,N_3040);
or U4390 (N_4390,N_3722,N_3813);
nor U4391 (N_4391,N_3237,N_3076);
or U4392 (N_4392,N_3619,N_3637);
and U4393 (N_4393,N_3362,N_3323);
nor U4394 (N_4394,N_3271,N_3552);
nand U4395 (N_4395,N_3179,N_3182);
and U4396 (N_4396,N_3893,N_3642);
nand U4397 (N_4397,N_3694,N_3808);
and U4398 (N_4398,N_3542,N_3173);
and U4399 (N_4399,N_3402,N_3119);
and U4400 (N_4400,N_3310,N_3023);
and U4401 (N_4401,N_3792,N_3785);
or U4402 (N_4402,N_3761,N_3047);
nand U4403 (N_4403,N_3661,N_3331);
nand U4404 (N_4404,N_3884,N_3670);
and U4405 (N_4405,N_3876,N_3246);
or U4406 (N_4406,N_3529,N_3338);
nand U4407 (N_4407,N_3583,N_3485);
and U4408 (N_4408,N_3254,N_3189);
or U4409 (N_4409,N_3850,N_3690);
or U4410 (N_4410,N_3603,N_3890);
nor U4411 (N_4411,N_3607,N_3365);
or U4412 (N_4412,N_3399,N_3692);
nor U4413 (N_4413,N_3332,N_3118);
nand U4414 (N_4414,N_3296,N_3388);
or U4415 (N_4415,N_3929,N_3109);
nor U4416 (N_4416,N_3130,N_3091);
nor U4417 (N_4417,N_3930,N_3474);
and U4418 (N_4418,N_3948,N_3746);
nand U4419 (N_4419,N_3375,N_3831);
xnor U4420 (N_4420,N_3847,N_3707);
or U4421 (N_4421,N_3217,N_3462);
or U4422 (N_4422,N_3231,N_3305);
or U4423 (N_4423,N_3174,N_3437);
and U4424 (N_4424,N_3548,N_3837);
and U4425 (N_4425,N_3963,N_3094);
or U4426 (N_4426,N_3232,N_3773);
nand U4427 (N_4427,N_3767,N_3343);
nor U4428 (N_4428,N_3735,N_3511);
or U4429 (N_4429,N_3533,N_3218);
or U4430 (N_4430,N_3460,N_3781);
or U4431 (N_4431,N_3723,N_3445);
or U4432 (N_4432,N_3630,N_3896);
nor U4433 (N_4433,N_3037,N_3814);
or U4434 (N_4434,N_3415,N_3081);
nor U4435 (N_4435,N_3032,N_3907);
nand U4436 (N_4436,N_3391,N_3137);
nand U4437 (N_4437,N_3976,N_3188);
or U4438 (N_4438,N_3629,N_3641);
and U4439 (N_4439,N_3617,N_3676);
nand U4440 (N_4440,N_3817,N_3659);
nor U4441 (N_4441,N_3162,N_3981);
nor U4442 (N_4442,N_3794,N_3300);
nor U4443 (N_4443,N_3251,N_3764);
nand U4444 (N_4444,N_3799,N_3318);
or U4445 (N_4445,N_3337,N_3075);
nor U4446 (N_4446,N_3523,N_3009);
xnor U4447 (N_4447,N_3560,N_3810);
and U4448 (N_4448,N_3392,N_3227);
xnor U4449 (N_4449,N_3631,N_3458);
and U4450 (N_4450,N_3845,N_3953);
nand U4451 (N_4451,N_3697,N_3497);
and U4452 (N_4452,N_3496,N_3592);
nand U4453 (N_4453,N_3446,N_3033);
nand U4454 (N_4454,N_3067,N_3803);
nor U4455 (N_4455,N_3656,N_3144);
and U4456 (N_4456,N_3531,N_3344);
xor U4457 (N_4457,N_3516,N_3054);
and U4458 (N_4458,N_3101,N_3741);
nand U4459 (N_4459,N_3580,N_3304);
or U4460 (N_4460,N_3681,N_3816);
nand U4461 (N_4461,N_3369,N_3361);
nand U4462 (N_4462,N_3367,N_3364);
nand U4463 (N_4463,N_3028,N_3328);
nor U4464 (N_4464,N_3085,N_3494);
or U4465 (N_4465,N_3280,N_3093);
or U4466 (N_4466,N_3242,N_3176);
nand U4467 (N_4467,N_3634,N_3204);
nor U4468 (N_4468,N_3775,N_3706);
nand U4469 (N_4469,N_3942,N_3099);
nor U4470 (N_4470,N_3186,N_3537);
xnor U4471 (N_4471,N_3864,N_3731);
nand U4472 (N_4472,N_3621,N_3684);
nand U4473 (N_4473,N_3389,N_3272);
nor U4474 (N_4474,N_3561,N_3606);
and U4475 (N_4475,N_3139,N_3420);
nor U4476 (N_4476,N_3053,N_3371);
nor U4477 (N_4477,N_3483,N_3973);
nand U4478 (N_4478,N_3400,N_3426);
nand U4479 (N_4479,N_3904,N_3124);
or U4480 (N_4480,N_3138,N_3498);
nand U4481 (N_4481,N_3441,N_3050);
nand U4482 (N_4482,N_3530,N_3200);
nor U4483 (N_4483,N_3083,N_3999);
nand U4484 (N_4484,N_3424,N_3786);
nor U4485 (N_4485,N_3882,N_3131);
nor U4486 (N_4486,N_3663,N_3063);
and U4487 (N_4487,N_3720,N_3266);
nand U4488 (N_4488,N_3917,N_3662);
xnor U4489 (N_4489,N_3765,N_3539);
nand U4490 (N_4490,N_3111,N_3313);
and U4491 (N_4491,N_3766,N_3084);
and U4492 (N_4492,N_3944,N_3971);
and U4493 (N_4493,N_3644,N_3372);
and U4494 (N_4494,N_3086,N_3527);
nand U4495 (N_4495,N_3576,N_3886);
or U4496 (N_4496,N_3862,N_3708);
and U4497 (N_4497,N_3448,N_3759);
or U4498 (N_4498,N_3208,N_3565);
nand U4499 (N_4499,N_3376,N_3443);
xnor U4500 (N_4500,N_3381,N_3299);
or U4501 (N_4501,N_3695,N_3639);
and U4502 (N_4502,N_3624,N_3713);
and U4503 (N_4503,N_3559,N_3716);
or U4504 (N_4504,N_3188,N_3458);
and U4505 (N_4505,N_3188,N_3802);
nor U4506 (N_4506,N_3848,N_3369);
nor U4507 (N_4507,N_3885,N_3383);
or U4508 (N_4508,N_3519,N_3325);
and U4509 (N_4509,N_3937,N_3888);
nor U4510 (N_4510,N_3946,N_3184);
and U4511 (N_4511,N_3416,N_3112);
and U4512 (N_4512,N_3965,N_3009);
or U4513 (N_4513,N_3984,N_3970);
nor U4514 (N_4514,N_3382,N_3276);
and U4515 (N_4515,N_3466,N_3458);
nor U4516 (N_4516,N_3206,N_3857);
nand U4517 (N_4517,N_3545,N_3922);
xor U4518 (N_4518,N_3771,N_3715);
nor U4519 (N_4519,N_3671,N_3017);
and U4520 (N_4520,N_3754,N_3264);
xnor U4521 (N_4521,N_3836,N_3593);
nand U4522 (N_4522,N_3326,N_3740);
and U4523 (N_4523,N_3212,N_3382);
nor U4524 (N_4524,N_3090,N_3713);
nand U4525 (N_4525,N_3766,N_3674);
or U4526 (N_4526,N_3837,N_3463);
or U4527 (N_4527,N_3098,N_3884);
nor U4528 (N_4528,N_3218,N_3226);
and U4529 (N_4529,N_3367,N_3693);
nor U4530 (N_4530,N_3733,N_3423);
xnor U4531 (N_4531,N_3716,N_3292);
nor U4532 (N_4532,N_3909,N_3385);
and U4533 (N_4533,N_3442,N_3958);
and U4534 (N_4534,N_3290,N_3539);
or U4535 (N_4535,N_3990,N_3008);
or U4536 (N_4536,N_3964,N_3497);
nand U4537 (N_4537,N_3292,N_3257);
nor U4538 (N_4538,N_3351,N_3132);
nor U4539 (N_4539,N_3759,N_3527);
nor U4540 (N_4540,N_3253,N_3262);
nor U4541 (N_4541,N_3926,N_3831);
or U4542 (N_4542,N_3700,N_3896);
nor U4543 (N_4543,N_3764,N_3394);
xor U4544 (N_4544,N_3398,N_3865);
nor U4545 (N_4545,N_3718,N_3587);
nor U4546 (N_4546,N_3182,N_3477);
or U4547 (N_4547,N_3393,N_3665);
and U4548 (N_4548,N_3080,N_3365);
nor U4549 (N_4549,N_3946,N_3337);
and U4550 (N_4550,N_3570,N_3994);
nand U4551 (N_4551,N_3917,N_3509);
or U4552 (N_4552,N_3086,N_3629);
and U4553 (N_4553,N_3476,N_3983);
nor U4554 (N_4554,N_3080,N_3644);
nand U4555 (N_4555,N_3761,N_3860);
or U4556 (N_4556,N_3220,N_3820);
nand U4557 (N_4557,N_3192,N_3099);
nand U4558 (N_4558,N_3359,N_3730);
and U4559 (N_4559,N_3362,N_3498);
nand U4560 (N_4560,N_3860,N_3921);
and U4561 (N_4561,N_3320,N_3531);
or U4562 (N_4562,N_3511,N_3081);
nor U4563 (N_4563,N_3296,N_3863);
nor U4564 (N_4564,N_3893,N_3734);
nor U4565 (N_4565,N_3292,N_3084);
nand U4566 (N_4566,N_3825,N_3790);
or U4567 (N_4567,N_3041,N_3361);
nor U4568 (N_4568,N_3249,N_3798);
or U4569 (N_4569,N_3937,N_3846);
nand U4570 (N_4570,N_3644,N_3465);
nor U4571 (N_4571,N_3030,N_3983);
and U4572 (N_4572,N_3336,N_3512);
or U4573 (N_4573,N_3479,N_3047);
nand U4574 (N_4574,N_3391,N_3944);
nand U4575 (N_4575,N_3712,N_3849);
and U4576 (N_4576,N_3629,N_3159);
nor U4577 (N_4577,N_3982,N_3959);
or U4578 (N_4578,N_3289,N_3447);
nand U4579 (N_4579,N_3596,N_3782);
nand U4580 (N_4580,N_3922,N_3734);
or U4581 (N_4581,N_3030,N_3677);
nand U4582 (N_4582,N_3606,N_3297);
xnor U4583 (N_4583,N_3987,N_3178);
and U4584 (N_4584,N_3240,N_3721);
xnor U4585 (N_4585,N_3248,N_3966);
nor U4586 (N_4586,N_3845,N_3477);
nand U4587 (N_4587,N_3253,N_3891);
or U4588 (N_4588,N_3178,N_3246);
nor U4589 (N_4589,N_3560,N_3595);
nand U4590 (N_4590,N_3733,N_3235);
or U4591 (N_4591,N_3075,N_3020);
or U4592 (N_4592,N_3887,N_3644);
or U4593 (N_4593,N_3859,N_3357);
nand U4594 (N_4594,N_3764,N_3175);
or U4595 (N_4595,N_3388,N_3714);
xor U4596 (N_4596,N_3492,N_3577);
or U4597 (N_4597,N_3558,N_3942);
xnor U4598 (N_4598,N_3469,N_3895);
nor U4599 (N_4599,N_3233,N_3373);
and U4600 (N_4600,N_3377,N_3396);
and U4601 (N_4601,N_3294,N_3058);
or U4602 (N_4602,N_3708,N_3247);
nand U4603 (N_4603,N_3850,N_3635);
nor U4604 (N_4604,N_3686,N_3473);
nor U4605 (N_4605,N_3569,N_3555);
nor U4606 (N_4606,N_3378,N_3828);
or U4607 (N_4607,N_3902,N_3925);
nor U4608 (N_4608,N_3330,N_3385);
nand U4609 (N_4609,N_3996,N_3427);
nor U4610 (N_4610,N_3769,N_3710);
xnor U4611 (N_4611,N_3436,N_3236);
nand U4612 (N_4612,N_3098,N_3453);
nand U4613 (N_4613,N_3323,N_3724);
xnor U4614 (N_4614,N_3635,N_3955);
nor U4615 (N_4615,N_3948,N_3774);
nand U4616 (N_4616,N_3306,N_3474);
nor U4617 (N_4617,N_3683,N_3458);
or U4618 (N_4618,N_3155,N_3493);
and U4619 (N_4619,N_3806,N_3580);
or U4620 (N_4620,N_3708,N_3220);
nor U4621 (N_4621,N_3230,N_3078);
and U4622 (N_4622,N_3132,N_3221);
nand U4623 (N_4623,N_3869,N_3086);
nor U4624 (N_4624,N_3864,N_3736);
and U4625 (N_4625,N_3012,N_3527);
nand U4626 (N_4626,N_3727,N_3349);
or U4627 (N_4627,N_3427,N_3422);
or U4628 (N_4628,N_3700,N_3799);
or U4629 (N_4629,N_3327,N_3075);
nor U4630 (N_4630,N_3256,N_3177);
and U4631 (N_4631,N_3590,N_3149);
nand U4632 (N_4632,N_3858,N_3808);
or U4633 (N_4633,N_3933,N_3592);
nand U4634 (N_4634,N_3730,N_3080);
nor U4635 (N_4635,N_3937,N_3660);
nand U4636 (N_4636,N_3638,N_3504);
nand U4637 (N_4637,N_3192,N_3847);
or U4638 (N_4638,N_3437,N_3062);
nand U4639 (N_4639,N_3263,N_3931);
nand U4640 (N_4640,N_3761,N_3349);
or U4641 (N_4641,N_3327,N_3573);
nor U4642 (N_4642,N_3628,N_3070);
nand U4643 (N_4643,N_3349,N_3274);
or U4644 (N_4644,N_3103,N_3890);
xnor U4645 (N_4645,N_3579,N_3201);
nand U4646 (N_4646,N_3145,N_3035);
and U4647 (N_4647,N_3377,N_3329);
nor U4648 (N_4648,N_3940,N_3571);
and U4649 (N_4649,N_3274,N_3961);
or U4650 (N_4650,N_3964,N_3015);
or U4651 (N_4651,N_3367,N_3030);
nand U4652 (N_4652,N_3247,N_3086);
or U4653 (N_4653,N_3443,N_3825);
and U4654 (N_4654,N_3988,N_3935);
and U4655 (N_4655,N_3931,N_3003);
or U4656 (N_4656,N_3943,N_3374);
or U4657 (N_4657,N_3125,N_3171);
nor U4658 (N_4658,N_3451,N_3374);
nand U4659 (N_4659,N_3321,N_3701);
and U4660 (N_4660,N_3055,N_3077);
nand U4661 (N_4661,N_3296,N_3280);
and U4662 (N_4662,N_3122,N_3818);
and U4663 (N_4663,N_3319,N_3678);
nand U4664 (N_4664,N_3817,N_3705);
xnor U4665 (N_4665,N_3425,N_3552);
nor U4666 (N_4666,N_3550,N_3874);
xnor U4667 (N_4667,N_3550,N_3868);
or U4668 (N_4668,N_3312,N_3886);
and U4669 (N_4669,N_3722,N_3552);
and U4670 (N_4670,N_3895,N_3289);
and U4671 (N_4671,N_3803,N_3946);
or U4672 (N_4672,N_3758,N_3948);
nand U4673 (N_4673,N_3681,N_3385);
nor U4674 (N_4674,N_3086,N_3252);
or U4675 (N_4675,N_3087,N_3738);
nor U4676 (N_4676,N_3629,N_3666);
nand U4677 (N_4677,N_3821,N_3384);
or U4678 (N_4678,N_3467,N_3113);
nor U4679 (N_4679,N_3660,N_3054);
or U4680 (N_4680,N_3634,N_3530);
and U4681 (N_4681,N_3309,N_3667);
xnor U4682 (N_4682,N_3064,N_3851);
nor U4683 (N_4683,N_3442,N_3503);
nand U4684 (N_4684,N_3464,N_3478);
nand U4685 (N_4685,N_3878,N_3480);
and U4686 (N_4686,N_3680,N_3239);
nand U4687 (N_4687,N_3428,N_3965);
nand U4688 (N_4688,N_3282,N_3996);
nor U4689 (N_4689,N_3204,N_3561);
and U4690 (N_4690,N_3396,N_3886);
and U4691 (N_4691,N_3418,N_3846);
nand U4692 (N_4692,N_3562,N_3444);
and U4693 (N_4693,N_3846,N_3763);
nor U4694 (N_4694,N_3262,N_3519);
or U4695 (N_4695,N_3794,N_3662);
nor U4696 (N_4696,N_3170,N_3007);
nand U4697 (N_4697,N_3405,N_3084);
or U4698 (N_4698,N_3986,N_3571);
and U4699 (N_4699,N_3837,N_3721);
nor U4700 (N_4700,N_3057,N_3158);
or U4701 (N_4701,N_3809,N_3207);
nand U4702 (N_4702,N_3556,N_3025);
or U4703 (N_4703,N_3790,N_3403);
or U4704 (N_4704,N_3915,N_3642);
nor U4705 (N_4705,N_3957,N_3160);
xnor U4706 (N_4706,N_3914,N_3999);
nor U4707 (N_4707,N_3414,N_3800);
nand U4708 (N_4708,N_3057,N_3742);
xnor U4709 (N_4709,N_3230,N_3845);
or U4710 (N_4710,N_3175,N_3428);
nand U4711 (N_4711,N_3732,N_3878);
and U4712 (N_4712,N_3838,N_3423);
nand U4713 (N_4713,N_3000,N_3417);
nor U4714 (N_4714,N_3431,N_3089);
or U4715 (N_4715,N_3193,N_3844);
nor U4716 (N_4716,N_3079,N_3887);
or U4717 (N_4717,N_3980,N_3391);
or U4718 (N_4718,N_3712,N_3989);
and U4719 (N_4719,N_3599,N_3512);
or U4720 (N_4720,N_3789,N_3492);
or U4721 (N_4721,N_3722,N_3235);
or U4722 (N_4722,N_3136,N_3015);
or U4723 (N_4723,N_3957,N_3915);
or U4724 (N_4724,N_3122,N_3779);
and U4725 (N_4725,N_3325,N_3403);
or U4726 (N_4726,N_3854,N_3929);
xor U4727 (N_4727,N_3323,N_3201);
or U4728 (N_4728,N_3733,N_3595);
xor U4729 (N_4729,N_3237,N_3566);
nand U4730 (N_4730,N_3015,N_3307);
nor U4731 (N_4731,N_3884,N_3828);
nor U4732 (N_4732,N_3238,N_3311);
or U4733 (N_4733,N_3161,N_3336);
or U4734 (N_4734,N_3860,N_3107);
xnor U4735 (N_4735,N_3526,N_3219);
nor U4736 (N_4736,N_3327,N_3159);
nand U4737 (N_4737,N_3678,N_3686);
nand U4738 (N_4738,N_3452,N_3908);
nor U4739 (N_4739,N_3684,N_3102);
nand U4740 (N_4740,N_3086,N_3340);
nor U4741 (N_4741,N_3673,N_3750);
or U4742 (N_4742,N_3595,N_3141);
nor U4743 (N_4743,N_3192,N_3631);
or U4744 (N_4744,N_3869,N_3050);
and U4745 (N_4745,N_3935,N_3071);
nor U4746 (N_4746,N_3384,N_3050);
or U4747 (N_4747,N_3415,N_3345);
nand U4748 (N_4748,N_3477,N_3626);
xor U4749 (N_4749,N_3740,N_3285);
nand U4750 (N_4750,N_3985,N_3507);
nor U4751 (N_4751,N_3008,N_3103);
or U4752 (N_4752,N_3439,N_3893);
and U4753 (N_4753,N_3521,N_3118);
xnor U4754 (N_4754,N_3595,N_3062);
or U4755 (N_4755,N_3593,N_3822);
or U4756 (N_4756,N_3980,N_3544);
and U4757 (N_4757,N_3179,N_3359);
nand U4758 (N_4758,N_3524,N_3772);
or U4759 (N_4759,N_3961,N_3908);
nor U4760 (N_4760,N_3393,N_3821);
or U4761 (N_4761,N_3313,N_3281);
nor U4762 (N_4762,N_3504,N_3175);
nor U4763 (N_4763,N_3955,N_3394);
or U4764 (N_4764,N_3931,N_3742);
nand U4765 (N_4765,N_3139,N_3658);
nand U4766 (N_4766,N_3309,N_3991);
and U4767 (N_4767,N_3889,N_3259);
nand U4768 (N_4768,N_3560,N_3535);
nor U4769 (N_4769,N_3963,N_3363);
nor U4770 (N_4770,N_3714,N_3888);
xnor U4771 (N_4771,N_3148,N_3171);
xor U4772 (N_4772,N_3907,N_3457);
and U4773 (N_4773,N_3438,N_3115);
nand U4774 (N_4774,N_3368,N_3813);
or U4775 (N_4775,N_3610,N_3983);
xor U4776 (N_4776,N_3509,N_3480);
nand U4777 (N_4777,N_3863,N_3636);
nand U4778 (N_4778,N_3406,N_3854);
xor U4779 (N_4779,N_3202,N_3104);
nand U4780 (N_4780,N_3501,N_3955);
or U4781 (N_4781,N_3362,N_3680);
xor U4782 (N_4782,N_3027,N_3795);
or U4783 (N_4783,N_3440,N_3222);
xor U4784 (N_4784,N_3733,N_3388);
and U4785 (N_4785,N_3986,N_3225);
nand U4786 (N_4786,N_3788,N_3018);
nand U4787 (N_4787,N_3369,N_3370);
nand U4788 (N_4788,N_3185,N_3093);
and U4789 (N_4789,N_3858,N_3615);
nand U4790 (N_4790,N_3535,N_3582);
and U4791 (N_4791,N_3178,N_3541);
nor U4792 (N_4792,N_3846,N_3063);
or U4793 (N_4793,N_3799,N_3820);
xor U4794 (N_4794,N_3546,N_3261);
nor U4795 (N_4795,N_3282,N_3592);
and U4796 (N_4796,N_3977,N_3979);
nor U4797 (N_4797,N_3292,N_3274);
nor U4798 (N_4798,N_3702,N_3624);
and U4799 (N_4799,N_3745,N_3807);
nand U4800 (N_4800,N_3509,N_3623);
and U4801 (N_4801,N_3887,N_3849);
nor U4802 (N_4802,N_3839,N_3170);
and U4803 (N_4803,N_3381,N_3457);
nor U4804 (N_4804,N_3756,N_3735);
or U4805 (N_4805,N_3137,N_3866);
or U4806 (N_4806,N_3193,N_3142);
nor U4807 (N_4807,N_3292,N_3473);
or U4808 (N_4808,N_3389,N_3912);
nand U4809 (N_4809,N_3009,N_3598);
or U4810 (N_4810,N_3158,N_3477);
nor U4811 (N_4811,N_3376,N_3032);
or U4812 (N_4812,N_3485,N_3191);
nor U4813 (N_4813,N_3704,N_3802);
or U4814 (N_4814,N_3842,N_3836);
or U4815 (N_4815,N_3997,N_3387);
or U4816 (N_4816,N_3042,N_3238);
or U4817 (N_4817,N_3007,N_3133);
or U4818 (N_4818,N_3927,N_3901);
or U4819 (N_4819,N_3677,N_3594);
or U4820 (N_4820,N_3790,N_3960);
nor U4821 (N_4821,N_3733,N_3814);
or U4822 (N_4822,N_3842,N_3796);
nand U4823 (N_4823,N_3006,N_3801);
nand U4824 (N_4824,N_3312,N_3558);
nor U4825 (N_4825,N_3403,N_3262);
nand U4826 (N_4826,N_3873,N_3178);
and U4827 (N_4827,N_3436,N_3566);
nor U4828 (N_4828,N_3462,N_3342);
xnor U4829 (N_4829,N_3634,N_3808);
or U4830 (N_4830,N_3617,N_3792);
nand U4831 (N_4831,N_3793,N_3374);
nor U4832 (N_4832,N_3712,N_3123);
or U4833 (N_4833,N_3576,N_3975);
nor U4834 (N_4834,N_3429,N_3244);
and U4835 (N_4835,N_3463,N_3481);
and U4836 (N_4836,N_3423,N_3289);
or U4837 (N_4837,N_3981,N_3438);
nor U4838 (N_4838,N_3850,N_3500);
or U4839 (N_4839,N_3111,N_3780);
or U4840 (N_4840,N_3962,N_3292);
nor U4841 (N_4841,N_3959,N_3811);
xnor U4842 (N_4842,N_3932,N_3950);
and U4843 (N_4843,N_3895,N_3184);
nand U4844 (N_4844,N_3063,N_3109);
nand U4845 (N_4845,N_3271,N_3157);
and U4846 (N_4846,N_3345,N_3610);
nor U4847 (N_4847,N_3528,N_3485);
or U4848 (N_4848,N_3262,N_3454);
and U4849 (N_4849,N_3631,N_3434);
and U4850 (N_4850,N_3912,N_3005);
or U4851 (N_4851,N_3722,N_3117);
xor U4852 (N_4852,N_3286,N_3265);
xor U4853 (N_4853,N_3874,N_3211);
nand U4854 (N_4854,N_3594,N_3104);
and U4855 (N_4855,N_3312,N_3874);
and U4856 (N_4856,N_3209,N_3424);
and U4857 (N_4857,N_3145,N_3508);
xor U4858 (N_4858,N_3803,N_3400);
nor U4859 (N_4859,N_3608,N_3953);
or U4860 (N_4860,N_3882,N_3392);
and U4861 (N_4861,N_3912,N_3940);
nand U4862 (N_4862,N_3685,N_3548);
nand U4863 (N_4863,N_3317,N_3261);
or U4864 (N_4864,N_3876,N_3668);
xor U4865 (N_4865,N_3358,N_3455);
or U4866 (N_4866,N_3442,N_3798);
and U4867 (N_4867,N_3704,N_3434);
nor U4868 (N_4868,N_3463,N_3855);
xnor U4869 (N_4869,N_3051,N_3601);
nand U4870 (N_4870,N_3573,N_3836);
or U4871 (N_4871,N_3535,N_3036);
and U4872 (N_4872,N_3219,N_3123);
and U4873 (N_4873,N_3348,N_3624);
and U4874 (N_4874,N_3241,N_3387);
and U4875 (N_4875,N_3503,N_3625);
nand U4876 (N_4876,N_3660,N_3138);
and U4877 (N_4877,N_3839,N_3809);
xnor U4878 (N_4878,N_3280,N_3670);
xnor U4879 (N_4879,N_3607,N_3323);
nand U4880 (N_4880,N_3460,N_3017);
or U4881 (N_4881,N_3434,N_3906);
nand U4882 (N_4882,N_3407,N_3688);
or U4883 (N_4883,N_3326,N_3865);
and U4884 (N_4884,N_3880,N_3168);
or U4885 (N_4885,N_3040,N_3742);
xnor U4886 (N_4886,N_3533,N_3957);
or U4887 (N_4887,N_3917,N_3520);
nor U4888 (N_4888,N_3041,N_3121);
nor U4889 (N_4889,N_3884,N_3296);
nor U4890 (N_4890,N_3012,N_3988);
or U4891 (N_4891,N_3301,N_3474);
or U4892 (N_4892,N_3708,N_3815);
xnor U4893 (N_4893,N_3441,N_3091);
nor U4894 (N_4894,N_3010,N_3573);
nand U4895 (N_4895,N_3100,N_3310);
nor U4896 (N_4896,N_3423,N_3544);
or U4897 (N_4897,N_3374,N_3992);
nor U4898 (N_4898,N_3462,N_3283);
nor U4899 (N_4899,N_3304,N_3104);
nand U4900 (N_4900,N_3374,N_3544);
or U4901 (N_4901,N_3938,N_3802);
nand U4902 (N_4902,N_3745,N_3225);
nand U4903 (N_4903,N_3340,N_3311);
nand U4904 (N_4904,N_3637,N_3583);
nand U4905 (N_4905,N_3725,N_3051);
nand U4906 (N_4906,N_3769,N_3716);
nand U4907 (N_4907,N_3951,N_3452);
nor U4908 (N_4908,N_3711,N_3304);
nand U4909 (N_4909,N_3361,N_3769);
nor U4910 (N_4910,N_3807,N_3400);
xor U4911 (N_4911,N_3852,N_3846);
or U4912 (N_4912,N_3284,N_3677);
and U4913 (N_4913,N_3074,N_3427);
nand U4914 (N_4914,N_3065,N_3412);
nand U4915 (N_4915,N_3411,N_3750);
nand U4916 (N_4916,N_3422,N_3989);
xnor U4917 (N_4917,N_3339,N_3085);
nand U4918 (N_4918,N_3116,N_3585);
nand U4919 (N_4919,N_3628,N_3951);
nand U4920 (N_4920,N_3675,N_3515);
and U4921 (N_4921,N_3423,N_3869);
nor U4922 (N_4922,N_3148,N_3188);
nor U4923 (N_4923,N_3606,N_3080);
xnor U4924 (N_4924,N_3436,N_3445);
and U4925 (N_4925,N_3662,N_3737);
and U4926 (N_4926,N_3140,N_3607);
nor U4927 (N_4927,N_3192,N_3404);
and U4928 (N_4928,N_3448,N_3052);
xnor U4929 (N_4929,N_3402,N_3365);
or U4930 (N_4930,N_3437,N_3143);
or U4931 (N_4931,N_3081,N_3720);
nand U4932 (N_4932,N_3316,N_3521);
and U4933 (N_4933,N_3234,N_3076);
or U4934 (N_4934,N_3241,N_3812);
nand U4935 (N_4935,N_3057,N_3220);
nand U4936 (N_4936,N_3163,N_3424);
nand U4937 (N_4937,N_3781,N_3076);
and U4938 (N_4938,N_3203,N_3796);
nand U4939 (N_4939,N_3985,N_3240);
and U4940 (N_4940,N_3571,N_3223);
nand U4941 (N_4941,N_3726,N_3189);
xor U4942 (N_4942,N_3471,N_3443);
nor U4943 (N_4943,N_3860,N_3631);
or U4944 (N_4944,N_3849,N_3962);
nor U4945 (N_4945,N_3931,N_3314);
nor U4946 (N_4946,N_3080,N_3527);
nor U4947 (N_4947,N_3294,N_3431);
and U4948 (N_4948,N_3160,N_3805);
nor U4949 (N_4949,N_3779,N_3735);
and U4950 (N_4950,N_3183,N_3785);
or U4951 (N_4951,N_3834,N_3229);
or U4952 (N_4952,N_3545,N_3774);
nand U4953 (N_4953,N_3893,N_3682);
or U4954 (N_4954,N_3985,N_3932);
or U4955 (N_4955,N_3304,N_3318);
xor U4956 (N_4956,N_3379,N_3839);
nand U4957 (N_4957,N_3538,N_3223);
nand U4958 (N_4958,N_3074,N_3070);
and U4959 (N_4959,N_3086,N_3445);
and U4960 (N_4960,N_3926,N_3486);
nor U4961 (N_4961,N_3994,N_3101);
nor U4962 (N_4962,N_3516,N_3018);
nand U4963 (N_4963,N_3205,N_3386);
and U4964 (N_4964,N_3071,N_3260);
nand U4965 (N_4965,N_3966,N_3648);
or U4966 (N_4966,N_3239,N_3263);
nand U4967 (N_4967,N_3696,N_3540);
or U4968 (N_4968,N_3536,N_3656);
or U4969 (N_4969,N_3722,N_3642);
xnor U4970 (N_4970,N_3544,N_3156);
or U4971 (N_4971,N_3138,N_3951);
or U4972 (N_4972,N_3079,N_3266);
xor U4973 (N_4973,N_3739,N_3244);
and U4974 (N_4974,N_3440,N_3124);
or U4975 (N_4975,N_3710,N_3167);
or U4976 (N_4976,N_3206,N_3021);
and U4977 (N_4977,N_3353,N_3366);
nor U4978 (N_4978,N_3314,N_3327);
or U4979 (N_4979,N_3956,N_3248);
or U4980 (N_4980,N_3039,N_3787);
or U4981 (N_4981,N_3597,N_3178);
nand U4982 (N_4982,N_3505,N_3556);
nor U4983 (N_4983,N_3295,N_3028);
nor U4984 (N_4984,N_3460,N_3741);
nor U4985 (N_4985,N_3072,N_3575);
nor U4986 (N_4986,N_3051,N_3696);
nand U4987 (N_4987,N_3070,N_3538);
nor U4988 (N_4988,N_3945,N_3190);
xnor U4989 (N_4989,N_3993,N_3257);
or U4990 (N_4990,N_3941,N_3903);
nor U4991 (N_4991,N_3581,N_3699);
or U4992 (N_4992,N_3149,N_3415);
nor U4993 (N_4993,N_3642,N_3527);
nand U4994 (N_4994,N_3288,N_3613);
nor U4995 (N_4995,N_3939,N_3727);
nand U4996 (N_4996,N_3035,N_3408);
or U4997 (N_4997,N_3826,N_3518);
xor U4998 (N_4998,N_3992,N_3770);
xnor U4999 (N_4999,N_3660,N_3574);
or U5000 (N_5000,N_4108,N_4902);
nor U5001 (N_5001,N_4097,N_4240);
and U5002 (N_5002,N_4104,N_4060);
and U5003 (N_5003,N_4632,N_4769);
or U5004 (N_5004,N_4347,N_4562);
and U5005 (N_5005,N_4956,N_4402);
xor U5006 (N_5006,N_4495,N_4684);
nand U5007 (N_5007,N_4563,N_4193);
or U5008 (N_5008,N_4688,N_4698);
and U5009 (N_5009,N_4690,N_4069);
nand U5010 (N_5010,N_4190,N_4901);
nor U5011 (N_5011,N_4815,N_4849);
nor U5012 (N_5012,N_4012,N_4460);
or U5013 (N_5013,N_4067,N_4145);
nor U5014 (N_5014,N_4597,N_4265);
or U5015 (N_5015,N_4057,N_4768);
xor U5016 (N_5016,N_4270,N_4055);
or U5017 (N_5017,N_4864,N_4619);
and U5018 (N_5018,N_4944,N_4788);
and U5019 (N_5019,N_4238,N_4940);
nand U5020 (N_5020,N_4878,N_4775);
xor U5021 (N_5021,N_4820,N_4388);
nor U5022 (N_5022,N_4842,N_4953);
and U5023 (N_5023,N_4628,N_4153);
nor U5024 (N_5024,N_4498,N_4365);
or U5025 (N_5025,N_4887,N_4089);
nand U5026 (N_5026,N_4242,N_4120);
or U5027 (N_5027,N_4152,N_4824);
nand U5028 (N_5028,N_4122,N_4435);
nor U5029 (N_5029,N_4269,N_4642);
and U5030 (N_5030,N_4750,N_4861);
nand U5031 (N_5031,N_4705,N_4056);
nor U5032 (N_5032,N_4657,N_4254);
nand U5033 (N_5033,N_4660,N_4349);
and U5034 (N_5034,N_4627,N_4149);
nand U5035 (N_5035,N_4214,N_4624);
nor U5036 (N_5036,N_4863,N_4724);
or U5037 (N_5037,N_4177,N_4356);
xor U5038 (N_5038,N_4150,N_4979);
or U5039 (N_5039,N_4276,N_4857);
xor U5040 (N_5040,N_4035,N_4751);
xor U5041 (N_5041,N_4507,N_4764);
and U5042 (N_5042,N_4047,N_4614);
nand U5043 (N_5043,N_4401,N_4653);
nor U5044 (N_5044,N_4667,N_4773);
nand U5045 (N_5045,N_4411,N_4034);
or U5046 (N_5046,N_4793,N_4123);
or U5047 (N_5047,N_4078,N_4294);
nor U5048 (N_5048,N_4701,N_4763);
or U5049 (N_5049,N_4519,N_4790);
and U5050 (N_5050,N_4397,N_4374);
nand U5051 (N_5051,N_4644,N_4704);
nor U5052 (N_5052,N_4364,N_4163);
nor U5053 (N_5053,N_4530,N_4168);
or U5054 (N_5054,N_4548,N_4101);
and U5055 (N_5055,N_4449,N_4283);
or U5056 (N_5056,N_4508,N_4175);
xor U5057 (N_5057,N_4219,N_4008);
and U5058 (N_5058,N_4187,N_4081);
xor U5059 (N_5059,N_4351,N_4129);
nor U5060 (N_5060,N_4327,N_4311);
or U5061 (N_5061,N_4394,N_4447);
xor U5062 (N_5062,N_4430,N_4522);
or U5063 (N_5063,N_4377,N_4165);
nand U5064 (N_5064,N_4231,N_4876);
nand U5065 (N_5065,N_4167,N_4247);
nor U5066 (N_5066,N_4074,N_4251);
or U5067 (N_5067,N_4299,N_4572);
nor U5068 (N_5068,N_4245,N_4837);
nor U5069 (N_5069,N_4531,N_4930);
nand U5070 (N_5070,N_4408,N_4604);
xor U5071 (N_5071,N_4516,N_4871);
and U5072 (N_5072,N_4023,N_4742);
xor U5073 (N_5073,N_4039,N_4072);
nor U5074 (N_5074,N_4528,N_4905);
nor U5075 (N_5075,N_4765,N_4180);
and U5076 (N_5076,N_4909,N_4969);
or U5077 (N_5077,N_4437,N_4752);
and U5078 (N_5078,N_4004,N_4179);
nand U5079 (N_5079,N_4770,N_4143);
nand U5080 (N_5080,N_4661,N_4256);
nand U5081 (N_5081,N_4418,N_4686);
nand U5082 (N_5082,N_4776,N_4346);
nor U5083 (N_5083,N_4564,N_4504);
and U5084 (N_5084,N_4094,N_4558);
or U5085 (N_5085,N_4221,N_4880);
xor U5086 (N_5086,N_4556,N_4225);
nor U5087 (N_5087,N_4307,N_4099);
nand U5088 (N_5088,N_4586,N_4048);
xor U5089 (N_5089,N_4199,N_4753);
or U5090 (N_5090,N_4259,N_4111);
nor U5091 (N_5091,N_4967,N_4345);
or U5092 (N_5092,N_4113,N_4471);
or U5093 (N_5093,N_4543,N_4220);
and U5094 (N_5094,N_4205,N_4869);
and U5095 (N_5095,N_4612,N_4816);
nor U5096 (N_5096,N_4466,N_4885);
nor U5097 (N_5097,N_4761,N_4234);
nor U5098 (N_5098,N_4469,N_4022);
nor U5099 (N_5099,N_4354,N_4695);
nand U5100 (N_5100,N_4798,N_4973);
nand U5101 (N_5101,N_4438,N_4479);
nand U5102 (N_5102,N_4319,N_4389);
or U5103 (N_5103,N_4313,N_4019);
nand U5104 (N_5104,N_4648,N_4856);
nor U5105 (N_5105,N_4808,N_4289);
or U5106 (N_5106,N_4159,N_4112);
xor U5107 (N_5107,N_4306,N_4706);
nand U5108 (N_5108,N_4791,N_4523);
nor U5109 (N_5109,N_4026,N_4981);
nor U5110 (N_5110,N_4710,N_4178);
nor U5111 (N_5111,N_4288,N_4441);
nand U5112 (N_5112,N_4410,N_4732);
nand U5113 (N_5113,N_4043,N_4779);
nor U5114 (N_5114,N_4384,N_4964);
or U5115 (N_5115,N_4813,N_4006);
nor U5116 (N_5116,N_4959,N_4188);
or U5117 (N_5117,N_4369,N_4325);
and U5118 (N_5118,N_4565,N_4772);
and U5119 (N_5119,N_4804,N_4566);
nor U5120 (N_5120,N_4229,N_4200);
and U5121 (N_5121,N_4756,N_4974);
xor U5122 (N_5122,N_4217,N_4865);
nand U5123 (N_5123,N_4593,N_4620);
and U5124 (N_5124,N_4223,N_4541);
nor U5125 (N_5125,N_4803,N_4841);
nand U5126 (N_5126,N_4680,N_4800);
and U5127 (N_5127,N_4016,N_4164);
nand U5128 (N_5128,N_4045,N_4456);
nor U5129 (N_5129,N_4392,N_4928);
nand U5130 (N_5130,N_4651,N_4198);
nand U5131 (N_5131,N_4420,N_4483);
or U5132 (N_5132,N_4128,N_4328);
nor U5133 (N_5133,N_4107,N_4414);
or U5134 (N_5134,N_4310,N_4204);
or U5135 (N_5135,N_4972,N_4540);
nor U5136 (N_5136,N_4577,N_4948);
nor U5137 (N_5137,N_4730,N_4239);
nor U5138 (N_5138,N_4598,N_4749);
and U5139 (N_5139,N_4296,N_4581);
and U5140 (N_5140,N_4966,N_4576);
and U5141 (N_5141,N_4098,N_4532);
nand U5142 (N_5142,N_4344,N_4396);
or U5143 (N_5143,N_4042,N_4362);
nand U5144 (N_5144,N_4000,N_4116);
or U5145 (N_5145,N_4774,N_4357);
xor U5146 (N_5146,N_4494,N_4372);
nor U5147 (N_5147,N_4213,N_4606);
nand U5148 (N_5148,N_4990,N_4692);
and U5149 (N_5149,N_4893,N_4064);
and U5150 (N_5150,N_4036,N_4427);
and U5151 (N_5151,N_4826,N_4912);
and U5152 (N_5152,N_4476,N_4124);
or U5153 (N_5153,N_4579,N_4637);
and U5154 (N_5154,N_4699,N_4434);
and U5155 (N_5155,N_4797,N_4907);
or U5156 (N_5156,N_4079,N_4485);
nor U5157 (N_5157,N_4809,N_4847);
xnor U5158 (N_5158,N_4984,N_4933);
nand U5159 (N_5159,N_4659,N_4819);
nand U5160 (N_5160,N_4118,N_4230);
nand U5161 (N_5161,N_4881,N_4119);
nor U5162 (N_5162,N_4324,N_4585);
nor U5163 (N_5163,N_4822,N_4400);
or U5164 (N_5164,N_4148,N_4802);
and U5165 (N_5165,N_4796,N_4271);
xnor U5166 (N_5166,N_4838,N_4649);
nand U5167 (N_5167,N_4810,N_4947);
nor U5168 (N_5168,N_4515,N_4601);
nor U5169 (N_5169,N_4812,N_4032);
nand U5170 (N_5170,N_4305,N_4656);
or U5171 (N_5171,N_4462,N_4925);
xor U5172 (N_5172,N_4058,N_4638);
xor U5173 (N_5173,N_4010,N_4158);
and U5174 (N_5174,N_4243,N_4664);
xnor U5175 (N_5175,N_4872,N_4169);
nor U5176 (N_5176,N_4370,N_4843);
nor U5177 (N_5177,N_4995,N_4350);
nor U5178 (N_5178,N_4040,N_4342);
or U5179 (N_5179,N_4708,N_4005);
or U5180 (N_5180,N_4255,N_4513);
and U5181 (N_5181,N_4147,N_4920);
and U5182 (N_5182,N_4465,N_4618);
nand U5183 (N_5183,N_4889,N_4714);
nor U5184 (N_5184,N_4201,N_4478);
or U5185 (N_5185,N_4286,N_4482);
and U5186 (N_5186,N_4105,N_4867);
and U5187 (N_5187,N_4671,N_4858);
or U5188 (N_5188,N_4718,N_4068);
and U5189 (N_5189,N_4801,N_4713);
nor U5190 (N_5190,N_4224,N_4899);
or U5191 (N_5191,N_4640,N_4212);
nor U5192 (N_5192,N_4962,N_4433);
or U5193 (N_5193,N_4102,N_4833);
or U5194 (N_5194,N_4918,N_4716);
nand U5195 (N_5195,N_4781,N_4183);
nand U5196 (N_5196,N_4115,N_4021);
or U5197 (N_5197,N_4358,N_4303);
xnor U5198 (N_5198,N_4567,N_4337);
nor U5199 (N_5199,N_4825,N_4759);
xor U5200 (N_5200,N_4983,N_4689);
nor U5201 (N_5201,N_4834,N_4828);
nand U5202 (N_5202,N_4279,N_4468);
or U5203 (N_5203,N_4831,N_4895);
nor U5204 (N_5204,N_4683,N_4840);
or U5205 (N_5205,N_4210,N_4676);
or U5206 (N_5206,N_4611,N_4549);
and U5207 (N_5207,N_4399,N_4375);
xnor U5208 (N_5208,N_4312,N_4237);
and U5209 (N_5209,N_4290,N_4302);
and U5210 (N_5210,N_4884,N_4189);
nor U5211 (N_5211,N_4156,N_4550);
and U5212 (N_5212,N_4323,N_4923);
and U5213 (N_5213,N_4052,N_4678);
nor U5214 (N_5214,N_4329,N_4547);
or U5215 (N_5215,N_4539,N_4429);
nand U5216 (N_5216,N_4154,N_4110);
nand U5217 (N_5217,N_4529,N_4870);
nor U5218 (N_5218,N_4295,N_4988);
nor U5219 (N_5219,N_4817,N_4343);
nand U5220 (N_5220,N_4709,N_4782);
nor U5221 (N_5221,N_4037,N_4246);
nand U5222 (N_5222,N_4961,N_4287);
and U5223 (N_5223,N_4075,N_4873);
and U5224 (N_5224,N_4317,N_4416);
and U5225 (N_5225,N_4053,N_4355);
and U5226 (N_5226,N_4426,N_4297);
xor U5227 (N_5227,N_4723,N_4157);
xor U5228 (N_5228,N_4274,N_4413);
nor U5229 (N_5229,N_4829,N_4398);
or U5230 (N_5230,N_4481,N_4600);
or U5231 (N_5231,N_4569,N_4551);
and U5232 (N_5232,N_4924,N_4268);
or U5233 (N_5233,N_4184,N_4202);
nor U5234 (N_5234,N_4298,N_4073);
and U5235 (N_5235,N_4971,N_4525);
xor U5236 (N_5236,N_4785,N_4376);
nand U5237 (N_5237,N_4077,N_4309);
or U5238 (N_5238,N_4011,N_4121);
nand U5239 (N_5239,N_4368,N_4636);
nand U5240 (N_5240,N_4352,N_4859);
nor U5241 (N_5241,N_4587,N_4645);
nor U5242 (N_5242,N_4561,N_4633);
and U5243 (N_5243,N_4996,N_4855);
nor U5244 (N_5244,N_4783,N_4314);
nor U5245 (N_5245,N_4146,N_4687);
nand U5246 (N_5246,N_4945,N_4677);
and U5247 (N_5247,N_4207,N_4758);
xnor U5248 (N_5248,N_4882,N_4291);
and U5249 (N_5249,N_4792,N_4087);
nor U5250 (N_5250,N_4919,N_4691);
or U5251 (N_5251,N_4062,N_4137);
or U5252 (N_5252,N_4707,N_4140);
nand U5253 (N_5253,N_4715,N_4521);
nor U5254 (N_5254,N_4737,N_4851);
and U5255 (N_5255,N_4135,N_4646);
nor U5256 (N_5256,N_4662,N_4703);
nand U5257 (N_5257,N_4949,N_4031);
and U5258 (N_5258,N_4748,N_4754);
and U5259 (N_5259,N_4589,N_4615);
or U5260 (N_5260,N_4736,N_4424);
nor U5261 (N_5261,N_4599,N_4711);
nor U5262 (N_5262,N_4407,N_4938);
nand U5263 (N_5263,N_4386,N_4139);
nor U5264 (N_5264,N_4332,N_4304);
or U5265 (N_5265,N_4832,N_4315);
nand U5266 (N_5266,N_4160,N_4109);
nand U5267 (N_5267,N_4162,N_4517);
or U5268 (N_5268,N_4100,N_4500);
nor U5269 (N_5269,N_4380,N_4951);
nor U5270 (N_5270,N_4131,N_4452);
nand U5271 (N_5271,N_4423,N_4744);
nand U5272 (N_5272,N_4806,N_4570);
and U5273 (N_5273,N_4574,N_4264);
or U5274 (N_5274,N_4341,N_4166);
and U5275 (N_5275,N_4070,N_4182);
nor U5276 (N_5276,N_4194,N_4729);
nor U5277 (N_5277,N_4061,N_4932);
xor U5278 (N_5278,N_4854,N_4827);
nand U5279 (N_5279,N_4621,N_4892);
nand U5280 (N_5280,N_4535,N_4029);
nand U5281 (N_5281,N_4088,N_4568);
nand U5282 (N_5282,N_4065,N_4852);
or U5283 (N_5283,N_4929,N_4927);
or U5284 (N_5284,N_4381,N_4499);
and U5285 (N_5285,N_4338,N_4248);
xnor U5286 (N_5286,N_4275,N_4063);
xor U5287 (N_5287,N_4382,N_4459);
xor U5288 (N_5288,N_4720,N_4244);
and U5289 (N_5289,N_4537,N_4717);
or U5290 (N_5290,N_4955,N_4954);
xnor U5291 (N_5291,N_4821,N_4883);
xor U5292 (N_5292,N_4473,N_4033);
nor U5293 (N_5293,N_4085,N_4127);
nor U5294 (N_5294,N_4554,N_4092);
nor U5295 (N_5295,N_4862,N_4650);
nor U5296 (N_5296,N_4898,N_4913);
or U5297 (N_5297,N_4669,N_4536);
xnor U5298 (N_5298,N_4719,N_4215);
or U5299 (N_5299,N_4181,N_4747);
nor U5300 (N_5300,N_4879,N_4987);
or U5301 (N_5301,N_4860,N_4836);
nor U5302 (N_5302,N_4968,N_4546);
and U5303 (N_5303,N_4890,N_4506);
or U5304 (N_5304,N_4524,N_4625);
xor U5305 (N_5305,N_4914,N_4675);
or U5306 (N_5306,N_4366,N_4629);
and U5307 (N_5307,N_4503,N_4226);
nor U5308 (N_5308,N_4450,N_4673);
nor U5309 (N_5309,N_4211,N_4480);
xor U5310 (N_5310,N_4915,N_4284);
nor U5311 (N_5311,N_4652,N_4527);
nor U5312 (N_5312,N_4745,N_4582);
nor U5313 (N_5313,N_4647,N_4038);
xnor U5314 (N_5314,N_4731,N_4455);
and U5315 (N_5315,N_4353,N_4963);
or U5316 (N_5316,N_4387,N_4335);
and U5317 (N_5317,N_4138,N_4931);
nor U5318 (N_5318,N_4257,N_4171);
and U5319 (N_5319,N_4518,N_4222);
nor U5320 (N_5320,N_4874,N_4446);
or U5321 (N_5321,N_4510,N_4475);
nand U5322 (N_5322,N_4330,N_4378);
nand U5323 (N_5323,N_4571,N_4333);
or U5324 (N_5324,N_4464,N_4934);
or U5325 (N_5325,N_4054,N_4786);
or U5326 (N_5326,N_4654,N_4976);
xor U5327 (N_5327,N_4958,N_4910);
and U5328 (N_5328,N_4007,N_4679);
nand U5329 (N_5329,N_4050,N_4367);
and U5330 (N_5330,N_4906,N_4084);
nand U5331 (N_5331,N_4639,N_4922);
and U5332 (N_5332,N_4144,N_4196);
nand U5333 (N_5333,N_4603,N_4682);
nor U5334 (N_5334,N_4845,N_4491);
nand U5335 (N_5335,N_4740,N_4383);
and U5336 (N_5336,N_4584,N_4970);
or U5337 (N_5337,N_4451,N_4106);
nor U5338 (N_5338,N_4114,N_4457);
or U5339 (N_5339,N_4273,N_4727);
nor U5340 (N_5340,N_4454,N_4025);
and U5341 (N_5341,N_4093,N_4939);
nand U5342 (N_5342,N_4590,N_4555);
or U5343 (N_5343,N_4320,N_4263);
nand U5344 (N_5344,N_4170,N_4300);
and U5345 (N_5345,N_4233,N_4900);
xnor U5346 (N_5346,N_4607,N_4935);
and U5347 (N_5347,N_4272,N_4440);
or U5348 (N_5348,N_4575,N_4493);
or U5349 (N_5349,N_4733,N_4681);
nor U5350 (N_5350,N_4693,N_4041);
nor U5351 (N_5351,N_4395,N_4404);
xnor U5352 (N_5352,N_4994,N_4608);
and U5353 (N_5353,N_4728,N_4743);
xor U5354 (N_5354,N_4066,N_4209);
nand U5355 (N_5355,N_4573,N_4839);
xnor U5356 (N_5356,N_4937,N_4755);
nor U5357 (N_5357,N_4818,N_4428);
or U5358 (N_5358,N_4028,N_4888);
and U5359 (N_5359,N_4942,N_4339);
nand U5360 (N_5360,N_4151,N_4557);
or U5361 (N_5361,N_4911,N_4674);
or U5362 (N_5362,N_4580,N_4002);
nor U5363 (N_5363,N_4197,N_4722);
or U5364 (N_5364,N_4293,N_4490);
nor U5365 (N_5365,N_4391,N_4331);
xnor U5366 (N_5366,N_4432,N_4095);
and U5367 (N_5367,N_4083,N_4076);
nor U5368 (N_5368,N_4236,N_4133);
or U5369 (N_5369,N_4908,N_4846);
and U5370 (N_5370,N_4014,N_4326);
nand U5371 (N_5371,N_4726,N_4795);
and U5372 (N_5372,N_4363,N_4439);
or U5373 (N_5373,N_4015,N_4321);
nor U5374 (N_5374,N_4393,N_4130);
and U5375 (N_5375,N_4174,N_4502);
xnor U5376 (N_5376,N_4721,N_4771);
nand U5377 (N_5377,N_4746,N_4278);
or U5378 (N_5378,N_4767,N_4497);
nor U5379 (N_5379,N_4477,N_4509);
nand U5380 (N_5380,N_4685,N_4991);
xor U5381 (N_5381,N_4448,N_4702);
nand U5382 (N_5382,N_4136,N_4616);
or U5383 (N_5383,N_4668,N_4534);
nor U5384 (N_5384,N_4916,N_4348);
nor U5385 (N_5385,N_4670,N_4725);
nor U5386 (N_5386,N_4020,N_4665);
or U5387 (N_5387,N_4672,N_4192);
nor U5388 (N_5388,N_4308,N_4917);
nor U5389 (N_5389,N_4617,N_4018);
xor U5390 (N_5390,N_4103,N_4978);
or U5391 (N_5391,N_4059,N_4866);
nor U5392 (N_5392,N_4361,N_4921);
nand U5393 (N_5393,N_4807,N_4488);
nand U5394 (N_5394,N_4186,N_4823);
nand U5395 (N_5395,N_4696,N_4003);
nand U5396 (N_5396,N_4596,N_4980);
and U5397 (N_5397,N_4700,N_4472);
or U5398 (N_5398,N_4626,N_4017);
or U5399 (N_5399,N_4301,N_4282);
xnor U5400 (N_5400,N_4583,N_4641);
and U5401 (N_5401,N_4185,N_4578);
or U5402 (N_5402,N_4142,N_4868);
or U5403 (N_5403,N_4712,N_4655);
nor U5404 (N_5404,N_4602,N_4850);
nand U5405 (N_5405,N_4371,N_4875);
and U5406 (N_5406,N_4340,N_4560);
nor U5407 (N_5407,N_4227,N_4206);
nand U5408 (N_5408,N_4336,N_4957);
xnor U5409 (N_5409,N_4780,N_4458);
and U5410 (N_5410,N_4195,N_4588);
or U5411 (N_5411,N_4634,N_4453);
nand U5412 (N_5412,N_4666,N_4258);
nor U5413 (N_5413,N_4533,N_4249);
or U5414 (N_5414,N_4986,N_4134);
xnor U5415 (N_5415,N_4373,N_4155);
or U5416 (N_5416,N_4425,N_4316);
nand U5417 (N_5417,N_4926,N_4082);
and U5418 (N_5418,N_4835,N_4463);
nor U5419 (N_5419,N_4250,N_4694);
xnor U5420 (N_5420,N_4741,N_4789);
xor U5421 (N_5421,N_4161,N_4993);
and U5422 (N_5422,N_4784,N_4762);
and U5423 (N_5423,N_4623,N_4894);
or U5424 (N_5424,N_4260,N_4760);
nand U5425 (N_5425,N_4431,N_4545);
xor U5426 (N_5426,N_4635,N_4663);
and U5427 (N_5427,N_4405,N_4191);
nor U5428 (N_5428,N_4252,N_4609);
and U5429 (N_5429,N_4992,N_4999);
nand U5430 (N_5430,N_4941,N_4390);
nor U5431 (N_5431,N_4266,N_4853);
and U5432 (N_5432,N_4496,N_4417);
nor U5433 (N_5433,N_4141,N_4044);
or U5434 (N_5434,N_4985,N_4126);
and U5435 (N_5435,N_4125,N_4975);
or U5436 (N_5436,N_4787,N_4897);
and U5437 (N_5437,N_4965,N_4794);
or U5438 (N_5438,N_4950,N_4071);
and U5439 (N_5439,N_4409,N_4232);
and U5440 (N_5440,N_4904,N_4591);
nor U5441 (N_5441,N_4610,N_4406);
nor U5442 (N_5442,N_4013,N_4086);
and U5443 (N_5443,N_4982,N_4622);
nand U5444 (N_5444,N_4415,N_4285);
and U5445 (N_5445,N_4412,N_4419);
or U5446 (N_5446,N_4511,N_4436);
or U5447 (N_5447,N_4989,N_4830);
or U5448 (N_5448,N_4896,N_4814);
and U5449 (N_5449,N_4461,N_4943);
nand U5450 (N_5450,N_4030,N_4592);
nand U5451 (N_5451,N_4051,N_4228);
nand U5452 (N_5452,N_4442,N_4738);
nor U5453 (N_5453,N_4757,N_4467);
nand U5454 (N_5454,N_4492,N_4844);
or U5455 (N_5455,N_4605,N_4172);
nand U5456 (N_5456,N_4281,N_4946);
or U5457 (N_5457,N_4552,N_4403);
and U5458 (N_5458,N_4277,N_4805);
or U5459 (N_5459,N_4280,N_4613);
and U5460 (N_5460,N_4261,N_4443);
xor U5461 (N_5461,N_4936,N_4080);
nand U5462 (N_5462,N_4090,N_4544);
nor U5463 (N_5463,N_4444,N_4262);
or U5464 (N_5464,N_4595,N_4735);
nand U5465 (N_5465,N_4631,N_4027);
or U5466 (N_5466,N_4322,N_4049);
xnor U5467 (N_5467,N_4360,N_4658);
xor U5468 (N_5468,N_4318,N_4766);
or U5469 (N_5469,N_4886,N_4643);
nor U5470 (N_5470,N_4777,N_4422);
nand U5471 (N_5471,N_4091,N_4484);
nand U5472 (N_5472,N_4903,N_4117);
nand U5473 (N_5473,N_4421,N_4514);
nor U5474 (N_5474,N_4216,N_4203);
xor U5475 (N_5475,N_4997,N_4998);
or U5476 (N_5476,N_4542,N_4891);
nor U5477 (N_5477,N_4526,N_4474);
nor U5478 (N_5478,N_4176,N_4173);
nand U5479 (N_5479,N_4253,N_4132);
or U5480 (N_5480,N_4009,N_4697);
or U5481 (N_5481,N_4538,N_4489);
nand U5482 (N_5482,N_4778,N_4512);
nand U5483 (N_5483,N_4734,N_4960);
nand U5484 (N_5484,N_4046,N_4952);
nand U5485 (N_5485,N_4024,N_4739);
nand U5486 (N_5486,N_4505,N_4267);
nand U5487 (N_5487,N_4594,N_4799);
nor U5488 (N_5488,N_4235,N_4001);
and U5489 (N_5489,N_4385,N_4559);
or U5490 (N_5490,N_4520,N_4553);
nand U5491 (N_5491,N_4811,N_4241);
and U5492 (N_5492,N_4445,N_4486);
xor U5493 (N_5493,N_4334,N_4630);
nor U5494 (N_5494,N_4096,N_4379);
nand U5495 (N_5495,N_4208,N_4470);
and U5496 (N_5496,N_4501,N_4877);
nand U5497 (N_5497,N_4292,N_4359);
or U5498 (N_5498,N_4977,N_4218);
nor U5499 (N_5499,N_4487,N_4848);
nand U5500 (N_5500,N_4175,N_4833);
nor U5501 (N_5501,N_4342,N_4154);
and U5502 (N_5502,N_4826,N_4063);
or U5503 (N_5503,N_4840,N_4868);
or U5504 (N_5504,N_4658,N_4496);
and U5505 (N_5505,N_4337,N_4928);
or U5506 (N_5506,N_4781,N_4727);
or U5507 (N_5507,N_4535,N_4855);
or U5508 (N_5508,N_4568,N_4792);
and U5509 (N_5509,N_4333,N_4372);
and U5510 (N_5510,N_4917,N_4714);
nor U5511 (N_5511,N_4634,N_4612);
and U5512 (N_5512,N_4913,N_4576);
xor U5513 (N_5513,N_4947,N_4930);
or U5514 (N_5514,N_4965,N_4570);
nor U5515 (N_5515,N_4283,N_4179);
nor U5516 (N_5516,N_4789,N_4443);
nor U5517 (N_5517,N_4963,N_4332);
and U5518 (N_5518,N_4135,N_4394);
nor U5519 (N_5519,N_4203,N_4944);
nor U5520 (N_5520,N_4090,N_4933);
or U5521 (N_5521,N_4195,N_4898);
nor U5522 (N_5522,N_4914,N_4443);
and U5523 (N_5523,N_4689,N_4120);
nand U5524 (N_5524,N_4691,N_4605);
xor U5525 (N_5525,N_4893,N_4645);
nand U5526 (N_5526,N_4528,N_4277);
or U5527 (N_5527,N_4986,N_4868);
and U5528 (N_5528,N_4057,N_4039);
and U5529 (N_5529,N_4819,N_4011);
and U5530 (N_5530,N_4678,N_4755);
xor U5531 (N_5531,N_4587,N_4927);
nand U5532 (N_5532,N_4888,N_4562);
xor U5533 (N_5533,N_4776,N_4827);
nor U5534 (N_5534,N_4316,N_4704);
nor U5535 (N_5535,N_4591,N_4844);
nor U5536 (N_5536,N_4434,N_4145);
and U5537 (N_5537,N_4651,N_4163);
nand U5538 (N_5538,N_4862,N_4473);
nand U5539 (N_5539,N_4793,N_4238);
or U5540 (N_5540,N_4764,N_4620);
nand U5541 (N_5541,N_4505,N_4813);
and U5542 (N_5542,N_4684,N_4271);
nand U5543 (N_5543,N_4228,N_4723);
and U5544 (N_5544,N_4658,N_4141);
xor U5545 (N_5545,N_4124,N_4313);
xnor U5546 (N_5546,N_4618,N_4037);
or U5547 (N_5547,N_4580,N_4604);
and U5548 (N_5548,N_4889,N_4268);
nand U5549 (N_5549,N_4326,N_4129);
or U5550 (N_5550,N_4680,N_4689);
nand U5551 (N_5551,N_4331,N_4453);
nor U5552 (N_5552,N_4078,N_4104);
nor U5553 (N_5553,N_4541,N_4510);
nor U5554 (N_5554,N_4110,N_4054);
and U5555 (N_5555,N_4988,N_4600);
nor U5556 (N_5556,N_4746,N_4116);
nor U5557 (N_5557,N_4022,N_4981);
or U5558 (N_5558,N_4725,N_4951);
nor U5559 (N_5559,N_4908,N_4727);
nor U5560 (N_5560,N_4243,N_4687);
or U5561 (N_5561,N_4789,N_4821);
nor U5562 (N_5562,N_4571,N_4057);
or U5563 (N_5563,N_4672,N_4822);
nor U5564 (N_5564,N_4014,N_4129);
or U5565 (N_5565,N_4743,N_4856);
and U5566 (N_5566,N_4138,N_4409);
or U5567 (N_5567,N_4695,N_4335);
nand U5568 (N_5568,N_4565,N_4286);
and U5569 (N_5569,N_4453,N_4096);
and U5570 (N_5570,N_4204,N_4132);
and U5571 (N_5571,N_4779,N_4842);
and U5572 (N_5572,N_4214,N_4136);
or U5573 (N_5573,N_4600,N_4715);
nor U5574 (N_5574,N_4129,N_4441);
nor U5575 (N_5575,N_4847,N_4941);
xnor U5576 (N_5576,N_4357,N_4618);
and U5577 (N_5577,N_4224,N_4959);
xnor U5578 (N_5578,N_4988,N_4456);
nand U5579 (N_5579,N_4412,N_4134);
and U5580 (N_5580,N_4693,N_4972);
and U5581 (N_5581,N_4448,N_4718);
or U5582 (N_5582,N_4410,N_4252);
and U5583 (N_5583,N_4287,N_4716);
and U5584 (N_5584,N_4449,N_4144);
or U5585 (N_5585,N_4867,N_4434);
or U5586 (N_5586,N_4736,N_4123);
nand U5587 (N_5587,N_4631,N_4686);
or U5588 (N_5588,N_4552,N_4379);
nor U5589 (N_5589,N_4299,N_4776);
and U5590 (N_5590,N_4547,N_4220);
and U5591 (N_5591,N_4638,N_4219);
and U5592 (N_5592,N_4530,N_4640);
and U5593 (N_5593,N_4638,N_4519);
nand U5594 (N_5594,N_4424,N_4296);
nand U5595 (N_5595,N_4838,N_4708);
or U5596 (N_5596,N_4812,N_4929);
or U5597 (N_5597,N_4786,N_4400);
nor U5598 (N_5598,N_4995,N_4760);
or U5599 (N_5599,N_4328,N_4580);
and U5600 (N_5600,N_4509,N_4709);
nand U5601 (N_5601,N_4957,N_4387);
or U5602 (N_5602,N_4377,N_4636);
or U5603 (N_5603,N_4954,N_4760);
nand U5604 (N_5604,N_4789,N_4774);
nor U5605 (N_5605,N_4774,N_4018);
xor U5606 (N_5606,N_4752,N_4730);
nand U5607 (N_5607,N_4225,N_4697);
and U5608 (N_5608,N_4575,N_4041);
nor U5609 (N_5609,N_4131,N_4447);
or U5610 (N_5610,N_4798,N_4689);
nor U5611 (N_5611,N_4006,N_4416);
nor U5612 (N_5612,N_4587,N_4634);
nand U5613 (N_5613,N_4621,N_4648);
nand U5614 (N_5614,N_4622,N_4108);
or U5615 (N_5615,N_4745,N_4545);
nor U5616 (N_5616,N_4906,N_4550);
nand U5617 (N_5617,N_4415,N_4267);
and U5618 (N_5618,N_4710,N_4711);
nor U5619 (N_5619,N_4113,N_4589);
xor U5620 (N_5620,N_4464,N_4841);
nand U5621 (N_5621,N_4979,N_4445);
and U5622 (N_5622,N_4196,N_4850);
and U5623 (N_5623,N_4291,N_4877);
nor U5624 (N_5624,N_4812,N_4622);
nor U5625 (N_5625,N_4644,N_4876);
xor U5626 (N_5626,N_4405,N_4443);
nor U5627 (N_5627,N_4918,N_4977);
and U5628 (N_5628,N_4508,N_4011);
nand U5629 (N_5629,N_4925,N_4424);
nand U5630 (N_5630,N_4076,N_4032);
or U5631 (N_5631,N_4447,N_4289);
xor U5632 (N_5632,N_4697,N_4252);
xor U5633 (N_5633,N_4665,N_4359);
nor U5634 (N_5634,N_4241,N_4910);
or U5635 (N_5635,N_4602,N_4432);
nand U5636 (N_5636,N_4473,N_4300);
or U5637 (N_5637,N_4445,N_4179);
xnor U5638 (N_5638,N_4155,N_4687);
and U5639 (N_5639,N_4382,N_4029);
and U5640 (N_5640,N_4752,N_4974);
or U5641 (N_5641,N_4899,N_4675);
xnor U5642 (N_5642,N_4554,N_4481);
nand U5643 (N_5643,N_4574,N_4130);
nand U5644 (N_5644,N_4278,N_4115);
nor U5645 (N_5645,N_4117,N_4515);
or U5646 (N_5646,N_4996,N_4864);
and U5647 (N_5647,N_4605,N_4963);
or U5648 (N_5648,N_4251,N_4540);
or U5649 (N_5649,N_4275,N_4937);
xor U5650 (N_5650,N_4867,N_4812);
or U5651 (N_5651,N_4956,N_4593);
or U5652 (N_5652,N_4492,N_4338);
xnor U5653 (N_5653,N_4119,N_4887);
and U5654 (N_5654,N_4270,N_4283);
nor U5655 (N_5655,N_4105,N_4525);
and U5656 (N_5656,N_4895,N_4998);
and U5657 (N_5657,N_4149,N_4753);
and U5658 (N_5658,N_4313,N_4444);
nand U5659 (N_5659,N_4864,N_4935);
nor U5660 (N_5660,N_4810,N_4779);
xor U5661 (N_5661,N_4982,N_4152);
nand U5662 (N_5662,N_4517,N_4576);
nand U5663 (N_5663,N_4789,N_4910);
nor U5664 (N_5664,N_4860,N_4678);
nand U5665 (N_5665,N_4938,N_4914);
and U5666 (N_5666,N_4196,N_4781);
nand U5667 (N_5667,N_4258,N_4038);
and U5668 (N_5668,N_4405,N_4208);
nand U5669 (N_5669,N_4412,N_4065);
or U5670 (N_5670,N_4444,N_4337);
nor U5671 (N_5671,N_4056,N_4458);
or U5672 (N_5672,N_4121,N_4556);
and U5673 (N_5673,N_4989,N_4522);
or U5674 (N_5674,N_4465,N_4048);
and U5675 (N_5675,N_4306,N_4278);
or U5676 (N_5676,N_4476,N_4355);
or U5677 (N_5677,N_4586,N_4435);
nand U5678 (N_5678,N_4218,N_4176);
nand U5679 (N_5679,N_4231,N_4680);
or U5680 (N_5680,N_4688,N_4310);
nor U5681 (N_5681,N_4383,N_4323);
nand U5682 (N_5682,N_4759,N_4997);
or U5683 (N_5683,N_4578,N_4194);
nor U5684 (N_5684,N_4671,N_4494);
nand U5685 (N_5685,N_4067,N_4513);
xnor U5686 (N_5686,N_4415,N_4567);
xor U5687 (N_5687,N_4101,N_4198);
and U5688 (N_5688,N_4959,N_4330);
nor U5689 (N_5689,N_4094,N_4058);
nor U5690 (N_5690,N_4316,N_4156);
nand U5691 (N_5691,N_4723,N_4060);
and U5692 (N_5692,N_4280,N_4077);
or U5693 (N_5693,N_4191,N_4002);
or U5694 (N_5694,N_4455,N_4534);
nor U5695 (N_5695,N_4107,N_4254);
nor U5696 (N_5696,N_4508,N_4533);
and U5697 (N_5697,N_4118,N_4856);
nand U5698 (N_5698,N_4793,N_4668);
nor U5699 (N_5699,N_4953,N_4485);
or U5700 (N_5700,N_4216,N_4010);
nand U5701 (N_5701,N_4255,N_4367);
and U5702 (N_5702,N_4456,N_4788);
or U5703 (N_5703,N_4781,N_4717);
nor U5704 (N_5704,N_4898,N_4093);
nand U5705 (N_5705,N_4037,N_4888);
nand U5706 (N_5706,N_4198,N_4369);
nand U5707 (N_5707,N_4180,N_4384);
nor U5708 (N_5708,N_4744,N_4856);
or U5709 (N_5709,N_4641,N_4775);
nor U5710 (N_5710,N_4190,N_4908);
and U5711 (N_5711,N_4357,N_4647);
xnor U5712 (N_5712,N_4371,N_4166);
xnor U5713 (N_5713,N_4249,N_4933);
or U5714 (N_5714,N_4345,N_4994);
nor U5715 (N_5715,N_4011,N_4780);
nand U5716 (N_5716,N_4954,N_4034);
nand U5717 (N_5717,N_4381,N_4140);
and U5718 (N_5718,N_4454,N_4266);
or U5719 (N_5719,N_4621,N_4373);
or U5720 (N_5720,N_4646,N_4104);
or U5721 (N_5721,N_4127,N_4583);
nand U5722 (N_5722,N_4470,N_4756);
nor U5723 (N_5723,N_4230,N_4138);
nor U5724 (N_5724,N_4660,N_4843);
nor U5725 (N_5725,N_4558,N_4691);
xnor U5726 (N_5726,N_4800,N_4545);
xor U5727 (N_5727,N_4733,N_4282);
xnor U5728 (N_5728,N_4305,N_4338);
xnor U5729 (N_5729,N_4887,N_4678);
or U5730 (N_5730,N_4024,N_4150);
nand U5731 (N_5731,N_4873,N_4469);
nand U5732 (N_5732,N_4687,N_4094);
or U5733 (N_5733,N_4474,N_4016);
nor U5734 (N_5734,N_4452,N_4920);
nor U5735 (N_5735,N_4250,N_4886);
nor U5736 (N_5736,N_4791,N_4939);
nor U5737 (N_5737,N_4148,N_4404);
xnor U5738 (N_5738,N_4958,N_4226);
or U5739 (N_5739,N_4853,N_4481);
nand U5740 (N_5740,N_4517,N_4859);
or U5741 (N_5741,N_4406,N_4190);
and U5742 (N_5742,N_4569,N_4842);
or U5743 (N_5743,N_4774,N_4411);
or U5744 (N_5744,N_4057,N_4851);
or U5745 (N_5745,N_4874,N_4410);
nor U5746 (N_5746,N_4886,N_4692);
nand U5747 (N_5747,N_4868,N_4140);
nor U5748 (N_5748,N_4002,N_4776);
or U5749 (N_5749,N_4847,N_4848);
nor U5750 (N_5750,N_4688,N_4058);
and U5751 (N_5751,N_4485,N_4934);
and U5752 (N_5752,N_4723,N_4863);
nand U5753 (N_5753,N_4648,N_4063);
nand U5754 (N_5754,N_4831,N_4096);
nand U5755 (N_5755,N_4248,N_4869);
nor U5756 (N_5756,N_4127,N_4163);
and U5757 (N_5757,N_4191,N_4576);
xnor U5758 (N_5758,N_4598,N_4910);
or U5759 (N_5759,N_4436,N_4641);
xor U5760 (N_5760,N_4365,N_4563);
nor U5761 (N_5761,N_4174,N_4701);
xor U5762 (N_5762,N_4614,N_4217);
or U5763 (N_5763,N_4773,N_4200);
and U5764 (N_5764,N_4377,N_4374);
and U5765 (N_5765,N_4628,N_4270);
nand U5766 (N_5766,N_4963,N_4369);
or U5767 (N_5767,N_4167,N_4395);
nor U5768 (N_5768,N_4302,N_4371);
and U5769 (N_5769,N_4607,N_4994);
nor U5770 (N_5770,N_4677,N_4622);
nor U5771 (N_5771,N_4801,N_4436);
or U5772 (N_5772,N_4094,N_4328);
xnor U5773 (N_5773,N_4207,N_4969);
or U5774 (N_5774,N_4038,N_4137);
or U5775 (N_5775,N_4112,N_4253);
and U5776 (N_5776,N_4727,N_4759);
nand U5777 (N_5777,N_4893,N_4974);
nand U5778 (N_5778,N_4526,N_4174);
and U5779 (N_5779,N_4748,N_4702);
xnor U5780 (N_5780,N_4095,N_4258);
nand U5781 (N_5781,N_4480,N_4584);
nand U5782 (N_5782,N_4852,N_4466);
nor U5783 (N_5783,N_4979,N_4854);
xor U5784 (N_5784,N_4873,N_4245);
and U5785 (N_5785,N_4390,N_4716);
and U5786 (N_5786,N_4480,N_4024);
nor U5787 (N_5787,N_4018,N_4732);
nand U5788 (N_5788,N_4171,N_4235);
nor U5789 (N_5789,N_4619,N_4566);
xnor U5790 (N_5790,N_4861,N_4699);
or U5791 (N_5791,N_4481,N_4065);
nor U5792 (N_5792,N_4779,N_4824);
nor U5793 (N_5793,N_4272,N_4027);
or U5794 (N_5794,N_4094,N_4951);
nand U5795 (N_5795,N_4483,N_4844);
or U5796 (N_5796,N_4910,N_4989);
or U5797 (N_5797,N_4097,N_4762);
and U5798 (N_5798,N_4096,N_4119);
nand U5799 (N_5799,N_4561,N_4131);
nor U5800 (N_5800,N_4488,N_4233);
nor U5801 (N_5801,N_4374,N_4682);
nand U5802 (N_5802,N_4514,N_4331);
and U5803 (N_5803,N_4916,N_4654);
nand U5804 (N_5804,N_4396,N_4805);
xnor U5805 (N_5805,N_4474,N_4022);
xor U5806 (N_5806,N_4874,N_4437);
nor U5807 (N_5807,N_4662,N_4766);
nor U5808 (N_5808,N_4777,N_4660);
nor U5809 (N_5809,N_4754,N_4994);
and U5810 (N_5810,N_4181,N_4188);
or U5811 (N_5811,N_4878,N_4931);
and U5812 (N_5812,N_4336,N_4713);
xor U5813 (N_5813,N_4271,N_4418);
or U5814 (N_5814,N_4864,N_4146);
nor U5815 (N_5815,N_4164,N_4630);
nor U5816 (N_5816,N_4148,N_4469);
or U5817 (N_5817,N_4309,N_4305);
nand U5818 (N_5818,N_4258,N_4552);
or U5819 (N_5819,N_4557,N_4301);
and U5820 (N_5820,N_4037,N_4195);
nand U5821 (N_5821,N_4229,N_4452);
nor U5822 (N_5822,N_4500,N_4191);
nand U5823 (N_5823,N_4271,N_4755);
or U5824 (N_5824,N_4561,N_4762);
nand U5825 (N_5825,N_4771,N_4380);
or U5826 (N_5826,N_4815,N_4929);
and U5827 (N_5827,N_4551,N_4633);
xor U5828 (N_5828,N_4251,N_4637);
nor U5829 (N_5829,N_4795,N_4674);
nand U5830 (N_5830,N_4266,N_4889);
nor U5831 (N_5831,N_4887,N_4479);
nor U5832 (N_5832,N_4372,N_4812);
and U5833 (N_5833,N_4487,N_4213);
and U5834 (N_5834,N_4932,N_4624);
and U5835 (N_5835,N_4265,N_4990);
nand U5836 (N_5836,N_4203,N_4472);
or U5837 (N_5837,N_4769,N_4292);
or U5838 (N_5838,N_4527,N_4295);
and U5839 (N_5839,N_4170,N_4828);
or U5840 (N_5840,N_4627,N_4482);
nand U5841 (N_5841,N_4939,N_4884);
or U5842 (N_5842,N_4603,N_4686);
or U5843 (N_5843,N_4446,N_4858);
or U5844 (N_5844,N_4853,N_4927);
nand U5845 (N_5845,N_4061,N_4134);
xor U5846 (N_5846,N_4949,N_4756);
and U5847 (N_5847,N_4006,N_4670);
nand U5848 (N_5848,N_4194,N_4502);
and U5849 (N_5849,N_4463,N_4148);
and U5850 (N_5850,N_4255,N_4685);
nand U5851 (N_5851,N_4674,N_4287);
nor U5852 (N_5852,N_4730,N_4086);
or U5853 (N_5853,N_4584,N_4051);
nor U5854 (N_5854,N_4193,N_4962);
or U5855 (N_5855,N_4545,N_4181);
or U5856 (N_5856,N_4380,N_4846);
nor U5857 (N_5857,N_4448,N_4660);
nor U5858 (N_5858,N_4067,N_4794);
nand U5859 (N_5859,N_4596,N_4553);
nor U5860 (N_5860,N_4276,N_4219);
nor U5861 (N_5861,N_4506,N_4367);
or U5862 (N_5862,N_4653,N_4334);
nor U5863 (N_5863,N_4325,N_4374);
or U5864 (N_5864,N_4024,N_4103);
nand U5865 (N_5865,N_4420,N_4388);
or U5866 (N_5866,N_4938,N_4730);
or U5867 (N_5867,N_4498,N_4319);
nor U5868 (N_5868,N_4120,N_4899);
nand U5869 (N_5869,N_4573,N_4163);
or U5870 (N_5870,N_4399,N_4810);
and U5871 (N_5871,N_4735,N_4409);
xor U5872 (N_5872,N_4088,N_4764);
nor U5873 (N_5873,N_4571,N_4477);
xor U5874 (N_5874,N_4965,N_4973);
and U5875 (N_5875,N_4388,N_4542);
nand U5876 (N_5876,N_4138,N_4141);
and U5877 (N_5877,N_4997,N_4022);
nand U5878 (N_5878,N_4774,N_4745);
and U5879 (N_5879,N_4585,N_4366);
or U5880 (N_5880,N_4561,N_4405);
and U5881 (N_5881,N_4157,N_4898);
nor U5882 (N_5882,N_4986,N_4506);
nor U5883 (N_5883,N_4933,N_4883);
and U5884 (N_5884,N_4221,N_4976);
nand U5885 (N_5885,N_4941,N_4513);
and U5886 (N_5886,N_4179,N_4138);
and U5887 (N_5887,N_4581,N_4114);
nand U5888 (N_5888,N_4064,N_4249);
nand U5889 (N_5889,N_4197,N_4043);
or U5890 (N_5890,N_4653,N_4433);
or U5891 (N_5891,N_4090,N_4700);
xor U5892 (N_5892,N_4792,N_4612);
nand U5893 (N_5893,N_4509,N_4414);
nor U5894 (N_5894,N_4197,N_4011);
nand U5895 (N_5895,N_4918,N_4811);
or U5896 (N_5896,N_4200,N_4994);
nor U5897 (N_5897,N_4320,N_4758);
and U5898 (N_5898,N_4154,N_4543);
nand U5899 (N_5899,N_4090,N_4101);
and U5900 (N_5900,N_4322,N_4812);
and U5901 (N_5901,N_4865,N_4612);
nor U5902 (N_5902,N_4774,N_4838);
and U5903 (N_5903,N_4895,N_4258);
nor U5904 (N_5904,N_4224,N_4463);
or U5905 (N_5905,N_4288,N_4345);
and U5906 (N_5906,N_4977,N_4985);
or U5907 (N_5907,N_4547,N_4211);
or U5908 (N_5908,N_4410,N_4663);
and U5909 (N_5909,N_4369,N_4629);
nor U5910 (N_5910,N_4608,N_4321);
nor U5911 (N_5911,N_4166,N_4053);
or U5912 (N_5912,N_4047,N_4176);
or U5913 (N_5913,N_4885,N_4413);
or U5914 (N_5914,N_4869,N_4755);
xor U5915 (N_5915,N_4393,N_4850);
or U5916 (N_5916,N_4657,N_4929);
xnor U5917 (N_5917,N_4826,N_4193);
or U5918 (N_5918,N_4865,N_4245);
nand U5919 (N_5919,N_4899,N_4777);
nand U5920 (N_5920,N_4396,N_4350);
or U5921 (N_5921,N_4996,N_4572);
or U5922 (N_5922,N_4059,N_4700);
or U5923 (N_5923,N_4586,N_4483);
or U5924 (N_5924,N_4460,N_4068);
nor U5925 (N_5925,N_4582,N_4980);
nor U5926 (N_5926,N_4974,N_4620);
nand U5927 (N_5927,N_4786,N_4002);
xnor U5928 (N_5928,N_4381,N_4131);
or U5929 (N_5929,N_4223,N_4293);
nand U5930 (N_5930,N_4733,N_4348);
and U5931 (N_5931,N_4595,N_4351);
nand U5932 (N_5932,N_4443,N_4795);
and U5933 (N_5933,N_4721,N_4391);
and U5934 (N_5934,N_4713,N_4553);
and U5935 (N_5935,N_4997,N_4436);
nand U5936 (N_5936,N_4130,N_4972);
nand U5937 (N_5937,N_4640,N_4613);
xor U5938 (N_5938,N_4290,N_4546);
or U5939 (N_5939,N_4708,N_4395);
and U5940 (N_5940,N_4233,N_4334);
xor U5941 (N_5941,N_4504,N_4717);
nand U5942 (N_5942,N_4432,N_4698);
nor U5943 (N_5943,N_4793,N_4752);
nor U5944 (N_5944,N_4865,N_4975);
or U5945 (N_5945,N_4915,N_4465);
and U5946 (N_5946,N_4473,N_4169);
nor U5947 (N_5947,N_4022,N_4297);
nor U5948 (N_5948,N_4220,N_4553);
nand U5949 (N_5949,N_4408,N_4310);
nand U5950 (N_5950,N_4120,N_4901);
xnor U5951 (N_5951,N_4090,N_4887);
nor U5952 (N_5952,N_4681,N_4482);
nor U5953 (N_5953,N_4071,N_4041);
and U5954 (N_5954,N_4684,N_4844);
nor U5955 (N_5955,N_4652,N_4999);
nand U5956 (N_5956,N_4954,N_4930);
and U5957 (N_5957,N_4308,N_4029);
and U5958 (N_5958,N_4008,N_4646);
nand U5959 (N_5959,N_4612,N_4255);
or U5960 (N_5960,N_4207,N_4268);
nor U5961 (N_5961,N_4670,N_4901);
and U5962 (N_5962,N_4862,N_4737);
nand U5963 (N_5963,N_4121,N_4038);
nor U5964 (N_5964,N_4647,N_4047);
xor U5965 (N_5965,N_4150,N_4741);
nand U5966 (N_5966,N_4889,N_4862);
or U5967 (N_5967,N_4885,N_4196);
nor U5968 (N_5968,N_4845,N_4181);
and U5969 (N_5969,N_4311,N_4582);
nand U5970 (N_5970,N_4564,N_4696);
and U5971 (N_5971,N_4533,N_4123);
or U5972 (N_5972,N_4874,N_4335);
nor U5973 (N_5973,N_4985,N_4688);
nand U5974 (N_5974,N_4410,N_4981);
or U5975 (N_5975,N_4511,N_4068);
xnor U5976 (N_5976,N_4320,N_4229);
or U5977 (N_5977,N_4800,N_4732);
nand U5978 (N_5978,N_4311,N_4679);
nor U5979 (N_5979,N_4746,N_4406);
or U5980 (N_5980,N_4945,N_4839);
or U5981 (N_5981,N_4220,N_4475);
or U5982 (N_5982,N_4192,N_4232);
and U5983 (N_5983,N_4765,N_4713);
and U5984 (N_5984,N_4853,N_4371);
nand U5985 (N_5985,N_4433,N_4691);
or U5986 (N_5986,N_4558,N_4656);
nand U5987 (N_5987,N_4284,N_4972);
nor U5988 (N_5988,N_4639,N_4174);
or U5989 (N_5989,N_4972,N_4106);
nand U5990 (N_5990,N_4546,N_4054);
and U5991 (N_5991,N_4265,N_4172);
nand U5992 (N_5992,N_4554,N_4837);
nand U5993 (N_5993,N_4387,N_4849);
and U5994 (N_5994,N_4630,N_4848);
nand U5995 (N_5995,N_4060,N_4024);
nand U5996 (N_5996,N_4556,N_4371);
nand U5997 (N_5997,N_4899,N_4122);
or U5998 (N_5998,N_4085,N_4454);
nand U5999 (N_5999,N_4464,N_4815);
nand U6000 (N_6000,N_5661,N_5976);
nor U6001 (N_6001,N_5488,N_5342);
nor U6002 (N_6002,N_5090,N_5256);
nand U6003 (N_6003,N_5613,N_5428);
and U6004 (N_6004,N_5222,N_5832);
nor U6005 (N_6005,N_5900,N_5260);
or U6006 (N_6006,N_5837,N_5277);
nor U6007 (N_6007,N_5359,N_5340);
or U6008 (N_6008,N_5162,N_5346);
and U6009 (N_6009,N_5586,N_5332);
nor U6010 (N_6010,N_5402,N_5907);
and U6011 (N_6011,N_5878,N_5110);
nor U6012 (N_6012,N_5377,N_5165);
nand U6013 (N_6013,N_5163,N_5019);
and U6014 (N_6014,N_5808,N_5128);
or U6015 (N_6015,N_5458,N_5489);
nand U6016 (N_6016,N_5047,N_5202);
nand U6017 (N_6017,N_5569,N_5461);
xor U6018 (N_6018,N_5008,N_5706);
and U6019 (N_6019,N_5963,N_5682);
nand U6020 (N_6020,N_5105,N_5379);
xor U6021 (N_6021,N_5732,N_5413);
or U6022 (N_6022,N_5739,N_5764);
or U6023 (N_6023,N_5447,N_5647);
nor U6024 (N_6024,N_5574,N_5628);
nand U6025 (N_6025,N_5931,N_5119);
nor U6026 (N_6026,N_5758,N_5098);
nand U6027 (N_6027,N_5812,N_5712);
nand U6028 (N_6028,N_5368,N_5212);
nor U6029 (N_6029,N_5376,N_5895);
and U6030 (N_6030,N_5085,N_5506);
and U6031 (N_6031,N_5692,N_5135);
nand U6032 (N_6032,N_5799,N_5022);
or U6033 (N_6033,N_5631,N_5834);
nor U6034 (N_6034,N_5152,N_5896);
or U6035 (N_6035,N_5718,N_5263);
nand U6036 (N_6036,N_5855,N_5276);
nand U6037 (N_6037,N_5564,N_5510);
or U6038 (N_6038,N_5906,N_5279);
xor U6039 (N_6039,N_5830,N_5897);
nand U6040 (N_6040,N_5169,N_5975);
and U6041 (N_6041,N_5054,N_5030);
and U6042 (N_6042,N_5171,N_5027);
and U6043 (N_6043,N_5814,N_5599);
nor U6044 (N_6044,N_5958,N_5088);
and U6045 (N_6045,N_5516,N_5549);
nor U6046 (N_6046,N_5203,N_5729);
and U6047 (N_6047,N_5410,N_5331);
nor U6048 (N_6048,N_5562,N_5534);
or U6049 (N_6049,N_5733,N_5343);
and U6050 (N_6050,N_5611,N_5716);
nor U6051 (N_6051,N_5490,N_5571);
xor U6052 (N_6052,N_5501,N_5172);
or U6053 (N_6053,N_5391,N_5939);
or U6054 (N_6054,N_5548,N_5318);
nor U6055 (N_6055,N_5969,N_5147);
and U6056 (N_6056,N_5092,N_5221);
nand U6057 (N_6057,N_5558,N_5587);
or U6058 (N_6058,N_5372,N_5794);
or U6059 (N_6059,N_5009,N_5483);
and U6060 (N_6060,N_5339,N_5590);
and U6061 (N_6061,N_5213,N_5151);
xnor U6062 (N_6062,N_5869,N_5679);
and U6063 (N_6063,N_5220,N_5018);
nor U6064 (N_6064,N_5528,N_5080);
and U6065 (N_6065,N_5580,N_5950);
and U6066 (N_6066,N_5772,N_5328);
nand U6067 (N_6067,N_5620,N_5125);
and U6068 (N_6068,N_5341,N_5782);
nand U6069 (N_6069,N_5797,N_5046);
nor U6070 (N_6070,N_5927,N_5314);
or U6071 (N_6071,N_5070,N_5435);
or U6072 (N_6072,N_5743,N_5420);
and U6073 (N_6073,N_5862,N_5703);
or U6074 (N_6074,N_5585,N_5633);
nand U6075 (N_6075,N_5068,N_5485);
nor U6076 (N_6076,N_5984,N_5042);
or U6077 (N_6077,N_5348,N_5638);
nand U6078 (N_6078,N_5871,N_5780);
nor U6079 (N_6079,N_5844,N_5186);
and U6080 (N_6080,N_5311,N_5236);
or U6081 (N_6081,N_5910,N_5595);
nor U6082 (N_6082,N_5394,N_5937);
xor U6083 (N_6083,N_5829,N_5330);
or U6084 (N_6084,N_5769,N_5416);
xnor U6085 (N_6085,N_5144,N_5544);
nand U6086 (N_6086,N_5185,N_5345);
nand U6087 (N_6087,N_5582,N_5691);
nor U6088 (N_6088,N_5879,N_5888);
and U6089 (N_6089,N_5655,N_5828);
xor U6090 (N_6090,N_5398,N_5541);
nor U6091 (N_6091,N_5892,N_5513);
nor U6092 (N_6092,N_5922,N_5473);
or U6093 (N_6093,N_5095,N_5014);
or U6094 (N_6094,N_5678,N_5167);
nor U6095 (N_6095,N_5563,N_5358);
xor U6096 (N_6096,N_5412,N_5781);
xnor U6097 (N_6097,N_5822,N_5357);
nand U6098 (N_6098,N_5217,N_5609);
or U6099 (N_6099,N_5320,N_5818);
or U6100 (N_6100,N_5974,N_5155);
and U6101 (N_6101,N_5324,N_5874);
nand U6102 (N_6102,N_5457,N_5384);
or U6103 (N_6103,N_5353,N_5460);
nor U6104 (N_6104,N_5048,N_5833);
or U6105 (N_6105,N_5920,N_5667);
or U6106 (N_6106,N_5934,N_5399);
nand U6107 (N_6107,N_5577,N_5454);
xnor U6108 (N_6108,N_5816,N_5850);
nand U6109 (N_6109,N_5056,N_5455);
or U6110 (N_6110,N_5363,N_5349);
or U6111 (N_6111,N_5545,N_5940);
nand U6112 (N_6112,N_5023,N_5658);
xnor U6113 (N_6113,N_5811,N_5946);
or U6114 (N_6114,N_5800,N_5366);
nor U6115 (N_6115,N_5573,N_5581);
and U6116 (N_6116,N_5004,N_5375);
or U6117 (N_6117,N_5676,N_5695);
and U6118 (N_6118,N_5329,N_5043);
or U6119 (N_6119,N_5124,N_5928);
and U6120 (N_6120,N_5744,N_5537);
nor U6121 (N_6121,N_5863,N_5189);
or U6122 (N_6122,N_5970,N_5193);
or U6123 (N_6123,N_5943,N_5861);
nand U6124 (N_6124,N_5941,N_5315);
nand U6125 (N_6125,N_5876,N_5400);
nor U6126 (N_6126,N_5336,N_5230);
nand U6127 (N_6127,N_5166,N_5396);
nor U6128 (N_6128,N_5710,N_5696);
and U6129 (N_6129,N_5350,N_5143);
nor U6130 (N_6130,N_5247,N_5326);
xor U6131 (N_6131,N_5737,N_5757);
nor U6132 (N_6132,N_5197,N_5267);
nand U6133 (N_6133,N_5069,N_5752);
and U6134 (N_6134,N_5999,N_5714);
and U6135 (N_6135,N_5231,N_5866);
or U6136 (N_6136,N_5264,N_5079);
or U6137 (N_6137,N_5351,N_5120);
and U6138 (N_6138,N_5687,N_5478);
nand U6139 (N_6139,N_5859,N_5983);
nand U6140 (N_6140,N_5444,N_5181);
nor U6141 (N_6141,N_5873,N_5148);
nand U6142 (N_6142,N_5005,N_5860);
nand U6143 (N_6143,N_5393,N_5037);
nand U6144 (N_6144,N_5530,N_5479);
xor U6145 (N_6145,N_5761,N_5664);
nand U6146 (N_6146,N_5292,N_5041);
nor U6147 (N_6147,N_5272,N_5310);
nand U6148 (N_6148,N_5001,N_5643);
or U6149 (N_6149,N_5367,N_5842);
xnor U6150 (N_6150,N_5361,N_5055);
xor U6151 (N_6151,N_5462,N_5028);
or U6152 (N_6152,N_5604,N_5034);
and U6153 (N_6153,N_5519,N_5547);
nand U6154 (N_6154,N_5387,N_5885);
nor U6155 (N_6155,N_5538,N_5497);
or U6156 (N_6156,N_5791,N_5076);
or U6157 (N_6157,N_5649,N_5415);
nor U6158 (N_6158,N_5550,N_5771);
or U6159 (N_6159,N_5887,N_5721);
or U6160 (N_6160,N_5319,N_5831);
and U6161 (N_6161,N_5565,N_5524);
nor U6162 (N_6162,N_5626,N_5918);
or U6163 (N_6163,N_5566,N_5235);
or U6164 (N_6164,N_5926,N_5734);
and U6165 (N_6165,N_5274,N_5347);
xnor U6166 (N_6166,N_5824,N_5698);
xnor U6167 (N_6167,N_5982,N_5917);
nor U6168 (N_6168,N_5551,N_5073);
nand U6169 (N_6169,N_5039,N_5126);
and U6170 (N_6170,N_5378,N_5063);
nor U6171 (N_6171,N_5841,N_5083);
and U6172 (N_6172,N_5190,N_5215);
or U6173 (N_6173,N_5759,N_5226);
or U6174 (N_6174,N_5060,N_5156);
and U6175 (N_6175,N_5094,N_5663);
or U6176 (N_6176,N_5188,N_5302);
or U6177 (N_6177,N_5443,N_5290);
nand U6178 (N_6178,N_5114,N_5559);
nor U6179 (N_6179,N_5209,N_5527);
xor U6180 (N_6180,N_5949,N_5770);
nand U6181 (N_6181,N_5645,N_5867);
nand U6182 (N_6182,N_5335,N_5921);
or U6183 (N_6183,N_5746,N_5715);
nor U6184 (N_6184,N_5919,N_5059);
and U6185 (N_6185,N_5945,N_5200);
nor U6186 (N_6186,N_5145,N_5262);
and U6187 (N_6187,N_5141,N_5291);
or U6188 (N_6188,N_5015,N_5321);
or U6189 (N_6189,N_5994,N_5623);
nor U6190 (N_6190,N_5929,N_5741);
or U6191 (N_6191,N_5817,N_5433);
or U6192 (N_6192,N_5865,N_5750);
or U6193 (N_6193,N_5726,N_5916);
or U6194 (N_6194,N_5751,N_5255);
nor U6195 (N_6195,N_5049,N_5825);
or U6196 (N_6196,N_5578,N_5334);
and U6197 (N_6197,N_5973,N_5904);
xnor U6198 (N_6198,N_5651,N_5567);
nand U6199 (N_6199,N_5270,N_5204);
xnor U6200 (N_6200,N_5498,N_5187);
nand U6201 (N_6201,N_5608,N_5293);
or U6202 (N_6202,N_5902,N_5074);
nor U6203 (N_6203,N_5851,N_5644);
and U6204 (N_6204,N_5838,N_5421);
nand U6205 (N_6205,N_5453,N_5370);
and U6206 (N_6206,N_5964,N_5522);
nor U6207 (N_6207,N_5300,N_5058);
or U6208 (N_6208,N_5621,N_5096);
nor U6209 (N_6209,N_5777,N_5542);
and U6210 (N_6210,N_5880,N_5669);
nor U6211 (N_6211,N_5438,N_5707);
and U6212 (N_6212,N_5081,N_5773);
nor U6213 (N_6213,N_5630,N_5536);
or U6214 (N_6214,N_5688,N_5077);
or U6215 (N_6215,N_5789,N_5680);
nand U6216 (N_6216,N_5670,N_5281);
and U6217 (N_6217,N_5052,N_5464);
or U6218 (N_6218,N_5675,N_5965);
nand U6219 (N_6219,N_5344,N_5507);
or U6220 (N_6220,N_5233,N_5955);
xnor U6221 (N_6221,N_5966,N_5295);
nand U6222 (N_6222,N_5409,N_5304);
nor U6223 (N_6223,N_5404,N_5557);
nand U6224 (N_6224,N_5252,N_5427);
or U6225 (N_6225,N_5445,N_5422);
nand U6226 (N_6226,N_5495,N_5803);
and U6227 (N_6227,N_5531,N_5561);
or U6228 (N_6228,N_5856,N_5423);
and U6229 (N_6229,N_5117,N_5529);
or U6230 (N_6230,N_5540,N_5603);
nor U6231 (N_6231,N_5191,N_5795);
and U6232 (N_6232,N_5634,N_5129);
nand U6233 (N_6233,N_5697,N_5360);
xnor U6234 (N_6234,N_5933,N_5210);
or U6235 (N_6235,N_5287,N_5783);
xor U6236 (N_6236,N_5891,N_5854);
or U6237 (N_6237,N_5442,N_5875);
nor U6238 (N_6238,N_5234,N_5686);
and U6239 (N_6239,N_5511,N_5901);
nand U6240 (N_6240,N_5286,N_5730);
nor U6241 (N_6241,N_5988,N_5660);
or U6242 (N_6242,N_5656,N_5753);
nand U6243 (N_6243,N_5952,N_5229);
and U6244 (N_6244,N_5813,N_5093);
xor U6245 (N_6245,N_5440,N_5767);
or U6246 (N_6246,N_5131,N_5257);
nand U6247 (N_6247,N_5748,N_5709);
or U6248 (N_6248,N_5877,N_5858);
nand U6249 (N_6249,N_5755,N_5665);
or U6250 (N_6250,N_5000,N_5239);
and U6251 (N_6251,N_5100,N_5199);
nor U6252 (N_6252,N_5806,N_5727);
nor U6253 (N_6253,N_5313,N_5543);
nand U6254 (N_6254,N_5177,N_5482);
nor U6255 (N_6255,N_5987,N_5108);
or U6256 (N_6256,N_5724,N_5990);
or U6257 (N_6257,N_5853,N_5371);
xor U6258 (N_6258,N_5639,N_5308);
xor U6259 (N_6259,N_5467,N_5477);
nand U6260 (N_6260,N_5790,N_5535);
nor U6261 (N_6261,N_5115,N_5184);
or U6262 (N_6262,N_5307,N_5884);
and U6263 (N_6263,N_5700,N_5352);
or U6264 (N_6264,N_5237,N_5006);
and U6265 (N_6265,N_5722,N_5521);
and U6266 (N_6266,N_5978,N_5451);
nand U6267 (N_6267,N_5798,N_5784);
and U6268 (N_6268,N_5406,N_5836);
or U6269 (N_6269,N_5130,N_5463);
and U6270 (N_6270,N_5020,N_5666);
xnor U6271 (N_6271,N_5429,N_5749);
nor U6272 (N_6272,N_5606,N_5299);
and U6273 (N_6273,N_5835,N_5240);
or U6274 (N_6274,N_5250,N_5972);
and U6275 (N_6275,N_5164,N_5652);
or U6276 (N_6276,N_5642,N_5882);
xor U6277 (N_6277,N_5801,N_5397);
nor U6278 (N_6278,N_5903,N_5881);
and U6279 (N_6279,N_5852,N_5820);
nor U6280 (N_6280,N_5207,N_5602);
nor U6281 (N_6281,N_5301,N_5066);
xor U6282 (N_6282,N_5011,N_5520);
nor U6283 (N_6283,N_5689,N_5954);
and U6284 (N_6284,N_5275,N_5839);
nand U6285 (N_6285,N_5512,N_5439);
nand U6286 (N_6286,N_5484,N_5157);
or U6287 (N_6287,N_5819,N_5364);
or U6288 (N_6288,N_5174,N_5807);
and U6289 (N_6289,N_5815,N_5981);
and U6290 (N_6290,N_5241,N_5909);
and U6291 (N_6291,N_5072,N_5296);
nand U6292 (N_6292,N_5116,N_5796);
nand U6293 (N_6293,N_5057,N_5168);
and U6294 (N_6294,N_5071,N_5102);
nor U6295 (N_6295,N_5673,N_5323);
or U6296 (N_6296,N_5723,N_5146);
xnor U6297 (N_6297,N_5554,N_5890);
or U6298 (N_6298,N_5133,N_5556);
nand U6299 (N_6299,N_5306,N_5893);
or U6300 (N_6300,N_5113,N_5754);
nor U6301 (N_6301,N_5078,N_5408);
and U6302 (N_6302,N_5786,N_5792);
nor U6303 (N_6303,N_5175,N_5826);
nor U6304 (N_6304,N_5635,N_5432);
and U6305 (N_6305,N_5594,N_5414);
nor U6306 (N_6306,N_5282,N_5154);
nor U6307 (N_6307,N_5003,N_5441);
or U6308 (N_6308,N_5742,N_5967);
or U6309 (N_6309,N_5224,N_5805);
or U6310 (N_6310,N_5469,N_5690);
and U6311 (N_6311,N_5123,N_5403);
nor U6312 (N_6312,N_5101,N_5762);
nor U6313 (N_6313,N_5061,N_5911);
and U6314 (N_6314,N_5244,N_5195);
nor U6315 (N_6315,N_5405,N_5338);
nor U6316 (N_6316,N_5327,N_5617);
nor U6317 (N_6317,N_5738,N_5238);
and U6318 (N_6318,N_5205,N_5596);
or U6319 (N_6319,N_5356,N_5614);
nand U6320 (N_6320,N_5486,N_5514);
nand U6321 (N_6321,N_5084,N_5864);
nand U6322 (N_6322,N_5389,N_5668);
nor U6323 (N_6323,N_5650,N_5646);
nand U6324 (N_6324,N_5024,N_5153);
xnor U6325 (N_6325,N_5021,N_5677);
nand U6326 (N_6326,N_5448,N_5476);
and U6327 (N_6327,N_5038,N_5555);
and U6328 (N_6328,N_5491,N_5745);
nand U6329 (N_6329,N_5708,N_5470);
xnor U6330 (N_6330,N_5846,N_5923);
and U6331 (N_6331,N_5390,N_5588);
and U6332 (N_6332,N_5474,N_5140);
or U6333 (N_6333,N_5459,N_5924);
nor U6334 (N_6334,N_5373,N_5546);
or U6335 (N_6335,N_5086,N_5434);
nor U6336 (N_6336,N_5870,N_5333);
nand U6337 (N_6337,N_5266,N_5278);
xor U6338 (N_6338,N_5572,N_5253);
or U6339 (N_6339,N_5763,N_5354);
and U6340 (N_6340,N_5273,N_5178);
and U6341 (N_6341,N_5849,N_5468);
or U6342 (N_6342,N_5713,N_5380);
and U6343 (N_6343,N_5449,N_5430);
xnor U6344 (N_6344,N_5627,N_5012);
nor U6345 (N_6345,N_5612,N_5089);
or U6346 (N_6346,N_5245,N_5418);
nor U6347 (N_6347,N_5930,N_5173);
or U6348 (N_6348,N_5201,N_5684);
and U6349 (N_6349,N_5465,N_5109);
nor U6350 (N_6350,N_5747,N_5064);
and U6351 (N_6351,N_5183,N_5383);
nor U6352 (N_6352,N_5913,N_5961);
xnor U6353 (N_6353,N_5509,N_5294);
nand U6354 (N_6354,N_5568,N_5775);
nand U6355 (N_6355,N_5297,N_5382);
and U6356 (N_6356,N_5993,N_5518);
nand U6357 (N_6357,N_5992,N_5158);
nor U6358 (N_6358,N_5525,N_5122);
nand U6359 (N_6359,N_5050,N_5539);
and U6360 (N_6360,N_5216,N_5065);
nor U6361 (N_6361,N_5425,N_5219);
xnor U6362 (N_6362,N_5471,N_5575);
and U6363 (N_6363,N_5087,N_5134);
or U6364 (N_6364,N_5305,N_5103);
xor U6365 (N_6365,N_5674,N_5446);
xnor U6366 (N_6366,N_5886,N_5127);
xor U6367 (N_6367,N_5194,N_5472);
nand U6368 (N_6368,N_5149,N_5728);
or U6369 (N_6369,N_5977,N_5091);
and U6370 (N_6370,N_5785,N_5960);
xor U6371 (N_6371,N_5456,N_5868);
and U6372 (N_6372,N_5840,N_5553);
and U6373 (N_6373,N_5533,N_5619);
nor U6374 (N_6374,N_5182,N_5283);
and U6375 (N_6375,N_5316,N_5788);
nor U6376 (N_6376,N_5899,N_5683);
and U6377 (N_6377,N_5589,N_5593);
nand U6378 (N_6378,N_5031,N_5914);
nand U6379 (N_6379,N_5637,N_5959);
and U6380 (N_6380,N_5419,N_5809);
nand U6381 (N_6381,N_5337,N_5610);
xnor U6382 (N_6382,N_5309,N_5317);
nand U6383 (N_6383,N_5107,N_5632);
or U6384 (N_6384,N_5082,N_5779);
and U6385 (N_6385,N_5436,N_5198);
or U6386 (N_6386,N_5289,N_5985);
nor U6387 (N_6387,N_5111,N_5223);
nor U6388 (N_6388,N_5312,N_5699);
nor U6389 (N_6389,N_5995,N_5179);
nand U6390 (N_6390,N_5925,N_5932);
nor U6391 (N_6391,N_5466,N_5325);
xnor U6392 (N_6392,N_5662,N_5225);
or U6393 (N_6393,N_5242,N_5261);
and U6394 (N_6394,N_5576,N_5942);
nand U6395 (N_6395,N_5979,N_5760);
nor U6396 (N_6396,N_5392,N_5810);
or U6397 (N_6397,N_5365,N_5249);
nand U6398 (N_6398,N_5615,N_5597);
and U6399 (N_6399,N_5618,N_5526);
nor U6400 (N_6400,N_5051,N_5025);
and U6401 (N_6401,N_5288,N_5654);
or U6402 (N_6402,N_5362,N_5936);
nor U6403 (N_6403,N_5139,N_5998);
and U6404 (N_6404,N_5957,N_5986);
or U6405 (N_6405,N_5374,N_5905);
nor U6406 (N_6406,N_5218,N_5997);
and U6407 (N_6407,N_5208,N_5912);
or U6408 (N_6408,N_5411,N_5417);
and U6409 (N_6409,N_5793,N_5246);
and U6410 (N_6410,N_5322,N_5160);
xor U6411 (N_6411,N_5685,N_5953);
nor U6412 (N_6412,N_5607,N_5598);
and U6413 (N_6413,N_5026,N_5505);
nand U6414 (N_6414,N_5502,N_5956);
nor U6415 (N_6415,N_5280,N_5872);
or U6416 (N_6416,N_5889,N_5681);
nand U6417 (N_6417,N_5176,N_5269);
nand U6418 (N_6418,N_5029,N_5132);
and U6419 (N_6419,N_5271,N_5017);
and U6420 (N_6420,N_5067,N_5731);
or U6421 (N_6421,N_5894,N_5487);
nor U6422 (N_6422,N_5258,N_5170);
nor U6423 (N_6423,N_5481,N_5496);
and U6424 (N_6424,N_5848,N_5648);
and U6425 (N_6425,N_5032,N_5035);
or U6426 (N_6426,N_5016,N_5494);
and U6427 (N_6427,N_5228,N_5898);
nand U6428 (N_6428,N_5180,N_5672);
nor U6429 (N_6429,N_5827,N_5659);
and U6430 (N_6430,N_5605,N_5044);
and U6431 (N_6431,N_5013,N_5591);
or U6432 (N_6432,N_5118,N_5500);
nand U6433 (N_6433,N_5138,N_5693);
nor U6434 (N_6434,N_5694,N_5104);
nor U6435 (N_6435,N_5989,N_5040);
or U6436 (N_6436,N_5385,N_5756);
xor U6437 (N_6437,N_5774,N_5475);
xnor U6438 (N_6438,N_5002,N_5584);
and U6439 (N_6439,N_5159,N_5823);
nor U6440 (N_6440,N_5150,N_5499);
nor U6441 (N_6441,N_5075,N_5381);
or U6442 (N_6442,N_5600,N_5915);
or U6443 (N_6443,N_5701,N_5935);
or U6444 (N_6444,N_5480,N_5388);
and U6445 (N_6445,N_5437,N_5980);
or U6446 (N_6446,N_5616,N_5948);
nand U6447 (N_6447,N_5369,N_5259);
nand U6448 (N_6448,N_5705,N_5450);
and U6449 (N_6449,N_5719,N_5883);
or U6450 (N_6450,N_5857,N_5211);
nor U6451 (N_6451,N_5702,N_5106);
or U6452 (N_6452,N_5640,N_5592);
or U6453 (N_6453,N_5493,N_5268);
xnor U6454 (N_6454,N_5007,N_5653);
or U6455 (N_6455,N_5625,N_5036);
nor U6456 (N_6456,N_5196,N_5962);
or U6457 (N_6457,N_5523,N_5503);
xor U6458 (N_6458,N_5424,N_5947);
and U6459 (N_6459,N_5161,N_5517);
or U6460 (N_6460,N_5515,N_5121);
nand U6461 (N_6461,N_5010,N_5601);
nand U6462 (N_6462,N_5355,N_5214);
nor U6463 (N_6463,N_5938,N_5227);
or U6464 (N_6464,N_5062,N_5532);
nor U6465 (N_6465,N_5192,N_5206);
nand U6466 (N_6466,N_5847,N_5508);
nand U6467 (N_6467,N_5431,N_5996);
nand U6468 (N_6468,N_5944,N_5778);
and U6469 (N_6469,N_5908,N_5704);
and U6470 (N_6470,N_5968,N_5395);
and U6471 (N_6471,N_5671,N_5265);
nor U6472 (N_6472,N_5622,N_5136);
nand U6473 (N_6473,N_5248,N_5401);
and U6474 (N_6474,N_5971,N_5787);
and U6475 (N_6475,N_5843,N_5636);
xor U6476 (N_6476,N_5776,N_5285);
nand U6477 (N_6477,N_5740,N_5232);
or U6478 (N_6478,N_5137,N_5492);
xor U6479 (N_6479,N_5804,N_5099);
and U6480 (N_6480,N_5711,N_5045);
nor U6481 (N_6481,N_5570,N_5629);
xor U6482 (N_6482,N_5951,N_5766);
or U6483 (N_6483,N_5142,N_5641);
nand U6484 (N_6484,N_5504,N_5720);
xnor U6485 (N_6485,N_5845,N_5717);
nor U6486 (N_6486,N_5112,N_5579);
nand U6487 (N_6487,N_5386,N_5251);
nor U6488 (N_6488,N_5560,N_5821);
nand U6489 (N_6489,N_5053,N_5768);
or U6490 (N_6490,N_5254,N_5298);
nand U6491 (N_6491,N_5284,N_5991);
nand U6492 (N_6492,N_5243,N_5735);
nor U6493 (N_6493,N_5765,N_5303);
or U6494 (N_6494,N_5552,N_5426);
or U6495 (N_6495,N_5802,N_5657);
nor U6496 (N_6496,N_5452,N_5624);
nand U6497 (N_6497,N_5033,N_5097);
nand U6498 (N_6498,N_5407,N_5725);
nand U6499 (N_6499,N_5736,N_5583);
or U6500 (N_6500,N_5156,N_5022);
nor U6501 (N_6501,N_5455,N_5338);
nand U6502 (N_6502,N_5042,N_5775);
or U6503 (N_6503,N_5237,N_5309);
xor U6504 (N_6504,N_5158,N_5369);
and U6505 (N_6505,N_5865,N_5671);
or U6506 (N_6506,N_5430,N_5251);
nand U6507 (N_6507,N_5083,N_5526);
or U6508 (N_6508,N_5682,N_5241);
or U6509 (N_6509,N_5731,N_5706);
nor U6510 (N_6510,N_5092,N_5176);
or U6511 (N_6511,N_5564,N_5891);
or U6512 (N_6512,N_5278,N_5946);
xnor U6513 (N_6513,N_5576,N_5678);
nor U6514 (N_6514,N_5823,N_5683);
or U6515 (N_6515,N_5535,N_5528);
xor U6516 (N_6516,N_5234,N_5510);
nor U6517 (N_6517,N_5050,N_5071);
or U6518 (N_6518,N_5198,N_5633);
and U6519 (N_6519,N_5018,N_5594);
xor U6520 (N_6520,N_5735,N_5410);
nand U6521 (N_6521,N_5186,N_5985);
and U6522 (N_6522,N_5944,N_5663);
or U6523 (N_6523,N_5899,N_5527);
xnor U6524 (N_6524,N_5614,N_5424);
and U6525 (N_6525,N_5702,N_5745);
xnor U6526 (N_6526,N_5388,N_5395);
or U6527 (N_6527,N_5648,N_5200);
or U6528 (N_6528,N_5693,N_5682);
nand U6529 (N_6529,N_5221,N_5283);
nand U6530 (N_6530,N_5607,N_5704);
nand U6531 (N_6531,N_5604,N_5383);
and U6532 (N_6532,N_5525,N_5386);
xor U6533 (N_6533,N_5001,N_5944);
or U6534 (N_6534,N_5948,N_5504);
or U6535 (N_6535,N_5896,N_5399);
nand U6536 (N_6536,N_5945,N_5783);
or U6537 (N_6537,N_5723,N_5498);
and U6538 (N_6538,N_5798,N_5484);
nor U6539 (N_6539,N_5969,N_5725);
and U6540 (N_6540,N_5452,N_5081);
and U6541 (N_6541,N_5140,N_5917);
nand U6542 (N_6542,N_5600,N_5254);
nand U6543 (N_6543,N_5540,N_5846);
nor U6544 (N_6544,N_5837,N_5151);
xor U6545 (N_6545,N_5755,N_5661);
xnor U6546 (N_6546,N_5109,N_5686);
and U6547 (N_6547,N_5296,N_5938);
and U6548 (N_6548,N_5774,N_5198);
nor U6549 (N_6549,N_5101,N_5611);
nor U6550 (N_6550,N_5490,N_5155);
or U6551 (N_6551,N_5036,N_5938);
nor U6552 (N_6552,N_5406,N_5027);
nand U6553 (N_6553,N_5550,N_5999);
xor U6554 (N_6554,N_5711,N_5666);
and U6555 (N_6555,N_5480,N_5770);
nand U6556 (N_6556,N_5863,N_5702);
nand U6557 (N_6557,N_5658,N_5845);
and U6558 (N_6558,N_5656,N_5820);
or U6559 (N_6559,N_5512,N_5558);
or U6560 (N_6560,N_5216,N_5369);
and U6561 (N_6561,N_5670,N_5259);
and U6562 (N_6562,N_5863,N_5506);
nor U6563 (N_6563,N_5310,N_5887);
nor U6564 (N_6564,N_5248,N_5619);
and U6565 (N_6565,N_5626,N_5430);
nand U6566 (N_6566,N_5748,N_5631);
xor U6567 (N_6567,N_5786,N_5328);
or U6568 (N_6568,N_5339,N_5455);
xor U6569 (N_6569,N_5076,N_5439);
nand U6570 (N_6570,N_5325,N_5087);
or U6571 (N_6571,N_5083,N_5090);
or U6572 (N_6572,N_5242,N_5030);
and U6573 (N_6573,N_5915,N_5163);
xnor U6574 (N_6574,N_5194,N_5489);
nor U6575 (N_6575,N_5053,N_5029);
nor U6576 (N_6576,N_5529,N_5834);
and U6577 (N_6577,N_5136,N_5103);
and U6578 (N_6578,N_5933,N_5560);
nor U6579 (N_6579,N_5262,N_5829);
and U6580 (N_6580,N_5806,N_5595);
and U6581 (N_6581,N_5328,N_5527);
xnor U6582 (N_6582,N_5220,N_5512);
and U6583 (N_6583,N_5388,N_5700);
nand U6584 (N_6584,N_5590,N_5852);
nor U6585 (N_6585,N_5804,N_5154);
or U6586 (N_6586,N_5965,N_5986);
or U6587 (N_6587,N_5322,N_5540);
nor U6588 (N_6588,N_5651,N_5334);
and U6589 (N_6589,N_5971,N_5442);
and U6590 (N_6590,N_5886,N_5158);
xnor U6591 (N_6591,N_5005,N_5323);
nor U6592 (N_6592,N_5696,N_5546);
and U6593 (N_6593,N_5946,N_5315);
and U6594 (N_6594,N_5952,N_5764);
nor U6595 (N_6595,N_5218,N_5246);
nand U6596 (N_6596,N_5603,N_5279);
nand U6597 (N_6597,N_5146,N_5972);
nor U6598 (N_6598,N_5022,N_5474);
xnor U6599 (N_6599,N_5686,N_5175);
and U6600 (N_6600,N_5138,N_5603);
xor U6601 (N_6601,N_5512,N_5262);
or U6602 (N_6602,N_5313,N_5729);
nor U6603 (N_6603,N_5872,N_5941);
nand U6604 (N_6604,N_5901,N_5966);
nor U6605 (N_6605,N_5222,N_5510);
and U6606 (N_6606,N_5844,N_5020);
and U6607 (N_6607,N_5780,N_5834);
xor U6608 (N_6608,N_5872,N_5710);
nand U6609 (N_6609,N_5745,N_5342);
or U6610 (N_6610,N_5759,N_5713);
or U6611 (N_6611,N_5027,N_5595);
xor U6612 (N_6612,N_5992,N_5629);
and U6613 (N_6613,N_5752,N_5457);
nand U6614 (N_6614,N_5498,N_5158);
xor U6615 (N_6615,N_5434,N_5540);
and U6616 (N_6616,N_5905,N_5620);
nor U6617 (N_6617,N_5664,N_5927);
and U6618 (N_6618,N_5030,N_5623);
or U6619 (N_6619,N_5556,N_5760);
or U6620 (N_6620,N_5146,N_5806);
xor U6621 (N_6621,N_5745,N_5498);
and U6622 (N_6622,N_5475,N_5367);
nand U6623 (N_6623,N_5927,N_5338);
or U6624 (N_6624,N_5861,N_5166);
and U6625 (N_6625,N_5474,N_5183);
nor U6626 (N_6626,N_5100,N_5654);
xor U6627 (N_6627,N_5195,N_5752);
nor U6628 (N_6628,N_5326,N_5625);
and U6629 (N_6629,N_5990,N_5535);
nor U6630 (N_6630,N_5984,N_5374);
nor U6631 (N_6631,N_5353,N_5610);
nor U6632 (N_6632,N_5783,N_5993);
or U6633 (N_6633,N_5177,N_5287);
nand U6634 (N_6634,N_5417,N_5467);
and U6635 (N_6635,N_5758,N_5234);
nand U6636 (N_6636,N_5706,N_5976);
or U6637 (N_6637,N_5817,N_5869);
or U6638 (N_6638,N_5900,N_5783);
nand U6639 (N_6639,N_5531,N_5300);
and U6640 (N_6640,N_5186,N_5617);
and U6641 (N_6641,N_5714,N_5854);
and U6642 (N_6642,N_5978,N_5789);
nand U6643 (N_6643,N_5623,N_5826);
and U6644 (N_6644,N_5062,N_5734);
nor U6645 (N_6645,N_5203,N_5232);
and U6646 (N_6646,N_5448,N_5849);
or U6647 (N_6647,N_5670,N_5100);
nor U6648 (N_6648,N_5220,N_5086);
xnor U6649 (N_6649,N_5567,N_5441);
and U6650 (N_6650,N_5380,N_5403);
or U6651 (N_6651,N_5544,N_5126);
nand U6652 (N_6652,N_5628,N_5338);
nand U6653 (N_6653,N_5495,N_5044);
nand U6654 (N_6654,N_5639,N_5090);
nand U6655 (N_6655,N_5701,N_5478);
nand U6656 (N_6656,N_5770,N_5931);
and U6657 (N_6657,N_5669,N_5523);
and U6658 (N_6658,N_5497,N_5998);
or U6659 (N_6659,N_5757,N_5297);
and U6660 (N_6660,N_5107,N_5563);
and U6661 (N_6661,N_5140,N_5542);
and U6662 (N_6662,N_5458,N_5617);
xnor U6663 (N_6663,N_5969,N_5004);
and U6664 (N_6664,N_5453,N_5592);
nand U6665 (N_6665,N_5400,N_5678);
nand U6666 (N_6666,N_5655,N_5480);
nor U6667 (N_6667,N_5286,N_5399);
or U6668 (N_6668,N_5665,N_5133);
or U6669 (N_6669,N_5805,N_5685);
xor U6670 (N_6670,N_5759,N_5809);
or U6671 (N_6671,N_5050,N_5799);
nor U6672 (N_6672,N_5417,N_5531);
and U6673 (N_6673,N_5501,N_5921);
nand U6674 (N_6674,N_5050,N_5405);
or U6675 (N_6675,N_5306,N_5951);
and U6676 (N_6676,N_5478,N_5591);
nand U6677 (N_6677,N_5775,N_5328);
or U6678 (N_6678,N_5012,N_5180);
or U6679 (N_6679,N_5736,N_5331);
and U6680 (N_6680,N_5641,N_5435);
and U6681 (N_6681,N_5321,N_5361);
nand U6682 (N_6682,N_5119,N_5593);
nor U6683 (N_6683,N_5654,N_5949);
xnor U6684 (N_6684,N_5802,N_5255);
and U6685 (N_6685,N_5551,N_5640);
xnor U6686 (N_6686,N_5851,N_5432);
xnor U6687 (N_6687,N_5173,N_5609);
or U6688 (N_6688,N_5500,N_5738);
xor U6689 (N_6689,N_5847,N_5861);
xnor U6690 (N_6690,N_5684,N_5489);
and U6691 (N_6691,N_5347,N_5005);
and U6692 (N_6692,N_5114,N_5475);
nor U6693 (N_6693,N_5647,N_5208);
or U6694 (N_6694,N_5135,N_5456);
nor U6695 (N_6695,N_5449,N_5903);
and U6696 (N_6696,N_5117,N_5581);
or U6697 (N_6697,N_5321,N_5916);
or U6698 (N_6698,N_5094,N_5140);
or U6699 (N_6699,N_5063,N_5143);
nor U6700 (N_6700,N_5943,N_5539);
nor U6701 (N_6701,N_5988,N_5167);
nand U6702 (N_6702,N_5529,N_5898);
and U6703 (N_6703,N_5961,N_5601);
and U6704 (N_6704,N_5999,N_5852);
nor U6705 (N_6705,N_5508,N_5515);
or U6706 (N_6706,N_5804,N_5062);
nor U6707 (N_6707,N_5092,N_5241);
and U6708 (N_6708,N_5759,N_5130);
nor U6709 (N_6709,N_5918,N_5233);
or U6710 (N_6710,N_5118,N_5613);
and U6711 (N_6711,N_5026,N_5854);
and U6712 (N_6712,N_5430,N_5391);
nand U6713 (N_6713,N_5313,N_5066);
nand U6714 (N_6714,N_5993,N_5885);
and U6715 (N_6715,N_5455,N_5813);
or U6716 (N_6716,N_5819,N_5334);
and U6717 (N_6717,N_5232,N_5165);
or U6718 (N_6718,N_5537,N_5032);
nand U6719 (N_6719,N_5620,N_5301);
nor U6720 (N_6720,N_5426,N_5960);
xnor U6721 (N_6721,N_5971,N_5906);
and U6722 (N_6722,N_5427,N_5319);
nand U6723 (N_6723,N_5345,N_5997);
nand U6724 (N_6724,N_5403,N_5447);
and U6725 (N_6725,N_5963,N_5112);
nor U6726 (N_6726,N_5927,N_5911);
and U6727 (N_6727,N_5033,N_5406);
nor U6728 (N_6728,N_5006,N_5208);
nor U6729 (N_6729,N_5772,N_5227);
or U6730 (N_6730,N_5716,N_5467);
nand U6731 (N_6731,N_5202,N_5731);
nand U6732 (N_6732,N_5122,N_5055);
and U6733 (N_6733,N_5919,N_5648);
or U6734 (N_6734,N_5719,N_5670);
and U6735 (N_6735,N_5957,N_5549);
xor U6736 (N_6736,N_5266,N_5876);
and U6737 (N_6737,N_5988,N_5342);
or U6738 (N_6738,N_5054,N_5052);
nor U6739 (N_6739,N_5395,N_5203);
xor U6740 (N_6740,N_5639,N_5364);
nor U6741 (N_6741,N_5572,N_5922);
nand U6742 (N_6742,N_5753,N_5063);
xnor U6743 (N_6743,N_5686,N_5618);
or U6744 (N_6744,N_5493,N_5460);
nand U6745 (N_6745,N_5245,N_5849);
and U6746 (N_6746,N_5249,N_5265);
and U6747 (N_6747,N_5989,N_5517);
and U6748 (N_6748,N_5019,N_5075);
nor U6749 (N_6749,N_5196,N_5605);
nor U6750 (N_6750,N_5334,N_5813);
xor U6751 (N_6751,N_5755,N_5587);
nor U6752 (N_6752,N_5301,N_5201);
or U6753 (N_6753,N_5141,N_5726);
or U6754 (N_6754,N_5824,N_5004);
nand U6755 (N_6755,N_5943,N_5626);
nor U6756 (N_6756,N_5677,N_5658);
xnor U6757 (N_6757,N_5473,N_5018);
xnor U6758 (N_6758,N_5038,N_5676);
nand U6759 (N_6759,N_5016,N_5249);
nand U6760 (N_6760,N_5274,N_5648);
or U6761 (N_6761,N_5853,N_5765);
or U6762 (N_6762,N_5192,N_5655);
xnor U6763 (N_6763,N_5409,N_5006);
or U6764 (N_6764,N_5116,N_5032);
nor U6765 (N_6765,N_5216,N_5965);
nor U6766 (N_6766,N_5208,N_5031);
nor U6767 (N_6767,N_5115,N_5204);
nand U6768 (N_6768,N_5032,N_5726);
and U6769 (N_6769,N_5768,N_5313);
or U6770 (N_6770,N_5533,N_5089);
or U6771 (N_6771,N_5253,N_5636);
nor U6772 (N_6772,N_5775,N_5486);
or U6773 (N_6773,N_5699,N_5756);
or U6774 (N_6774,N_5383,N_5250);
or U6775 (N_6775,N_5765,N_5496);
and U6776 (N_6776,N_5874,N_5848);
nor U6777 (N_6777,N_5828,N_5644);
and U6778 (N_6778,N_5341,N_5980);
nand U6779 (N_6779,N_5737,N_5193);
or U6780 (N_6780,N_5168,N_5756);
or U6781 (N_6781,N_5345,N_5599);
and U6782 (N_6782,N_5484,N_5458);
or U6783 (N_6783,N_5297,N_5210);
nand U6784 (N_6784,N_5007,N_5477);
and U6785 (N_6785,N_5693,N_5626);
and U6786 (N_6786,N_5489,N_5539);
and U6787 (N_6787,N_5806,N_5162);
or U6788 (N_6788,N_5580,N_5022);
or U6789 (N_6789,N_5715,N_5157);
and U6790 (N_6790,N_5764,N_5289);
xor U6791 (N_6791,N_5199,N_5670);
and U6792 (N_6792,N_5449,N_5830);
or U6793 (N_6793,N_5934,N_5813);
xor U6794 (N_6794,N_5995,N_5402);
nand U6795 (N_6795,N_5074,N_5743);
and U6796 (N_6796,N_5124,N_5347);
xnor U6797 (N_6797,N_5429,N_5416);
nor U6798 (N_6798,N_5626,N_5802);
nor U6799 (N_6799,N_5338,N_5216);
nor U6800 (N_6800,N_5673,N_5728);
or U6801 (N_6801,N_5125,N_5739);
and U6802 (N_6802,N_5173,N_5302);
nand U6803 (N_6803,N_5480,N_5571);
nand U6804 (N_6804,N_5368,N_5195);
or U6805 (N_6805,N_5725,N_5192);
or U6806 (N_6806,N_5625,N_5680);
nor U6807 (N_6807,N_5427,N_5945);
or U6808 (N_6808,N_5088,N_5917);
nor U6809 (N_6809,N_5474,N_5687);
nor U6810 (N_6810,N_5018,N_5002);
nor U6811 (N_6811,N_5008,N_5731);
nand U6812 (N_6812,N_5920,N_5410);
nor U6813 (N_6813,N_5121,N_5451);
or U6814 (N_6814,N_5417,N_5199);
nand U6815 (N_6815,N_5816,N_5234);
or U6816 (N_6816,N_5674,N_5192);
xnor U6817 (N_6817,N_5343,N_5011);
xnor U6818 (N_6818,N_5002,N_5554);
or U6819 (N_6819,N_5054,N_5500);
nand U6820 (N_6820,N_5058,N_5059);
xor U6821 (N_6821,N_5581,N_5325);
and U6822 (N_6822,N_5398,N_5166);
nand U6823 (N_6823,N_5361,N_5856);
nand U6824 (N_6824,N_5947,N_5721);
nor U6825 (N_6825,N_5341,N_5097);
xnor U6826 (N_6826,N_5903,N_5357);
nor U6827 (N_6827,N_5429,N_5098);
or U6828 (N_6828,N_5519,N_5922);
nor U6829 (N_6829,N_5629,N_5316);
nand U6830 (N_6830,N_5197,N_5463);
and U6831 (N_6831,N_5344,N_5063);
nand U6832 (N_6832,N_5382,N_5741);
or U6833 (N_6833,N_5338,N_5783);
and U6834 (N_6834,N_5195,N_5973);
nand U6835 (N_6835,N_5340,N_5065);
nor U6836 (N_6836,N_5227,N_5671);
xor U6837 (N_6837,N_5874,N_5151);
and U6838 (N_6838,N_5541,N_5994);
nand U6839 (N_6839,N_5427,N_5454);
nand U6840 (N_6840,N_5267,N_5020);
or U6841 (N_6841,N_5036,N_5973);
nand U6842 (N_6842,N_5238,N_5446);
xor U6843 (N_6843,N_5024,N_5398);
or U6844 (N_6844,N_5604,N_5025);
nor U6845 (N_6845,N_5170,N_5156);
nor U6846 (N_6846,N_5832,N_5997);
or U6847 (N_6847,N_5283,N_5588);
nor U6848 (N_6848,N_5168,N_5242);
nand U6849 (N_6849,N_5532,N_5257);
nand U6850 (N_6850,N_5801,N_5348);
xnor U6851 (N_6851,N_5092,N_5037);
nor U6852 (N_6852,N_5941,N_5437);
and U6853 (N_6853,N_5791,N_5859);
nor U6854 (N_6854,N_5248,N_5316);
or U6855 (N_6855,N_5456,N_5719);
nand U6856 (N_6856,N_5917,N_5703);
nor U6857 (N_6857,N_5074,N_5036);
nand U6858 (N_6858,N_5215,N_5234);
nand U6859 (N_6859,N_5403,N_5998);
or U6860 (N_6860,N_5718,N_5032);
nor U6861 (N_6861,N_5562,N_5843);
nor U6862 (N_6862,N_5801,N_5970);
nand U6863 (N_6863,N_5849,N_5474);
and U6864 (N_6864,N_5885,N_5117);
nand U6865 (N_6865,N_5929,N_5286);
or U6866 (N_6866,N_5569,N_5677);
or U6867 (N_6867,N_5809,N_5194);
or U6868 (N_6868,N_5389,N_5340);
and U6869 (N_6869,N_5144,N_5519);
nand U6870 (N_6870,N_5520,N_5223);
nor U6871 (N_6871,N_5339,N_5874);
nor U6872 (N_6872,N_5404,N_5825);
nor U6873 (N_6873,N_5939,N_5634);
nand U6874 (N_6874,N_5095,N_5800);
nand U6875 (N_6875,N_5896,N_5497);
or U6876 (N_6876,N_5259,N_5188);
nand U6877 (N_6877,N_5658,N_5965);
or U6878 (N_6878,N_5384,N_5568);
nor U6879 (N_6879,N_5827,N_5315);
and U6880 (N_6880,N_5156,N_5448);
or U6881 (N_6881,N_5564,N_5778);
or U6882 (N_6882,N_5747,N_5957);
nor U6883 (N_6883,N_5044,N_5358);
nor U6884 (N_6884,N_5701,N_5623);
nor U6885 (N_6885,N_5231,N_5122);
and U6886 (N_6886,N_5089,N_5842);
nor U6887 (N_6887,N_5159,N_5384);
nor U6888 (N_6888,N_5800,N_5059);
and U6889 (N_6889,N_5683,N_5618);
and U6890 (N_6890,N_5945,N_5512);
and U6891 (N_6891,N_5321,N_5211);
or U6892 (N_6892,N_5390,N_5365);
and U6893 (N_6893,N_5213,N_5649);
or U6894 (N_6894,N_5146,N_5069);
and U6895 (N_6895,N_5932,N_5588);
or U6896 (N_6896,N_5523,N_5326);
xor U6897 (N_6897,N_5715,N_5942);
or U6898 (N_6898,N_5530,N_5600);
nand U6899 (N_6899,N_5035,N_5996);
and U6900 (N_6900,N_5318,N_5383);
xor U6901 (N_6901,N_5193,N_5903);
nor U6902 (N_6902,N_5254,N_5166);
nor U6903 (N_6903,N_5012,N_5239);
nor U6904 (N_6904,N_5986,N_5401);
or U6905 (N_6905,N_5050,N_5015);
and U6906 (N_6906,N_5310,N_5593);
xor U6907 (N_6907,N_5269,N_5079);
or U6908 (N_6908,N_5965,N_5706);
and U6909 (N_6909,N_5076,N_5632);
and U6910 (N_6910,N_5944,N_5814);
xor U6911 (N_6911,N_5577,N_5500);
nor U6912 (N_6912,N_5662,N_5549);
or U6913 (N_6913,N_5390,N_5663);
and U6914 (N_6914,N_5383,N_5004);
and U6915 (N_6915,N_5613,N_5943);
nor U6916 (N_6916,N_5071,N_5804);
nor U6917 (N_6917,N_5868,N_5955);
and U6918 (N_6918,N_5961,N_5904);
nand U6919 (N_6919,N_5124,N_5029);
or U6920 (N_6920,N_5520,N_5268);
and U6921 (N_6921,N_5946,N_5455);
nor U6922 (N_6922,N_5226,N_5300);
or U6923 (N_6923,N_5283,N_5236);
nor U6924 (N_6924,N_5632,N_5021);
nor U6925 (N_6925,N_5906,N_5316);
and U6926 (N_6926,N_5519,N_5341);
or U6927 (N_6927,N_5419,N_5269);
xor U6928 (N_6928,N_5383,N_5815);
or U6929 (N_6929,N_5727,N_5523);
nor U6930 (N_6930,N_5849,N_5370);
and U6931 (N_6931,N_5721,N_5426);
xnor U6932 (N_6932,N_5219,N_5814);
nand U6933 (N_6933,N_5741,N_5194);
and U6934 (N_6934,N_5334,N_5031);
and U6935 (N_6935,N_5189,N_5708);
nand U6936 (N_6936,N_5167,N_5056);
or U6937 (N_6937,N_5208,N_5750);
xor U6938 (N_6938,N_5929,N_5723);
nor U6939 (N_6939,N_5133,N_5908);
nand U6940 (N_6940,N_5902,N_5363);
xor U6941 (N_6941,N_5240,N_5445);
or U6942 (N_6942,N_5733,N_5476);
nand U6943 (N_6943,N_5587,N_5969);
and U6944 (N_6944,N_5781,N_5902);
xnor U6945 (N_6945,N_5699,N_5177);
nand U6946 (N_6946,N_5895,N_5076);
xor U6947 (N_6947,N_5190,N_5060);
nor U6948 (N_6948,N_5240,N_5776);
nor U6949 (N_6949,N_5932,N_5229);
or U6950 (N_6950,N_5724,N_5344);
nand U6951 (N_6951,N_5853,N_5578);
nor U6952 (N_6952,N_5665,N_5864);
nand U6953 (N_6953,N_5589,N_5565);
or U6954 (N_6954,N_5349,N_5865);
nand U6955 (N_6955,N_5224,N_5842);
xnor U6956 (N_6956,N_5716,N_5299);
nand U6957 (N_6957,N_5331,N_5348);
xor U6958 (N_6958,N_5212,N_5538);
or U6959 (N_6959,N_5285,N_5792);
or U6960 (N_6960,N_5654,N_5270);
nand U6961 (N_6961,N_5389,N_5810);
or U6962 (N_6962,N_5845,N_5619);
or U6963 (N_6963,N_5575,N_5754);
and U6964 (N_6964,N_5485,N_5090);
nand U6965 (N_6965,N_5255,N_5240);
xor U6966 (N_6966,N_5447,N_5282);
xnor U6967 (N_6967,N_5544,N_5109);
nor U6968 (N_6968,N_5181,N_5058);
and U6969 (N_6969,N_5257,N_5756);
or U6970 (N_6970,N_5256,N_5202);
xnor U6971 (N_6971,N_5713,N_5684);
or U6972 (N_6972,N_5347,N_5959);
or U6973 (N_6973,N_5756,N_5595);
xor U6974 (N_6974,N_5776,N_5712);
and U6975 (N_6975,N_5703,N_5837);
nand U6976 (N_6976,N_5164,N_5903);
or U6977 (N_6977,N_5358,N_5204);
and U6978 (N_6978,N_5709,N_5658);
and U6979 (N_6979,N_5875,N_5053);
nor U6980 (N_6980,N_5648,N_5325);
nor U6981 (N_6981,N_5349,N_5772);
or U6982 (N_6982,N_5880,N_5186);
nand U6983 (N_6983,N_5482,N_5234);
nand U6984 (N_6984,N_5969,N_5449);
xor U6985 (N_6985,N_5974,N_5706);
xor U6986 (N_6986,N_5593,N_5427);
nand U6987 (N_6987,N_5893,N_5796);
nand U6988 (N_6988,N_5420,N_5164);
nand U6989 (N_6989,N_5056,N_5233);
and U6990 (N_6990,N_5487,N_5137);
nor U6991 (N_6991,N_5841,N_5466);
or U6992 (N_6992,N_5039,N_5395);
and U6993 (N_6993,N_5427,N_5610);
nor U6994 (N_6994,N_5447,N_5648);
and U6995 (N_6995,N_5982,N_5123);
nor U6996 (N_6996,N_5417,N_5534);
and U6997 (N_6997,N_5168,N_5740);
or U6998 (N_6998,N_5288,N_5186);
xor U6999 (N_6999,N_5867,N_5173);
nand U7000 (N_7000,N_6079,N_6644);
and U7001 (N_7001,N_6062,N_6169);
nor U7002 (N_7002,N_6792,N_6496);
xnor U7003 (N_7003,N_6696,N_6107);
nand U7004 (N_7004,N_6879,N_6040);
and U7005 (N_7005,N_6574,N_6605);
and U7006 (N_7006,N_6474,N_6695);
or U7007 (N_7007,N_6916,N_6177);
and U7008 (N_7008,N_6816,N_6170);
nor U7009 (N_7009,N_6687,N_6338);
xnor U7010 (N_7010,N_6835,N_6093);
nand U7011 (N_7011,N_6602,N_6502);
or U7012 (N_7012,N_6274,N_6821);
nor U7013 (N_7013,N_6822,N_6128);
and U7014 (N_7014,N_6343,N_6701);
or U7015 (N_7015,N_6830,N_6264);
nor U7016 (N_7016,N_6453,N_6796);
nand U7017 (N_7017,N_6889,N_6568);
nand U7018 (N_7018,N_6771,N_6967);
nor U7019 (N_7019,N_6087,N_6313);
and U7020 (N_7020,N_6371,N_6194);
nor U7021 (N_7021,N_6447,N_6206);
nand U7022 (N_7022,N_6965,N_6509);
or U7023 (N_7023,N_6524,N_6640);
or U7024 (N_7024,N_6323,N_6305);
and U7025 (N_7025,N_6270,N_6489);
xor U7026 (N_7026,N_6384,N_6347);
and U7027 (N_7027,N_6849,N_6482);
and U7028 (N_7028,N_6829,N_6892);
nor U7029 (N_7029,N_6272,N_6478);
or U7030 (N_7030,N_6787,N_6232);
or U7031 (N_7031,N_6205,N_6240);
nand U7032 (N_7032,N_6633,N_6464);
or U7033 (N_7033,N_6863,N_6077);
nand U7034 (N_7034,N_6656,N_6690);
or U7035 (N_7035,N_6257,N_6675);
and U7036 (N_7036,N_6426,N_6480);
nand U7037 (N_7037,N_6679,N_6424);
and U7038 (N_7038,N_6488,N_6880);
nand U7039 (N_7039,N_6363,N_6623);
nand U7040 (N_7040,N_6642,N_6777);
nand U7041 (N_7041,N_6058,N_6824);
or U7042 (N_7042,N_6418,N_6613);
or U7043 (N_7043,N_6462,N_6708);
nor U7044 (N_7044,N_6068,N_6537);
or U7045 (N_7045,N_6033,N_6684);
nand U7046 (N_7046,N_6969,N_6666);
xnor U7047 (N_7047,N_6491,N_6584);
nor U7048 (N_7048,N_6731,N_6794);
or U7049 (N_7049,N_6331,N_6097);
or U7050 (N_7050,N_6667,N_6922);
nor U7051 (N_7051,N_6229,N_6858);
nand U7052 (N_7052,N_6985,N_6799);
xnor U7053 (N_7053,N_6050,N_6555);
and U7054 (N_7054,N_6452,N_6939);
and U7055 (N_7055,N_6336,N_6645);
xor U7056 (N_7056,N_6844,N_6903);
or U7057 (N_7057,N_6944,N_6127);
and U7058 (N_7058,N_6597,N_6108);
and U7059 (N_7059,N_6410,N_6357);
nand U7060 (N_7060,N_6089,N_6990);
and U7061 (N_7061,N_6560,N_6899);
or U7062 (N_7062,N_6102,N_6070);
nand U7063 (N_7063,N_6484,N_6303);
nor U7064 (N_7064,N_6664,N_6519);
nand U7065 (N_7065,N_6398,N_6373);
nand U7066 (N_7066,N_6795,N_6700);
nor U7067 (N_7067,N_6628,N_6974);
nor U7068 (N_7068,N_6578,N_6199);
and U7069 (N_7069,N_6278,N_6571);
nand U7070 (N_7070,N_6736,N_6273);
xnor U7071 (N_7071,N_6988,N_6707);
and U7072 (N_7072,N_6119,N_6222);
nand U7073 (N_7073,N_6387,N_6327);
and U7074 (N_7074,N_6254,N_6359);
or U7075 (N_7075,N_6786,N_6505);
and U7076 (N_7076,N_6122,N_6607);
xor U7077 (N_7077,N_6504,N_6562);
nor U7078 (N_7078,N_6643,N_6814);
nand U7079 (N_7079,N_6325,N_6860);
or U7080 (N_7080,N_6782,N_6789);
nand U7081 (N_7081,N_6724,N_6296);
nand U7082 (N_7082,N_6351,N_6167);
or U7083 (N_7083,N_6685,N_6023);
nor U7084 (N_7084,N_6246,N_6266);
nor U7085 (N_7085,N_6900,N_6295);
or U7086 (N_7086,N_6015,N_6412);
or U7087 (N_7087,N_6815,N_6963);
nand U7088 (N_7088,N_6495,N_6737);
and U7089 (N_7089,N_6702,N_6051);
nand U7090 (N_7090,N_6111,N_6012);
or U7091 (N_7091,N_6928,N_6590);
and U7092 (N_7092,N_6554,N_6465);
xnor U7093 (N_7093,N_6201,N_6671);
nand U7094 (N_7094,N_6970,N_6804);
xnor U7095 (N_7095,N_6636,N_6181);
nor U7096 (N_7096,N_6791,N_6923);
xnor U7097 (N_7097,N_6297,N_6376);
and U7098 (N_7098,N_6759,N_6365);
and U7099 (N_7099,N_6385,N_6676);
and U7100 (N_7100,N_6711,N_6224);
nor U7101 (N_7101,N_6971,N_6742);
xnor U7102 (N_7102,N_6219,N_6168);
and U7103 (N_7103,N_6510,N_6419);
nand U7104 (N_7104,N_6031,N_6896);
or U7105 (N_7105,N_6917,N_6277);
nand U7106 (N_7106,N_6751,N_6790);
and U7107 (N_7107,N_6958,N_6984);
nand U7108 (N_7108,N_6330,N_6120);
nand U7109 (N_7109,N_6216,N_6226);
nand U7110 (N_7110,N_6150,N_6755);
and U7111 (N_7111,N_6907,N_6801);
nand U7112 (N_7112,N_6714,N_6723);
and U7113 (N_7113,N_6692,N_6008);
xnor U7114 (N_7114,N_6542,N_6959);
nand U7115 (N_7115,N_6839,N_6318);
nor U7116 (N_7116,N_6573,N_6115);
or U7117 (N_7117,N_6601,N_6655);
and U7118 (N_7118,N_6680,N_6867);
nor U7119 (N_7119,N_6648,N_6874);
nor U7120 (N_7120,N_6556,N_6641);
nand U7121 (N_7121,N_6720,N_6469);
nor U7122 (N_7122,N_6457,N_6503);
nand U7123 (N_7123,N_6173,N_6533);
xnor U7124 (N_7124,N_6352,N_6856);
nor U7125 (N_7125,N_6481,N_6287);
nor U7126 (N_7126,N_6069,N_6951);
nand U7127 (N_7127,N_6187,N_6261);
nor U7128 (N_7128,N_6448,N_6218);
and U7129 (N_7129,N_6490,N_6629);
nand U7130 (N_7130,N_6995,N_6615);
nor U7131 (N_7131,N_6933,N_6250);
nor U7132 (N_7132,N_6299,N_6048);
nor U7133 (N_7133,N_6081,N_6611);
nand U7134 (N_7134,N_6779,N_6800);
or U7135 (N_7135,N_6483,N_6151);
and U7136 (N_7136,N_6603,N_6783);
nand U7137 (N_7137,N_6432,N_6761);
nor U7138 (N_7138,N_6258,N_6178);
nor U7139 (N_7139,N_6019,N_6911);
or U7140 (N_7140,N_6583,N_6831);
or U7141 (N_7141,N_6434,N_6414);
or U7142 (N_7142,N_6757,N_6072);
or U7143 (N_7143,N_6091,N_6339);
or U7144 (N_7144,N_6189,N_6227);
nand U7145 (N_7145,N_6064,N_6084);
nand U7146 (N_7146,N_6871,N_6565);
or U7147 (N_7147,N_6972,N_6683);
xnor U7148 (N_7148,N_6172,N_6857);
nand U7149 (N_7149,N_6054,N_6516);
or U7150 (N_7150,N_6765,N_6756);
nor U7151 (N_7151,N_6999,N_6047);
nor U7152 (N_7152,N_6739,N_6677);
xnor U7153 (N_7153,N_6924,N_6383);
or U7154 (N_7154,N_6421,N_6750);
nand U7155 (N_7155,N_6709,N_6989);
nand U7156 (N_7156,N_6842,N_6598);
nand U7157 (N_7157,N_6329,N_6520);
and U7158 (N_7158,N_6029,N_6214);
nand U7159 (N_7159,N_6293,N_6957);
or U7160 (N_7160,N_6785,N_6838);
nand U7161 (N_7161,N_6112,N_6852);
or U7162 (N_7162,N_6076,N_6877);
nand U7163 (N_7163,N_6302,N_6859);
nor U7164 (N_7164,N_6725,N_6698);
nor U7165 (N_7165,N_6500,N_6833);
nand U7166 (N_7166,N_6143,N_6596);
and U7167 (N_7167,N_6397,N_6847);
nand U7168 (N_7168,N_6909,N_6139);
or U7169 (N_7169,N_6651,N_6362);
or U7170 (N_7170,N_6234,N_6895);
or U7171 (N_7171,N_6620,N_6300);
or U7172 (N_7172,N_6522,N_6818);
or U7173 (N_7173,N_6841,N_6646);
or U7174 (N_7174,N_6773,N_6126);
xor U7175 (N_7175,N_6016,N_6380);
nand U7176 (N_7176,N_6007,N_6512);
and U7177 (N_7177,N_6514,N_6055);
nand U7178 (N_7178,N_6658,N_6441);
nand U7179 (N_7179,N_6389,N_6836);
xor U7180 (N_7180,N_6271,N_6553);
xnor U7181 (N_7181,N_6558,N_6003);
nand U7182 (N_7182,N_6886,N_6890);
or U7183 (N_7183,N_6834,N_6024);
and U7184 (N_7184,N_6211,N_6057);
nand U7185 (N_7185,N_6088,N_6121);
xnor U7186 (N_7186,N_6105,N_6766);
and U7187 (N_7187,N_6797,N_6987);
nor U7188 (N_7188,N_6570,N_6592);
or U7189 (N_7189,N_6027,N_6445);
nand U7190 (N_7190,N_6672,N_6668);
or U7191 (N_7191,N_6103,N_6255);
nand U7192 (N_7192,N_6098,N_6728);
and U7193 (N_7193,N_6021,N_6733);
xnor U7194 (N_7194,N_6950,N_6501);
nor U7195 (N_7195,N_6322,N_6547);
or U7196 (N_7196,N_6165,N_6523);
nor U7197 (N_7197,N_6936,N_6735);
and U7198 (N_7198,N_6861,N_6017);
or U7199 (N_7199,N_6065,N_6964);
xnor U7200 (N_7200,N_6061,N_6355);
xor U7201 (N_7201,N_6925,N_6037);
or U7202 (N_7202,N_6334,N_6026);
nor U7203 (N_7203,N_6321,N_6080);
nand U7204 (N_7204,N_6941,N_6993);
and U7205 (N_7205,N_6022,N_6036);
nand U7206 (N_7206,N_6231,N_6914);
and U7207 (N_7207,N_6073,N_6606);
or U7208 (N_7208,N_6203,N_6328);
and U7209 (N_7209,N_6030,N_6530);
nor U7210 (N_7210,N_6154,N_6808);
and U7211 (N_7211,N_6499,N_6180);
or U7212 (N_7212,N_6525,N_6146);
xnor U7213 (N_7213,N_6375,N_6832);
nand U7214 (N_7214,N_6968,N_6552);
nand U7215 (N_7215,N_6979,N_6193);
and U7216 (N_7216,N_6546,N_6973);
nand U7217 (N_7217,N_6279,N_6541);
or U7218 (N_7218,N_6043,N_6588);
or U7219 (N_7219,N_6772,N_6018);
nand U7220 (N_7220,N_6534,N_6210);
and U7221 (N_7221,N_6768,N_6652);
and U7222 (N_7222,N_6446,N_6475);
or U7223 (N_7223,N_6353,N_6550);
or U7224 (N_7224,N_6837,N_6497);
xnor U7225 (N_7225,N_6309,N_6114);
nor U7226 (N_7226,N_6282,N_6083);
and U7227 (N_7227,N_6721,N_6265);
or U7228 (N_7228,N_6780,N_6631);
and U7229 (N_7229,N_6585,N_6152);
or U7230 (N_7230,N_6955,N_6479);
nor U7231 (N_7231,N_6594,N_6345);
and U7232 (N_7232,N_6747,N_6090);
or U7233 (N_7233,N_6576,N_6401);
nand U7234 (N_7234,N_6809,N_6171);
or U7235 (N_7235,N_6106,N_6075);
xor U7236 (N_7236,N_6511,N_6186);
nand U7237 (N_7237,N_6729,N_6204);
or U7238 (N_7238,N_6249,N_6360);
or U7239 (N_7239,N_6798,N_6506);
and U7240 (N_7240,N_6937,N_6622);
and U7241 (N_7241,N_6619,N_6316);
and U7242 (N_7242,N_6776,N_6044);
and U7243 (N_7243,N_6011,N_6307);
nand U7244 (N_7244,N_6208,N_6716);
or U7245 (N_7245,N_6630,N_6025);
or U7246 (N_7246,N_6314,N_6415);
and U7247 (N_7247,N_6241,N_6634);
nand U7248 (N_7248,N_6758,N_6392);
nand U7249 (N_7249,N_6245,N_6196);
and U7250 (N_7250,N_6366,N_6819);
xor U7251 (N_7251,N_6134,N_6734);
nor U7252 (N_7252,N_6096,N_6388);
and U7253 (N_7253,N_6095,N_6148);
nand U7254 (N_7254,N_6540,N_6348);
nand U7255 (N_7255,N_6133,N_6678);
and U7256 (N_7256,N_6324,N_6650);
and U7257 (N_7257,N_6932,N_6461);
and U7258 (N_7258,N_6191,N_6717);
nand U7259 (N_7259,N_6034,N_6846);
or U7260 (N_7260,N_6929,N_6660);
nand U7261 (N_7261,N_6346,N_6869);
and U7262 (N_7262,N_6252,N_6649);
or U7263 (N_7263,N_6545,N_6269);
nor U7264 (N_7264,N_6913,N_6748);
nand U7265 (N_7265,N_6153,N_6010);
and U7266 (N_7266,N_6082,N_6209);
nand U7267 (N_7267,N_6212,N_6940);
xor U7268 (N_7268,N_6100,N_6865);
xnor U7269 (N_7269,N_6367,N_6673);
and U7270 (N_7270,N_6086,N_6866);
or U7271 (N_7271,N_6333,N_6637);
or U7272 (N_7272,N_6223,N_6752);
nand U7273 (N_7273,N_6404,N_6099);
nand U7274 (N_7274,N_6727,N_6635);
nor U7275 (N_7275,N_6060,N_6456);
or U7276 (N_7276,N_6812,N_6551);
nand U7277 (N_7277,N_6740,N_6848);
nor U7278 (N_7278,N_6450,N_6532);
or U7279 (N_7279,N_6290,N_6123);
nand U7280 (N_7280,N_6626,N_6774);
nor U7281 (N_7281,N_6342,N_6920);
nor U7282 (N_7282,N_6429,N_6732);
nor U7283 (N_7283,N_6810,N_6382);
or U7284 (N_7284,N_6921,N_6719);
nor U7285 (N_7285,N_6425,N_6942);
xor U7286 (N_7286,N_6136,N_6039);
and U7287 (N_7287,N_6268,N_6986);
or U7288 (N_7288,N_6315,N_6820);
or U7289 (N_7289,N_6286,N_6919);
and U7290 (N_7290,N_6473,N_6827);
and U7291 (N_7291,N_6369,N_6195);
nor U7292 (N_7292,N_6291,N_6624);
nand U7293 (N_7293,N_6283,N_6947);
xnor U7294 (N_7294,N_6710,N_6374);
or U7295 (N_7295,N_6217,N_6312);
nand U7296 (N_7296,N_6579,N_6443);
nor U7297 (N_7297,N_6788,N_6674);
and U7298 (N_7298,N_6663,N_6354);
and U7299 (N_7299,N_6236,N_6528);
and U7300 (N_7300,N_6966,N_6625);
or U7301 (N_7301,N_6306,N_6915);
nor U7302 (N_7302,N_6926,N_6310);
and U7303 (N_7303,N_6686,N_6982);
or U7304 (N_7304,N_6851,N_6433);
and U7305 (N_7305,N_6960,N_6904);
nand U7306 (N_7306,N_6862,N_6697);
nand U7307 (N_7307,N_6991,N_6507);
nand U7308 (N_7308,N_6014,N_6164);
or U7309 (N_7309,N_6332,N_6517);
nand U7310 (N_7310,N_6317,N_6581);
and U7311 (N_7311,N_6416,N_6349);
and U7312 (N_7312,N_6372,N_6681);
nor U7313 (N_7313,N_6163,N_6341);
nor U7314 (N_7314,N_6162,N_6370);
nand U7315 (N_7315,N_6364,N_6763);
nor U7316 (N_7316,N_6378,N_6535);
or U7317 (N_7317,N_6140,N_6001);
and U7318 (N_7318,N_6670,N_6141);
nor U7319 (N_7319,N_6912,N_6400);
nor U7320 (N_7320,N_6092,N_6067);
nor U7321 (N_7321,N_6161,N_6233);
xor U7322 (N_7322,N_6399,N_6130);
nand U7323 (N_7323,N_6391,N_6992);
and U7324 (N_7324,N_6221,N_6753);
nand U7325 (N_7325,N_6361,N_6888);
nand U7326 (N_7326,N_6237,N_6803);
and U7327 (N_7327,N_6045,N_6052);
nand U7328 (N_7328,N_6459,N_6595);
nand U7329 (N_7329,N_6730,N_6543);
nor U7330 (N_7330,N_6248,N_6049);
nand U7331 (N_7331,N_6449,N_6854);
and U7332 (N_7332,N_6826,N_6807);
nor U7333 (N_7333,N_6840,N_6174);
nor U7334 (N_7334,N_6632,N_6132);
and U7335 (N_7335,N_6669,N_6215);
and U7336 (N_7336,N_6427,N_6770);
and U7337 (N_7337,N_6104,N_6238);
or U7338 (N_7338,N_6954,N_6393);
or U7339 (N_7339,N_6428,N_6407);
nor U7340 (N_7340,N_6653,N_6129);
nand U7341 (N_7341,N_6580,N_6745);
and U7342 (N_7342,N_6706,N_6591);
nand U7343 (N_7343,N_6976,N_6567);
xnor U7344 (N_7344,N_6110,N_6396);
or U7345 (N_7345,N_6587,N_6949);
and U7346 (N_7346,N_6875,N_6998);
or U7347 (N_7347,N_6402,N_6262);
or U7348 (N_7348,N_6131,N_6013);
nor U7349 (N_7349,N_6775,N_6781);
xor U7350 (N_7350,N_6616,N_6486);
nor U7351 (N_7351,N_6028,N_6891);
or U7352 (N_7352,N_6124,N_6438);
nand U7353 (N_7353,N_6593,N_6572);
nor U7354 (N_7354,N_6508,N_6526);
xnor U7355 (N_7355,N_6485,N_6157);
and U7356 (N_7356,N_6935,N_6557);
or U7357 (N_7357,N_6539,N_6627);
nand U7358 (N_7358,N_6559,N_6873);
or U7359 (N_7359,N_6894,N_6767);
nand U7360 (N_7360,N_6147,N_6467);
nand U7361 (N_7361,N_6778,N_6882);
nand U7362 (N_7362,N_6487,N_6665);
nor U7363 (N_7363,N_6952,N_6056);
xnor U7364 (N_7364,N_6741,N_6138);
or U7365 (N_7365,N_6319,N_6845);
nor U7366 (N_7366,N_6413,N_6905);
nor U7367 (N_7367,N_6358,N_6403);
or U7368 (N_7368,N_6864,N_6498);
or U7369 (N_7369,N_6116,N_6244);
and U7370 (N_7370,N_6762,N_6769);
xor U7371 (N_7371,N_6053,N_6183);
nand U7372 (N_7372,N_6032,N_6561);
and U7373 (N_7373,N_6586,N_6004);
nor U7374 (N_7374,N_6137,N_6997);
nor U7375 (N_7375,N_6298,N_6609);
or U7376 (N_7376,N_6604,N_6908);
or U7377 (N_7377,N_6197,N_6326);
nand U7378 (N_7378,N_6843,N_6078);
nand U7379 (N_7379,N_6292,N_6005);
and U7380 (N_7380,N_6294,N_6704);
or U7381 (N_7381,N_6887,N_6884);
or U7382 (N_7382,N_6718,N_6149);
nand U7383 (N_7383,N_6145,N_6125);
or U7384 (N_7384,N_6454,N_6430);
nor U7385 (N_7385,N_6872,N_6823);
nand U7386 (N_7386,N_6320,N_6198);
and U7387 (N_7387,N_6538,N_6142);
nor U7388 (N_7388,N_6893,N_6420);
nand U7389 (N_7389,N_6943,N_6117);
or U7390 (N_7390,N_6746,N_6423);
and U7391 (N_7391,N_6182,N_6417);
nand U7392 (N_7392,N_6460,N_6647);
or U7393 (N_7393,N_6529,N_6868);
nand U7394 (N_7394,N_6876,N_6945);
xnor U7395 (N_7395,N_6442,N_6806);
and U7396 (N_7396,N_6377,N_6682);
nor U7397 (N_7397,N_6304,N_6308);
nand U7398 (N_7398,N_6379,N_6536);
or U7399 (N_7399,N_6749,N_6094);
xnor U7400 (N_7400,N_6492,N_6458);
nor U7401 (N_7401,N_6589,N_6337);
nand U7402 (N_7402,N_6738,N_6694);
xnor U7403 (N_7403,N_6621,N_6251);
nand U7404 (N_7404,N_6437,N_6531);
nand U7405 (N_7405,N_6811,N_6703);
or U7406 (N_7406,N_6513,N_6190);
nand U7407 (N_7407,N_6439,N_6962);
xor U7408 (N_7408,N_6978,N_6247);
and U7409 (N_7409,N_6466,N_6828);
or U7410 (N_7410,N_6109,N_6156);
nor U7411 (N_7411,N_6135,N_6563);
and U7412 (N_7412,N_6994,N_6118);
xor U7413 (N_7413,N_6657,N_6406);
nand U7414 (N_7414,N_6395,N_6996);
or U7415 (N_7415,N_6870,N_6267);
and U7416 (N_7416,N_6661,N_6948);
nand U7417 (N_7417,N_6639,N_6085);
nor U7418 (N_7418,N_6038,N_6722);
and U7419 (N_7419,N_6144,N_6662);
nor U7420 (N_7420,N_6927,N_6898);
nor U7421 (N_7421,N_6220,N_6242);
and U7422 (N_7422,N_6235,N_6000);
nor U7423 (N_7423,N_6793,N_6243);
or U7424 (N_7424,N_6521,N_6638);
nand U7425 (N_7425,N_6980,N_6202);
nand U7426 (N_7426,N_6975,N_6693);
or U7427 (N_7427,N_6689,N_6910);
nor U7428 (N_7428,N_6356,N_6101);
and U7429 (N_7429,N_6712,N_6906);
or U7430 (N_7430,N_6515,N_6158);
or U7431 (N_7431,N_6784,N_6897);
and U7432 (N_7432,N_6066,N_6825);
nor U7433 (N_7433,N_6760,N_6472);
nor U7434 (N_7434,N_6444,N_6471);
and U7435 (N_7435,N_6608,N_6956);
nand U7436 (N_7436,N_6435,N_6582);
or U7437 (N_7437,N_6569,N_6059);
nand U7438 (N_7438,N_6176,N_6113);
nor U7439 (N_7439,N_6184,N_6744);
xnor U7440 (N_7440,N_6207,N_6311);
and U7441 (N_7441,N_6159,N_6654);
and U7442 (N_7442,N_6881,N_6411);
nand U7443 (N_7443,N_6046,N_6726);
and U7444 (N_7444,N_6276,N_6805);
nor U7445 (N_7445,N_6188,N_6850);
and U7446 (N_7446,N_6883,N_6009);
nand U7447 (N_7447,N_6063,N_6228);
nor U7448 (N_7448,N_6549,N_6409);
and U7449 (N_7449,N_6288,N_6600);
and U7450 (N_7450,N_6691,N_6885);
or U7451 (N_7451,N_6179,N_6853);
nor U7452 (N_7452,N_6225,N_6577);
and U7453 (N_7453,N_6213,N_6934);
nor U7454 (N_7454,N_6548,N_6953);
and U7455 (N_7455,N_6335,N_6350);
and U7456 (N_7456,N_6688,N_6041);
nor U7457 (N_7457,N_6239,N_6155);
xor U7458 (N_7458,N_6470,N_6301);
nor U7459 (N_7459,N_6817,N_6946);
nor U7460 (N_7460,N_6494,N_6192);
and U7461 (N_7461,N_6699,N_6284);
and U7462 (N_7462,N_6476,N_6042);
or U7463 (N_7463,N_6566,N_6381);
nor U7464 (N_7464,N_6918,N_6263);
and U7465 (N_7465,N_6451,N_6575);
nor U7466 (N_7466,N_6659,N_6340);
and U7467 (N_7467,N_6422,N_6931);
nor U7468 (N_7468,N_6901,N_6006);
or U7469 (N_7469,N_6518,N_6617);
or U7470 (N_7470,N_6166,N_6705);
and U7471 (N_7471,N_6071,N_6275);
xor U7472 (N_7472,N_6390,N_6431);
nand U7473 (N_7473,N_6408,N_6436);
and U7474 (N_7474,N_6527,N_6493);
nor U7475 (N_7475,N_6855,N_6280);
xnor U7476 (N_7476,N_6256,N_6764);
or U7477 (N_7477,N_6961,N_6200);
nor U7478 (N_7478,N_6405,N_6618);
nor U7479 (N_7479,N_6564,N_6368);
xor U7480 (N_7480,N_6285,N_6614);
and U7481 (N_7481,N_6878,N_6468);
and U7482 (N_7482,N_6610,N_6230);
nand U7483 (N_7483,N_6455,N_6983);
nor U7484 (N_7484,N_6175,N_6259);
and U7485 (N_7485,N_6715,N_6981);
or U7486 (N_7486,N_6160,N_6002);
or U7487 (N_7487,N_6440,N_6185);
nor U7488 (N_7488,N_6260,N_6281);
nor U7489 (N_7489,N_6599,N_6253);
or U7490 (N_7490,N_6463,N_6802);
nand U7491 (N_7491,N_6035,N_6902);
xnor U7492 (N_7492,N_6612,N_6938);
or U7493 (N_7493,N_6477,N_6743);
or U7494 (N_7494,N_6344,N_6074);
nor U7495 (N_7495,N_6977,N_6394);
and U7496 (N_7496,N_6754,N_6713);
nand U7497 (N_7497,N_6289,N_6544);
nand U7498 (N_7498,N_6930,N_6020);
nor U7499 (N_7499,N_6386,N_6813);
or U7500 (N_7500,N_6536,N_6042);
and U7501 (N_7501,N_6114,N_6549);
nor U7502 (N_7502,N_6141,N_6647);
or U7503 (N_7503,N_6097,N_6955);
nor U7504 (N_7504,N_6409,N_6890);
nor U7505 (N_7505,N_6926,N_6272);
nor U7506 (N_7506,N_6462,N_6207);
nand U7507 (N_7507,N_6437,N_6235);
nor U7508 (N_7508,N_6176,N_6920);
xnor U7509 (N_7509,N_6209,N_6013);
and U7510 (N_7510,N_6281,N_6188);
nand U7511 (N_7511,N_6749,N_6737);
nand U7512 (N_7512,N_6131,N_6640);
nand U7513 (N_7513,N_6738,N_6068);
nand U7514 (N_7514,N_6829,N_6683);
nor U7515 (N_7515,N_6442,N_6953);
and U7516 (N_7516,N_6691,N_6957);
nor U7517 (N_7517,N_6401,N_6179);
and U7518 (N_7518,N_6794,N_6591);
and U7519 (N_7519,N_6909,N_6933);
or U7520 (N_7520,N_6006,N_6509);
nor U7521 (N_7521,N_6458,N_6295);
and U7522 (N_7522,N_6567,N_6710);
nor U7523 (N_7523,N_6844,N_6390);
nand U7524 (N_7524,N_6314,N_6424);
or U7525 (N_7525,N_6225,N_6437);
and U7526 (N_7526,N_6979,N_6177);
and U7527 (N_7527,N_6637,N_6465);
xor U7528 (N_7528,N_6238,N_6360);
or U7529 (N_7529,N_6839,N_6593);
nor U7530 (N_7530,N_6519,N_6093);
nand U7531 (N_7531,N_6085,N_6980);
xnor U7532 (N_7532,N_6655,N_6097);
and U7533 (N_7533,N_6811,N_6620);
xnor U7534 (N_7534,N_6828,N_6709);
nand U7535 (N_7535,N_6043,N_6919);
nand U7536 (N_7536,N_6404,N_6400);
and U7537 (N_7537,N_6265,N_6011);
nor U7538 (N_7538,N_6207,N_6000);
and U7539 (N_7539,N_6417,N_6919);
nand U7540 (N_7540,N_6466,N_6294);
or U7541 (N_7541,N_6016,N_6391);
nand U7542 (N_7542,N_6331,N_6953);
nand U7543 (N_7543,N_6235,N_6689);
nor U7544 (N_7544,N_6384,N_6901);
or U7545 (N_7545,N_6432,N_6527);
nand U7546 (N_7546,N_6103,N_6831);
xor U7547 (N_7547,N_6583,N_6111);
and U7548 (N_7548,N_6676,N_6396);
nand U7549 (N_7549,N_6633,N_6404);
nand U7550 (N_7550,N_6312,N_6660);
nor U7551 (N_7551,N_6581,N_6549);
nor U7552 (N_7552,N_6108,N_6860);
nand U7553 (N_7553,N_6832,N_6924);
and U7554 (N_7554,N_6983,N_6427);
nor U7555 (N_7555,N_6620,N_6837);
and U7556 (N_7556,N_6851,N_6412);
or U7557 (N_7557,N_6665,N_6531);
nand U7558 (N_7558,N_6618,N_6351);
nand U7559 (N_7559,N_6126,N_6709);
nor U7560 (N_7560,N_6395,N_6766);
nor U7561 (N_7561,N_6181,N_6769);
nand U7562 (N_7562,N_6498,N_6351);
and U7563 (N_7563,N_6235,N_6005);
nand U7564 (N_7564,N_6291,N_6904);
and U7565 (N_7565,N_6671,N_6155);
and U7566 (N_7566,N_6739,N_6333);
or U7567 (N_7567,N_6195,N_6966);
and U7568 (N_7568,N_6703,N_6615);
xor U7569 (N_7569,N_6484,N_6010);
and U7570 (N_7570,N_6682,N_6942);
xor U7571 (N_7571,N_6322,N_6782);
and U7572 (N_7572,N_6921,N_6321);
nor U7573 (N_7573,N_6778,N_6687);
and U7574 (N_7574,N_6070,N_6090);
nor U7575 (N_7575,N_6158,N_6448);
nand U7576 (N_7576,N_6632,N_6380);
or U7577 (N_7577,N_6442,N_6779);
and U7578 (N_7578,N_6195,N_6128);
xnor U7579 (N_7579,N_6468,N_6590);
nand U7580 (N_7580,N_6748,N_6404);
and U7581 (N_7581,N_6256,N_6748);
nor U7582 (N_7582,N_6848,N_6633);
nand U7583 (N_7583,N_6395,N_6631);
xnor U7584 (N_7584,N_6505,N_6043);
or U7585 (N_7585,N_6484,N_6109);
nor U7586 (N_7586,N_6199,N_6959);
nor U7587 (N_7587,N_6294,N_6524);
nor U7588 (N_7588,N_6865,N_6331);
or U7589 (N_7589,N_6295,N_6155);
nand U7590 (N_7590,N_6777,N_6435);
xor U7591 (N_7591,N_6445,N_6788);
nand U7592 (N_7592,N_6974,N_6874);
nor U7593 (N_7593,N_6906,N_6024);
xnor U7594 (N_7594,N_6691,N_6716);
xnor U7595 (N_7595,N_6976,N_6728);
nor U7596 (N_7596,N_6237,N_6276);
nor U7597 (N_7597,N_6144,N_6324);
nor U7598 (N_7598,N_6040,N_6508);
xnor U7599 (N_7599,N_6105,N_6476);
and U7600 (N_7600,N_6977,N_6015);
or U7601 (N_7601,N_6027,N_6822);
nor U7602 (N_7602,N_6407,N_6092);
and U7603 (N_7603,N_6932,N_6311);
and U7604 (N_7604,N_6435,N_6176);
nor U7605 (N_7605,N_6675,N_6460);
or U7606 (N_7606,N_6701,N_6044);
or U7607 (N_7607,N_6659,N_6011);
xnor U7608 (N_7608,N_6696,N_6970);
xnor U7609 (N_7609,N_6832,N_6934);
xnor U7610 (N_7610,N_6074,N_6458);
and U7611 (N_7611,N_6288,N_6389);
nor U7612 (N_7612,N_6737,N_6897);
nand U7613 (N_7613,N_6915,N_6754);
nor U7614 (N_7614,N_6469,N_6443);
or U7615 (N_7615,N_6116,N_6844);
or U7616 (N_7616,N_6103,N_6993);
nand U7617 (N_7617,N_6981,N_6140);
nand U7618 (N_7618,N_6112,N_6094);
or U7619 (N_7619,N_6646,N_6311);
nor U7620 (N_7620,N_6376,N_6835);
nand U7621 (N_7621,N_6414,N_6241);
nand U7622 (N_7622,N_6305,N_6654);
nor U7623 (N_7623,N_6770,N_6383);
and U7624 (N_7624,N_6767,N_6409);
nor U7625 (N_7625,N_6332,N_6390);
and U7626 (N_7626,N_6347,N_6722);
and U7627 (N_7627,N_6104,N_6613);
and U7628 (N_7628,N_6568,N_6594);
or U7629 (N_7629,N_6104,N_6664);
nor U7630 (N_7630,N_6348,N_6353);
nand U7631 (N_7631,N_6895,N_6753);
nand U7632 (N_7632,N_6271,N_6589);
nor U7633 (N_7633,N_6100,N_6646);
and U7634 (N_7634,N_6166,N_6272);
nand U7635 (N_7635,N_6325,N_6502);
or U7636 (N_7636,N_6731,N_6109);
nor U7637 (N_7637,N_6435,N_6257);
or U7638 (N_7638,N_6961,N_6380);
nand U7639 (N_7639,N_6311,N_6606);
or U7640 (N_7640,N_6008,N_6210);
nor U7641 (N_7641,N_6244,N_6231);
and U7642 (N_7642,N_6808,N_6834);
nand U7643 (N_7643,N_6864,N_6591);
or U7644 (N_7644,N_6563,N_6749);
or U7645 (N_7645,N_6051,N_6924);
or U7646 (N_7646,N_6926,N_6102);
nor U7647 (N_7647,N_6239,N_6153);
nand U7648 (N_7648,N_6453,N_6859);
or U7649 (N_7649,N_6420,N_6109);
or U7650 (N_7650,N_6639,N_6543);
nand U7651 (N_7651,N_6194,N_6111);
and U7652 (N_7652,N_6876,N_6342);
nor U7653 (N_7653,N_6967,N_6585);
or U7654 (N_7654,N_6584,N_6315);
or U7655 (N_7655,N_6918,N_6447);
xnor U7656 (N_7656,N_6981,N_6619);
and U7657 (N_7657,N_6946,N_6987);
or U7658 (N_7658,N_6762,N_6627);
nand U7659 (N_7659,N_6611,N_6743);
nor U7660 (N_7660,N_6229,N_6736);
or U7661 (N_7661,N_6676,N_6613);
nor U7662 (N_7662,N_6102,N_6201);
nor U7663 (N_7663,N_6221,N_6428);
xnor U7664 (N_7664,N_6870,N_6530);
and U7665 (N_7665,N_6881,N_6568);
and U7666 (N_7666,N_6212,N_6282);
xnor U7667 (N_7667,N_6459,N_6456);
and U7668 (N_7668,N_6049,N_6081);
nor U7669 (N_7669,N_6621,N_6362);
and U7670 (N_7670,N_6133,N_6514);
nand U7671 (N_7671,N_6905,N_6288);
and U7672 (N_7672,N_6624,N_6640);
and U7673 (N_7673,N_6099,N_6794);
xor U7674 (N_7674,N_6730,N_6715);
or U7675 (N_7675,N_6481,N_6486);
xnor U7676 (N_7676,N_6371,N_6560);
and U7677 (N_7677,N_6448,N_6152);
and U7678 (N_7678,N_6086,N_6360);
or U7679 (N_7679,N_6344,N_6231);
or U7680 (N_7680,N_6621,N_6823);
and U7681 (N_7681,N_6033,N_6666);
nand U7682 (N_7682,N_6390,N_6625);
nand U7683 (N_7683,N_6648,N_6130);
nand U7684 (N_7684,N_6587,N_6656);
and U7685 (N_7685,N_6867,N_6945);
and U7686 (N_7686,N_6925,N_6753);
or U7687 (N_7687,N_6121,N_6816);
nor U7688 (N_7688,N_6342,N_6761);
or U7689 (N_7689,N_6200,N_6712);
nand U7690 (N_7690,N_6872,N_6534);
and U7691 (N_7691,N_6736,N_6808);
nand U7692 (N_7692,N_6183,N_6869);
nand U7693 (N_7693,N_6446,N_6934);
and U7694 (N_7694,N_6039,N_6510);
xor U7695 (N_7695,N_6855,N_6336);
or U7696 (N_7696,N_6492,N_6370);
nand U7697 (N_7697,N_6061,N_6592);
xor U7698 (N_7698,N_6318,N_6665);
nand U7699 (N_7699,N_6933,N_6832);
and U7700 (N_7700,N_6509,N_6223);
and U7701 (N_7701,N_6930,N_6494);
nor U7702 (N_7702,N_6534,N_6909);
and U7703 (N_7703,N_6492,N_6459);
nand U7704 (N_7704,N_6885,N_6472);
nor U7705 (N_7705,N_6758,N_6491);
nor U7706 (N_7706,N_6613,N_6422);
nor U7707 (N_7707,N_6295,N_6875);
nor U7708 (N_7708,N_6835,N_6522);
nand U7709 (N_7709,N_6968,N_6205);
xor U7710 (N_7710,N_6151,N_6078);
and U7711 (N_7711,N_6566,N_6849);
nor U7712 (N_7712,N_6192,N_6048);
nor U7713 (N_7713,N_6084,N_6858);
and U7714 (N_7714,N_6297,N_6448);
or U7715 (N_7715,N_6761,N_6391);
xnor U7716 (N_7716,N_6014,N_6827);
nand U7717 (N_7717,N_6632,N_6535);
and U7718 (N_7718,N_6280,N_6927);
nand U7719 (N_7719,N_6945,N_6515);
and U7720 (N_7720,N_6111,N_6936);
and U7721 (N_7721,N_6083,N_6892);
nand U7722 (N_7722,N_6450,N_6765);
and U7723 (N_7723,N_6492,N_6799);
xnor U7724 (N_7724,N_6042,N_6605);
or U7725 (N_7725,N_6515,N_6944);
and U7726 (N_7726,N_6375,N_6202);
nand U7727 (N_7727,N_6327,N_6712);
nor U7728 (N_7728,N_6344,N_6181);
nand U7729 (N_7729,N_6118,N_6467);
nand U7730 (N_7730,N_6585,N_6175);
nor U7731 (N_7731,N_6879,N_6381);
xnor U7732 (N_7732,N_6880,N_6518);
or U7733 (N_7733,N_6380,N_6002);
and U7734 (N_7734,N_6563,N_6163);
nor U7735 (N_7735,N_6974,N_6043);
nor U7736 (N_7736,N_6907,N_6574);
or U7737 (N_7737,N_6494,N_6948);
nand U7738 (N_7738,N_6345,N_6590);
or U7739 (N_7739,N_6424,N_6727);
or U7740 (N_7740,N_6391,N_6616);
and U7741 (N_7741,N_6141,N_6774);
xnor U7742 (N_7742,N_6834,N_6123);
and U7743 (N_7743,N_6735,N_6512);
nand U7744 (N_7744,N_6544,N_6900);
nand U7745 (N_7745,N_6558,N_6740);
or U7746 (N_7746,N_6152,N_6805);
and U7747 (N_7747,N_6045,N_6130);
and U7748 (N_7748,N_6448,N_6319);
xnor U7749 (N_7749,N_6356,N_6328);
nand U7750 (N_7750,N_6706,N_6637);
nor U7751 (N_7751,N_6204,N_6754);
xnor U7752 (N_7752,N_6601,N_6765);
xnor U7753 (N_7753,N_6514,N_6374);
nor U7754 (N_7754,N_6585,N_6798);
and U7755 (N_7755,N_6454,N_6173);
and U7756 (N_7756,N_6436,N_6503);
nand U7757 (N_7757,N_6984,N_6616);
nor U7758 (N_7758,N_6791,N_6702);
nor U7759 (N_7759,N_6956,N_6724);
nand U7760 (N_7760,N_6446,N_6606);
nor U7761 (N_7761,N_6510,N_6897);
or U7762 (N_7762,N_6330,N_6350);
and U7763 (N_7763,N_6508,N_6074);
xor U7764 (N_7764,N_6178,N_6371);
nor U7765 (N_7765,N_6417,N_6454);
nand U7766 (N_7766,N_6578,N_6123);
or U7767 (N_7767,N_6385,N_6821);
nor U7768 (N_7768,N_6804,N_6576);
nor U7769 (N_7769,N_6316,N_6732);
and U7770 (N_7770,N_6053,N_6236);
and U7771 (N_7771,N_6448,N_6906);
xor U7772 (N_7772,N_6901,N_6152);
nor U7773 (N_7773,N_6127,N_6301);
nor U7774 (N_7774,N_6629,N_6697);
nand U7775 (N_7775,N_6513,N_6834);
nor U7776 (N_7776,N_6488,N_6178);
nor U7777 (N_7777,N_6260,N_6780);
nand U7778 (N_7778,N_6966,N_6093);
and U7779 (N_7779,N_6933,N_6594);
xnor U7780 (N_7780,N_6784,N_6150);
nand U7781 (N_7781,N_6140,N_6210);
nand U7782 (N_7782,N_6960,N_6085);
or U7783 (N_7783,N_6896,N_6302);
nor U7784 (N_7784,N_6275,N_6152);
or U7785 (N_7785,N_6699,N_6175);
or U7786 (N_7786,N_6175,N_6469);
nor U7787 (N_7787,N_6480,N_6029);
nor U7788 (N_7788,N_6874,N_6861);
or U7789 (N_7789,N_6047,N_6293);
nand U7790 (N_7790,N_6422,N_6232);
nor U7791 (N_7791,N_6468,N_6288);
and U7792 (N_7792,N_6006,N_6418);
xnor U7793 (N_7793,N_6545,N_6276);
and U7794 (N_7794,N_6219,N_6196);
nor U7795 (N_7795,N_6722,N_6101);
or U7796 (N_7796,N_6153,N_6608);
or U7797 (N_7797,N_6023,N_6249);
nand U7798 (N_7798,N_6238,N_6468);
or U7799 (N_7799,N_6196,N_6405);
nor U7800 (N_7800,N_6909,N_6482);
xnor U7801 (N_7801,N_6971,N_6678);
nand U7802 (N_7802,N_6486,N_6157);
nor U7803 (N_7803,N_6138,N_6348);
nand U7804 (N_7804,N_6222,N_6862);
nand U7805 (N_7805,N_6439,N_6919);
or U7806 (N_7806,N_6093,N_6160);
and U7807 (N_7807,N_6526,N_6567);
xor U7808 (N_7808,N_6657,N_6351);
and U7809 (N_7809,N_6202,N_6708);
nand U7810 (N_7810,N_6894,N_6327);
and U7811 (N_7811,N_6679,N_6018);
and U7812 (N_7812,N_6751,N_6586);
nor U7813 (N_7813,N_6553,N_6537);
nand U7814 (N_7814,N_6094,N_6237);
nor U7815 (N_7815,N_6823,N_6984);
or U7816 (N_7816,N_6414,N_6351);
xnor U7817 (N_7817,N_6255,N_6054);
nand U7818 (N_7818,N_6585,N_6557);
nand U7819 (N_7819,N_6513,N_6371);
nand U7820 (N_7820,N_6886,N_6279);
xnor U7821 (N_7821,N_6933,N_6901);
and U7822 (N_7822,N_6876,N_6966);
or U7823 (N_7823,N_6652,N_6163);
or U7824 (N_7824,N_6245,N_6538);
or U7825 (N_7825,N_6262,N_6248);
nor U7826 (N_7826,N_6705,N_6058);
nor U7827 (N_7827,N_6954,N_6672);
nor U7828 (N_7828,N_6240,N_6524);
or U7829 (N_7829,N_6299,N_6924);
nand U7830 (N_7830,N_6129,N_6014);
nor U7831 (N_7831,N_6021,N_6131);
or U7832 (N_7832,N_6320,N_6984);
nor U7833 (N_7833,N_6262,N_6546);
and U7834 (N_7834,N_6023,N_6328);
or U7835 (N_7835,N_6535,N_6563);
nor U7836 (N_7836,N_6344,N_6873);
nand U7837 (N_7837,N_6489,N_6706);
or U7838 (N_7838,N_6408,N_6197);
nand U7839 (N_7839,N_6277,N_6350);
or U7840 (N_7840,N_6389,N_6949);
nor U7841 (N_7841,N_6498,N_6304);
nor U7842 (N_7842,N_6155,N_6072);
nor U7843 (N_7843,N_6553,N_6782);
and U7844 (N_7844,N_6286,N_6646);
nand U7845 (N_7845,N_6144,N_6049);
nand U7846 (N_7846,N_6995,N_6232);
xor U7847 (N_7847,N_6077,N_6350);
or U7848 (N_7848,N_6225,N_6135);
xnor U7849 (N_7849,N_6138,N_6010);
or U7850 (N_7850,N_6795,N_6267);
nor U7851 (N_7851,N_6707,N_6426);
nand U7852 (N_7852,N_6647,N_6458);
nor U7853 (N_7853,N_6773,N_6954);
nor U7854 (N_7854,N_6175,N_6637);
or U7855 (N_7855,N_6379,N_6089);
xnor U7856 (N_7856,N_6055,N_6650);
xnor U7857 (N_7857,N_6598,N_6666);
nor U7858 (N_7858,N_6292,N_6145);
or U7859 (N_7859,N_6594,N_6321);
and U7860 (N_7860,N_6873,N_6824);
nor U7861 (N_7861,N_6413,N_6540);
xor U7862 (N_7862,N_6735,N_6320);
xnor U7863 (N_7863,N_6336,N_6303);
and U7864 (N_7864,N_6283,N_6454);
nor U7865 (N_7865,N_6608,N_6708);
or U7866 (N_7866,N_6080,N_6988);
xnor U7867 (N_7867,N_6143,N_6226);
or U7868 (N_7868,N_6248,N_6865);
or U7869 (N_7869,N_6184,N_6761);
nor U7870 (N_7870,N_6890,N_6388);
or U7871 (N_7871,N_6390,N_6898);
nor U7872 (N_7872,N_6659,N_6003);
and U7873 (N_7873,N_6158,N_6537);
or U7874 (N_7874,N_6093,N_6330);
nor U7875 (N_7875,N_6471,N_6105);
and U7876 (N_7876,N_6689,N_6060);
and U7877 (N_7877,N_6381,N_6813);
nor U7878 (N_7878,N_6145,N_6559);
nor U7879 (N_7879,N_6044,N_6152);
or U7880 (N_7880,N_6403,N_6912);
and U7881 (N_7881,N_6541,N_6999);
nor U7882 (N_7882,N_6748,N_6693);
and U7883 (N_7883,N_6249,N_6552);
nor U7884 (N_7884,N_6309,N_6018);
and U7885 (N_7885,N_6517,N_6744);
and U7886 (N_7886,N_6078,N_6137);
nand U7887 (N_7887,N_6245,N_6024);
xnor U7888 (N_7888,N_6416,N_6782);
and U7889 (N_7889,N_6425,N_6794);
nor U7890 (N_7890,N_6985,N_6464);
and U7891 (N_7891,N_6443,N_6942);
nand U7892 (N_7892,N_6730,N_6675);
or U7893 (N_7893,N_6162,N_6228);
and U7894 (N_7894,N_6350,N_6369);
nand U7895 (N_7895,N_6387,N_6148);
xnor U7896 (N_7896,N_6348,N_6141);
or U7897 (N_7897,N_6410,N_6206);
nor U7898 (N_7898,N_6053,N_6645);
and U7899 (N_7899,N_6624,N_6762);
nand U7900 (N_7900,N_6335,N_6212);
and U7901 (N_7901,N_6274,N_6855);
or U7902 (N_7902,N_6523,N_6160);
nand U7903 (N_7903,N_6749,N_6370);
nor U7904 (N_7904,N_6902,N_6368);
nand U7905 (N_7905,N_6106,N_6438);
or U7906 (N_7906,N_6551,N_6796);
nor U7907 (N_7907,N_6153,N_6303);
or U7908 (N_7908,N_6139,N_6878);
and U7909 (N_7909,N_6029,N_6271);
xnor U7910 (N_7910,N_6239,N_6381);
xnor U7911 (N_7911,N_6126,N_6804);
nand U7912 (N_7912,N_6879,N_6130);
or U7913 (N_7913,N_6487,N_6337);
or U7914 (N_7914,N_6809,N_6875);
xor U7915 (N_7915,N_6016,N_6972);
and U7916 (N_7916,N_6570,N_6061);
and U7917 (N_7917,N_6963,N_6847);
nand U7918 (N_7918,N_6382,N_6198);
nor U7919 (N_7919,N_6922,N_6708);
xnor U7920 (N_7920,N_6974,N_6281);
and U7921 (N_7921,N_6842,N_6861);
or U7922 (N_7922,N_6958,N_6216);
and U7923 (N_7923,N_6575,N_6825);
nand U7924 (N_7924,N_6006,N_6863);
nor U7925 (N_7925,N_6267,N_6083);
nand U7926 (N_7926,N_6080,N_6649);
xnor U7927 (N_7927,N_6941,N_6762);
and U7928 (N_7928,N_6172,N_6356);
and U7929 (N_7929,N_6653,N_6305);
and U7930 (N_7930,N_6765,N_6475);
nor U7931 (N_7931,N_6601,N_6519);
xor U7932 (N_7932,N_6748,N_6369);
or U7933 (N_7933,N_6734,N_6148);
or U7934 (N_7934,N_6764,N_6386);
nor U7935 (N_7935,N_6553,N_6554);
and U7936 (N_7936,N_6847,N_6887);
and U7937 (N_7937,N_6088,N_6688);
and U7938 (N_7938,N_6980,N_6781);
or U7939 (N_7939,N_6889,N_6767);
xor U7940 (N_7940,N_6036,N_6232);
nand U7941 (N_7941,N_6379,N_6106);
and U7942 (N_7942,N_6294,N_6059);
nand U7943 (N_7943,N_6041,N_6470);
nor U7944 (N_7944,N_6380,N_6304);
and U7945 (N_7945,N_6570,N_6289);
nor U7946 (N_7946,N_6088,N_6455);
xnor U7947 (N_7947,N_6983,N_6358);
nor U7948 (N_7948,N_6274,N_6537);
or U7949 (N_7949,N_6074,N_6423);
nor U7950 (N_7950,N_6607,N_6195);
and U7951 (N_7951,N_6544,N_6821);
xor U7952 (N_7952,N_6686,N_6594);
xor U7953 (N_7953,N_6454,N_6089);
nand U7954 (N_7954,N_6554,N_6891);
nor U7955 (N_7955,N_6352,N_6149);
and U7956 (N_7956,N_6890,N_6623);
or U7957 (N_7957,N_6992,N_6842);
or U7958 (N_7958,N_6474,N_6778);
and U7959 (N_7959,N_6529,N_6539);
xnor U7960 (N_7960,N_6121,N_6217);
and U7961 (N_7961,N_6776,N_6838);
nand U7962 (N_7962,N_6285,N_6802);
nand U7963 (N_7963,N_6619,N_6249);
nand U7964 (N_7964,N_6960,N_6559);
nor U7965 (N_7965,N_6528,N_6721);
and U7966 (N_7966,N_6267,N_6241);
or U7967 (N_7967,N_6490,N_6059);
or U7968 (N_7968,N_6822,N_6650);
and U7969 (N_7969,N_6903,N_6803);
nor U7970 (N_7970,N_6892,N_6480);
nor U7971 (N_7971,N_6900,N_6595);
nand U7972 (N_7972,N_6638,N_6409);
or U7973 (N_7973,N_6741,N_6896);
nand U7974 (N_7974,N_6200,N_6422);
or U7975 (N_7975,N_6905,N_6755);
xnor U7976 (N_7976,N_6699,N_6373);
nand U7977 (N_7977,N_6866,N_6699);
and U7978 (N_7978,N_6038,N_6253);
nor U7979 (N_7979,N_6417,N_6607);
and U7980 (N_7980,N_6221,N_6308);
nor U7981 (N_7981,N_6029,N_6264);
nor U7982 (N_7982,N_6202,N_6911);
and U7983 (N_7983,N_6962,N_6456);
nor U7984 (N_7984,N_6428,N_6571);
and U7985 (N_7985,N_6643,N_6092);
and U7986 (N_7986,N_6017,N_6621);
and U7987 (N_7987,N_6876,N_6262);
xnor U7988 (N_7988,N_6213,N_6876);
nand U7989 (N_7989,N_6775,N_6721);
nand U7990 (N_7990,N_6259,N_6091);
nand U7991 (N_7991,N_6535,N_6363);
nand U7992 (N_7992,N_6632,N_6391);
nor U7993 (N_7993,N_6122,N_6192);
nor U7994 (N_7994,N_6943,N_6698);
or U7995 (N_7995,N_6421,N_6249);
nor U7996 (N_7996,N_6416,N_6891);
nand U7997 (N_7997,N_6924,N_6452);
xnor U7998 (N_7998,N_6456,N_6132);
or U7999 (N_7999,N_6512,N_6211);
or U8000 (N_8000,N_7322,N_7949);
nand U8001 (N_8001,N_7639,N_7951);
nand U8002 (N_8002,N_7017,N_7994);
or U8003 (N_8003,N_7962,N_7769);
nor U8004 (N_8004,N_7521,N_7021);
xnor U8005 (N_8005,N_7064,N_7016);
and U8006 (N_8006,N_7301,N_7798);
nand U8007 (N_8007,N_7065,N_7572);
and U8008 (N_8008,N_7472,N_7445);
nand U8009 (N_8009,N_7265,N_7595);
nor U8010 (N_8010,N_7508,N_7709);
xnor U8011 (N_8011,N_7050,N_7434);
xor U8012 (N_8012,N_7402,N_7598);
nor U8013 (N_8013,N_7297,N_7259);
nand U8014 (N_8014,N_7840,N_7924);
and U8015 (N_8015,N_7992,N_7466);
or U8016 (N_8016,N_7929,N_7523);
or U8017 (N_8017,N_7602,N_7827);
xnor U8018 (N_8018,N_7770,N_7063);
nor U8019 (N_8019,N_7309,N_7708);
and U8020 (N_8020,N_7323,N_7990);
and U8021 (N_8021,N_7348,N_7435);
or U8022 (N_8022,N_7078,N_7055);
or U8023 (N_8023,N_7652,N_7889);
nand U8024 (N_8024,N_7628,N_7220);
nor U8025 (N_8025,N_7554,N_7496);
nor U8026 (N_8026,N_7288,N_7387);
and U8027 (N_8027,N_7395,N_7796);
nor U8028 (N_8028,N_7237,N_7773);
and U8029 (N_8029,N_7275,N_7597);
nor U8030 (N_8030,N_7742,N_7933);
xnor U8031 (N_8031,N_7683,N_7306);
and U8032 (N_8032,N_7056,N_7191);
xnor U8033 (N_8033,N_7745,N_7583);
or U8034 (N_8034,N_7379,N_7541);
nand U8035 (N_8035,N_7299,N_7406);
xnor U8036 (N_8036,N_7231,N_7932);
and U8037 (N_8037,N_7083,N_7669);
nor U8038 (N_8038,N_7898,N_7548);
or U8039 (N_8039,N_7151,N_7535);
or U8040 (N_8040,N_7824,N_7490);
xor U8041 (N_8041,N_7673,N_7945);
nor U8042 (N_8042,N_7678,N_7650);
nor U8043 (N_8043,N_7319,N_7431);
nand U8044 (N_8044,N_7833,N_7041);
nor U8045 (N_8045,N_7978,N_7640);
and U8046 (N_8046,N_7218,N_7117);
nand U8047 (N_8047,N_7426,N_7555);
and U8048 (N_8048,N_7152,N_7953);
nor U8049 (N_8049,N_7396,N_7410);
nand U8050 (N_8050,N_7080,N_7736);
and U8051 (N_8051,N_7852,N_7760);
nor U8052 (N_8052,N_7418,N_7748);
and U8053 (N_8053,N_7140,N_7293);
nand U8054 (N_8054,N_7251,N_7329);
or U8055 (N_8055,N_7966,N_7529);
nor U8056 (N_8056,N_7776,N_7453);
nand U8057 (N_8057,N_7812,N_7473);
and U8058 (N_8058,N_7834,N_7592);
or U8059 (N_8059,N_7458,N_7260);
or U8060 (N_8060,N_7757,N_7782);
and U8061 (N_8061,N_7278,N_7113);
and U8062 (N_8062,N_7412,N_7980);
xor U8063 (N_8063,N_7003,N_7871);
nand U8064 (N_8064,N_7882,N_7741);
nor U8065 (N_8065,N_7784,N_7333);
nor U8066 (N_8066,N_7921,N_7764);
nand U8067 (N_8067,N_7486,N_7235);
or U8068 (N_8068,N_7034,N_7934);
nand U8069 (N_8069,N_7906,N_7802);
nand U8070 (N_8070,N_7897,N_7352);
or U8071 (N_8071,N_7847,N_7677);
nor U8072 (N_8072,N_7522,N_7343);
and U8073 (N_8073,N_7586,N_7858);
and U8074 (N_8074,N_7312,N_7607);
or U8075 (N_8075,N_7698,N_7681);
nor U8076 (N_8076,N_7032,N_7038);
nand U8077 (N_8077,N_7591,N_7877);
nor U8078 (N_8078,N_7706,N_7112);
or U8079 (N_8079,N_7720,N_7403);
nor U8080 (N_8080,N_7285,N_7666);
xor U8081 (N_8081,N_7066,N_7984);
or U8082 (N_8082,N_7327,N_7242);
nor U8083 (N_8083,N_7208,N_7726);
nor U8084 (N_8084,N_7665,N_7226);
nand U8085 (N_8085,N_7539,N_7713);
nor U8086 (N_8086,N_7731,N_7828);
nand U8087 (N_8087,N_7605,N_7927);
xor U8088 (N_8088,N_7789,N_7613);
or U8089 (N_8089,N_7059,N_7289);
or U8090 (N_8090,N_7389,N_7623);
and U8091 (N_8091,N_7023,N_7479);
nand U8092 (N_8092,N_7717,N_7991);
nor U8093 (N_8093,N_7097,N_7621);
nand U8094 (N_8094,N_7475,N_7918);
xnor U8095 (N_8095,N_7361,N_7845);
nor U8096 (N_8096,N_7631,N_7230);
and U8097 (N_8097,N_7714,N_7753);
xor U8098 (N_8098,N_7244,N_7452);
nand U8099 (N_8099,N_7855,N_7502);
and U8100 (N_8100,N_7779,N_7813);
nand U8101 (N_8101,N_7762,N_7162);
xnor U8102 (N_8102,N_7822,N_7200);
and U8103 (N_8103,N_7353,N_7675);
xnor U8104 (N_8104,N_7381,N_7965);
or U8105 (N_8105,N_7946,N_7691);
nand U8106 (N_8106,N_7892,N_7792);
nand U8107 (N_8107,N_7635,N_7136);
nor U8108 (N_8108,N_7212,N_7817);
or U8109 (N_8109,N_7545,N_7421);
nand U8110 (N_8110,N_7380,N_7103);
nand U8111 (N_8111,N_7729,N_7108);
nand U8112 (N_8112,N_7931,N_7443);
or U8113 (N_8113,N_7517,N_7245);
nand U8114 (N_8114,N_7912,N_7777);
and U8115 (N_8115,N_7718,N_7193);
nand U8116 (N_8116,N_7414,N_7542);
or U8117 (N_8117,N_7254,N_7077);
and U8118 (N_8118,N_7916,N_7975);
nand U8119 (N_8119,N_7651,N_7759);
nand U8120 (N_8120,N_7331,N_7186);
or U8121 (N_8121,N_7207,N_7600);
or U8122 (N_8122,N_7175,N_7154);
nand U8123 (N_8123,N_7612,N_7314);
nand U8124 (N_8124,N_7087,N_7001);
or U8125 (N_8125,N_7483,N_7660);
or U8126 (N_8126,N_7095,N_7608);
or U8127 (N_8127,N_7981,N_7560);
nand U8128 (N_8128,N_7205,N_7375);
nand U8129 (N_8129,N_7716,N_7819);
and U8130 (N_8130,N_7227,N_7470);
nor U8131 (N_8131,N_7754,N_7866);
nand U8132 (N_8132,N_7659,N_7843);
or U8133 (N_8133,N_7519,N_7494);
or U8134 (N_8134,N_7724,N_7126);
xnor U8135 (N_8135,N_7577,N_7030);
nor U8136 (N_8136,N_7766,N_7197);
nor U8137 (N_8137,N_7585,N_7328);
and U8138 (N_8138,N_7463,N_7184);
nor U8139 (N_8139,N_7619,N_7841);
nand U8140 (N_8140,N_7336,N_7446);
nor U8141 (N_8141,N_7895,N_7582);
nor U8142 (N_8142,N_7570,N_7401);
xor U8143 (N_8143,N_7450,N_7310);
nor U8144 (N_8144,N_7225,N_7068);
xnor U8145 (N_8145,N_7250,N_7477);
nor U8146 (N_8146,N_7524,N_7642);
nand U8147 (N_8147,N_7223,N_7124);
nand U8148 (N_8148,N_7861,N_7498);
nand U8149 (N_8149,N_7354,N_7697);
or U8150 (N_8150,N_7940,N_7509);
or U8151 (N_8151,N_7578,N_7537);
nor U8152 (N_8152,N_7143,N_7057);
nand U8153 (N_8153,N_7604,N_7547);
xnor U8154 (N_8154,N_7376,N_7688);
or U8155 (N_8155,N_7211,N_7388);
nor U8156 (N_8156,N_7132,N_7177);
or U8157 (N_8157,N_7657,N_7100);
or U8158 (N_8158,N_7772,N_7611);
and U8159 (N_8159,N_7625,N_7090);
nand U8160 (N_8160,N_7295,N_7526);
or U8161 (N_8161,N_7894,N_7195);
nand U8162 (N_8162,N_7025,N_7181);
nand U8163 (N_8163,N_7674,N_7262);
and U8164 (N_8164,N_7854,N_7165);
xor U8165 (N_8165,N_7734,N_7829);
nor U8166 (N_8166,N_7864,N_7495);
nor U8167 (N_8167,N_7385,N_7000);
nor U8168 (N_8168,N_7010,N_7174);
xor U8169 (N_8169,N_7944,N_7727);
and U8170 (N_8170,N_7672,N_7499);
and U8171 (N_8171,N_7648,N_7298);
xor U8172 (N_8172,N_7093,N_7455);
nand U8173 (N_8173,N_7420,N_7169);
nor U8174 (N_8174,N_7964,N_7974);
nand U8175 (N_8175,N_7115,N_7166);
and U8176 (N_8176,N_7071,N_7255);
nor U8177 (N_8177,N_7249,N_7007);
xnor U8178 (N_8178,N_7771,N_7922);
nand U8179 (N_8179,N_7042,N_7082);
nand U8180 (N_8180,N_7930,N_7416);
or U8181 (N_8181,N_7860,N_7950);
and U8182 (N_8182,N_7576,N_7755);
xnor U8183 (N_8183,N_7735,N_7024);
nand U8184 (N_8184,N_7324,N_7890);
or U8185 (N_8185,N_7948,N_7926);
nor U8186 (N_8186,N_7656,N_7638);
nand U8187 (N_8187,N_7317,N_7969);
and U8188 (N_8188,N_7270,N_7682);
nand U8189 (N_8189,N_7601,N_7913);
xor U8190 (N_8190,N_7842,N_7531);
nor U8191 (N_8191,N_7500,N_7559);
or U8192 (N_8192,N_7125,N_7196);
and U8193 (N_8193,N_7334,N_7456);
nand U8194 (N_8194,N_7147,N_7012);
or U8195 (N_8195,N_7355,N_7911);
and U8196 (N_8196,N_7627,N_7510);
and U8197 (N_8197,N_7616,N_7359);
or U8198 (N_8198,N_7590,N_7234);
and U8199 (N_8199,N_7955,N_7337);
or U8200 (N_8200,N_7549,N_7422);
nor U8201 (N_8201,N_7763,N_7002);
nand U8202 (N_8202,N_7960,N_7091);
and U8203 (N_8203,N_7814,N_7867);
nor U8204 (N_8204,N_7561,N_7914);
nand U8205 (N_8205,N_7971,N_7935);
xor U8206 (N_8206,N_7344,N_7037);
nor U8207 (N_8207,N_7179,N_7869);
nand U8208 (N_8208,N_7409,N_7504);
and U8209 (N_8209,N_7051,N_7909);
and U8210 (N_8210,N_7340,N_7893);
nor U8211 (N_8211,N_7768,N_7680);
and U8212 (N_8212,N_7345,N_7111);
nor U8213 (N_8213,N_7272,N_7655);
and U8214 (N_8214,N_7138,N_7367);
xnor U8215 (N_8215,N_7743,N_7269);
or U8216 (N_8216,N_7120,N_7332);
and U8217 (N_8217,N_7865,N_7139);
and U8218 (N_8218,N_7228,N_7941);
and U8219 (N_8219,N_7313,N_7569);
nor U8220 (N_8220,N_7121,N_7905);
nand U8221 (N_8221,N_7690,N_7505);
nand U8222 (N_8222,N_7214,N_7687);
nand U8223 (N_8223,N_7807,N_7923);
and U8224 (N_8224,N_7471,N_7316);
nand U8225 (N_8225,N_7821,N_7788);
nor U8226 (N_8226,N_7527,N_7074);
and U8227 (N_8227,N_7398,N_7543);
xnor U8228 (N_8228,N_7052,N_7610);
and U8229 (N_8229,N_7979,N_7280);
or U8230 (N_8230,N_7116,N_7982);
and U8231 (N_8231,N_7808,N_7127);
or U8232 (N_8232,N_7844,N_7694);
and U8233 (N_8233,N_7049,N_7469);
or U8234 (N_8234,N_7099,N_7746);
nor U8235 (N_8235,N_7967,N_7263);
and U8236 (N_8236,N_7029,N_7315);
and U8237 (N_8237,N_7624,N_7973);
nor U8238 (N_8238,N_7054,N_7062);
xnor U8239 (N_8239,N_7781,N_7036);
and U8240 (N_8240,N_7557,N_7928);
or U8241 (N_8241,N_7141,N_7378);
and U8242 (N_8242,N_7031,N_7185);
or U8243 (N_8243,N_7558,N_7837);
nor U8244 (N_8244,N_7404,N_7160);
or U8245 (N_8245,N_7119,N_7210);
and U8246 (N_8246,N_7791,N_7904);
nor U8247 (N_8247,N_7252,N_7073);
and U8248 (N_8248,N_7287,N_7851);
nor U8249 (N_8249,N_7663,N_7647);
nand U8250 (N_8250,N_7849,N_7302);
nand U8251 (N_8251,N_7530,N_7303);
and U8252 (N_8252,N_7863,N_7008);
xnor U8253 (N_8253,N_7723,N_7581);
nor U8254 (N_8254,N_7146,N_7887);
nand U8255 (N_8255,N_7831,N_7085);
and U8256 (N_8256,N_7879,N_7474);
xor U8257 (N_8257,N_7862,N_7571);
or U8258 (N_8258,N_7325,N_7711);
xor U8259 (N_8259,N_7256,N_7544);
xor U8260 (N_8260,N_7615,N_7240);
nand U8261 (N_8261,N_7579,N_7465);
nand U8262 (N_8262,N_7084,N_7968);
nor U8263 (N_8263,N_7460,N_7556);
nand U8264 (N_8264,N_7067,N_7538);
xor U8265 (N_8265,N_7342,N_7751);
and U8266 (N_8266,N_7804,N_7761);
nand U8267 (N_8267,N_7506,N_7920);
nand U8268 (N_8268,N_7492,N_7149);
xor U8269 (N_8269,N_7487,N_7565);
nand U8270 (N_8270,N_7999,N_7489);
xor U8271 (N_8271,N_7229,N_7820);
nor U8272 (N_8272,N_7187,N_7109);
xnor U8273 (N_8273,N_7366,N_7907);
and U8274 (N_8274,N_7518,N_7338);
and U8275 (N_8275,N_7171,N_7462);
or U8276 (N_8276,N_7296,N_7936);
nor U8277 (N_8277,N_7917,N_7850);
nor U8278 (N_8278,N_7566,N_7370);
nor U8279 (N_8279,N_7159,N_7995);
xnor U8280 (N_8280,N_7956,N_7341);
and U8281 (N_8281,N_7092,N_7192);
or U8282 (N_8282,N_7550,N_7070);
nand U8283 (N_8283,N_7176,N_7189);
and U8284 (N_8284,N_7069,N_7374);
nor U8285 (N_8285,N_7428,N_7636);
nand U8286 (N_8286,N_7730,N_7400);
nand U8287 (N_8287,N_7253,N_7292);
and U8288 (N_8288,N_7134,N_7805);
or U8289 (N_8289,N_7880,N_7747);
xnor U8290 (N_8290,N_7977,N_7397);
nand U8291 (N_8291,N_7876,N_7279);
nor U8292 (N_8292,N_7096,N_7019);
xor U8293 (N_8293,N_7178,N_7075);
xor U8294 (N_8294,N_7986,N_7204);
and U8295 (N_8295,N_7365,N_7721);
nand U8296 (N_8296,N_7157,N_7028);
or U8297 (N_8297,N_7161,N_7006);
nor U8298 (N_8298,N_7238,N_7998);
nand U8299 (N_8299,N_7321,N_7908);
nand U8300 (N_8300,N_7511,N_7167);
nand U8301 (N_8301,N_7649,N_7993);
or U8302 (N_8302,N_7142,N_7732);
xor U8303 (N_8303,N_7394,N_7744);
and U8304 (N_8304,N_7749,N_7386);
or U8305 (N_8305,N_7305,N_7653);
xnor U8306 (N_8306,N_7358,N_7806);
or U8307 (N_8307,N_7679,N_7009);
and U8308 (N_8308,N_7294,N_7015);
nand U8309 (N_8309,N_7221,N_7739);
and U8310 (N_8310,N_7122,N_7795);
and U8311 (N_8311,N_7183,N_7020);
nand U8312 (N_8312,N_7430,N_7444);
and U8313 (N_8313,N_7290,N_7970);
nor U8314 (N_8314,N_7939,N_7481);
nand U8315 (N_8315,N_7419,N_7818);
or U8316 (N_8316,N_7988,N_7780);
nand U8317 (N_8317,N_7372,N_7670);
nand U8318 (N_8318,N_7765,N_7239);
and U8319 (N_8319,N_7201,N_7552);
or U8320 (N_8320,N_7079,N_7058);
nand U8321 (N_8321,N_7282,N_7035);
nand U8322 (N_8322,N_7232,N_7740);
nor U8323 (N_8323,N_7872,N_7133);
nor U8324 (N_8324,N_7213,N_7696);
nand U8325 (N_8325,N_7098,N_7704);
nand U8326 (N_8326,N_7947,N_7130);
or U8327 (N_8327,N_7589,N_7884);
and U8328 (N_8328,N_7567,N_7883);
nand U8329 (N_8329,N_7150,N_7432);
nand U8330 (N_8330,N_7281,N_7826);
or U8331 (N_8331,N_7300,N_7040);
nor U8332 (N_8332,N_7241,N_7026);
and U8333 (N_8333,N_7686,N_7836);
nor U8334 (N_8334,N_7362,N_7144);
nor U8335 (N_8335,N_7188,N_7942);
and U8336 (N_8336,N_7919,N_7667);
and U8337 (N_8337,N_7902,N_7573);
and U8338 (N_8338,N_7137,N_7107);
or U8339 (N_8339,N_7209,N_7580);
and U8340 (N_8340,N_7832,N_7658);
nand U8341 (N_8341,N_7086,N_7039);
nor U8342 (N_8342,N_7369,N_7702);
and U8343 (N_8343,N_7901,N_7447);
nand U8344 (N_8344,N_7163,N_7417);
and U8345 (N_8345,N_7507,N_7047);
nand U8346 (N_8346,N_7158,N_7614);
nand U8347 (N_8347,N_7425,N_7712);
nand U8348 (N_8348,N_7393,N_7399);
nor U8349 (N_8349,N_7004,N_7534);
or U8350 (N_8350,N_7785,N_7013);
nor U8351 (N_8351,N_7439,N_7596);
nand U8352 (N_8352,N_7963,N_7110);
xnor U8353 (N_8353,N_7273,N_7533);
nor U8354 (N_8354,N_7692,N_7794);
xnor U8355 (N_8355,N_7118,N_7493);
nor U8356 (N_8356,N_7816,N_7258);
nor U8357 (N_8357,N_7643,N_7170);
nand U8358 (N_8358,N_7043,N_7457);
xnor U8359 (N_8359,N_7335,N_7484);
xor U8360 (N_8360,N_7587,N_7985);
and U8361 (N_8361,N_7875,N_7634);
nand U8362 (N_8362,N_7976,N_7476);
nor U8363 (N_8363,N_7349,N_7276);
or U8364 (N_8364,N_7286,N_7801);
and U8365 (N_8365,N_7206,N_7436);
nand U8366 (N_8366,N_7793,N_7046);
nand U8367 (N_8367,N_7266,N_7383);
xor U8368 (N_8368,N_7027,N_7856);
and U8369 (N_8369,N_7180,N_7488);
and U8370 (N_8370,N_7267,N_7937);
nor U8371 (N_8371,N_7996,N_7553);
or U8372 (N_8372,N_7878,N_7684);
and U8373 (N_8373,N_7224,N_7903);
nand U8374 (N_8374,N_7705,N_7609);
nor U8375 (N_8375,N_7815,N_7528);
and U8376 (N_8376,N_7899,N_7076);
nand U8377 (N_8377,N_7954,N_7629);
and U8378 (N_8378,N_7800,N_7148);
nand U8379 (N_8379,N_7440,N_7584);
nand U8380 (N_8380,N_7128,N_7859);
nor U8381 (N_8381,N_7774,N_7390);
or U8382 (N_8382,N_7733,N_7786);
nor U8383 (N_8383,N_7599,N_7664);
xnor U8384 (N_8384,N_7646,N_7671);
or U8385 (N_8385,N_7215,N_7236);
and U8386 (N_8386,N_7373,N_7464);
or U8387 (N_8387,N_7449,N_7459);
nor U8388 (N_8388,N_7896,N_7501);
or U8389 (N_8389,N_7536,N_7448);
and U8390 (N_8390,N_7233,N_7797);
and U8391 (N_8391,N_7405,N_7392);
nor U8392 (N_8392,N_7825,N_7513);
and U8393 (N_8393,N_7810,N_7377);
nand U8394 (N_8394,N_7088,N_7881);
nand U8395 (N_8395,N_7482,N_7364);
or U8396 (N_8396,N_7384,N_7198);
and U8397 (N_8397,N_7268,N_7018);
nor U8398 (N_8398,N_7952,N_7532);
nand U8399 (N_8399,N_7594,N_7514);
or U8400 (N_8400,N_7283,N_7438);
or U8401 (N_8401,N_7168,N_7958);
xor U8402 (N_8402,N_7216,N_7371);
nand U8403 (N_8403,N_7617,N_7943);
or U8404 (N_8404,N_7676,N_7005);
and U8405 (N_8405,N_7997,N_7710);
and U8406 (N_8406,N_7645,N_7382);
nor U8407 (N_8407,N_7853,N_7131);
or U8408 (N_8408,N_7407,N_7308);
nor U8409 (N_8409,N_7222,N_7756);
or U8410 (N_8410,N_7467,N_7105);
or U8411 (N_8411,N_7830,N_7106);
and U8412 (N_8412,N_7846,N_7516);
nor U8413 (N_8413,N_7081,N_7715);
nor U8414 (N_8414,N_7891,N_7987);
or U8415 (N_8415,N_7520,N_7622);
nor U8416 (N_8416,N_7767,N_7790);
nor U8417 (N_8417,N_7357,N_7102);
and U8418 (N_8418,N_7783,N_7699);
nor U8419 (N_8419,N_7423,N_7938);
nand U8420 (N_8420,N_7060,N_7722);
xnor U8421 (N_8421,N_7022,N_7391);
xnor U8422 (N_8422,N_7045,N_7546);
xor U8423 (N_8423,N_7989,N_7194);
or U8424 (N_8424,N_7155,N_7114);
nand U8425 (N_8425,N_7424,N_7202);
nand U8426 (N_8426,N_7330,N_7503);
nor U8427 (N_8427,N_7261,N_7351);
nor U8428 (N_8428,N_7011,N_7568);
and U8429 (N_8429,N_7983,N_7874);
xnor U8430 (N_8430,N_7641,N_7562);
and U8431 (N_8431,N_7803,N_7632);
or U8432 (N_8432,N_7491,N_7247);
nand U8433 (N_8433,N_7700,N_7811);
or U8434 (N_8434,N_7606,N_7701);
or U8435 (N_8435,N_7129,N_7787);
nor U8436 (N_8436,N_7123,N_7274);
nor U8437 (N_8437,N_7725,N_7429);
nor U8438 (N_8438,N_7512,N_7662);
nand U8439 (N_8439,N_7689,N_7630);
or U8440 (N_8440,N_7307,N_7101);
and U8441 (N_8441,N_7441,N_7618);
nand U8442 (N_8442,N_7551,N_7173);
xor U8443 (N_8443,N_7360,N_7271);
nand U8444 (N_8444,N_7728,N_7593);
and U8445 (N_8445,N_7693,N_7053);
xnor U8446 (N_8446,N_7437,N_7750);
or U8447 (N_8447,N_7873,N_7048);
nor U8448 (N_8448,N_7442,N_7304);
nor U8449 (N_8449,N_7809,N_7823);
and U8450 (N_8450,N_7915,N_7661);
nand U8451 (N_8451,N_7540,N_7094);
xor U8452 (N_8452,N_7775,N_7644);
or U8453 (N_8453,N_7277,N_7654);
and U8454 (N_8454,N_7468,N_7243);
nand U8455 (N_8455,N_7014,N_7668);
and U8456 (N_8456,N_7415,N_7199);
and U8457 (N_8457,N_7707,N_7203);
nand U8458 (N_8458,N_7145,N_7326);
nor U8459 (N_8459,N_7413,N_7888);
nand U8460 (N_8460,N_7284,N_7311);
xor U8461 (N_8461,N_7190,N_7972);
and U8462 (N_8462,N_7172,N_7156);
xnor U8463 (N_8463,N_7320,N_7219);
and U8464 (N_8464,N_7838,N_7427);
or U8465 (N_8465,N_7703,N_7291);
and U8466 (N_8466,N_7497,N_7044);
nand U8467 (N_8467,N_7835,N_7870);
and U8468 (N_8468,N_7574,N_7563);
xor U8469 (N_8469,N_7695,N_7339);
and U8470 (N_8470,N_7356,N_7478);
nand U8471 (N_8471,N_7182,N_7164);
nor U8472 (N_8472,N_7719,N_7153);
nor U8473 (N_8473,N_7433,N_7368);
nor U8474 (N_8474,N_7217,N_7868);
nand U8475 (N_8475,N_7525,N_7839);
nor U8476 (N_8476,N_7485,N_7104);
nor U8477 (N_8477,N_7885,N_7461);
or U8478 (N_8478,N_7347,N_7061);
nand U8479 (N_8479,N_7248,N_7633);
nor U8480 (N_8480,N_7318,N_7959);
or U8481 (N_8481,N_7515,N_7454);
nand U8482 (N_8482,N_7363,N_7886);
nand U8483 (N_8483,N_7564,N_7072);
and U8484 (N_8484,N_7961,N_7778);
or U8485 (N_8485,N_7089,N_7857);
nand U8486 (N_8486,N_7799,N_7737);
or U8487 (N_8487,N_7350,N_7264);
and U8488 (N_8488,N_7758,N_7910);
xor U8489 (N_8489,N_7588,N_7738);
nand U8490 (N_8490,N_7346,N_7033);
nor U8491 (N_8491,N_7575,N_7752);
or U8492 (N_8492,N_7257,N_7620);
nor U8493 (N_8493,N_7848,N_7626);
nand U8494 (N_8494,N_7451,N_7685);
or U8495 (N_8495,N_7900,N_7411);
or U8496 (N_8496,N_7135,N_7246);
nor U8497 (N_8497,N_7603,N_7637);
and U8498 (N_8498,N_7925,N_7480);
nand U8499 (N_8499,N_7957,N_7408);
xnor U8500 (N_8500,N_7518,N_7427);
nor U8501 (N_8501,N_7731,N_7299);
nand U8502 (N_8502,N_7277,N_7241);
xnor U8503 (N_8503,N_7882,N_7641);
and U8504 (N_8504,N_7277,N_7934);
and U8505 (N_8505,N_7861,N_7500);
nor U8506 (N_8506,N_7420,N_7886);
nor U8507 (N_8507,N_7359,N_7360);
or U8508 (N_8508,N_7406,N_7588);
nor U8509 (N_8509,N_7688,N_7801);
or U8510 (N_8510,N_7118,N_7175);
or U8511 (N_8511,N_7747,N_7380);
or U8512 (N_8512,N_7748,N_7853);
nand U8513 (N_8513,N_7314,N_7404);
nand U8514 (N_8514,N_7767,N_7922);
or U8515 (N_8515,N_7412,N_7758);
nand U8516 (N_8516,N_7757,N_7206);
nor U8517 (N_8517,N_7997,N_7260);
nor U8518 (N_8518,N_7104,N_7209);
or U8519 (N_8519,N_7859,N_7632);
xor U8520 (N_8520,N_7114,N_7996);
or U8521 (N_8521,N_7586,N_7791);
nand U8522 (N_8522,N_7335,N_7245);
and U8523 (N_8523,N_7719,N_7564);
nand U8524 (N_8524,N_7948,N_7958);
and U8525 (N_8525,N_7140,N_7475);
xnor U8526 (N_8526,N_7766,N_7607);
and U8527 (N_8527,N_7307,N_7574);
and U8528 (N_8528,N_7853,N_7229);
or U8529 (N_8529,N_7816,N_7508);
or U8530 (N_8530,N_7308,N_7699);
xnor U8531 (N_8531,N_7376,N_7398);
nand U8532 (N_8532,N_7570,N_7954);
and U8533 (N_8533,N_7061,N_7025);
or U8534 (N_8534,N_7999,N_7996);
nor U8535 (N_8535,N_7776,N_7465);
nand U8536 (N_8536,N_7878,N_7706);
or U8537 (N_8537,N_7821,N_7104);
nor U8538 (N_8538,N_7964,N_7168);
and U8539 (N_8539,N_7584,N_7359);
nand U8540 (N_8540,N_7545,N_7887);
or U8541 (N_8541,N_7401,N_7142);
or U8542 (N_8542,N_7997,N_7740);
or U8543 (N_8543,N_7682,N_7794);
or U8544 (N_8544,N_7470,N_7084);
nand U8545 (N_8545,N_7061,N_7096);
and U8546 (N_8546,N_7619,N_7251);
nor U8547 (N_8547,N_7370,N_7310);
nor U8548 (N_8548,N_7818,N_7563);
or U8549 (N_8549,N_7698,N_7847);
xnor U8550 (N_8550,N_7356,N_7016);
or U8551 (N_8551,N_7055,N_7666);
nand U8552 (N_8552,N_7298,N_7487);
or U8553 (N_8553,N_7410,N_7676);
or U8554 (N_8554,N_7928,N_7197);
or U8555 (N_8555,N_7728,N_7837);
or U8556 (N_8556,N_7005,N_7122);
nand U8557 (N_8557,N_7131,N_7065);
nand U8558 (N_8558,N_7276,N_7368);
and U8559 (N_8559,N_7128,N_7785);
nand U8560 (N_8560,N_7996,N_7803);
nor U8561 (N_8561,N_7348,N_7402);
and U8562 (N_8562,N_7239,N_7180);
or U8563 (N_8563,N_7566,N_7721);
and U8564 (N_8564,N_7166,N_7643);
nor U8565 (N_8565,N_7649,N_7083);
nand U8566 (N_8566,N_7593,N_7326);
or U8567 (N_8567,N_7408,N_7620);
nor U8568 (N_8568,N_7368,N_7490);
and U8569 (N_8569,N_7716,N_7732);
nor U8570 (N_8570,N_7790,N_7862);
or U8571 (N_8571,N_7489,N_7388);
nor U8572 (N_8572,N_7881,N_7754);
and U8573 (N_8573,N_7404,N_7622);
and U8574 (N_8574,N_7600,N_7954);
or U8575 (N_8575,N_7419,N_7402);
or U8576 (N_8576,N_7284,N_7027);
nor U8577 (N_8577,N_7993,N_7997);
nand U8578 (N_8578,N_7196,N_7981);
and U8579 (N_8579,N_7090,N_7716);
nor U8580 (N_8580,N_7225,N_7658);
or U8581 (N_8581,N_7236,N_7121);
or U8582 (N_8582,N_7614,N_7309);
or U8583 (N_8583,N_7327,N_7281);
xnor U8584 (N_8584,N_7061,N_7927);
or U8585 (N_8585,N_7423,N_7217);
nor U8586 (N_8586,N_7359,N_7296);
nor U8587 (N_8587,N_7410,N_7471);
nor U8588 (N_8588,N_7371,N_7642);
nor U8589 (N_8589,N_7914,N_7664);
nor U8590 (N_8590,N_7385,N_7497);
and U8591 (N_8591,N_7050,N_7482);
nor U8592 (N_8592,N_7251,N_7117);
or U8593 (N_8593,N_7751,N_7626);
nor U8594 (N_8594,N_7720,N_7780);
nor U8595 (N_8595,N_7935,N_7166);
xnor U8596 (N_8596,N_7648,N_7120);
xnor U8597 (N_8597,N_7993,N_7782);
or U8598 (N_8598,N_7200,N_7164);
nand U8599 (N_8599,N_7790,N_7623);
nor U8600 (N_8600,N_7674,N_7337);
nor U8601 (N_8601,N_7430,N_7487);
nor U8602 (N_8602,N_7680,N_7723);
nand U8603 (N_8603,N_7223,N_7034);
nor U8604 (N_8604,N_7519,N_7475);
or U8605 (N_8605,N_7439,N_7052);
and U8606 (N_8606,N_7855,N_7877);
nor U8607 (N_8607,N_7240,N_7481);
nor U8608 (N_8608,N_7947,N_7805);
nor U8609 (N_8609,N_7677,N_7873);
or U8610 (N_8610,N_7590,N_7849);
nor U8611 (N_8611,N_7732,N_7330);
and U8612 (N_8612,N_7973,N_7440);
nor U8613 (N_8613,N_7901,N_7330);
nand U8614 (N_8614,N_7995,N_7542);
or U8615 (N_8615,N_7854,N_7052);
nor U8616 (N_8616,N_7474,N_7548);
or U8617 (N_8617,N_7370,N_7974);
nor U8618 (N_8618,N_7564,N_7053);
nand U8619 (N_8619,N_7134,N_7631);
and U8620 (N_8620,N_7835,N_7360);
nor U8621 (N_8621,N_7024,N_7653);
and U8622 (N_8622,N_7107,N_7165);
nand U8623 (N_8623,N_7446,N_7783);
and U8624 (N_8624,N_7959,N_7495);
nand U8625 (N_8625,N_7768,N_7682);
nand U8626 (N_8626,N_7484,N_7917);
nor U8627 (N_8627,N_7774,N_7615);
nor U8628 (N_8628,N_7804,N_7011);
nand U8629 (N_8629,N_7308,N_7710);
xnor U8630 (N_8630,N_7640,N_7966);
xnor U8631 (N_8631,N_7041,N_7609);
and U8632 (N_8632,N_7310,N_7920);
nand U8633 (N_8633,N_7974,N_7160);
and U8634 (N_8634,N_7977,N_7678);
or U8635 (N_8635,N_7354,N_7178);
nor U8636 (N_8636,N_7061,N_7976);
and U8637 (N_8637,N_7560,N_7002);
nand U8638 (N_8638,N_7293,N_7569);
and U8639 (N_8639,N_7619,N_7495);
xor U8640 (N_8640,N_7550,N_7475);
and U8641 (N_8641,N_7539,N_7570);
or U8642 (N_8642,N_7438,N_7298);
and U8643 (N_8643,N_7152,N_7818);
and U8644 (N_8644,N_7440,N_7434);
xor U8645 (N_8645,N_7457,N_7488);
nand U8646 (N_8646,N_7418,N_7383);
and U8647 (N_8647,N_7191,N_7505);
and U8648 (N_8648,N_7797,N_7077);
or U8649 (N_8649,N_7221,N_7297);
nand U8650 (N_8650,N_7375,N_7597);
or U8651 (N_8651,N_7075,N_7354);
nand U8652 (N_8652,N_7129,N_7144);
nor U8653 (N_8653,N_7626,N_7142);
or U8654 (N_8654,N_7146,N_7024);
or U8655 (N_8655,N_7142,N_7640);
nor U8656 (N_8656,N_7844,N_7148);
nor U8657 (N_8657,N_7003,N_7952);
nor U8658 (N_8658,N_7246,N_7767);
nand U8659 (N_8659,N_7560,N_7063);
nor U8660 (N_8660,N_7313,N_7225);
and U8661 (N_8661,N_7448,N_7855);
nor U8662 (N_8662,N_7155,N_7819);
nor U8663 (N_8663,N_7562,N_7245);
and U8664 (N_8664,N_7107,N_7045);
nand U8665 (N_8665,N_7395,N_7136);
and U8666 (N_8666,N_7266,N_7711);
nor U8667 (N_8667,N_7795,N_7371);
or U8668 (N_8668,N_7655,N_7819);
nand U8669 (N_8669,N_7631,N_7216);
or U8670 (N_8670,N_7310,N_7327);
or U8671 (N_8671,N_7351,N_7181);
nor U8672 (N_8672,N_7173,N_7235);
or U8673 (N_8673,N_7668,N_7005);
and U8674 (N_8674,N_7830,N_7952);
nor U8675 (N_8675,N_7520,N_7923);
or U8676 (N_8676,N_7346,N_7046);
or U8677 (N_8677,N_7701,N_7799);
or U8678 (N_8678,N_7791,N_7671);
and U8679 (N_8679,N_7330,N_7905);
nand U8680 (N_8680,N_7168,N_7085);
and U8681 (N_8681,N_7791,N_7556);
nor U8682 (N_8682,N_7293,N_7900);
or U8683 (N_8683,N_7917,N_7671);
and U8684 (N_8684,N_7835,N_7033);
xnor U8685 (N_8685,N_7006,N_7875);
or U8686 (N_8686,N_7686,N_7458);
nand U8687 (N_8687,N_7345,N_7942);
xor U8688 (N_8688,N_7950,N_7889);
and U8689 (N_8689,N_7708,N_7052);
or U8690 (N_8690,N_7361,N_7585);
or U8691 (N_8691,N_7974,N_7496);
xnor U8692 (N_8692,N_7658,N_7520);
and U8693 (N_8693,N_7844,N_7583);
and U8694 (N_8694,N_7944,N_7062);
or U8695 (N_8695,N_7711,N_7721);
or U8696 (N_8696,N_7130,N_7064);
nor U8697 (N_8697,N_7214,N_7104);
nor U8698 (N_8698,N_7385,N_7370);
xor U8699 (N_8699,N_7845,N_7454);
and U8700 (N_8700,N_7380,N_7026);
nand U8701 (N_8701,N_7970,N_7991);
xnor U8702 (N_8702,N_7743,N_7200);
nand U8703 (N_8703,N_7857,N_7730);
nand U8704 (N_8704,N_7222,N_7500);
and U8705 (N_8705,N_7229,N_7137);
nor U8706 (N_8706,N_7134,N_7456);
xnor U8707 (N_8707,N_7386,N_7486);
nor U8708 (N_8708,N_7849,N_7869);
or U8709 (N_8709,N_7921,N_7272);
nor U8710 (N_8710,N_7196,N_7186);
or U8711 (N_8711,N_7599,N_7918);
nand U8712 (N_8712,N_7527,N_7110);
and U8713 (N_8713,N_7436,N_7211);
nand U8714 (N_8714,N_7010,N_7596);
or U8715 (N_8715,N_7766,N_7507);
nor U8716 (N_8716,N_7805,N_7461);
nor U8717 (N_8717,N_7166,N_7601);
nand U8718 (N_8718,N_7393,N_7229);
xnor U8719 (N_8719,N_7990,N_7236);
or U8720 (N_8720,N_7177,N_7811);
or U8721 (N_8721,N_7000,N_7350);
or U8722 (N_8722,N_7310,N_7893);
or U8723 (N_8723,N_7357,N_7955);
nor U8724 (N_8724,N_7056,N_7600);
and U8725 (N_8725,N_7221,N_7547);
and U8726 (N_8726,N_7158,N_7080);
or U8727 (N_8727,N_7488,N_7035);
xor U8728 (N_8728,N_7700,N_7575);
nor U8729 (N_8729,N_7939,N_7133);
nand U8730 (N_8730,N_7755,N_7222);
or U8731 (N_8731,N_7791,N_7107);
nand U8732 (N_8732,N_7129,N_7581);
nand U8733 (N_8733,N_7939,N_7271);
or U8734 (N_8734,N_7479,N_7308);
and U8735 (N_8735,N_7083,N_7276);
nor U8736 (N_8736,N_7007,N_7065);
and U8737 (N_8737,N_7477,N_7671);
or U8738 (N_8738,N_7122,N_7775);
and U8739 (N_8739,N_7759,N_7400);
nor U8740 (N_8740,N_7937,N_7292);
nor U8741 (N_8741,N_7612,N_7419);
or U8742 (N_8742,N_7508,N_7900);
and U8743 (N_8743,N_7949,N_7754);
and U8744 (N_8744,N_7288,N_7319);
or U8745 (N_8745,N_7376,N_7270);
xnor U8746 (N_8746,N_7353,N_7244);
nor U8747 (N_8747,N_7727,N_7811);
or U8748 (N_8748,N_7635,N_7794);
or U8749 (N_8749,N_7136,N_7843);
nor U8750 (N_8750,N_7492,N_7588);
or U8751 (N_8751,N_7787,N_7307);
nor U8752 (N_8752,N_7141,N_7603);
nor U8753 (N_8753,N_7463,N_7248);
and U8754 (N_8754,N_7509,N_7941);
or U8755 (N_8755,N_7305,N_7141);
or U8756 (N_8756,N_7554,N_7821);
nand U8757 (N_8757,N_7075,N_7141);
nor U8758 (N_8758,N_7612,N_7095);
nor U8759 (N_8759,N_7325,N_7189);
and U8760 (N_8760,N_7086,N_7403);
xor U8761 (N_8761,N_7059,N_7255);
or U8762 (N_8762,N_7639,N_7474);
nor U8763 (N_8763,N_7364,N_7526);
xor U8764 (N_8764,N_7051,N_7459);
xnor U8765 (N_8765,N_7835,N_7907);
or U8766 (N_8766,N_7269,N_7676);
nand U8767 (N_8767,N_7102,N_7218);
or U8768 (N_8768,N_7900,N_7850);
and U8769 (N_8769,N_7338,N_7266);
and U8770 (N_8770,N_7708,N_7096);
or U8771 (N_8771,N_7767,N_7415);
and U8772 (N_8772,N_7025,N_7035);
nand U8773 (N_8773,N_7355,N_7530);
nand U8774 (N_8774,N_7886,N_7858);
nand U8775 (N_8775,N_7685,N_7132);
xor U8776 (N_8776,N_7388,N_7095);
and U8777 (N_8777,N_7002,N_7105);
or U8778 (N_8778,N_7614,N_7658);
or U8779 (N_8779,N_7882,N_7306);
and U8780 (N_8780,N_7936,N_7760);
xnor U8781 (N_8781,N_7978,N_7975);
nand U8782 (N_8782,N_7250,N_7270);
nand U8783 (N_8783,N_7746,N_7065);
and U8784 (N_8784,N_7144,N_7600);
nor U8785 (N_8785,N_7852,N_7882);
nor U8786 (N_8786,N_7422,N_7194);
nor U8787 (N_8787,N_7695,N_7817);
and U8788 (N_8788,N_7514,N_7164);
and U8789 (N_8789,N_7472,N_7732);
and U8790 (N_8790,N_7704,N_7970);
nand U8791 (N_8791,N_7849,N_7096);
and U8792 (N_8792,N_7152,N_7199);
nor U8793 (N_8793,N_7716,N_7117);
xnor U8794 (N_8794,N_7026,N_7826);
nor U8795 (N_8795,N_7551,N_7216);
xor U8796 (N_8796,N_7456,N_7832);
nor U8797 (N_8797,N_7575,N_7321);
and U8798 (N_8798,N_7249,N_7998);
or U8799 (N_8799,N_7265,N_7661);
xnor U8800 (N_8800,N_7288,N_7909);
or U8801 (N_8801,N_7871,N_7541);
and U8802 (N_8802,N_7083,N_7262);
or U8803 (N_8803,N_7759,N_7054);
or U8804 (N_8804,N_7660,N_7028);
nand U8805 (N_8805,N_7250,N_7352);
or U8806 (N_8806,N_7265,N_7499);
or U8807 (N_8807,N_7189,N_7535);
nor U8808 (N_8808,N_7683,N_7455);
and U8809 (N_8809,N_7836,N_7848);
or U8810 (N_8810,N_7020,N_7311);
xnor U8811 (N_8811,N_7567,N_7037);
nand U8812 (N_8812,N_7216,N_7622);
xor U8813 (N_8813,N_7501,N_7078);
or U8814 (N_8814,N_7777,N_7405);
and U8815 (N_8815,N_7867,N_7556);
nor U8816 (N_8816,N_7003,N_7824);
nor U8817 (N_8817,N_7786,N_7111);
and U8818 (N_8818,N_7963,N_7427);
nand U8819 (N_8819,N_7323,N_7984);
nor U8820 (N_8820,N_7539,N_7778);
or U8821 (N_8821,N_7968,N_7758);
nor U8822 (N_8822,N_7667,N_7094);
or U8823 (N_8823,N_7722,N_7222);
or U8824 (N_8824,N_7096,N_7336);
or U8825 (N_8825,N_7894,N_7953);
nand U8826 (N_8826,N_7304,N_7410);
nand U8827 (N_8827,N_7018,N_7815);
and U8828 (N_8828,N_7035,N_7424);
or U8829 (N_8829,N_7810,N_7777);
nor U8830 (N_8830,N_7490,N_7350);
and U8831 (N_8831,N_7863,N_7484);
or U8832 (N_8832,N_7675,N_7865);
nand U8833 (N_8833,N_7102,N_7524);
xor U8834 (N_8834,N_7734,N_7421);
nand U8835 (N_8835,N_7226,N_7174);
or U8836 (N_8836,N_7494,N_7064);
xor U8837 (N_8837,N_7503,N_7045);
nand U8838 (N_8838,N_7888,N_7714);
or U8839 (N_8839,N_7899,N_7948);
nand U8840 (N_8840,N_7583,N_7582);
xor U8841 (N_8841,N_7046,N_7598);
or U8842 (N_8842,N_7312,N_7749);
nand U8843 (N_8843,N_7947,N_7495);
nand U8844 (N_8844,N_7305,N_7542);
nand U8845 (N_8845,N_7302,N_7408);
and U8846 (N_8846,N_7848,N_7239);
or U8847 (N_8847,N_7612,N_7368);
or U8848 (N_8848,N_7305,N_7096);
nand U8849 (N_8849,N_7271,N_7631);
and U8850 (N_8850,N_7995,N_7369);
and U8851 (N_8851,N_7696,N_7257);
xor U8852 (N_8852,N_7600,N_7734);
or U8853 (N_8853,N_7838,N_7163);
nand U8854 (N_8854,N_7988,N_7767);
or U8855 (N_8855,N_7895,N_7812);
nor U8856 (N_8856,N_7123,N_7501);
nand U8857 (N_8857,N_7339,N_7123);
xor U8858 (N_8858,N_7239,N_7884);
nand U8859 (N_8859,N_7061,N_7315);
nand U8860 (N_8860,N_7210,N_7743);
or U8861 (N_8861,N_7205,N_7123);
and U8862 (N_8862,N_7758,N_7135);
xnor U8863 (N_8863,N_7112,N_7643);
nand U8864 (N_8864,N_7066,N_7980);
and U8865 (N_8865,N_7571,N_7195);
nand U8866 (N_8866,N_7361,N_7684);
nand U8867 (N_8867,N_7561,N_7049);
or U8868 (N_8868,N_7168,N_7893);
or U8869 (N_8869,N_7551,N_7510);
xnor U8870 (N_8870,N_7319,N_7976);
nor U8871 (N_8871,N_7791,N_7154);
nor U8872 (N_8872,N_7017,N_7545);
nor U8873 (N_8873,N_7702,N_7426);
nor U8874 (N_8874,N_7230,N_7975);
and U8875 (N_8875,N_7466,N_7538);
xnor U8876 (N_8876,N_7696,N_7033);
or U8877 (N_8877,N_7552,N_7683);
nor U8878 (N_8878,N_7352,N_7525);
nand U8879 (N_8879,N_7054,N_7675);
or U8880 (N_8880,N_7492,N_7209);
nand U8881 (N_8881,N_7674,N_7021);
and U8882 (N_8882,N_7433,N_7553);
nor U8883 (N_8883,N_7460,N_7035);
and U8884 (N_8884,N_7977,N_7234);
and U8885 (N_8885,N_7370,N_7535);
nor U8886 (N_8886,N_7323,N_7887);
nor U8887 (N_8887,N_7554,N_7991);
nor U8888 (N_8888,N_7070,N_7100);
nand U8889 (N_8889,N_7951,N_7696);
nand U8890 (N_8890,N_7590,N_7389);
or U8891 (N_8891,N_7395,N_7964);
and U8892 (N_8892,N_7596,N_7957);
xnor U8893 (N_8893,N_7628,N_7983);
and U8894 (N_8894,N_7292,N_7969);
nor U8895 (N_8895,N_7175,N_7622);
or U8896 (N_8896,N_7506,N_7065);
or U8897 (N_8897,N_7876,N_7017);
or U8898 (N_8898,N_7217,N_7522);
or U8899 (N_8899,N_7679,N_7041);
nand U8900 (N_8900,N_7473,N_7732);
nor U8901 (N_8901,N_7285,N_7775);
nor U8902 (N_8902,N_7658,N_7197);
nand U8903 (N_8903,N_7604,N_7175);
and U8904 (N_8904,N_7548,N_7278);
or U8905 (N_8905,N_7531,N_7782);
and U8906 (N_8906,N_7363,N_7275);
or U8907 (N_8907,N_7981,N_7824);
or U8908 (N_8908,N_7724,N_7138);
or U8909 (N_8909,N_7317,N_7489);
and U8910 (N_8910,N_7252,N_7499);
or U8911 (N_8911,N_7728,N_7565);
and U8912 (N_8912,N_7367,N_7045);
nand U8913 (N_8913,N_7460,N_7743);
or U8914 (N_8914,N_7705,N_7126);
and U8915 (N_8915,N_7228,N_7433);
or U8916 (N_8916,N_7576,N_7068);
and U8917 (N_8917,N_7249,N_7215);
or U8918 (N_8918,N_7631,N_7603);
nor U8919 (N_8919,N_7528,N_7262);
nor U8920 (N_8920,N_7483,N_7384);
or U8921 (N_8921,N_7654,N_7580);
and U8922 (N_8922,N_7755,N_7728);
nand U8923 (N_8923,N_7476,N_7945);
or U8924 (N_8924,N_7620,N_7078);
or U8925 (N_8925,N_7142,N_7201);
xor U8926 (N_8926,N_7626,N_7257);
and U8927 (N_8927,N_7429,N_7220);
and U8928 (N_8928,N_7355,N_7004);
nor U8929 (N_8929,N_7181,N_7049);
nand U8930 (N_8930,N_7258,N_7560);
nand U8931 (N_8931,N_7904,N_7611);
or U8932 (N_8932,N_7957,N_7177);
nand U8933 (N_8933,N_7509,N_7279);
nand U8934 (N_8934,N_7208,N_7496);
and U8935 (N_8935,N_7926,N_7476);
xnor U8936 (N_8936,N_7735,N_7530);
and U8937 (N_8937,N_7649,N_7511);
nand U8938 (N_8938,N_7355,N_7286);
and U8939 (N_8939,N_7489,N_7827);
nor U8940 (N_8940,N_7343,N_7888);
xor U8941 (N_8941,N_7393,N_7071);
or U8942 (N_8942,N_7774,N_7499);
nand U8943 (N_8943,N_7860,N_7742);
nand U8944 (N_8944,N_7354,N_7543);
nand U8945 (N_8945,N_7519,N_7074);
and U8946 (N_8946,N_7557,N_7424);
or U8947 (N_8947,N_7695,N_7664);
xor U8948 (N_8948,N_7283,N_7348);
nand U8949 (N_8949,N_7154,N_7983);
and U8950 (N_8950,N_7836,N_7490);
xor U8951 (N_8951,N_7200,N_7965);
nor U8952 (N_8952,N_7198,N_7619);
nor U8953 (N_8953,N_7660,N_7064);
or U8954 (N_8954,N_7071,N_7939);
nand U8955 (N_8955,N_7248,N_7036);
or U8956 (N_8956,N_7270,N_7614);
nor U8957 (N_8957,N_7229,N_7179);
nor U8958 (N_8958,N_7147,N_7583);
or U8959 (N_8959,N_7842,N_7489);
or U8960 (N_8960,N_7486,N_7695);
or U8961 (N_8961,N_7799,N_7212);
xor U8962 (N_8962,N_7374,N_7743);
or U8963 (N_8963,N_7236,N_7175);
xnor U8964 (N_8964,N_7811,N_7882);
and U8965 (N_8965,N_7540,N_7797);
or U8966 (N_8966,N_7441,N_7115);
xnor U8967 (N_8967,N_7162,N_7193);
and U8968 (N_8968,N_7130,N_7193);
nor U8969 (N_8969,N_7451,N_7164);
nor U8970 (N_8970,N_7228,N_7682);
nand U8971 (N_8971,N_7405,N_7958);
or U8972 (N_8972,N_7608,N_7599);
nor U8973 (N_8973,N_7179,N_7167);
and U8974 (N_8974,N_7310,N_7894);
xor U8975 (N_8975,N_7465,N_7840);
nand U8976 (N_8976,N_7765,N_7179);
nor U8977 (N_8977,N_7965,N_7878);
nor U8978 (N_8978,N_7051,N_7366);
nand U8979 (N_8979,N_7071,N_7499);
and U8980 (N_8980,N_7619,N_7097);
and U8981 (N_8981,N_7006,N_7841);
or U8982 (N_8982,N_7134,N_7040);
nand U8983 (N_8983,N_7669,N_7448);
or U8984 (N_8984,N_7956,N_7724);
or U8985 (N_8985,N_7287,N_7450);
nand U8986 (N_8986,N_7919,N_7603);
nor U8987 (N_8987,N_7703,N_7870);
or U8988 (N_8988,N_7766,N_7425);
xnor U8989 (N_8989,N_7163,N_7681);
nor U8990 (N_8990,N_7004,N_7344);
nand U8991 (N_8991,N_7149,N_7137);
nor U8992 (N_8992,N_7805,N_7854);
nand U8993 (N_8993,N_7372,N_7101);
xnor U8994 (N_8994,N_7900,N_7817);
and U8995 (N_8995,N_7613,N_7044);
and U8996 (N_8996,N_7882,N_7102);
nand U8997 (N_8997,N_7279,N_7769);
nor U8998 (N_8998,N_7762,N_7403);
and U8999 (N_8999,N_7802,N_7157);
nor U9000 (N_9000,N_8107,N_8797);
nor U9001 (N_9001,N_8702,N_8517);
nor U9002 (N_9002,N_8201,N_8653);
nand U9003 (N_9003,N_8471,N_8903);
or U9004 (N_9004,N_8084,N_8985);
nor U9005 (N_9005,N_8256,N_8499);
or U9006 (N_9006,N_8624,N_8464);
nand U9007 (N_9007,N_8675,N_8351);
nand U9008 (N_9008,N_8595,N_8053);
nand U9009 (N_9009,N_8699,N_8161);
nor U9010 (N_9010,N_8440,N_8576);
nor U9011 (N_9011,N_8852,N_8063);
or U9012 (N_9012,N_8924,N_8183);
xnor U9013 (N_9013,N_8844,N_8661);
nand U9014 (N_9014,N_8268,N_8825);
nor U9015 (N_9015,N_8111,N_8211);
or U9016 (N_9016,N_8424,N_8663);
and U9017 (N_9017,N_8950,N_8771);
nand U9018 (N_9018,N_8807,N_8745);
nand U9019 (N_9019,N_8796,N_8008);
or U9020 (N_9020,N_8850,N_8441);
nor U9021 (N_9021,N_8848,N_8033);
and U9022 (N_9022,N_8735,N_8393);
nor U9023 (N_9023,N_8960,N_8536);
nor U9024 (N_9024,N_8504,N_8698);
xor U9025 (N_9025,N_8181,N_8946);
nor U9026 (N_9026,N_8120,N_8388);
nand U9027 (N_9027,N_8235,N_8336);
nor U9028 (N_9028,N_8673,N_8737);
and U9029 (N_9029,N_8124,N_8944);
and U9030 (N_9030,N_8882,N_8206);
or U9031 (N_9031,N_8414,N_8831);
or U9032 (N_9032,N_8748,N_8380);
nor U9033 (N_9033,N_8971,N_8701);
xnor U9034 (N_9034,N_8671,N_8563);
nand U9035 (N_9035,N_8812,N_8788);
and U9036 (N_9036,N_8587,N_8872);
xor U9037 (N_9037,N_8939,N_8695);
nor U9038 (N_9038,N_8945,N_8011);
nor U9039 (N_9039,N_8606,N_8876);
and U9040 (N_9040,N_8453,N_8109);
or U9041 (N_9041,N_8479,N_8794);
and U9042 (N_9042,N_8209,N_8190);
and U9043 (N_9043,N_8976,N_8878);
nand U9044 (N_9044,N_8058,N_8870);
nor U9045 (N_9045,N_8472,N_8954);
or U9046 (N_9046,N_8941,N_8288);
xor U9047 (N_9047,N_8935,N_8961);
nor U9048 (N_9048,N_8460,N_8833);
nand U9049 (N_9049,N_8205,N_8400);
and U9050 (N_9050,N_8880,N_8834);
nand U9051 (N_9051,N_8358,N_8384);
or U9052 (N_9052,N_8591,N_8173);
or U9053 (N_9053,N_8719,N_8118);
xor U9054 (N_9054,N_8616,N_8317);
nand U9055 (N_9055,N_8943,N_8168);
xnor U9056 (N_9056,N_8476,N_8710);
and U9057 (N_9057,N_8247,N_8642);
and U9058 (N_9058,N_8095,N_8327);
and U9059 (N_9059,N_8886,N_8895);
or U9060 (N_9060,N_8319,N_8708);
or U9061 (N_9061,N_8601,N_8417);
nand U9062 (N_9062,N_8324,N_8607);
nand U9063 (N_9063,N_8902,N_8717);
or U9064 (N_9064,N_8864,N_8530);
nand U9065 (N_9065,N_8128,N_8592);
nand U9066 (N_9066,N_8805,N_8314);
nand U9067 (N_9067,N_8552,N_8223);
and U9068 (N_9068,N_8192,N_8066);
and U9069 (N_9069,N_8547,N_8559);
nor U9070 (N_9070,N_8619,N_8044);
or U9071 (N_9071,N_8691,N_8622);
nor U9072 (N_9072,N_8693,N_8134);
nand U9073 (N_9073,N_8186,N_8936);
nand U9074 (N_9074,N_8222,N_8052);
nand U9075 (N_9075,N_8605,N_8694);
nand U9076 (N_9076,N_8277,N_8610);
nor U9077 (N_9077,N_8260,N_8838);
and U9078 (N_9078,N_8979,N_8059);
and U9079 (N_9079,N_8625,N_8697);
nand U9080 (N_9080,N_8357,N_8915);
nand U9081 (N_9081,N_8275,N_8258);
or U9082 (N_9082,N_8801,N_8230);
xor U9083 (N_9083,N_8113,N_8993);
nand U9084 (N_9084,N_8366,N_8452);
and U9085 (N_9085,N_8396,N_8569);
and U9086 (N_9086,N_8135,N_8637);
or U9087 (N_9087,N_8767,N_8104);
nor U9088 (N_9088,N_8980,N_8332);
nand U9089 (N_9089,N_8855,N_8254);
or U9090 (N_9090,N_8212,N_8392);
and U9091 (N_9091,N_8076,N_8662);
nand U9092 (N_9092,N_8437,N_8297);
nand U9093 (N_9093,N_8543,N_8024);
and U9094 (N_9094,N_8463,N_8740);
or U9095 (N_9095,N_8583,N_8974);
nor U9096 (N_9096,N_8139,N_8656);
and U9097 (N_9097,N_8474,N_8567);
nand U9098 (N_9098,N_8784,N_8928);
xnor U9099 (N_9099,N_8473,N_8466);
nor U9100 (N_9100,N_8395,N_8813);
nand U9101 (N_9101,N_8225,N_8588);
or U9102 (N_9102,N_8165,N_8612);
nand U9103 (N_9103,N_8753,N_8454);
xor U9104 (N_9104,N_8712,N_8204);
nor U9105 (N_9105,N_8199,N_8436);
and U9106 (N_9106,N_8892,N_8132);
nand U9107 (N_9107,N_8506,N_8420);
or U9108 (N_9108,N_8761,N_8166);
xor U9109 (N_9109,N_8023,N_8611);
or U9110 (N_9110,N_8434,N_8615);
and U9111 (N_9111,N_8861,N_8713);
nand U9112 (N_9112,N_8545,N_8500);
or U9113 (N_9113,N_8450,N_8816);
nor U9114 (N_9114,N_8746,N_8550);
or U9115 (N_9115,N_8425,N_8343);
and U9116 (N_9116,N_8034,N_8514);
xor U9117 (N_9117,N_8185,N_8913);
xor U9118 (N_9118,N_8187,N_8069);
and U9119 (N_9119,N_8683,N_8065);
and U9120 (N_9120,N_8951,N_8240);
nor U9121 (N_9121,N_8233,N_8786);
or U9122 (N_9122,N_8129,N_8724);
or U9123 (N_9123,N_8178,N_8540);
nand U9124 (N_9124,N_8074,N_8660);
nand U9125 (N_9125,N_8692,N_8362);
and U9126 (N_9126,N_8339,N_8546);
nand U9127 (N_9127,N_8755,N_8217);
xor U9128 (N_9128,N_8732,N_8854);
or U9129 (N_9129,N_8887,N_8346);
nand U9130 (N_9130,N_8459,N_8598);
or U9131 (N_9131,N_8325,N_8604);
or U9132 (N_9132,N_8981,N_8992);
or U9133 (N_9133,N_8893,N_8435);
nand U9134 (N_9134,N_8681,N_8197);
nor U9135 (N_9135,N_8176,N_8342);
nand U9136 (N_9136,N_8729,N_8068);
nor U9137 (N_9137,N_8394,N_8940);
nor U9138 (N_9138,N_8221,N_8018);
or U9139 (N_9139,N_8775,N_8078);
nand U9140 (N_9140,N_8064,N_8937);
xnor U9141 (N_9141,N_8766,N_8012);
or U9142 (N_9142,N_8734,N_8808);
or U9143 (N_9143,N_8010,N_8196);
nand U9144 (N_9144,N_8868,N_8883);
nand U9145 (N_9145,N_8207,N_8410);
or U9146 (N_9146,N_8110,N_8597);
and U9147 (N_9147,N_8073,N_8029);
nand U9148 (N_9148,N_8641,N_8818);
nor U9149 (N_9149,N_8482,N_8926);
nor U9150 (N_9150,N_8898,N_8492);
nand U9151 (N_9151,N_8635,N_8665);
or U9152 (N_9152,N_8997,N_8050);
nand U9153 (N_9153,N_8412,N_8518);
or U9154 (N_9154,N_8909,N_8820);
nand U9155 (N_9155,N_8016,N_8035);
nand U9156 (N_9156,N_8401,N_8933);
or U9157 (N_9157,N_8080,N_8251);
or U9158 (N_9158,N_8707,N_8005);
or U9159 (N_9159,N_8790,N_8776);
and U9160 (N_9160,N_8741,N_8930);
nand U9161 (N_9161,N_8842,N_8000);
nor U9162 (N_9162,N_8925,N_8285);
and U9163 (N_9163,N_8274,N_8823);
nand U9164 (N_9164,N_8041,N_8977);
or U9165 (N_9165,N_8756,N_8533);
or U9166 (N_9166,N_8573,N_8894);
and U9167 (N_9167,N_8220,N_8231);
and U9168 (N_9168,N_8562,N_8731);
xnor U9169 (N_9169,N_8851,N_8374);
nand U9170 (N_9170,N_8305,N_8269);
or U9171 (N_9171,N_8791,N_8955);
nor U9172 (N_9172,N_8426,N_8966);
nand U9173 (N_9173,N_8371,N_8914);
and U9174 (N_9174,N_8502,N_8525);
nor U9175 (N_9175,N_8867,N_8302);
nor U9176 (N_9176,N_8389,N_8811);
and U9177 (N_9177,N_8363,N_8989);
or U9178 (N_9178,N_8633,N_8070);
or U9179 (N_9179,N_8089,N_8709);
nand U9180 (N_9180,N_8164,N_8609);
and U9181 (N_9181,N_8227,N_8157);
xor U9182 (N_9182,N_8520,N_8310);
nand U9183 (N_9183,N_8077,N_8793);
or U9184 (N_9184,N_8809,N_8272);
or U9185 (N_9185,N_8037,N_8350);
and U9186 (N_9186,N_8154,N_8246);
nor U9187 (N_9187,N_8379,N_8055);
nand U9188 (N_9188,N_8579,N_8398);
and U9189 (N_9189,N_8590,N_8096);
or U9190 (N_9190,N_8087,N_8524);
or U9191 (N_9191,N_8382,N_8334);
nand U9192 (N_9192,N_8326,N_8081);
nand U9193 (N_9193,N_8083,N_8983);
nor U9194 (N_9194,N_8248,N_8323);
nor U9195 (N_9195,N_8564,N_8172);
and U9196 (N_9196,N_8744,N_8853);
or U9197 (N_9197,N_8758,N_8099);
and U9198 (N_9198,N_8191,N_8022);
nand U9199 (N_9199,N_8581,N_8743);
and U9200 (N_9200,N_8904,N_8690);
nand U9201 (N_9201,N_8787,N_8458);
or U9202 (N_9202,N_8515,N_8542);
or U9203 (N_9203,N_8079,N_8281);
or U9204 (N_9204,N_8726,N_8534);
xnor U9205 (N_9205,N_8650,N_8210);
xnor U9206 (N_9206,N_8193,N_8969);
xor U9207 (N_9207,N_8341,N_8652);
nor U9208 (N_9208,N_8723,N_8535);
xnor U9209 (N_9209,N_8042,N_8860);
nand U9210 (N_9210,N_8602,N_8521);
nand U9211 (N_9211,N_8369,N_8447);
and U9212 (N_9212,N_8301,N_8762);
or U9213 (N_9213,N_8431,N_8760);
or U9214 (N_9214,N_8575,N_8102);
nor U9215 (N_9215,N_8017,N_8307);
nand U9216 (N_9216,N_8802,N_8299);
nor U9217 (N_9217,N_8718,N_8910);
nand U9218 (N_9218,N_8501,N_8555);
nand U9219 (N_9219,N_8965,N_8705);
and U9220 (N_9220,N_8122,N_8330);
nor U9221 (N_9221,N_8188,N_8040);
xor U9222 (N_9222,N_8649,N_8169);
and U9223 (N_9223,N_8028,N_8238);
xor U9224 (N_9224,N_8832,N_8287);
nand U9225 (N_9225,N_8978,N_8027);
nand U9226 (N_9226,N_8179,N_8742);
nor U9227 (N_9227,N_8489,N_8090);
nor U9228 (N_9228,N_8556,N_8048);
nand U9229 (N_9229,N_8510,N_8901);
xor U9230 (N_9230,N_8483,N_8086);
nand U9231 (N_9231,N_8075,N_8266);
and U9232 (N_9232,N_8145,N_8045);
nand U9233 (N_9233,N_8614,N_8337);
nand U9234 (N_9234,N_8177,N_8770);
and U9235 (N_9235,N_8331,N_8988);
nand U9236 (N_9236,N_8531,N_8121);
nand U9237 (N_9237,N_8202,N_8214);
or U9238 (N_9238,N_8255,N_8144);
or U9239 (N_9239,N_8640,N_8779);
and U9240 (N_9240,N_8561,N_8627);
nand U9241 (N_9241,N_8194,N_8329);
nor U9242 (N_9242,N_8998,N_8123);
and U9243 (N_9243,N_8752,N_8948);
or U9244 (N_9244,N_8728,N_8047);
nand U9245 (N_9245,N_8383,N_8421);
and U9246 (N_9246,N_8780,N_8162);
or U9247 (N_9247,N_8956,N_8490);
and U9248 (N_9248,N_8405,N_8439);
nand U9249 (N_9249,N_8934,N_8413);
nor U9250 (N_9250,N_8427,N_8879);
nor U9251 (N_9251,N_8171,N_8964);
nor U9252 (N_9252,N_8685,N_8824);
or U9253 (N_9253,N_8320,N_8491);
and U9254 (N_9254,N_8657,N_8513);
or U9255 (N_9255,N_8494,N_8344);
nor U9256 (N_9256,N_8647,N_8630);
nand U9257 (N_9257,N_8585,N_8608);
or U9258 (N_9258,N_8278,N_8865);
xnor U9259 (N_9259,N_8829,N_8303);
or U9260 (N_9260,N_8676,N_8242);
nor U9261 (N_9261,N_8658,N_8432);
or U9262 (N_9262,N_8101,N_8313);
xnor U9263 (N_9263,N_8486,N_8250);
or U9264 (N_9264,N_8443,N_8749);
nor U9265 (N_9265,N_8270,N_8409);
nand U9266 (N_9266,N_8714,N_8727);
xor U9267 (N_9267,N_8907,N_8236);
nand U9268 (N_9268,N_8105,N_8519);
nand U9269 (N_9269,N_8666,N_8803);
nor U9270 (N_9270,N_8406,N_8528);
nor U9271 (N_9271,N_8019,N_8373);
nor U9272 (N_9272,N_8725,N_8733);
and U9273 (N_9273,N_8001,N_8416);
and U9274 (N_9274,N_8548,N_8408);
nor U9275 (N_9275,N_8826,N_8309);
nor U9276 (N_9276,N_8335,N_8419);
nor U9277 (N_9277,N_8284,N_8982);
nor U9278 (N_9278,N_8036,N_8365);
and U9279 (N_9279,N_8461,N_8487);
nand U9280 (N_9280,N_8234,N_8043);
nand U9281 (N_9281,N_8991,N_8815);
or U9282 (N_9282,N_8891,N_8228);
and U9283 (N_9283,N_8574,N_8446);
and U9284 (N_9284,N_8912,N_8137);
and U9285 (N_9285,N_8999,N_8237);
nor U9286 (N_9286,N_8908,N_8271);
and U9287 (N_9287,N_8088,N_8679);
and U9288 (N_9288,N_8468,N_8821);
nor U9289 (N_9289,N_8859,N_8376);
or U9290 (N_9290,N_8814,N_8557);
nor U9291 (N_9291,N_8160,N_8368);
and U9292 (N_9292,N_8094,N_8208);
or U9293 (N_9293,N_8031,N_8298);
nor U9294 (N_9294,N_8817,N_8798);
and U9295 (N_9295,N_8115,N_8152);
or U9296 (N_9296,N_8198,N_8819);
and U9297 (N_9297,N_8021,N_8032);
nand U9298 (N_9298,N_8577,N_8539);
nor U9299 (N_9299,N_8906,N_8738);
or U9300 (N_9300,N_8578,N_8167);
or U9301 (N_9301,N_8163,N_8843);
or U9302 (N_9302,N_8617,N_8927);
nor U9303 (N_9303,N_8847,N_8566);
nor U9304 (N_9304,N_8387,N_8153);
nor U9305 (N_9305,N_8062,N_8835);
nand U9306 (N_9306,N_8618,N_8958);
nor U9307 (N_9307,N_8862,N_8311);
xor U9308 (N_9308,N_8899,N_8026);
nor U9309 (N_9309,N_8498,N_8804);
or U9310 (N_9310,N_8216,N_8554);
and U9311 (N_9311,N_8551,N_8952);
or U9312 (N_9312,N_8252,N_8783);
nor U9313 (N_9313,N_8768,N_8493);
or U9314 (N_9314,N_8594,N_8004);
or U9315 (N_9315,N_8651,N_8478);
nand U9316 (N_9316,N_8736,N_8863);
or U9317 (N_9317,N_8318,N_8621);
and U9318 (N_9318,N_8512,N_8565);
nor U9319 (N_9319,N_8159,N_8990);
nor U9320 (N_9320,N_8570,N_8480);
nor U9321 (N_9321,N_8112,N_8837);
and U9322 (N_9322,N_8182,N_8349);
nor U9323 (N_9323,N_8232,N_8968);
nand U9324 (N_9324,N_8340,N_8131);
and U9325 (N_9325,N_8774,N_8503);
nand U9326 (N_9326,N_8149,N_8025);
nand U9327 (N_9327,N_8664,N_8264);
nand U9328 (N_9328,N_8778,N_8655);
nand U9329 (N_9329,N_8792,N_8315);
or U9330 (N_9330,N_8856,N_8529);
and U9331 (N_9331,N_8537,N_8677);
nor U9332 (N_9332,N_8259,N_8747);
nor U9333 (N_9333,N_8639,N_8923);
and U9334 (N_9334,N_8972,N_8789);
nor U9335 (N_9335,N_8423,N_8060);
nand U9336 (N_9336,N_8987,N_8049);
nand U9337 (N_9337,N_8253,N_8527);
or U9338 (N_9338,N_8082,N_8397);
or U9339 (N_9339,N_8477,N_8553);
nor U9340 (N_9340,N_8688,N_8359);
nand U9341 (N_9341,N_8444,N_8411);
nor U9342 (N_9342,N_8241,N_8888);
nor U9343 (N_9343,N_8293,N_8455);
or U9344 (N_9344,N_8385,N_8377);
or U9345 (N_9345,N_8549,N_8184);
or U9346 (N_9346,N_8875,N_8629);
or U9347 (N_9347,N_8626,N_8457);
and U9348 (N_9348,N_8496,N_8356);
nand U9349 (N_9349,N_8292,N_8881);
or U9350 (N_9350,N_8481,N_8245);
nand U9351 (N_9351,N_8684,N_8739);
nand U9352 (N_9352,N_8061,N_8143);
nand U9353 (N_9353,N_8680,N_8922);
nor U9354 (N_9354,N_8263,N_8715);
or U9355 (N_9355,N_8919,N_8433);
nand U9356 (N_9356,N_8039,N_8636);
or U9357 (N_9357,N_8051,N_8404);
and U9358 (N_9358,N_8646,N_8703);
or U9359 (N_9359,N_8704,N_8013);
and U9360 (N_9360,N_8957,N_8345);
and U9361 (N_9361,N_8103,N_8038);
nand U9362 (N_9362,N_8097,N_8781);
nand U9363 (N_9363,N_8106,N_8386);
xnor U9364 (N_9364,N_8189,N_8800);
and U9365 (N_9365,N_8507,N_8905);
or U9366 (N_9366,N_8670,N_8568);
and U9367 (N_9367,N_8361,N_8773);
nor U9368 (N_9368,N_8422,N_8003);
nand U9369 (N_9369,N_8352,N_8827);
nand U9370 (N_9370,N_8721,N_8828);
or U9371 (N_9371,N_8151,N_8582);
or U9372 (N_9372,N_8975,N_8469);
nand U9373 (N_9373,N_8402,N_8219);
and U9374 (N_9374,N_8322,N_8126);
xor U9375 (N_9375,N_8226,N_8890);
or U9376 (N_9376,N_8257,N_8644);
nand U9377 (N_9377,N_8140,N_8092);
or U9378 (N_9378,N_8866,N_8584);
nand U9379 (N_9379,N_8449,N_8200);
nor U9380 (N_9380,N_8456,N_8795);
nand U9381 (N_9381,N_8757,N_8261);
and U9382 (N_9382,N_8429,N_8764);
or U9383 (N_9383,N_8338,N_8072);
or U9384 (N_9384,N_8917,N_8858);
nand U9385 (N_9385,N_8030,N_8942);
and U9386 (N_9386,N_8628,N_8117);
nand U9387 (N_9387,N_8716,N_8295);
xnor U9388 (N_9388,N_8215,N_8959);
and U9389 (N_9389,N_8884,N_8526);
nand U9390 (N_9390,N_8470,N_8996);
or U9391 (N_9391,N_8654,N_8672);
nand U9392 (N_9392,N_8390,N_8720);
nor U9393 (N_9393,N_8874,N_8438);
nand U9394 (N_9394,N_8130,N_8054);
xnor U9395 (N_9395,N_8071,N_8696);
or U9396 (N_9396,N_8857,N_8623);
nand U9397 (N_9397,N_8462,N_8170);
nor U9398 (N_9398,N_8754,N_8015);
and U9399 (N_9399,N_8378,N_8967);
or U9400 (N_9400,N_8505,N_8931);
nor U9401 (N_9401,N_8283,N_8180);
or U9402 (N_9402,N_8348,N_8667);
and U9403 (N_9403,N_8391,N_8306);
and U9404 (N_9404,N_8750,N_8007);
and U9405 (N_9405,N_8229,N_8511);
and U9406 (N_9406,N_8497,N_8290);
nand U9407 (N_9407,N_8632,N_8769);
and U9408 (N_9408,N_8638,N_8218);
and U9409 (N_9409,N_8294,N_8304);
xnor U9410 (N_9410,N_8648,N_8643);
nor U9411 (N_9411,N_8114,N_8586);
xor U9412 (N_9412,N_8845,N_8687);
nor U9413 (N_9413,N_8372,N_8949);
and U9414 (N_9414,N_8836,N_8355);
nand U9415 (N_9415,N_8620,N_8484);
or U9416 (N_9416,N_8249,N_8243);
and U9417 (N_9417,N_8407,N_8485);
nand U9418 (N_9418,N_8929,N_8428);
nor U9419 (N_9419,N_8475,N_8634);
or U9420 (N_9420,N_8150,N_8279);
nor U9421 (N_9421,N_8116,N_8100);
or U9422 (N_9422,N_8347,N_8125);
or U9423 (N_9423,N_8158,N_8763);
and U9424 (N_9424,N_8785,N_8267);
and U9425 (N_9425,N_8451,N_8014);
nand U9426 (N_9426,N_8085,N_8333);
or U9427 (N_9427,N_8846,N_8889);
nor U9428 (N_9428,N_8544,N_8495);
and U9429 (N_9429,N_8286,N_8289);
and U9430 (N_9430,N_8448,N_8599);
nor U9431 (N_9431,N_8668,N_8678);
and U9432 (N_9432,N_8921,N_8669);
or U9433 (N_9433,N_8174,N_8354);
and U9434 (N_9434,N_8175,N_8146);
and U9435 (N_9435,N_8541,N_8532);
or U9436 (N_9436,N_8156,N_8488);
and U9437 (N_9437,N_8686,N_8963);
and U9438 (N_9438,N_8415,N_8869);
or U9439 (N_9439,N_8580,N_8558);
or U9440 (N_9440,N_8572,N_8986);
nand U9441 (N_9441,N_8994,N_8002);
and U9442 (N_9442,N_8830,N_8142);
or U9443 (N_9443,N_8953,N_8706);
nand U9444 (N_9444,N_8896,N_8467);
and U9445 (N_9445,N_8689,N_8300);
nor U9446 (N_9446,N_8508,N_8445);
xnor U9447 (N_9447,N_8631,N_8155);
and U9448 (N_9448,N_8516,N_8730);
xnor U9449 (N_9449,N_8932,N_8213);
nand U9450 (N_9450,N_8920,N_8296);
xor U9451 (N_9451,N_8885,N_8522);
nor U9452 (N_9452,N_8375,N_8136);
and U9453 (N_9453,N_8900,N_8119);
xnor U9454 (N_9454,N_8316,N_8674);
or U9455 (N_9455,N_8765,N_8938);
or U9456 (N_9456,N_8962,N_8841);
nor U9457 (N_9457,N_8806,N_8593);
nand U9458 (N_9458,N_8321,N_8418);
xor U9459 (N_9459,N_8006,N_8984);
nor U9460 (N_9460,N_8916,N_8877);
and U9461 (N_9461,N_8589,N_8273);
nand U9462 (N_9462,N_8777,N_8810);
nor U9463 (N_9463,N_8442,N_8147);
nor U9464 (N_9464,N_8108,N_8364);
or U9465 (N_9465,N_8312,N_8141);
xnor U9466 (N_9466,N_8093,N_8571);
and U9467 (N_9467,N_8839,N_8308);
nor U9468 (N_9468,N_8523,N_8148);
nor U9469 (N_9469,N_8603,N_8711);
nand U9470 (N_9470,N_8067,N_8224);
nor U9471 (N_9471,N_8403,N_8822);
nand U9472 (N_9472,N_8328,N_8020);
and U9473 (N_9473,N_8897,N_8360);
nand U9474 (N_9474,N_8367,N_8613);
or U9475 (N_9475,N_8509,N_8918);
and U9476 (N_9476,N_8947,N_8009);
nand U9477 (N_9477,N_8133,N_8282);
and U9478 (N_9478,N_8138,N_8873);
or U9479 (N_9479,N_8722,N_8645);
and U9480 (N_9480,N_8195,N_8659);
xnor U9481 (N_9481,N_8995,N_8973);
nor U9482 (N_9482,N_8276,N_8262);
and U9483 (N_9483,N_8370,N_8381);
and U9484 (N_9484,N_8759,N_8970);
nor U9485 (N_9485,N_8353,N_8399);
and U9486 (N_9486,N_8239,N_8280);
and U9487 (N_9487,N_8751,N_8046);
xor U9488 (N_9488,N_8871,N_8465);
nor U9489 (N_9489,N_8560,N_8057);
nor U9490 (N_9490,N_8538,N_8682);
nand U9491 (N_9491,N_8799,N_8782);
nor U9492 (N_9492,N_8244,N_8091);
xor U9493 (N_9493,N_8265,N_8772);
and U9494 (N_9494,N_8127,N_8291);
xnor U9495 (N_9495,N_8849,N_8056);
nand U9496 (N_9496,N_8700,N_8596);
or U9497 (N_9497,N_8840,N_8600);
and U9498 (N_9498,N_8098,N_8911);
nor U9499 (N_9499,N_8203,N_8430);
nor U9500 (N_9500,N_8510,N_8749);
and U9501 (N_9501,N_8590,N_8856);
or U9502 (N_9502,N_8790,N_8235);
or U9503 (N_9503,N_8734,N_8211);
nand U9504 (N_9504,N_8383,N_8622);
nand U9505 (N_9505,N_8486,N_8310);
and U9506 (N_9506,N_8222,N_8033);
nand U9507 (N_9507,N_8906,N_8532);
and U9508 (N_9508,N_8727,N_8167);
nand U9509 (N_9509,N_8385,N_8583);
or U9510 (N_9510,N_8931,N_8965);
nor U9511 (N_9511,N_8098,N_8418);
and U9512 (N_9512,N_8494,N_8603);
or U9513 (N_9513,N_8493,N_8196);
or U9514 (N_9514,N_8922,N_8554);
nand U9515 (N_9515,N_8037,N_8127);
or U9516 (N_9516,N_8402,N_8759);
xor U9517 (N_9517,N_8107,N_8574);
nor U9518 (N_9518,N_8853,N_8496);
nand U9519 (N_9519,N_8021,N_8942);
nand U9520 (N_9520,N_8554,N_8959);
nand U9521 (N_9521,N_8045,N_8057);
nand U9522 (N_9522,N_8941,N_8508);
or U9523 (N_9523,N_8914,N_8253);
nor U9524 (N_9524,N_8430,N_8519);
nand U9525 (N_9525,N_8288,N_8014);
nor U9526 (N_9526,N_8838,N_8841);
xnor U9527 (N_9527,N_8892,N_8193);
nand U9528 (N_9528,N_8057,N_8076);
nand U9529 (N_9529,N_8431,N_8146);
and U9530 (N_9530,N_8623,N_8089);
or U9531 (N_9531,N_8770,N_8721);
and U9532 (N_9532,N_8225,N_8265);
or U9533 (N_9533,N_8191,N_8308);
nor U9534 (N_9534,N_8592,N_8420);
nor U9535 (N_9535,N_8633,N_8736);
or U9536 (N_9536,N_8205,N_8477);
nand U9537 (N_9537,N_8720,N_8454);
and U9538 (N_9538,N_8144,N_8422);
and U9539 (N_9539,N_8249,N_8694);
nand U9540 (N_9540,N_8522,N_8807);
nor U9541 (N_9541,N_8645,N_8377);
nand U9542 (N_9542,N_8834,N_8018);
nor U9543 (N_9543,N_8257,N_8402);
nor U9544 (N_9544,N_8285,N_8113);
and U9545 (N_9545,N_8724,N_8745);
nand U9546 (N_9546,N_8374,N_8537);
and U9547 (N_9547,N_8078,N_8480);
xnor U9548 (N_9548,N_8521,N_8184);
nor U9549 (N_9549,N_8890,N_8858);
nor U9550 (N_9550,N_8580,N_8956);
nor U9551 (N_9551,N_8441,N_8203);
or U9552 (N_9552,N_8689,N_8865);
and U9553 (N_9553,N_8167,N_8446);
or U9554 (N_9554,N_8250,N_8591);
nand U9555 (N_9555,N_8632,N_8136);
nor U9556 (N_9556,N_8265,N_8179);
nand U9557 (N_9557,N_8562,N_8658);
or U9558 (N_9558,N_8089,N_8301);
or U9559 (N_9559,N_8185,N_8916);
nand U9560 (N_9560,N_8441,N_8595);
nor U9561 (N_9561,N_8864,N_8104);
and U9562 (N_9562,N_8439,N_8389);
nor U9563 (N_9563,N_8027,N_8320);
nand U9564 (N_9564,N_8267,N_8448);
nand U9565 (N_9565,N_8276,N_8235);
and U9566 (N_9566,N_8122,N_8919);
nor U9567 (N_9567,N_8633,N_8256);
and U9568 (N_9568,N_8900,N_8366);
nor U9569 (N_9569,N_8216,N_8176);
nor U9570 (N_9570,N_8305,N_8192);
xnor U9571 (N_9571,N_8278,N_8931);
and U9572 (N_9572,N_8374,N_8652);
nand U9573 (N_9573,N_8992,N_8431);
and U9574 (N_9574,N_8739,N_8963);
and U9575 (N_9575,N_8746,N_8397);
nor U9576 (N_9576,N_8171,N_8079);
xnor U9577 (N_9577,N_8090,N_8984);
or U9578 (N_9578,N_8719,N_8006);
and U9579 (N_9579,N_8518,N_8697);
or U9580 (N_9580,N_8716,N_8774);
nor U9581 (N_9581,N_8248,N_8685);
nor U9582 (N_9582,N_8006,N_8665);
xnor U9583 (N_9583,N_8521,N_8700);
or U9584 (N_9584,N_8969,N_8201);
xnor U9585 (N_9585,N_8607,N_8649);
nand U9586 (N_9586,N_8471,N_8468);
and U9587 (N_9587,N_8656,N_8741);
and U9588 (N_9588,N_8355,N_8881);
and U9589 (N_9589,N_8565,N_8478);
nor U9590 (N_9590,N_8529,N_8659);
xor U9591 (N_9591,N_8238,N_8778);
and U9592 (N_9592,N_8257,N_8661);
and U9593 (N_9593,N_8312,N_8052);
nor U9594 (N_9594,N_8423,N_8864);
or U9595 (N_9595,N_8473,N_8479);
xor U9596 (N_9596,N_8620,N_8622);
xor U9597 (N_9597,N_8638,N_8777);
xnor U9598 (N_9598,N_8338,N_8238);
and U9599 (N_9599,N_8254,N_8714);
and U9600 (N_9600,N_8391,N_8575);
and U9601 (N_9601,N_8616,N_8451);
nor U9602 (N_9602,N_8631,N_8651);
xor U9603 (N_9603,N_8925,N_8146);
nand U9604 (N_9604,N_8857,N_8841);
or U9605 (N_9605,N_8011,N_8213);
or U9606 (N_9606,N_8716,N_8102);
or U9607 (N_9607,N_8957,N_8006);
nand U9608 (N_9608,N_8599,N_8000);
and U9609 (N_9609,N_8424,N_8176);
and U9610 (N_9610,N_8676,N_8225);
nand U9611 (N_9611,N_8170,N_8505);
or U9612 (N_9612,N_8108,N_8188);
xnor U9613 (N_9613,N_8027,N_8767);
and U9614 (N_9614,N_8070,N_8899);
and U9615 (N_9615,N_8136,N_8371);
or U9616 (N_9616,N_8332,N_8716);
and U9617 (N_9617,N_8388,N_8711);
xor U9618 (N_9618,N_8280,N_8711);
nand U9619 (N_9619,N_8051,N_8403);
and U9620 (N_9620,N_8260,N_8586);
nor U9621 (N_9621,N_8100,N_8824);
and U9622 (N_9622,N_8161,N_8546);
and U9623 (N_9623,N_8424,N_8435);
and U9624 (N_9624,N_8804,N_8513);
and U9625 (N_9625,N_8261,N_8570);
xnor U9626 (N_9626,N_8600,N_8336);
nand U9627 (N_9627,N_8619,N_8253);
or U9628 (N_9628,N_8733,N_8326);
and U9629 (N_9629,N_8404,N_8853);
and U9630 (N_9630,N_8715,N_8360);
nor U9631 (N_9631,N_8742,N_8510);
nor U9632 (N_9632,N_8646,N_8667);
and U9633 (N_9633,N_8231,N_8452);
xor U9634 (N_9634,N_8477,N_8347);
or U9635 (N_9635,N_8522,N_8972);
nor U9636 (N_9636,N_8561,N_8776);
nand U9637 (N_9637,N_8359,N_8677);
nor U9638 (N_9638,N_8742,N_8570);
nand U9639 (N_9639,N_8565,N_8602);
nand U9640 (N_9640,N_8081,N_8529);
or U9641 (N_9641,N_8378,N_8457);
nand U9642 (N_9642,N_8628,N_8634);
or U9643 (N_9643,N_8994,N_8631);
nand U9644 (N_9644,N_8888,N_8849);
nand U9645 (N_9645,N_8509,N_8841);
and U9646 (N_9646,N_8027,N_8474);
and U9647 (N_9647,N_8141,N_8735);
xnor U9648 (N_9648,N_8729,N_8905);
or U9649 (N_9649,N_8976,N_8264);
or U9650 (N_9650,N_8918,N_8744);
or U9651 (N_9651,N_8830,N_8807);
and U9652 (N_9652,N_8133,N_8089);
nand U9653 (N_9653,N_8035,N_8244);
nor U9654 (N_9654,N_8534,N_8370);
nor U9655 (N_9655,N_8887,N_8658);
nand U9656 (N_9656,N_8838,N_8626);
nand U9657 (N_9657,N_8704,N_8925);
nor U9658 (N_9658,N_8544,N_8911);
nand U9659 (N_9659,N_8901,N_8195);
and U9660 (N_9660,N_8425,N_8003);
nand U9661 (N_9661,N_8899,N_8183);
nand U9662 (N_9662,N_8885,N_8852);
or U9663 (N_9663,N_8511,N_8566);
nor U9664 (N_9664,N_8730,N_8169);
nor U9665 (N_9665,N_8556,N_8336);
xnor U9666 (N_9666,N_8468,N_8287);
or U9667 (N_9667,N_8766,N_8713);
nor U9668 (N_9668,N_8234,N_8271);
and U9669 (N_9669,N_8369,N_8505);
nor U9670 (N_9670,N_8784,N_8040);
xor U9671 (N_9671,N_8701,N_8838);
nor U9672 (N_9672,N_8475,N_8707);
and U9673 (N_9673,N_8685,N_8355);
xor U9674 (N_9674,N_8045,N_8134);
nor U9675 (N_9675,N_8485,N_8053);
and U9676 (N_9676,N_8876,N_8714);
nor U9677 (N_9677,N_8547,N_8397);
or U9678 (N_9678,N_8354,N_8314);
xnor U9679 (N_9679,N_8442,N_8433);
and U9680 (N_9680,N_8039,N_8482);
nand U9681 (N_9681,N_8393,N_8144);
and U9682 (N_9682,N_8239,N_8454);
and U9683 (N_9683,N_8326,N_8313);
nor U9684 (N_9684,N_8862,N_8491);
and U9685 (N_9685,N_8686,N_8858);
nand U9686 (N_9686,N_8871,N_8830);
and U9687 (N_9687,N_8131,N_8522);
and U9688 (N_9688,N_8271,N_8927);
and U9689 (N_9689,N_8525,N_8333);
nor U9690 (N_9690,N_8882,N_8953);
and U9691 (N_9691,N_8977,N_8755);
or U9692 (N_9692,N_8359,N_8958);
nand U9693 (N_9693,N_8353,N_8701);
nor U9694 (N_9694,N_8185,N_8144);
xor U9695 (N_9695,N_8678,N_8997);
nor U9696 (N_9696,N_8519,N_8715);
or U9697 (N_9697,N_8734,N_8455);
nor U9698 (N_9698,N_8438,N_8456);
or U9699 (N_9699,N_8217,N_8067);
and U9700 (N_9700,N_8282,N_8270);
or U9701 (N_9701,N_8446,N_8712);
xor U9702 (N_9702,N_8371,N_8041);
nor U9703 (N_9703,N_8900,N_8662);
and U9704 (N_9704,N_8835,N_8035);
xor U9705 (N_9705,N_8764,N_8321);
nand U9706 (N_9706,N_8999,N_8789);
nand U9707 (N_9707,N_8875,N_8656);
or U9708 (N_9708,N_8166,N_8839);
nor U9709 (N_9709,N_8696,N_8388);
nor U9710 (N_9710,N_8208,N_8846);
nand U9711 (N_9711,N_8742,N_8638);
and U9712 (N_9712,N_8603,N_8696);
nor U9713 (N_9713,N_8245,N_8165);
or U9714 (N_9714,N_8400,N_8885);
and U9715 (N_9715,N_8831,N_8843);
and U9716 (N_9716,N_8332,N_8601);
or U9717 (N_9717,N_8210,N_8842);
nor U9718 (N_9718,N_8325,N_8985);
nand U9719 (N_9719,N_8802,N_8617);
nor U9720 (N_9720,N_8121,N_8654);
nand U9721 (N_9721,N_8672,N_8279);
or U9722 (N_9722,N_8778,N_8496);
nor U9723 (N_9723,N_8800,N_8967);
nand U9724 (N_9724,N_8674,N_8100);
or U9725 (N_9725,N_8427,N_8787);
xnor U9726 (N_9726,N_8090,N_8302);
or U9727 (N_9727,N_8175,N_8908);
or U9728 (N_9728,N_8743,N_8731);
nand U9729 (N_9729,N_8036,N_8475);
and U9730 (N_9730,N_8174,N_8050);
or U9731 (N_9731,N_8822,N_8101);
or U9732 (N_9732,N_8037,N_8530);
or U9733 (N_9733,N_8294,N_8272);
and U9734 (N_9734,N_8959,N_8370);
or U9735 (N_9735,N_8506,N_8076);
nand U9736 (N_9736,N_8580,N_8517);
nor U9737 (N_9737,N_8898,N_8427);
nor U9738 (N_9738,N_8011,N_8786);
and U9739 (N_9739,N_8240,N_8912);
nor U9740 (N_9740,N_8588,N_8370);
nand U9741 (N_9741,N_8838,N_8310);
and U9742 (N_9742,N_8037,N_8150);
or U9743 (N_9743,N_8927,N_8555);
and U9744 (N_9744,N_8641,N_8719);
nor U9745 (N_9745,N_8636,N_8477);
nand U9746 (N_9746,N_8895,N_8615);
nor U9747 (N_9747,N_8903,N_8306);
or U9748 (N_9748,N_8088,N_8503);
nor U9749 (N_9749,N_8742,N_8099);
or U9750 (N_9750,N_8544,N_8476);
nor U9751 (N_9751,N_8526,N_8810);
and U9752 (N_9752,N_8480,N_8094);
or U9753 (N_9753,N_8066,N_8928);
nand U9754 (N_9754,N_8190,N_8195);
or U9755 (N_9755,N_8635,N_8149);
nor U9756 (N_9756,N_8235,N_8555);
or U9757 (N_9757,N_8116,N_8614);
nand U9758 (N_9758,N_8793,N_8416);
nor U9759 (N_9759,N_8931,N_8523);
or U9760 (N_9760,N_8609,N_8276);
xnor U9761 (N_9761,N_8026,N_8193);
nor U9762 (N_9762,N_8128,N_8706);
and U9763 (N_9763,N_8290,N_8163);
or U9764 (N_9764,N_8908,N_8230);
xnor U9765 (N_9765,N_8715,N_8563);
xnor U9766 (N_9766,N_8607,N_8154);
and U9767 (N_9767,N_8316,N_8046);
nand U9768 (N_9768,N_8644,N_8249);
nor U9769 (N_9769,N_8714,N_8485);
nand U9770 (N_9770,N_8883,N_8428);
and U9771 (N_9771,N_8360,N_8602);
nand U9772 (N_9772,N_8509,N_8468);
nand U9773 (N_9773,N_8318,N_8367);
xor U9774 (N_9774,N_8757,N_8598);
nand U9775 (N_9775,N_8337,N_8022);
and U9776 (N_9776,N_8001,N_8321);
and U9777 (N_9777,N_8915,N_8800);
and U9778 (N_9778,N_8668,N_8653);
and U9779 (N_9779,N_8979,N_8862);
xor U9780 (N_9780,N_8811,N_8656);
nand U9781 (N_9781,N_8155,N_8869);
xor U9782 (N_9782,N_8574,N_8736);
or U9783 (N_9783,N_8452,N_8317);
and U9784 (N_9784,N_8029,N_8433);
nor U9785 (N_9785,N_8828,N_8023);
nor U9786 (N_9786,N_8283,N_8104);
xor U9787 (N_9787,N_8804,N_8139);
nor U9788 (N_9788,N_8076,N_8850);
and U9789 (N_9789,N_8157,N_8394);
nand U9790 (N_9790,N_8488,N_8821);
or U9791 (N_9791,N_8292,N_8150);
or U9792 (N_9792,N_8183,N_8248);
and U9793 (N_9793,N_8187,N_8157);
nor U9794 (N_9794,N_8098,N_8718);
nor U9795 (N_9795,N_8809,N_8731);
and U9796 (N_9796,N_8555,N_8502);
or U9797 (N_9797,N_8402,N_8096);
nand U9798 (N_9798,N_8005,N_8201);
or U9799 (N_9799,N_8727,N_8705);
nand U9800 (N_9800,N_8236,N_8277);
and U9801 (N_9801,N_8798,N_8714);
or U9802 (N_9802,N_8386,N_8989);
and U9803 (N_9803,N_8341,N_8673);
or U9804 (N_9804,N_8012,N_8283);
xnor U9805 (N_9805,N_8156,N_8556);
or U9806 (N_9806,N_8101,N_8325);
and U9807 (N_9807,N_8125,N_8946);
nor U9808 (N_9808,N_8151,N_8032);
and U9809 (N_9809,N_8038,N_8412);
nand U9810 (N_9810,N_8672,N_8271);
nand U9811 (N_9811,N_8989,N_8953);
nand U9812 (N_9812,N_8243,N_8503);
nor U9813 (N_9813,N_8404,N_8327);
nand U9814 (N_9814,N_8695,N_8151);
nand U9815 (N_9815,N_8351,N_8222);
nor U9816 (N_9816,N_8477,N_8154);
nand U9817 (N_9817,N_8074,N_8685);
or U9818 (N_9818,N_8583,N_8366);
or U9819 (N_9819,N_8669,N_8861);
nor U9820 (N_9820,N_8303,N_8854);
and U9821 (N_9821,N_8945,N_8409);
xor U9822 (N_9822,N_8458,N_8102);
nand U9823 (N_9823,N_8594,N_8840);
nand U9824 (N_9824,N_8001,N_8936);
nand U9825 (N_9825,N_8109,N_8954);
nand U9826 (N_9826,N_8803,N_8127);
nor U9827 (N_9827,N_8188,N_8370);
nor U9828 (N_9828,N_8812,N_8922);
nand U9829 (N_9829,N_8456,N_8652);
nor U9830 (N_9830,N_8713,N_8515);
nor U9831 (N_9831,N_8949,N_8497);
nor U9832 (N_9832,N_8952,N_8505);
nand U9833 (N_9833,N_8530,N_8414);
and U9834 (N_9834,N_8275,N_8464);
nor U9835 (N_9835,N_8836,N_8803);
nor U9836 (N_9836,N_8934,N_8945);
nor U9837 (N_9837,N_8954,N_8158);
nor U9838 (N_9838,N_8352,N_8059);
and U9839 (N_9839,N_8622,N_8898);
nand U9840 (N_9840,N_8613,N_8694);
and U9841 (N_9841,N_8151,N_8578);
and U9842 (N_9842,N_8834,N_8012);
nor U9843 (N_9843,N_8258,N_8828);
or U9844 (N_9844,N_8090,N_8149);
nand U9845 (N_9845,N_8770,N_8510);
xnor U9846 (N_9846,N_8625,N_8321);
nand U9847 (N_9847,N_8476,N_8190);
and U9848 (N_9848,N_8227,N_8782);
nor U9849 (N_9849,N_8364,N_8177);
and U9850 (N_9850,N_8978,N_8268);
nand U9851 (N_9851,N_8580,N_8978);
and U9852 (N_9852,N_8109,N_8936);
nor U9853 (N_9853,N_8825,N_8755);
nand U9854 (N_9854,N_8353,N_8667);
nor U9855 (N_9855,N_8704,N_8396);
and U9856 (N_9856,N_8459,N_8284);
or U9857 (N_9857,N_8754,N_8455);
xor U9858 (N_9858,N_8092,N_8372);
nor U9859 (N_9859,N_8902,N_8926);
and U9860 (N_9860,N_8857,N_8497);
or U9861 (N_9861,N_8378,N_8228);
and U9862 (N_9862,N_8956,N_8912);
and U9863 (N_9863,N_8820,N_8463);
xor U9864 (N_9864,N_8751,N_8847);
or U9865 (N_9865,N_8925,N_8399);
nand U9866 (N_9866,N_8914,N_8145);
and U9867 (N_9867,N_8006,N_8602);
and U9868 (N_9868,N_8050,N_8396);
nand U9869 (N_9869,N_8511,N_8458);
or U9870 (N_9870,N_8115,N_8955);
nand U9871 (N_9871,N_8272,N_8812);
and U9872 (N_9872,N_8086,N_8638);
nor U9873 (N_9873,N_8020,N_8446);
xor U9874 (N_9874,N_8093,N_8226);
nand U9875 (N_9875,N_8077,N_8250);
nor U9876 (N_9876,N_8294,N_8345);
or U9877 (N_9877,N_8484,N_8775);
nor U9878 (N_9878,N_8311,N_8944);
nor U9879 (N_9879,N_8490,N_8494);
nand U9880 (N_9880,N_8717,N_8856);
nor U9881 (N_9881,N_8605,N_8059);
or U9882 (N_9882,N_8004,N_8698);
or U9883 (N_9883,N_8432,N_8852);
nor U9884 (N_9884,N_8106,N_8662);
nand U9885 (N_9885,N_8507,N_8155);
nand U9886 (N_9886,N_8784,N_8555);
nor U9887 (N_9887,N_8584,N_8194);
xor U9888 (N_9888,N_8921,N_8897);
and U9889 (N_9889,N_8191,N_8630);
and U9890 (N_9890,N_8437,N_8933);
xnor U9891 (N_9891,N_8583,N_8378);
nand U9892 (N_9892,N_8767,N_8680);
xnor U9893 (N_9893,N_8824,N_8583);
or U9894 (N_9894,N_8356,N_8299);
or U9895 (N_9895,N_8765,N_8536);
nand U9896 (N_9896,N_8965,N_8421);
nand U9897 (N_9897,N_8988,N_8721);
and U9898 (N_9898,N_8154,N_8553);
or U9899 (N_9899,N_8503,N_8738);
or U9900 (N_9900,N_8128,N_8496);
nor U9901 (N_9901,N_8193,N_8062);
and U9902 (N_9902,N_8965,N_8625);
nand U9903 (N_9903,N_8609,N_8320);
and U9904 (N_9904,N_8378,N_8109);
and U9905 (N_9905,N_8646,N_8670);
and U9906 (N_9906,N_8412,N_8683);
and U9907 (N_9907,N_8199,N_8176);
nand U9908 (N_9908,N_8820,N_8124);
nand U9909 (N_9909,N_8829,N_8098);
nand U9910 (N_9910,N_8188,N_8517);
nor U9911 (N_9911,N_8790,N_8719);
nand U9912 (N_9912,N_8971,N_8236);
nand U9913 (N_9913,N_8806,N_8229);
nand U9914 (N_9914,N_8692,N_8591);
xor U9915 (N_9915,N_8823,N_8635);
nor U9916 (N_9916,N_8683,N_8164);
nand U9917 (N_9917,N_8259,N_8989);
nor U9918 (N_9918,N_8324,N_8293);
xnor U9919 (N_9919,N_8656,N_8962);
or U9920 (N_9920,N_8607,N_8202);
nand U9921 (N_9921,N_8056,N_8321);
nor U9922 (N_9922,N_8680,N_8786);
nand U9923 (N_9923,N_8388,N_8319);
nand U9924 (N_9924,N_8005,N_8862);
nor U9925 (N_9925,N_8616,N_8698);
nand U9926 (N_9926,N_8724,N_8472);
and U9927 (N_9927,N_8462,N_8399);
nand U9928 (N_9928,N_8728,N_8422);
nand U9929 (N_9929,N_8257,N_8967);
and U9930 (N_9930,N_8710,N_8899);
nand U9931 (N_9931,N_8923,N_8326);
or U9932 (N_9932,N_8911,N_8455);
or U9933 (N_9933,N_8221,N_8347);
xor U9934 (N_9934,N_8430,N_8630);
or U9935 (N_9935,N_8261,N_8710);
xnor U9936 (N_9936,N_8081,N_8513);
nor U9937 (N_9937,N_8911,N_8049);
and U9938 (N_9938,N_8343,N_8930);
nor U9939 (N_9939,N_8272,N_8171);
or U9940 (N_9940,N_8408,N_8374);
nor U9941 (N_9941,N_8586,N_8424);
nor U9942 (N_9942,N_8160,N_8253);
and U9943 (N_9943,N_8334,N_8251);
nor U9944 (N_9944,N_8572,N_8523);
or U9945 (N_9945,N_8264,N_8016);
or U9946 (N_9946,N_8790,N_8839);
or U9947 (N_9947,N_8645,N_8538);
nand U9948 (N_9948,N_8618,N_8960);
and U9949 (N_9949,N_8196,N_8238);
nor U9950 (N_9950,N_8853,N_8560);
nand U9951 (N_9951,N_8078,N_8892);
or U9952 (N_9952,N_8173,N_8883);
nor U9953 (N_9953,N_8866,N_8505);
or U9954 (N_9954,N_8588,N_8047);
or U9955 (N_9955,N_8585,N_8426);
nor U9956 (N_9956,N_8469,N_8594);
or U9957 (N_9957,N_8873,N_8409);
or U9958 (N_9958,N_8013,N_8966);
nand U9959 (N_9959,N_8535,N_8777);
and U9960 (N_9960,N_8473,N_8671);
nand U9961 (N_9961,N_8071,N_8525);
or U9962 (N_9962,N_8227,N_8547);
nor U9963 (N_9963,N_8614,N_8813);
and U9964 (N_9964,N_8878,N_8617);
nor U9965 (N_9965,N_8733,N_8088);
and U9966 (N_9966,N_8482,N_8712);
nor U9967 (N_9967,N_8555,N_8868);
nor U9968 (N_9968,N_8469,N_8331);
and U9969 (N_9969,N_8470,N_8235);
and U9970 (N_9970,N_8520,N_8768);
nor U9971 (N_9971,N_8821,N_8024);
nor U9972 (N_9972,N_8196,N_8795);
nor U9973 (N_9973,N_8571,N_8689);
nand U9974 (N_9974,N_8682,N_8149);
or U9975 (N_9975,N_8207,N_8197);
and U9976 (N_9976,N_8338,N_8208);
nor U9977 (N_9977,N_8122,N_8299);
and U9978 (N_9978,N_8933,N_8097);
nor U9979 (N_9979,N_8719,N_8290);
nor U9980 (N_9980,N_8709,N_8500);
and U9981 (N_9981,N_8066,N_8039);
nand U9982 (N_9982,N_8001,N_8793);
and U9983 (N_9983,N_8862,N_8635);
nand U9984 (N_9984,N_8428,N_8696);
nor U9985 (N_9985,N_8007,N_8917);
and U9986 (N_9986,N_8189,N_8567);
nand U9987 (N_9987,N_8695,N_8862);
or U9988 (N_9988,N_8844,N_8812);
or U9989 (N_9989,N_8991,N_8137);
and U9990 (N_9990,N_8128,N_8072);
nand U9991 (N_9991,N_8739,N_8887);
or U9992 (N_9992,N_8940,N_8749);
xnor U9993 (N_9993,N_8742,N_8320);
or U9994 (N_9994,N_8671,N_8348);
or U9995 (N_9995,N_8649,N_8106);
and U9996 (N_9996,N_8479,N_8632);
or U9997 (N_9997,N_8174,N_8991);
and U9998 (N_9998,N_8049,N_8805);
nand U9999 (N_9999,N_8765,N_8547);
xor UO_0 (O_0,N_9997,N_9789);
nand UO_1 (O_1,N_9173,N_9960);
nor UO_2 (O_2,N_9659,N_9594);
nand UO_3 (O_3,N_9549,N_9236);
and UO_4 (O_4,N_9274,N_9810);
nor UO_5 (O_5,N_9668,N_9928);
nor UO_6 (O_6,N_9673,N_9772);
or UO_7 (O_7,N_9692,N_9033);
and UO_8 (O_8,N_9003,N_9342);
xor UO_9 (O_9,N_9022,N_9749);
or UO_10 (O_10,N_9219,N_9848);
nor UO_11 (O_11,N_9183,N_9199);
nor UO_12 (O_12,N_9311,N_9457);
or UO_13 (O_13,N_9462,N_9717);
and UO_14 (O_14,N_9374,N_9017);
or UO_15 (O_15,N_9840,N_9704);
and UO_16 (O_16,N_9460,N_9028);
nor UO_17 (O_17,N_9043,N_9114);
xor UO_18 (O_18,N_9417,N_9331);
nor UO_19 (O_19,N_9349,N_9925);
or UO_20 (O_20,N_9228,N_9874);
nor UO_21 (O_21,N_9786,N_9634);
or UO_22 (O_22,N_9011,N_9646);
xnor UO_23 (O_23,N_9871,N_9447);
or UO_24 (O_24,N_9888,N_9841);
nand UO_25 (O_25,N_9034,N_9525);
and UO_26 (O_26,N_9446,N_9718);
nor UO_27 (O_27,N_9843,N_9314);
and UO_28 (O_28,N_9640,N_9522);
or UO_29 (O_29,N_9320,N_9651);
and UO_30 (O_30,N_9328,N_9542);
or UO_31 (O_31,N_9935,N_9357);
nand UO_32 (O_32,N_9152,N_9687);
and UO_33 (O_33,N_9852,N_9790);
or UO_34 (O_34,N_9570,N_9279);
nor UO_35 (O_35,N_9067,N_9587);
or UO_36 (O_36,N_9760,N_9260);
or UO_37 (O_37,N_9965,N_9423);
nor UO_38 (O_38,N_9834,N_9283);
or UO_39 (O_39,N_9915,N_9376);
nand UO_40 (O_40,N_9861,N_9978);
and UO_41 (O_41,N_9176,N_9050);
and UO_42 (O_42,N_9383,N_9139);
or UO_43 (O_43,N_9675,N_9591);
nor UO_44 (O_44,N_9637,N_9577);
or UO_45 (O_45,N_9348,N_9102);
and UO_46 (O_46,N_9459,N_9837);
or UO_47 (O_47,N_9836,N_9911);
nand UO_48 (O_48,N_9905,N_9649);
nor UO_49 (O_49,N_9906,N_9481);
nand UO_50 (O_50,N_9574,N_9647);
nor UO_51 (O_51,N_9268,N_9652);
xnor UO_52 (O_52,N_9338,N_9739);
xnor UO_53 (O_53,N_9742,N_9509);
or UO_54 (O_54,N_9293,N_9734);
and UO_55 (O_55,N_9927,N_9347);
nor UO_56 (O_56,N_9444,N_9467);
nor UO_57 (O_57,N_9100,N_9166);
xnor UO_58 (O_58,N_9977,N_9626);
xor UO_59 (O_59,N_9958,N_9341);
nor UO_60 (O_60,N_9014,N_9711);
nor UO_61 (O_61,N_9614,N_9916);
nor UO_62 (O_62,N_9396,N_9878);
or UO_63 (O_63,N_9815,N_9390);
and UO_64 (O_64,N_9060,N_9126);
xor UO_65 (O_65,N_9974,N_9129);
and UO_66 (O_66,N_9572,N_9294);
or UO_67 (O_67,N_9719,N_9002);
xor UO_68 (O_68,N_9024,N_9650);
and UO_69 (O_69,N_9197,N_9732);
or UO_70 (O_70,N_9846,N_9431);
nand UO_71 (O_71,N_9523,N_9451);
and UO_72 (O_72,N_9504,N_9681);
nand UO_73 (O_73,N_9812,N_9910);
nand UO_74 (O_74,N_9330,N_9220);
and UO_75 (O_75,N_9486,N_9241);
xor UO_76 (O_76,N_9370,N_9122);
nor UO_77 (O_77,N_9606,N_9566);
nor UO_78 (O_78,N_9146,N_9098);
nor UO_79 (O_79,N_9356,N_9086);
nand UO_80 (O_80,N_9669,N_9271);
xnor UO_81 (O_81,N_9720,N_9365);
and UO_82 (O_82,N_9782,N_9585);
nand UO_83 (O_83,N_9078,N_9691);
and UO_84 (O_84,N_9121,N_9496);
xnor UO_85 (O_85,N_9829,N_9851);
or UO_86 (O_86,N_9391,N_9855);
and UO_87 (O_87,N_9619,N_9821);
nand UO_88 (O_88,N_9303,N_9252);
or UO_89 (O_89,N_9027,N_9420);
xnor UO_90 (O_90,N_9477,N_9571);
xor UO_91 (O_91,N_9545,N_9339);
nor UO_92 (O_92,N_9699,N_9666);
nor UO_93 (O_93,N_9218,N_9991);
and UO_94 (O_94,N_9985,N_9941);
nand UO_95 (O_95,N_9913,N_9520);
nor UO_96 (O_96,N_9546,N_9018);
or UO_97 (O_97,N_9233,N_9180);
nor UO_98 (O_98,N_9528,N_9979);
nand UO_99 (O_99,N_9280,N_9893);
nand UO_100 (O_100,N_9601,N_9072);
nand UO_101 (O_101,N_9042,N_9517);
or UO_102 (O_102,N_9230,N_9285);
or UO_103 (O_103,N_9982,N_9284);
nor UO_104 (O_104,N_9748,N_9111);
or UO_105 (O_105,N_9468,N_9278);
and UO_106 (O_106,N_9456,N_9701);
or UO_107 (O_107,N_9209,N_9149);
and UO_108 (O_108,N_9151,N_9275);
nand UO_109 (O_109,N_9682,N_9804);
and UO_110 (O_110,N_9108,N_9992);
and UO_111 (O_111,N_9671,N_9531);
and UO_112 (O_112,N_9883,N_9707);
or UO_113 (O_113,N_9886,N_9296);
nor UO_114 (O_114,N_9784,N_9377);
nor UO_115 (O_115,N_9071,N_9793);
and UO_116 (O_116,N_9565,N_9696);
nand UO_117 (O_117,N_9697,N_9205);
and UO_118 (O_118,N_9973,N_9448);
and UO_119 (O_119,N_9737,N_9224);
nand UO_120 (O_120,N_9094,N_9360);
xor UO_121 (O_121,N_9740,N_9074);
nor UO_122 (O_122,N_9187,N_9505);
nand UO_123 (O_123,N_9493,N_9385);
nor UO_124 (O_124,N_9966,N_9632);
nand UO_125 (O_125,N_9990,N_9381);
nor UO_126 (O_126,N_9140,N_9947);
nor UO_127 (O_127,N_9788,N_9196);
nor UO_128 (O_128,N_9487,N_9475);
nor UO_129 (O_129,N_9195,N_9970);
nand UO_130 (O_130,N_9324,N_9488);
and UO_131 (O_131,N_9787,N_9639);
xor UO_132 (O_132,N_9256,N_9138);
nand UO_133 (O_133,N_9511,N_9688);
or UO_134 (O_134,N_9779,N_9471);
and UO_135 (O_135,N_9313,N_9708);
nor UO_136 (O_136,N_9246,N_9052);
nor UO_137 (O_137,N_9576,N_9750);
nor UO_138 (O_138,N_9802,N_9445);
or UO_139 (O_139,N_9744,N_9474);
or UO_140 (O_140,N_9845,N_9534);
nor UO_141 (O_141,N_9627,N_9590);
or UO_142 (O_142,N_9610,N_9255);
nor UO_143 (O_143,N_9858,N_9876);
or UO_144 (O_144,N_9679,N_9604);
nand UO_145 (O_145,N_9473,N_9062);
and UO_146 (O_146,N_9579,N_9661);
or UO_147 (O_147,N_9729,N_9560);
or UO_148 (O_148,N_9461,N_9118);
nor UO_149 (O_149,N_9856,N_9388);
and UO_150 (O_150,N_9521,N_9235);
xor UO_151 (O_151,N_9794,N_9269);
or UO_152 (O_152,N_9117,N_9115);
or UO_153 (O_153,N_9956,N_9880);
or UO_154 (O_154,N_9434,N_9158);
or UO_155 (O_155,N_9077,N_9645);
and UO_156 (O_156,N_9103,N_9045);
xnor UO_157 (O_157,N_9367,N_9380);
nor UO_158 (O_158,N_9919,N_9685);
and UO_159 (O_159,N_9409,N_9144);
xnor UO_160 (O_160,N_9148,N_9055);
or UO_161 (O_161,N_9624,N_9395);
or UO_162 (O_162,N_9999,N_9672);
or UO_163 (O_163,N_9405,N_9818);
or UO_164 (O_164,N_9684,N_9472);
or UO_165 (O_165,N_9644,N_9502);
xor UO_166 (O_166,N_9896,N_9286);
or UO_167 (O_167,N_9642,N_9184);
xor UO_168 (O_168,N_9948,N_9512);
or UO_169 (O_169,N_9809,N_9242);
and UO_170 (O_170,N_9070,N_9245);
nand UO_171 (O_171,N_9301,N_9312);
nor UO_172 (O_172,N_9427,N_9993);
xor UO_173 (O_173,N_9581,N_9706);
or UO_174 (O_174,N_9305,N_9657);
nand UO_175 (O_175,N_9860,N_9690);
xor UO_176 (O_176,N_9930,N_9325);
nand UO_177 (O_177,N_9389,N_9302);
or UO_178 (O_178,N_9082,N_9101);
nor UO_179 (O_179,N_9298,N_9145);
or UO_180 (O_180,N_9938,N_9617);
nand UO_181 (O_181,N_9902,N_9127);
nand UO_182 (O_182,N_9253,N_9518);
or UO_183 (O_183,N_9605,N_9698);
or UO_184 (O_184,N_9636,N_9728);
nand UO_185 (O_185,N_9232,N_9559);
and UO_186 (O_186,N_9163,N_9250);
nand UO_187 (O_187,N_9819,N_9498);
nand UO_188 (O_188,N_9125,N_9863);
and UO_189 (O_189,N_9934,N_9227);
nor UO_190 (O_190,N_9988,N_9808);
nor UO_191 (O_191,N_9214,N_9020);
and UO_192 (O_192,N_9774,N_9937);
and UO_193 (O_193,N_9226,N_9393);
and UO_194 (O_194,N_9641,N_9375);
and UO_195 (O_195,N_9678,N_9693);
nor UO_196 (O_196,N_9484,N_9048);
nand UO_197 (O_197,N_9709,N_9827);
and UO_198 (O_198,N_9894,N_9918);
xnor UO_199 (O_199,N_9746,N_9695);
xnor UO_200 (O_200,N_9010,N_9519);
nor UO_201 (O_201,N_9004,N_9000);
or UO_202 (O_202,N_9854,N_9986);
xor UO_203 (O_203,N_9954,N_9398);
or UO_204 (O_204,N_9607,N_9862);
nor UO_205 (O_205,N_9038,N_9142);
and UO_206 (O_206,N_9914,N_9277);
nor UO_207 (O_207,N_9623,N_9191);
nand UO_208 (O_208,N_9318,N_9066);
and UO_209 (O_209,N_9217,N_9713);
nor UO_210 (O_210,N_9628,N_9677);
nand UO_211 (O_211,N_9552,N_9160);
xnor UO_212 (O_212,N_9442,N_9508);
nor UO_213 (O_213,N_9538,N_9154);
nand UO_214 (O_214,N_9676,N_9539);
nand UO_215 (O_215,N_9814,N_9130);
xnor UO_216 (O_216,N_9440,N_9540);
and UO_217 (O_217,N_9295,N_9363);
or UO_218 (O_218,N_9785,N_9135);
nor UO_219 (O_219,N_9105,N_9767);
and UO_220 (O_220,N_9537,N_9795);
and UO_221 (O_221,N_9109,N_9890);
or UO_222 (O_222,N_9733,N_9306);
nand UO_223 (O_223,N_9407,N_9482);
nand UO_224 (O_224,N_9562,N_9007);
and UO_225 (O_225,N_9912,N_9612);
xor UO_226 (O_226,N_9797,N_9063);
nand UO_227 (O_227,N_9200,N_9247);
nand UO_228 (O_228,N_9813,N_9806);
nand UO_229 (O_229,N_9575,N_9929);
nand UO_230 (O_230,N_9736,N_9611);
and UO_231 (O_231,N_9037,N_9238);
nand UO_232 (O_232,N_9476,N_9332);
nand UO_233 (O_233,N_9944,N_9506);
nor UO_234 (O_234,N_9408,N_9132);
nor UO_235 (O_235,N_9887,N_9454);
and UO_236 (O_236,N_9384,N_9006);
and UO_237 (O_237,N_9198,N_9157);
or UO_238 (O_238,N_9485,N_9465);
nand UO_239 (O_239,N_9258,N_9625);
nand UO_240 (O_240,N_9942,N_9656);
and UO_241 (O_241,N_9980,N_9541);
nor UO_242 (O_242,N_9621,N_9399);
nor UO_243 (O_243,N_9207,N_9831);
nor UO_244 (O_244,N_9583,N_9291);
and UO_245 (O_245,N_9382,N_9658);
and UO_246 (O_246,N_9175,N_9470);
and UO_247 (O_247,N_9922,N_9087);
nor UO_248 (O_248,N_9620,N_9327);
nand UO_249 (O_249,N_9188,N_9865);
or UO_250 (O_250,N_9240,N_9853);
or UO_251 (O_251,N_9609,N_9613);
and UO_252 (O_252,N_9364,N_9346);
and UO_253 (O_253,N_9753,N_9174);
and UO_254 (O_254,N_9273,N_9875);
nor UO_255 (O_255,N_9397,N_9436);
and UO_256 (O_256,N_9563,N_9449);
nor UO_257 (O_257,N_9901,N_9113);
and UO_258 (O_258,N_9595,N_9780);
or UO_259 (O_259,N_9768,N_9680);
xor UO_260 (O_260,N_9297,N_9165);
or UO_261 (O_261,N_9859,N_9439);
xor UO_262 (O_262,N_9081,N_9730);
nand UO_263 (O_263,N_9532,N_9257);
nor UO_264 (O_264,N_9016,N_9317);
and UO_265 (O_265,N_9403,N_9618);
and UO_266 (O_266,N_9336,N_9172);
and UO_267 (O_267,N_9694,N_9047);
or UO_268 (O_268,N_9820,N_9653);
nand UO_269 (O_269,N_9603,N_9769);
xor UO_270 (O_270,N_9764,N_9839);
nand UO_271 (O_271,N_9091,N_9833);
nor UO_272 (O_272,N_9757,N_9061);
nor UO_273 (O_273,N_9872,N_9869);
or UO_274 (O_274,N_9097,N_9478);
nand UO_275 (O_275,N_9288,N_9358);
nor UO_276 (O_276,N_9727,N_9259);
and UO_277 (O_277,N_9355,N_9322);
or UO_278 (O_278,N_9029,N_9190);
and UO_279 (O_279,N_9775,N_9394);
nand UO_280 (O_280,N_9321,N_9128);
and UO_281 (O_281,N_9410,N_9781);
and UO_282 (O_282,N_9501,N_9580);
nor UO_283 (O_283,N_9281,N_9326);
nor UO_284 (O_284,N_9073,N_9044);
or UO_285 (O_285,N_9527,N_9971);
nor UO_286 (O_286,N_9714,N_9892);
nand UO_287 (O_287,N_9307,N_9369);
nor UO_288 (O_288,N_9805,N_9400);
and UO_289 (O_289,N_9137,N_9134);
nand UO_290 (O_290,N_9756,N_9084);
nor UO_291 (O_291,N_9304,N_9968);
xor UO_292 (O_292,N_9438,N_9012);
xnor UO_293 (O_293,N_9529,N_9556);
and UO_294 (O_294,N_9582,N_9558);
xor UO_295 (O_295,N_9939,N_9530);
xor UO_296 (O_296,N_9169,N_9089);
nor UO_297 (O_297,N_9870,N_9555);
nor UO_298 (O_298,N_9674,N_9231);
or UO_299 (O_299,N_9751,N_9334);
xor UO_300 (O_300,N_9263,N_9243);
and UO_301 (O_301,N_9368,N_9287);
and UO_302 (O_302,N_9013,N_9867);
or UO_303 (O_303,N_9588,N_9026);
or UO_304 (O_304,N_9994,N_9616);
and UO_305 (O_305,N_9879,N_9093);
and UO_306 (O_306,N_9497,N_9608);
and UO_307 (O_307,N_9762,N_9435);
and UO_308 (O_308,N_9664,N_9510);
nand UO_309 (O_309,N_9857,N_9201);
xor UO_310 (O_310,N_9755,N_9747);
nor UO_311 (O_311,N_9957,N_9386);
nand UO_312 (O_312,N_9904,N_9466);
or UO_313 (O_313,N_9758,N_9340);
or UO_314 (O_314,N_9526,N_9424);
nand UO_315 (O_315,N_9513,N_9335);
and UO_316 (O_316,N_9112,N_9412);
xor UO_317 (O_317,N_9453,N_9725);
and UO_318 (O_318,N_9310,N_9107);
nand UO_319 (O_319,N_9773,N_9898);
nor UO_320 (O_320,N_9864,N_9907);
nand UO_321 (O_321,N_9343,N_9373);
and UO_322 (O_322,N_9500,N_9547);
nand UO_323 (O_323,N_9212,N_9766);
or UO_324 (O_324,N_9299,N_9266);
nor UO_325 (O_325,N_9463,N_9602);
and UO_326 (O_326,N_9244,N_9437);
and UO_327 (O_327,N_9031,N_9975);
and UO_328 (O_328,N_9761,N_9536);
nor UO_329 (O_329,N_9554,N_9503);
nand UO_330 (O_330,N_9079,N_9792);
nor UO_331 (O_331,N_9983,N_9203);
nor UO_332 (O_332,N_9933,N_9164);
and UO_333 (O_333,N_9159,N_9741);
xor UO_334 (O_334,N_9516,N_9705);
xor UO_335 (O_335,N_9884,N_9300);
xor UO_336 (O_336,N_9450,N_9036);
nor UO_337 (O_337,N_9700,N_9202);
and UO_338 (O_338,N_9359,N_9249);
xnor UO_339 (O_339,N_9216,N_9800);
nor UO_340 (O_340,N_9835,N_9080);
nor UO_341 (O_341,N_9032,N_9229);
nor UO_342 (O_342,N_9830,N_9458);
nand UO_343 (O_343,N_9589,N_9251);
and UO_344 (O_344,N_9309,N_9411);
xor UO_345 (O_345,N_9593,N_9168);
xor UO_346 (O_346,N_9262,N_9239);
nand UO_347 (O_347,N_9738,N_9936);
nand UO_348 (O_348,N_9660,N_9561);
or UO_349 (O_349,N_9989,N_9945);
or UO_350 (O_350,N_9670,N_9655);
nor UO_351 (O_351,N_9881,N_9816);
or UO_352 (O_352,N_9065,N_9025);
nor UO_353 (O_353,N_9131,N_9019);
and UO_354 (O_354,N_9584,N_9123);
or UO_355 (O_355,N_9931,N_9972);
xor UO_356 (O_356,N_9432,N_9665);
nand UO_357 (O_357,N_9254,N_9596);
or UO_358 (O_358,N_9054,N_9419);
nand UO_359 (O_359,N_9030,N_9564);
nor UO_360 (O_360,N_9119,N_9801);
nor UO_361 (O_361,N_9282,N_9726);
nand UO_362 (O_362,N_9351,N_9039);
and UO_363 (O_363,N_9177,N_9599);
or UO_364 (O_364,N_9426,N_9413);
and UO_365 (O_365,N_9452,N_9551);
nor UO_366 (O_366,N_9223,N_9807);
and UO_367 (O_367,N_9323,N_9959);
and UO_368 (O_368,N_9068,N_9008);
nand UO_369 (O_369,N_9631,N_9569);
nand UO_370 (O_370,N_9686,N_9416);
nor UO_371 (O_371,N_9663,N_9316);
nor UO_372 (O_372,N_9237,N_9156);
nand UO_373 (O_373,N_9104,N_9885);
or UO_374 (O_374,N_9362,N_9735);
and UO_375 (O_375,N_9133,N_9425);
nor UO_376 (O_376,N_9832,N_9791);
and UO_377 (O_377,N_9897,N_9315);
nor UO_378 (O_378,N_9361,N_9194);
and UO_379 (O_379,N_9041,N_9514);
nand UO_380 (O_380,N_9162,N_9290);
or UO_381 (O_381,N_9076,N_9265);
nand UO_382 (O_382,N_9868,N_9882);
and UO_383 (O_383,N_9120,N_9329);
xor UO_384 (O_384,N_9096,N_9058);
nand UO_385 (O_385,N_9703,N_9206);
nor UO_386 (O_386,N_9745,N_9548);
nor UO_387 (O_387,N_9951,N_9147);
or UO_388 (O_388,N_9005,N_9193);
nand UO_389 (O_389,N_9056,N_9192);
or UO_390 (O_390,N_9629,N_9778);
nor UO_391 (O_391,N_9415,N_9981);
nor UO_392 (O_392,N_9181,N_9850);
xor UO_393 (O_393,N_9143,N_9721);
or UO_394 (O_394,N_9387,N_9333);
nand UO_395 (O_395,N_9900,N_9889);
xnor UO_396 (O_396,N_9917,N_9507);
and UO_397 (O_397,N_9568,N_9185);
xor UO_398 (O_398,N_9689,N_9578);
nor UO_399 (O_399,N_9213,N_9155);
nand UO_400 (O_400,N_9150,N_9754);
and UO_401 (O_401,N_9178,N_9702);
nor UO_402 (O_402,N_9515,N_9350);
nor UO_403 (O_403,N_9354,N_9838);
nand UO_404 (O_404,N_9116,N_9844);
or UO_405 (O_405,N_9492,N_9998);
nand UO_406 (O_406,N_9035,N_9489);
nor UO_407 (O_407,N_9464,N_9828);
or UO_408 (O_408,N_9001,N_9811);
and UO_409 (O_409,N_9204,N_9099);
nor UO_410 (O_410,N_9716,N_9171);
or UO_411 (O_411,N_9866,N_9428);
nor UO_412 (O_412,N_9783,N_9963);
nand UO_413 (O_413,N_9996,N_9987);
nand UO_414 (O_414,N_9633,N_9479);
nand UO_415 (O_415,N_9480,N_9319);
or UO_416 (O_416,N_9049,N_9490);
and UO_417 (O_417,N_9345,N_9270);
nand UO_418 (O_418,N_9776,N_9952);
and UO_419 (O_419,N_9352,N_9847);
and UO_420 (O_420,N_9976,N_9940);
nand UO_421 (O_421,N_9946,N_9524);
or UO_422 (O_422,N_9234,N_9095);
nor UO_423 (O_423,N_9635,N_9943);
or UO_424 (O_424,N_9189,N_9378);
or UO_425 (O_425,N_9494,N_9110);
nor UO_426 (O_426,N_9553,N_9731);
or UO_427 (O_427,N_9153,N_9923);
nand UO_428 (O_428,N_9069,N_9995);
or UO_429 (O_429,N_9124,N_9433);
nand UO_430 (O_430,N_9372,N_9950);
or UO_431 (O_431,N_9215,N_9088);
nand UO_432 (O_432,N_9170,N_9418);
nor UO_433 (O_433,N_9822,N_9873);
nand UO_434 (O_434,N_9483,N_9429);
and UO_435 (O_435,N_9495,N_9877);
or UO_436 (O_436,N_9899,N_9292);
nand UO_437 (O_437,N_9353,N_9366);
and UO_438 (O_438,N_9961,N_9763);
nand UO_439 (O_439,N_9092,N_9722);
or UO_440 (O_440,N_9926,N_9908);
or UO_441 (O_441,N_9752,N_9799);
nand UO_442 (O_442,N_9046,N_9337);
nand UO_443 (O_443,N_9955,N_9499);
nor UO_444 (O_444,N_9909,N_9075);
or UO_445 (O_445,N_9535,N_9264);
nand UO_446 (O_446,N_9825,N_9040);
and UO_447 (O_447,N_9964,N_9622);
or UO_448 (O_448,N_9712,N_9106);
nand UO_449 (O_449,N_9064,N_9225);
nor UO_450 (O_450,N_9683,N_9550);
and UO_451 (O_451,N_9969,N_9422);
and UO_452 (O_452,N_9598,N_9638);
or UO_453 (O_453,N_9021,N_9267);
or UO_454 (O_454,N_9289,N_9059);
and UO_455 (O_455,N_9272,N_9803);
nor UO_456 (O_456,N_9404,N_9765);
nor UO_457 (O_457,N_9724,N_9573);
or UO_458 (O_458,N_9441,N_9891);
nand UO_459 (O_459,N_9557,N_9932);
nor UO_460 (O_460,N_9469,N_9308);
or UO_461 (O_461,N_9167,N_9743);
nand UO_462 (O_462,N_9085,N_9600);
nor UO_463 (O_463,N_9491,N_9715);
nor UO_464 (O_464,N_9015,N_9222);
nand UO_465 (O_465,N_9210,N_9371);
or UO_466 (O_466,N_9083,N_9903);
or UO_467 (O_467,N_9920,N_9051);
nand UO_468 (O_468,N_9009,N_9406);
or UO_469 (O_469,N_9824,N_9895);
and UO_470 (O_470,N_9344,N_9953);
xor UO_471 (O_471,N_9967,N_9261);
nor UO_472 (O_472,N_9842,N_9161);
nor UO_473 (O_473,N_9023,N_9796);
and UO_474 (O_474,N_9455,N_9592);
nand UO_475 (O_475,N_9248,N_9777);
xor UO_476 (O_476,N_9379,N_9544);
or UO_477 (O_477,N_9533,N_9392);
and UO_478 (O_478,N_9141,N_9276);
nand UO_479 (O_479,N_9136,N_9962);
or UO_480 (O_480,N_9543,N_9401);
xor UO_481 (O_481,N_9654,N_9211);
or UO_482 (O_482,N_9182,N_9402);
and UO_483 (O_483,N_9924,N_9759);
or UO_484 (O_484,N_9771,N_9817);
and UO_485 (O_485,N_9823,N_9723);
or UO_486 (O_486,N_9648,N_9949);
nand UO_487 (O_487,N_9615,N_9826);
and UO_488 (O_488,N_9443,N_9179);
nor UO_489 (O_489,N_9798,N_9643);
or UO_490 (O_490,N_9053,N_9662);
or UO_491 (O_491,N_9090,N_9630);
nor UO_492 (O_492,N_9057,N_9921);
nor UO_493 (O_493,N_9770,N_9567);
and UO_494 (O_494,N_9208,N_9597);
and UO_495 (O_495,N_9849,N_9667);
nand UO_496 (O_496,N_9186,N_9414);
or UO_497 (O_497,N_9984,N_9710);
or UO_498 (O_498,N_9586,N_9421);
nand UO_499 (O_499,N_9221,N_9430);
and UO_500 (O_500,N_9449,N_9020);
nand UO_501 (O_501,N_9159,N_9393);
xnor UO_502 (O_502,N_9297,N_9905);
nand UO_503 (O_503,N_9377,N_9836);
nor UO_504 (O_504,N_9183,N_9763);
nor UO_505 (O_505,N_9794,N_9539);
and UO_506 (O_506,N_9586,N_9232);
nor UO_507 (O_507,N_9561,N_9158);
nor UO_508 (O_508,N_9376,N_9499);
nand UO_509 (O_509,N_9336,N_9052);
nand UO_510 (O_510,N_9787,N_9067);
and UO_511 (O_511,N_9841,N_9263);
nor UO_512 (O_512,N_9819,N_9043);
nand UO_513 (O_513,N_9732,N_9967);
nand UO_514 (O_514,N_9155,N_9866);
nor UO_515 (O_515,N_9588,N_9684);
nand UO_516 (O_516,N_9807,N_9239);
or UO_517 (O_517,N_9875,N_9498);
or UO_518 (O_518,N_9699,N_9466);
nor UO_519 (O_519,N_9740,N_9281);
nor UO_520 (O_520,N_9815,N_9494);
nor UO_521 (O_521,N_9103,N_9776);
nor UO_522 (O_522,N_9911,N_9504);
and UO_523 (O_523,N_9132,N_9956);
nand UO_524 (O_524,N_9781,N_9059);
nor UO_525 (O_525,N_9626,N_9077);
or UO_526 (O_526,N_9544,N_9454);
and UO_527 (O_527,N_9022,N_9223);
or UO_528 (O_528,N_9808,N_9053);
and UO_529 (O_529,N_9629,N_9860);
xnor UO_530 (O_530,N_9996,N_9653);
nor UO_531 (O_531,N_9261,N_9767);
nor UO_532 (O_532,N_9728,N_9739);
xnor UO_533 (O_533,N_9393,N_9591);
or UO_534 (O_534,N_9443,N_9920);
xnor UO_535 (O_535,N_9859,N_9940);
or UO_536 (O_536,N_9407,N_9486);
nor UO_537 (O_537,N_9996,N_9763);
nor UO_538 (O_538,N_9461,N_9340);
and UO_539 (O_539,N_9188,N_9612);
or UO_540 (O_540,N_9282,N_9514);
or UO_541 (O_541,N_9735,N_9244);
and UO_542 (O_542,N_9652,N_9429);
or UO_543 (O_543,N_9561,N_9760);
or UO_544 (O_544,N_9083,N_9293);
and UO_545 (O_545,N_9016,N_9612);
nand UO_546 (O_546,N_9828,N_9756);
xor UO_547 (O_547,N_9206,N_9569);
nand UO_548 (O_548,N_9610,N_9739);
and UO_549 (O_549,N_9096,N_9685);
nand UO_550 (O_550,N_9271,N_9856);
nand UO_551 (O_551,N_9441,N_9605);
xnor UO_552 (O_552,N_9296,N_9852);
or UO_553 (O_553,N_9116,N_9696);
and UO_554 (O_554,N_9460,N_9200);
nand UO_555 (O_555,N_9056,N_9226);
xnor UO_556 (O_556,N_9501,N_9534);
and UO_557 (O_557,N_9886,N_9761);
nand UO_558 (O_558,N_9897,N_9137);
and UO_559 (O_559,N_9310,N_9264);
and UO_560 (O_560,N_9504,N_9479);
or UO_561 (O_561,N_9459,N_9217);
nor UO_562 (O_562,N_9991,N_9126);
nand UO_563 (O_563,N_9201,N_9689);
and UO_564 (O_564,N_9088,N_9882);
nand UO_565 (O_565,N_9371,N_9411);
and UO_566 (O_566,N_9050,N_9095);
or UO_567 (O_567,N_9832,N_9747);
and UO_568 (O_568,N_9001,N_9955);
and UO_569 (O_569,N_9218,N_9787);
xnor UO_570 (O_570,N_9869,N_9129);
or UO_571 (O_571,N_9698,N_9807);
xnor UO_572 (O_572,N_9580,N_9702);
or UO_573 (O_573,N_9454,N_9644);
xor UO_574 (O_574,N_9020,N_9179);
xnor UO_575 (O_575,N_9216,N_9554);
or UO_576 (O_576,N_9697,N_9041);
or UO_577 (O_577,N_9871,N_9094);
nor UO_578 (O_578,N_9006,N_9172);
nor UO_579 (O_579,N_9490,N_9047);
or UO_580 (O_580,N_9262,N_9602);
or UO_581 (O_581,N_9390,N_9908);
or UO_582 (O_582,N_9661,N_9456);
nand UO_583 (O_583,N_9236,N_9118);
and UO_584 (O_584,N_9299,N_9470);
nand UO_585 (O_585,N_9184,N_9825);
nand UO_586 (O_586,N_9312,N_9482);
or UO_587 (O_587,N_9154,N_9465);
and UO_588 (O_588,N_9487,N_9372);
and UO_589 (O_589,N_9468,N_9627);
nor UO_590 (O_590,N_9633,N_9122);
nand UO_591 (O_591,N_9339,N_9833);
or UO_592 (O_592,N_9657,N_9988);
xor UO_593 (O_593,N_9383,N_9157);
xnor UO_594 (O_594,N_9794,N_9320);
nand UO_595 (O_595,N_9936,N_9658);
or UO_596 (O_596,N_9423,N_9378);
nand UO_597 (O_597,N_9874,N_9743);
xnor UO_598 (O_598,N_9036,N_9864);
and UO_599 (O_599,N_9083,N_9044);
and UO_600 (O_600,N_9475,N_9626);
or UO_601 (O_601,N_9517,N_9068);
nor UO_602 (O_602,N_9305,N_9351);
nor UO_603 (O_603,N_9337,N_9722);
and UO_604 (O_604,N_9742,N_9820);
nor UO_605 (O_605,N_9492,N_9428);
nor UO_606 (O_606,N_9031,N_9962);
and UO_607 (O_607,N_9427,N_9683);
xnor UO_608 (O_608,N_9037,N_9639);
nor UO_609 (O_609,N_9032,N_9548);
and UO_610 (O_610,N_9946,N_9662);
or UO_611 (O_611,N_9299,N_9571);
or UO_612 (O_612,N_9631,N_9981);
nor UO_613 (O_613,N_9055,N_9450);
xor UO_614 (O_614,N_9231,N_9211);
and UO_615 (O_615,N_9875,N_9845);
or UO_616 (O_616,N_9293,N_9904);
xor UO_617 (O_617,N_9503,N_9473);
or UO_618 (O_618,N_9070,N_9013);
or UO_619 (O_619,N_9417,N_9601);
and UO_620 (O_620,N_9702,N_9062);
and UO_621 (O_621,N_9218,N_9890);
nor UO_622 (O_622,N_9682,N_9965);
and UO_623 (O_623,N_9926,N_9666);
xnor UO_624 (O_624,N_9952,N_9033);
nand UO_625 (O_625,N_9145,N_9231);
or UO_626 (O_626,N_9411,N_9489);
and UO_627 (O_627,N_9536,N_9387);
nor UO_628 (O_628,N_9133,N_9117);
and UO_629 (O_629,N_9483,N_9262);
xnor UO_630 (O_630,N_9765,N_9844);
and UO_631 (O_631,N_9447,N_9563);
or UO_632 (O_632,N_9429,N_9874);
nand UO_633 (O_633,N_9636,N_9709);
or UO_634 (O_634,N_9641,N_9723);
nor UO_635 (O_635,N_9952,N_9282);
nor UO_636 (O_636,N_9744,N_9792);
nor UO_637 (O_637,N_9332,N_9136);
xnor UO_638 (O_638,N_9396,N_9485);
xor UO_639 (O_639,N_9609,N_9488);
xor UO_640 (O_640,N_9453,N_9404);
and UO_641 (O_641,N_9221,N_9737);
and UO_642 (O_642,N_9652,N_9887);
nand UO_643 (O_643,N_9327,N_9564);
or UO_644 (O_644,N_9233,N_9100);
nor UO_645 (O_645,N_9703,N_9751);
or UO_646 (O_646,N_9866,N_9818);
nand UO_647 (O_647,N_9579,N_9684);
nor UO_648 (O_648,N_9801,N_9365);
nor UO_649 (O_649,N_9055,N_9351);
xnor UO_650 (O_650,N_9053,N_9495);
nand UO_651 (O_651,N_9051,N_9571);
and UO_652 (O_652,N_9662,N_9527);
nor UO_653 (O_653,N_9789,N_9817);
nor UO_654 (O_654,N_9947,N_9330);
or UO_655 (O_655,N_9442,N_9891);
or UO_656 (O_656,N_9892,N_9852);
nand UO_657 (O_657,N_9791,N_9944);
and UO_658 (O_658,N_9954,N_9513);
or UO_659 (O_659,N_9445,N_9328);
nor UO_660 (O_660,N_9862,N_9693);
nor UO_661 (O_661,N_9471,N_9527);
nand UO_662 (O_662,N_9050,N_9122);
or UO_663 (O_663,N_9923,N_9744);
and UO_664 (O_664,N_9024,N_9222);
or UO_665 (O_665,N_9407,N_9830);
or UO_666 (O_666,N_9935,N_9420);
or UO_667 (O_667,N_9003,N_9793);
and UO_668 (O_668,N_9691,N_9481);
nor UO_669 (O_669,N_9523,N_9468);
or UO_670 (O_670,N_9558,N_9116);
xor UO_671 (O_671,N_9789,N_9926);
nor UO_672 (O_672,N_9227,N_9434);
nand UO_673 (O_673,N_9965,N_9362);
nor UO_674 (O_674,N_9963,N_9730);
nor UO_675 (O_675,N_9338,N_9965);
nor UO_676 (O_676,N_9669,N_9435);
or UO_677 (O_677,N_9754,N_9259);
xor UO_678 (O_678,N_9231,N_9381);
and UO_679 (O_679,N_9197,N_9481);
or UO_680 (O_680,N_9361,N_9755);
and UO_681 (O_681,N_9504,N_9757);
and UO_682 (O_682,N_9507,N_9792);
nand UO_683 (O_683,N_9291,N_9963);
or UO_684 (O_684,N_9527,N_9891);
and UO_685 (O_685,N_9574,N_9415);
or UO_686 (O_686,N_9157,N_9739);
nor UO_687 (O_687,N_9281,N_9622);
and UO_688 (O_688,N_9915,N_9906);
or UO_689 (O_689,N_9174,N_9342);
nor UO_690 (O_690,N_9512,N_9152);
nor UO_691 (O_691,N_9044,N_9175);
xnor UO_692 (O_692,N_9273,N_9749);
xor UO_693 (O_693,N_9744,N_9401);
and UO_694 (O_694,N_9427,N_9342);
and UO_695 (O_695,N_9541,N_9674);
and UO_696 (O_696,N_9085,N_9370);
nand UO_697 (O_697,N_9855,N_9581);
xnor UO_698 (O_698,N_9312,N_9617);
and UO_699 (O_699,N_9613,N_9030);
and UO_700 (O_700,N_9680,N_9655);
nand UO_701 (O_701,N_9755,N_9589);
nand UO_702 (O_702,N_9334,N_9119);
or UO_703 (O_703,N_9998,N_9884);
xnor UO_704 (O_704,N_9379,N_9337);
or UO_705 (O_705,N_9493,N_9773);
and UO_706 (O_706,N_9516,N_9431);
nand UO_707 (O_707,N_9837,N_9805);
nor UO_708 (O_708,N_9817,N_9490);
or UO_709 (O_709,N_9570,N_9594);
or UO_710 (O_710,N_9249,N_9854);
nor UO_711 (O_711,N_9896,N_9144);
and UO_712 (O_712,N_9349,N_9167);
and UO_713 (O_713,N_9193,N_9560);
or UO_714 (O_714,N_9030,N_9047);
xnor UO_715 (O_715,N_9117,N_9710);
and UO_716 (O_716,N_9955,N_9204);
xor UO_717 (O_717,N_9518,N_9625);
nor UO_718 (O_718,N_9016,N_9846);
and UO_719 (O_719,N_9095,N_9153);
or UO_720 (O_720,N_9805,N_9821);
nand UO_721 (O_721,N_9612,N_9541);
and UO_722 (O_722,N_9689,N_9666);
nor UO_723 (O_723,N_9358,N_9665);
or UO_724 (O_724,N_9259,N_9583);
nand UO_725 (O_725,N_9610,N_9685);
and UO_726 (O_726,N_9665,N_9352);
or UO_727 (O_727,N_9873,N_9080);
nand UO_728 (O_728,N_9172,N_9182);
or UO_729 (O_729,N_9836,N_9666);
or UO_730 (O_730,N_9355,N_9432);
nor UO_731 (O_731,N_9923,N_9271);
or UO_732 (O_732,N_9400,N_9956);
nand UO_733 (O_733,N_9482,N_9769);
nor UO_734 (O_734,N_9542,N_9629);
and UO_735 (O_735,N_9319,N_9596);
and UO_736 (O_736,N_9886,N_9757);
xor UO_737 (O_737,N_9284,N_9673);
nor UO_738 (O_738,N_9394,N_9355);
nor UO_739 (O_739,N_9758,N_9205);
and UO_740 (O_740,N_9983,N_9510);
nand UO_741 (O_741,N_9251,N_9289);
nor UO_742 (O_742,N_9106,N_9601);
or UO_743 (O_743,N_9990,N_9789);
or UO_744 (O_744,N_9627,N_9327);
xnor UO_745 (O_745,N_9114,N_9720);
and UO_746 (O_746,N_9432,N_9865);
xnor UO_747 (O_747,N_9239,N_9257);
nand UO_748 (O_748,N_9963,N_9450);
nor UO_749 (O_749,N_9023,N_9812);
nor UO_750 (O_750,N_9195,N_9235);
and UO_751 (O_751,N_9686,N_9089);
and UO_752 (O_752,N_9540,N_9180);
or UO_753 (O_753,N_9991,N_9755);
nor UO_754 (O_754,N_9497,N_9064);
nand UO_755 (O_755,N_9396,N_9993);
nor UO_756 (O_756,N_9526,N_9750);
nand UO_757 (O_757,N_9161,N_9638);
nor UO_758 (O_758,N_9371,N_9807);
and UO_759 (O_759,N_9487,N_9284);
or UO_760 (O_760,N_9958,N_9849);
or UO_761 (O_761,N_9326,N_9082);
xnor UO_762 (O_762,N_9377,N_9114);
nor UO_763 (O_763,N_9046,N_9093);
or UO_764 (O_764,N_9153,N_9551);
or UO_765 (O_765,N_9836,N_9723);
nor UO_766 (O_766,N_9518,N_9312);
and UO_767 (O_767,N_9962,N_9155);
nor UO_768 (O_768,N_9746,N_9838);
nor UO_769 (O_769,N_9685,N_9275);
or UO_770 (O_770,N_9899,N_9077);
or UO_771 (O_771,N_9261,N_9729);
or UO_772 (O_772,N_9018,N_9060);
nand UO_773 (O_773,N_9900,N_9818);
or UO_774 (O_774,N_9693,N_9686);
nand UO_775 (O_775,N_9618,N_9900);
or UO_776 (O_776,N_9139,N_9529);
and UO_777 (O_777,N_9988,N_9996);
or UO_778 (O_778,N_9937,N_9154);
and UO_779 (O_779,N_9773,N_9903);
and UO_780 (O_780,N_9224,N_9419);
nand UO_781 (O_781,N_9856,N_9888);
and UO_782 (O_782,N_9380,N_9132);
nand UO_783 (O_783,N_9595,N_9040);
nor UO_784 (O_784,N_9184,N_9643);
nor UO_785 (O_785,N_9861,N_9605);
nand UO_786 (O_786,N_9021,N_9064);
nand UO_787 (O_787,N_9561,N_9140);
nor UO_788 (O_788,N_9535,N_9164);
nor UO_789 (O_789,N_9283,N_9130);
nand UO_790 (O_790,N_9033,N_9724);
or UO_791 (O_791,N_9461,N_9078);
or UO_792 (O_792,N_9098,N_9629);
nor UO_793 (O_793,N_9345,N_9758);
xnor UO_794 (O_794,N_9926,N_9642);
nand UO_795 (O_795,N_9515,N_9871);
and UO_796 (O_796,N_9904,N_9835);
or UO_797 (O_797,N_9076,N_9548);
nand UO_798 (O_798,N_9288,N_9193);
and UO_799 (O_799,N_9877,N_9335);
or UO_800 (O_800,N_9567,N_9686);
and UO_801 (O_801,N_9268,N_9473);
or UO_802 (O_802,N_9967,N_9624);
or UO_803 (O_803,N_9601,N_9182);
nand UO_804 (O_804,N_9448,N_9933);
or UO_805 (O_805,N_9594,N_9741);
nor UO_806 (O_806,N_9597,N_9340);
nand UO_807 (O_807,N_9395,N_9146);
nand UO_808 (O_808,N_9123,N_9543);
nand UO_809 (O_809,N_9996,N_9813);
nand UO_810 (O_810,N_9875,N_9185);
nor UO_811 (O_811,N_9054,N_9163);
and UO_812 (O_812,N_9720,N_9265);
nand UO_813 (O_813,N_9973,N_9450);
or UO_814 (O_814,N_9565,N_9864);
and UO_815 (O_815,N_9753,N_9524);
xor UO_816 (O_816,N_9932,N_9654);
nor UO_817 (O_817,N_9514,N_9334);
xnor UO_818 (O_818,N_9460,N_9457);
and UO_819 (O_819,N_9452,N_9470);
nand UO_820 (O_820,N_9051,N_9120);
nor UO_821 (O_821,N_9838,N_9923);
nand UO_822 (O_822,N_9788,N_9164);
or UO_823 (O_823,N_9024,N_9804);
nor UO_824 (O_824,N_9126,N_9711);
nand UO_825 (O_825,N_9013,N_9102);
or UO_826 (O_826,N_9119,N_9858);
nand UO_827 (O_827,N_9079,N_9723);
nor UO_828 (O_828,N_9924,N_9518);
nand UO_829 (O_829,N_9042,N_9453);
or UO_830 (O_830,N_9392,N_9490);
or UO_831 (O_831,N_9010,N_9026);
or UO_832 (O_832,N_9208,N_9446);
nand UO_833 (O_833,N_9353,N_9691);
nand UO_834 (O_834,N_9243,N_9013);
and UO_835 (O_835,N_9619,N_9393);
or UO_836 (O_836,N_9199,N_9159);
and UO_837 (O_837,N_9302,N_9222);
nor UO_838 (O_838,N_9234,N_9680);
or UO_839 (O_839,N_9242,N_9039);
nor UO_840 (O_840,N_9176,N_9798);
and UO_841 (O_841,N_9549,N_9280);
and UO_842 (O_842,N_9486,N_9171);
nor UO_843 (O_843,N_9393,N_9058);
or UO_844 (O_844,N_9720,N_9552);
and UO_845 (O_845,N_9005,N_9358);
or UO_846 (O_846,N_9182,N_9996);
and UO_847 (O_847,N_9713,N_9089);
or UO_848 (O_848,N_9030,N_9688);
or UO_849 (O_849,N_9701,N_9686);
nor UO_850 (O_850,N_9395,N_9837);
nor UO_851 (O_851,N_9226,N_9860);
or UO_852 (O_852,N_9309,N_9545);
or UO_853 (O_853,N_9034,N_9045);
xnor UO_854 (O_854,N_9300,N_9736);
or UO_855 (O_855,N_9882,N_9713);
or UO_856 (O_856,N_9277,N_9363);
and UO_857 (O_857,N_9932,N_9360);
or UO_858 (O_858,N_9932,N_9964);
nand UO_859 (O_859,N_9865,N_9861);
xor UO_860 (O_860,N_9214,N_9821);
nor UO_861 (O_861,N_9150,N_9050);
and UO_862 (O_862,N_9906,N_9977);
nor UO_863 (O_863,N_9967,N_9830);
nand UO_864 (O_864,N_9191,N_9315);
or UO_865 (O_865,N_9956,N_9410);
and UO_866 (O_866,N_9186,N_9825);
or UO_867 (O_867,N_9975,N_9874);
nor UO_868 (O_868,N_9148,N_9630);
or UO_869 (O_869,N_9759,N_9782);
or UO_870 (O_870,N_9257,N_9334);
nand UO_871 (O_871,N_9371,N_9725);
nand UO_872 (O_872,N_9938,N_9606);
and UO_873 (O_873,N_9241,N_9745);
or UO_874 (O_874,N_9970,N_9622);
and UO_875 (O_875,N_9472,N_9326);
xnor UO_876 (O_876,N_9918,N_9558);
xnor UO_877 (O_877,N_9327,N_9251);
nor UO_878 (O_878,N_9607,N_9445);
and UO_879 (O_879,N_9498,N_9017);
xor UO_880 (O_880,N_9907,N_9981);
nand UO_881 (O_881,N_9746,N_9159);
nor UO_882 (O_882,N_9536,N_9328);
or UO_883 (O_883,N_9904,N_9828);
nand UO_884 (O_884,N_9254,N_9567);
or UO_885 (O_885,N_9882,N_9446);
nand UO_886 (O_886,N_9244,N_9698);
xor UO_887 (O_887,N_9683,N_9028);
nor UO_888 (O_888,N_9970,N_9545);
or UO_889 (O_889,N_9572,N_9015);
nor UO_890 (O_890,N_9812,N_9946);
or UO_891 (O_891,N_9259,N_9337);
and UO_892 (O_892,N_9076,N_9043);
nor UO_893 (O_893,N_9282,N_9169);
or UO_894 (O_894,N_9844,N_9374);
and UO_895 (O_895,N_9778,N_9338);
or UO_896 (O_896,N_9256,N_9356);
and UO_897 (O_897,N_9393,N_9782);
xnor UO_898 (O_898,N_9184,N_9713);
or UO_899 (O_899,N_9168,N_9427);
and UO_900 (O_900,N_9770,N_9049);
or UO_901 (O_901,N_9913,N_9944);
or UO_902 (O_902,N_9414,N_9967);
or UO_903 (O_903,N_9841,N_9847);
or UO_904 (O_904,N_9857,N_9137);
or UO_905 (O_905,N_9405,N_9564);
and UO_906 (O_906,N_9506,N_9414);
and UO_907 (O_907,N_9482,N_9326);
nand UO_908 (O_908,N_9452,N_9457);
or UO_909 (O_909,N_9094,N_9338);
nand UO_910 (O_910,N_9038,N_9474);
nor UO_911 (O_911,N_9745,N_9307);
nor UO_912 (O_912,N_9665,N_9766);
and UO_913 (O_913,N_9451,N_9168);
nand UO_914 (O_914,N_9543,N_9151);
or UO_915 (O_915,N_9730,N_9435);
nand UO_916 (O_916,N_9250,N_9192);
nand UO_917 (O_917,N_9145,N_9591);
and UO_918 (O_918,N_9162,N_9526);
nand UO_919 (O_919,N_9909,N_9256);
nor UO_920 (O_920,N_9269,N_9312);
and UO_921 (O_921,N_9536,N_9383);
nand UO_922 (O_922,N_9382,N_9756);
xor UO_923 (O_923,N_9761,N_9209);
nor UO_924 (O_924,N_9000,N_9954);
nand UO_925 (O_925,N_9735,N_9030);
xor UO_926 (O_926,N_9140,N_9134);
nand UO_927 (O_927,N_9948,N_9169);
xnor UO_928 (O_928,N_9621,N_9174);
nor UO_929 (O_929,N_9776,N_9090);
nor UO_930 (O_930,N_9783,N_9413);
or UO_931 (O_931,N_9568,N_9773);
nor UO_932 (O_932,N_9363,N_9118);
nor UO_933 (O_933,N_9318,N_9572);
nor UO_934 (O_934,N_9269,N_9982);
and UO_935 (O_935,N_9690,N_9404);
nand UO_936 (O_936,N_9832,N_9009);
nand UO_937 (O_937,N_9488,N_9000);
and UO_938 (O_938,N_9397,N_9780);
xnor UO_939 (O_939,N_9700,N_9842);
nor UO_940 (O_940,N_9630,N_9596);
or UO_941 (O_941,N_9044,N_9828);
nor UO_942 (O_942,N_9923,N_9074);
nor UO_943 (O_943,N_9004,N_9305);
or UO_944 (O_944,N_9106,N_9947);
nand UO_945 (O_945,N_9373,N_9510);
nand UO_946 (O_946,N_9631,N_9095);
and UO_947 (O_947,N_9752,N_9771);
xor UO_948 (O_948,N_9015,N_9085);
nor UO_949 (O_949,N_9630,N_9699);
nand UO_950 (O_950,N_9452,N_9715);
nand UO_951 (O_951,N_9622,N_9403);
or UO_952 (O_952,N_9679,N_9796);
nor UO_953 (O_953,N_9368,N_9709);
nor UO_954 (O_954,N_9524,N_9553);
nor UO_955 (O_955,N_9271,N_9467);
nand UO_956 (O_956,N_9263,N_9192);
nand UO_957 (O_957,N_9206,N_9857);
or UO_958 (O_958,N_9492,N_9795);
and UO_959 (O_959,N_9917,N_9944);
nor UO_960 (O_960,N_9481,N_9292);
or UO_961 (O_961,N_9356,N_9466);
xor UO_962 (O_962,N_9230,N_9956);
and UO_963 (O_963,N_9747,N_9362);
nor UO_964 (O_964,N_9632,N_9780);
nor UO_965 (O_965,N_9776,N_9618);
and UO_966 (O_966,N_9368,N_9129);
nor UO_967 (O_967,N_9149,N_9125);
nand UO_968 (O_968,N_9529,N_9499);
and UO_969 (O_969,N_9527,N_9153);
or UO_970 (O_970,N_9004,N_9051);
and UO_971 (O_971,N_9756,N_9129);
nor UO_972 (O_972,N_9655,N_9651);
nand UO_973 (O_973,N_9501,N_9136);
nor UO_974 (O_974,N_9448,N_9084);
nor UO_975 (O_975,N_9721,N_9170);
or UO_976 (O_976,N_9746,N_9946);
xor UO_977 (O_977,N_9920,N_9323);
xnor UO_978 (O_978,N_9838,N_9373);
nand UO_979 (O_979,N_9678,N_9097);
nor UO_980 (O_980,N_9401,N_9903);
or UO_981 (O_981,N_9343,N_9251);
nand UO_982 (O_982,N_9734,N_9631);
nand UO_983 (O_983,N_9512,N_9385);
xor UO_984 (O_984,N_9014,N_9137);
or UO_985 (O_985,N_9834,N_9524);
xor UO_986 (O_986,N_9995,N_9045);
or UO_987 (O_987,N_9455,N_9125);
nor UO_988 (O_988,N_9890,N_9989);
nor UO_989 (O_989,N_9529,N_9924);
nand UO_990 (O_990,N_9874,N_9408);
or UO_991 (O_991,N_9906,N_9664);
xnor UO_992 (O_992,N_9463,N_9595);
nor UO_993 (O_993,N_9701,N_9849);
or UO_994 (O_994,N_9430,N_9244);
and UO_995 (O_995,N_9973,N_9039);
or UO_996 (O_996,N_9492,N_9627);
and UO_997 (O_997,N_9750,N_9870);
nand UO_998 (O_998,N_9801,N_9273);
nor UO_999 (O_999,N_9309,N_9128);
and UO_1000 (O_1000,N_9842,N_9921);
or UO_1001 (O_1001,N_9220,N_9286);
nand UO_1002 (O_1002,N_9451,N_9669);
nand UO_1003 (O_1003,N_9826,N_9487);
and UO_1004 (O_1004,N_9460,N_9808);
or UO_1005 (O_1005,N_9802,N_9951);
nand UO_1006 (O_1006,N_9749,N_9562);
or UO_1007 (O_1007,N_9355,N_9846);
nor UO_1008 (O_1008,N_9334,N_9536);
nand UO_1009 (O_1009,N_9812,N_9622);
or UO_1010 (O_1010,N_9330,N_9449);
nor UO_1011 (O_1011,N_9227,N_9753);
nor UO_1012 (O_1012,N_9227,N_9002);
nand UO_1013 (O_1013,N_9138,N_9931);
nor UO_1014 (O_1014,N_9517,N_9470);
or UO_1015 (O_1015,N_9497,N_9380);
nor UO_1016 (O_1016,N_9265,N_9696);
and UO_1017 (O_1017,N_9605,N_9638);
nand UO_1018 (O_1018,N_9719,N_9247);
and UO_1019 (O_1019,N_9477,N_9843);
xor UO_1020 (O_1020,N_9850,N_9598);
nand UO_1021 (O_1021,N_9328,N_9663);
nor UO_1022 (O_1022,N_9352,N_9714);
nor UO_1023 (O_1023,N_9157,N_9345);
or UO_1024 (O_1024,N_9060,N_9767);
nand UO_1025 (O_1025,N_9828,N_9167);
nor UO_1026 (O_1026,N_9449,N_9942);
xor UO_1027 (O_1027,N_9292,N_9144);
and UO_1028 (O_1028,N_9726,N_9851);
or UO_1029 (O_1029,N_9340,N_9850);
nand UO_1030 (O_1030,N_9079,N_9871);
xnor UO_1031 (O_1031,N_9395,N_9928);
nor UO_1032 (O_1032,N_9779,N_9447);
and UO_1033 (O_1033,N_9812,N_9114);
nor UO_1034 (O_1034,N_9467,N_9156);
xnor UO_1035 (O_1035,N_9975,N_9679);
and UO_1036 (O_1036,N_9408,N_9258);
nand UO_1037 (O_1037,N_9931,N_9160);
nand UO_1038 (O_1038,N_9783,N_9686);
nand UO_1039 (O_1039,N_9133,N_9663);
or UO_1040 (O_1040,N_9366,N_9253);
nor UO_1041 (O_1041,N_9924,N_9292);
and UO_1042 (O_1042,N_9690,N_9224);
nand UO_1043 (O_1043,N_9587,N_9326);
nor UO_1044 (O_1044,N_9153,N_9927);
and UO_1045 (O_1045,N_9364,N_9361);
and UO_1046 (O_1046,N_9035,N_9236);
and UO_1047 (O_1047,N_9930,N_9211);
nor UO_1048 (O_1048,N_9136,N_9019);
xnor UO_1049 (O_1049,N_9649,N_9650);
and UO_1050 (O_1050,N_9310,N_9419);
nor UO_1051 (O_1051,N_9765,N_9109);
nand UO_1052 (O_1052,N_9922,N_9442);
nor UO_1053 (O_1053,N_9173,N_9883);
nand UO_1054 (O_1054,N_9604,N_9570);
nor UO_1055 (O_1055,N_9535,N_9515);
and UO_1056 (O_1056,N_9837,N_9414);
nand UO_1057 (O_1057,N_9388,N_9404);
nor UO_1058 (O_1058,N_9832,N_9758);
nor UO_1059 (O_1059,N_9162,N_9998);
nand UO_1060 (O_1060,N_9524,N_9894);
nor UO_1061 (O_1061,N_9381,N_9372);
or UO_1062 (O_1062,N_9419,N_9028);
and UO_1063 (O_1063,N_9037,N_9516);
nand UO_1064 (O_1064,N_9114,N_9586);
or UO_1065 (O_1065,N_9339,N_9594);
nand UO_1066 (O_1066,N_9220,N_9130);
or UO_1067 (O_1067,N_9024,N_9814);
nor UO_1068 (O_1068,N_9637,N_9306);
and UO_1069 (O_1069,N_9495,N_9781);
and UO_1070 (O_1070,N_9125,N_9736);
or UO_1071 (O_1071,N_9064,N_9858);
nor UO_1072 (O_1072,N_9910,N_9027);
nor UO_1073 (O_1073,N_9901,N_9301);
nor UO_1074 (O_1074,N_9982,N_9833);
nand UO_1075 (O_1075,N_9429,N_9577);
nor UO_1076 (O_1076,N_9133,N_9235);
or UO_1077 (O_1077,N_9931,N_9830);
nor UO_1078 (O_1078,N_9987,N_9877);
nor UO_1079 (O_1079,N_9078,N_9405);
and UO_1080 (O_1080,N_9033,N_9903);
nor UO_1081 (O_1081,N_9366,N_9922);
and UO_1082 (O_1082,N_9794,N_9756);
nor UO_1083 (O_1083,N_9536,N_9594);
nand UO_1084 (O_1084,N_9145,N_9191);
nand UO_1085 (O_1085,N_9280,N_9283);
nand UO_1086 (O_1086,N_9871,N_9722);
nor UO_1087 (O_1087,N_9040,N_9946);
and UO_1088 (O_1088,N_9551,N_9895);
or UO_1089 (O_1089,N_9533,N_9266);
or UO_1090 (O_1090,N_9108,N_9450);
or UO_1091 (O_1091,N_9006,N_9920);
or UO_1092 (O_1092,N_9066,N_9309);
nor UO_1093 (O_1093,N_9731,N_9415);
xor UO_1094 (O_1094,N_9690,N_9247);
nor UO_1095 (O_1095,N_9610,N_9818);
nor UO_1096 (O_1096,N_9424,N_9126);
nor UO_1097 (O_1097,N_9608,N_9802);
nand UO_1098 (O_1098,N_9997,N_9037);
nor UO_1099 (O_1099,N_9139,N_9966);
nor UO_1100 (O_1100,N_9149,N_9952);
or UO_1101 (O_1101,N_9065,N_9490);
or UO_1102 (O_1102,N_9497,N_9869);
nor UO_1103 (O_1103,N_9527,N_9811);
nor UO_1104 (O_1104,N_9637,N_9773);
or UO_1105 (O_1105,N_9508,N_9732);
or UO_1106 (O_1106,N_9538,N_9898);
nand UO_1107 (O_1107,N_9947,N_9781);
and UO_1108 (O_1108,N_9706,N_9310);
nor UO_1109 (O_1109,N_9839,N_9312);
nor UO_1110 (O_1110,N_9695,N_9209);
and UO_1111 (O_1111,N_9831,N_9225);
xor UO_1112 (O_1112,N_9453,N_9727);
nor UO_1113 (O_1113,N_9570,N_9350);
xor UO_1114 (O_1114,N_9919,N_9826);
nand UO_1115 (O_1115,N_9606,N_9101);
nor UO_1116 (O_1116,N_9909,N_9900);
nand UO_1117 (O_1117,N_9512,N_9641);
and UO_1118 (O_1118,N_9969,N_9834);
or UO_1119 (O_1119,N_9224,N_9707);
and UO_1120 (O_1120,N_9231,N_9861);
nor UO_1121 (O_1121,N_9919,N_9847);
nand UO_1122 (O_1122,N_9726,N_9272);
nor UO_1123 (O_1123,N_9640,N_9768);
and UO_1124 (O_1124,N_9363,N_9745);
and UO_1125 (O_1125,N_9904,N_9237);
or UO_1126 (O_1126,N_9635,N_9534);
or UO_1127 (O_1127,N_9192,N_9863);
nand UO_1128 (O_1128,N_9659,N_9520);
xnor UO_1129 (O_1129,N_9184,N_9033);
nand UO_1130 (O_1130,N_9556,N_9454);
nor UO_1131 (O_1131,N_9325,N_9266);
and UO_1132 (O_1132,N_9839,N_9954);
or UO_1133 (O_1133,N_9987,N_9119);
and UO_1134 (O_1134,N_9139,N_9534);
nand UO_1135 (O_1135,N_9169,N_9301);
nand UO_1136 (O_1136,N_9341,N_9708);
nand UO_1137 (O_1137,N_9352,N_9511);
and UO_1138 (O_1138,N_9611,N_9907);
nand UO_1139 (O_1139,N_9970,N_9919);
nand UO_1140 (O_1140,N_9285,N_9166);
nor UO_1141 (O_1141,N_9369,N_9160);
nor UO_1142 (O_1142,N_9584,N_9479);
and UO_1143 (O_1143,N_9523,N_9116);
and UO_1144 (O_1144,N_9001,N_9066);
or UO_1145 (O_1145,N_9859,N_9580);
nor UO_1146 (O_1146,N_9645,N_9939);
or UO_1147 (O_1147,N_9776,N_9653);
nand UO_1148 (O_1148,N_9594,N_9711);
nor UO_1149 (O_1149,N_9166,N_9793);
xnor UO_1150 (O_1150,N_9432,N_9962);
nor UO_1151 (O_1151,N_9813,N_9552);
nor UO_1152 (O_1152,N_9665,N_9790);
nor UO_1153 (O_1153,N_9674,N_9011);
nor UO_1154 (O_1154,N_9367,N_9570);
nor UO_1155 (O_1155,N_9754,N_9984);
nor UO_1156 (O_1156,N_9267,N_9803);
nor UO_1157 (O_1157,N_9403,N_9526);
nor UO_1158 (O_1158,N_9034,N_9370);
nand UO_1159 (O_1159,N_9204,N_9128);
nor UO_1160 (O_1160,N_9887,N_9991);
and UO_1161 (O_1161,N_9174,N_9372);
nand UO_1162 (O_1162,N_9054,N_9602);
nand UO_1163 (O_1163,N_9070,N_9944);
and UO_1164 (O_1164,N_9915,N_9745);
nor UO_1165 (O_1165,N_9914,N_9567);
or UO_1166 (O_1166,N_9747,N_9818);
nor UO_1167 (O_1167,N_9734,N_9558);
nor UO_1168 (O_1168,N_9339,N_9025);
or UO_1169 (O_1169,N_9057,N_9068);
nand UO_1170 (O_1170,N_9296,N_9694);
and UO_1171 (O_1171,N_9303,N_9422);
nor UO_1172 (O_1172,N_9311,N_9536);
and UO_1173 (O_1173,N_9290,N_9311);
nor UO_1174 (O_1174,N_9804,N_9990);
or UO_1175 (O_1175,N_9224,N_9853);
and UO_1176 (O_1176,N_9132,N_9021);
nand UO_1177 (O_1177,N_9477,N_9957);
and UO_1178 (O_1178,N_9016,N_9112);
xor UO_1179 (O_1179,N_9988,N_9475);
nor UO_1180 (O_1180,N_9016,N_9926);
and UO_1181 (O_1181,N_9901,N_9789);
xor UO_1182 (O_1182,N_9917,N_9152);
nor UO_1183 (O_1183,N_9754,N_9704);
and UO_1184 (O_1184,N_9941,N_9394);
xor UO_1185 (O_1185,N_9975,N_9685);
xnor UO_1186 (O_1186,N_9584,N_9259);
nand UO_1187 (O_1187,N_9443,N_9458);
nand UO_1188 (O_1188,N_9790,N_9206);
xnor UO_1189 (O_1189,N_9630,N_9975);
nand UO_1190 (O_1190,N_9579,N_9682);
nand UO_1191 (O_1191,N_9023,N_9845);
and UO_1192 (O_1192,N_9677,N_9752);
nand UO_1193 (O_1193,N_9135,N_9110);
xor UO_1194 (O_1194,N_9426,N_9971);
and UO_1195 (O_1195,N_9879,N_9152);
and UO_1196 (O_1196,N_9997,N_9283);
nand UO_1197 (O_1197,N_9005,N_9295);
or UO_1198 (O_1198,N_9617,N_9606);
nand UO_1199 (O_1199,N_9155,N_9233);
or UO_1200 (O_1200,N_9842,N_9408);
and UO_1201 (O_1201,N_9631,N_9599);
and UO_1202 (O_1202,N_9471,N_9945);
nand UO_1203 (O_1203,N_9743,N_9005);
nor UO_1204 (O_1204,N_9604,N_9650);
nor UO_1205 (O_1205,N_9464,N_9177);
nor UO_1206 (O_1206,N_9475,N_9665);
and UO_1207 (O_1207,N_9104,N_9380);
or UO_1208 (O_1208,N_9461,N_9302);
nor UO_1209 (O_1209,N_9626,N_9064);
nand UO_1210 (O_1210,N_9866,N_9399);
nand UO_1211 (O_1211,N_9179,N_9673);
or UO_1212 (O_1212,N_9210,N_9390);
nand UO_1213 (O_1213,N_9706,N_9298);
or UO_1214 (O_1214,N_9405,N_9797);
nor UO_1215 (O_1215,N_9908,N_9254);
nand UO_1216 (O_1216,N_9116,N_9247);
xor UO_1217 (O_1217,N_9367,N_9163);
nor UO_1218 (O_1218,N_9402,N_9935);
and UO_1219 (O_1219,N_9000,N_9301);
nand UO_1220 (O_1220,N_9679,N_9783);
and UO_1221 (O_1221,N_9295,N_9055);
nand UO_1222 (O_1222,N_9084,N_9009);
or UO_1223 (O_1223,N_9494,N_9836);
xor UO_1224 (O_1224,N_9859,N_9756);
or UO_1225 (O_1225,N_9612,N_9882);
nand UO_1226 (O_1226,N_9529,N_9361);
nor UO_1227 (O_1227,N_9596,N_9274);
and UO_1228 (O_1228,N_9285,N_9942);
nand UO_1229 (O_1229,N_9923,N_9414);
xor UO_1230 (O_1230,N_9866,N_9599);
or UO_1231 (O_1231,N_9438,N_9873);
xnor UO_1232 (O_1232,N_9462,N_9759);
nor UO_1233 (O_1233,N_9278,N_9079);
nand UO_1234 (O_1234,N_9585,N_9647);
nand UO_1235 (O_1235,N_9425,N_9600);
nand UO_1236 (O_1236,N_9676,N_9097);
and UO_1237 (O_1237,N_9710,N_9817);
nor UO_1238 (O_1238,N_9155,N_9231);
and UO_1239 (O_1239,N_9648,N_9177);
or UO_1240 (O_1240,N_9459,N_9272);
and UO_1241 (O_1241,N_9705,N_9362);
nand UO_1242 (O_1242,N_9983,N_9623);
and UO_1243 (O_1243,N_9644,N_9612);
or UO_1244 (O_1244,N_9656,N_9951);
or UO_1245 (O_1245,N_9132,N_9221);
and UO_1246 (O_1246,N_9249,N_9108);
or UO_1247 (O_1247,N_9780,N_9854);
and UO_1248 (O_1248,N_9449,N_9906);
nor UO_1249 (O_1249,N_9166,N_9701);
nor UO_1250 (O_1250,N_9947,N_9223);
nand UO_1251 (O_1251,N_9919,N_9821);
nand UO_1252 (O_1252,N_9971,N_9198);
and UO_1253 (O_1253,N_9096,N_9345);
nor UO_1254 (O_1254,N_9994,N_9893);
nor UO_1255 (O_1255,N_9459,N_9867);
or UO_1256 (O_1256,N_9817,N_9561);
or UO_1257 (O_1257,N_9534,N_9235);
or UO_1258 (O_1258,N_9247,N_9466);
nand UO_1259 (O_1259,N_9908,N_9611);
or UO_1260 (O_1260,N_9787,N_9958);
nand UO_1261 (O_1261,N_9554,N_9141);
and UO_1262 (O_1262,N_9805,N_9173);
and UO_1263 (O_1263,N_9544,N_9989);
and UO_1264 (O_1264,N_9115,N_9305);
nor UO_1265 (O_1265,N_9362,N_9511);
xor UO_1266 (O_1266,N_9571,N_9232);
nor UO_1267 (O_1267,N_9084,N_9313);
and UO_1268 (O_1268,N_9249,N_9024);
nor UO_1269 (O_1269,N_9839,N_9673);
nand UO_1270 (O_1270,N_9296,N_9700);
or UO_1271 (O_1271,N_9191,N_9350);
and UO_1272 (O_1272,N_9180,N_9981);
nor UO_1273 (O_1273,N_9191,N_9843);
or UO_1274 (O_1274,N_9028,N_9584);
or UO_1275 (O_1275,N_9289,N_9632);
nor UO_1276 (O_1276,N_9098,N_9774);
nor UO_1277 (O_1277,N_9565,N_9261);
nor UO_1278 (O_1278,N_9514,N_9993);
nor UO_1279 (O_1279,N_9665,N_9982);
nor UO_1280 (O_1280,N_9078,N_9672);
xor UO_1281 (O_1281,N_9349,N_9482);
and UO_1282 (O_1282,N_9453,N_9977);
nand UO_1283 (O_1283,N_9044,N_9209);
nor UO_1284 (O_1284,N_9257,N_9190);
or UO_1285 (O_1285,N_9199,N_9764);
and UO_1286 (O_1286,N_9356,N_9564);
or UO_1287 (O_1287,N_9247,N_9585);
nor UO_1288 (O_1288,N_9715,N_9051);
nor UO_1289 (O_1289,N_9390,N_9583);
nand UO_1290 (O_1290,N_9088,N_9993);
or UO_1291 (O_1291,N_9997,N_9787);
and UO_1292 (O_1292,N_9505,N_9036);
and UO_1293 (O_1293,N_9546,N_9182);
nand UO_1294 (O_1294,N_9189,N_9963);
nor UO_1295 (O_1295,N_9486,N_9254);
nor UO_1296 (O_1296,N_9250,N_9776);
and UO_1297 (O_1297,N_9799,N_9923);
nand UO_1298 (O_1298,N_9400,N_9030);
and UO_1299 (O_1299,N_9520,N_9263);
and UO_1300 (O_1300,N_9683,N_9502);
nor UO_1301 (O_1301,N_9666,N_9428);
nand UO_1302 (O_1302,N_9545,N_9512);
nor UO_1303 (O_1303,N_9876,N_9037);
nand UO_1304 (O_1304,N_9563,N_9411);
xnor UO_1305 (O_1305,N_9498,N_9934);
nand UO_1306 (O_1306,N_9601,N_9445);
or UO_1307 (O_1307,N_9881,N_9167);
nor UO_1308 (O_1308,N_9726,N_9461);
and UO_1309 (O_1309,N_9408,N_9336);
and UO_1310 (O_1310,N_9584,N_9280);
and UO_1311 (O_1311,N_9139,N_9293);
and UO_1312 (O_1312,N_9444,N_9616);
and UO_1313 (O_1313,N_9497,N_9371);
nand UO_1314 (O_1314,N_9143,N_9998);
nand UO_1315 (O_1315,N_9399,N_9773);
or UO_1316 (O_1316,N_9899,N_9394);
and UO_1317 (O_1317,N_9495,N_9642);
and UO_1318 (O_1318,N_9961,N_9660);
or UO_1319 (O_1319,N_9090,N_9018);
nand UO_1320 (O_1320,N_9234,N_9419);
nor UO_1321 (O_1321,N_9734,N_9213);
or UO_1322 (O_1322,N_9237,N_9115);
or UO_1323 (O_1323,N_9022,N_9780);
and UO_1324 (O_1324,N_9849,N_9905);
xnor UO_1325 (O_1325,N_9618,N_9061);
or UO_1326 (O_1326,N_9216,N_9396);
nor UO_1327 (O_1327,N_9330,N_9633);
nor UO_1328 (O_1328,N_9831,N_9413);
nand UO_1329 (O_1329,N_9197,N_9223);
nand UO_1330 (O_1330,N_9846,N_9716);
or UO_1331 (O_1331,N_9366,N_9149);
or UO_1332 (O_1332,N_9015,N_9699);
and UO_1333 (O_1333,N_9112,N_9278);
nor UO_1334 (O_1334,N_9519,N_9779);
nor UO_1335 (O_1335,N_9169,N_9907);
and UO_1336 (O_1336,N_9256,N_9422);
nor UO_1337 (O_1337,N_9010,N_9886);
and UO_1338 (O_1338,N_9419,N_9962);
nor UO_1339 (O_1339,N_9874,N_9972);
nor UO_1340 (O_1340,N_9146,N_9579);
or UO_1341 (O_1341,N_9437,N_9492);
xnor UO_1342 (O_1342,N_9113,N_9724);
and UO_1343 (O_1343,N_9677,N_9781);
and UO_1344 (O_1344,N_9650,N_9186);
or UO_1345 (O_1345,N_9675,N_9822);
or UO_1346 (O_1346,N_9970,N_9553);
nand UO_1347 (O_1347,N_9605,N_9702);
nor UO_1348 (O_1348,N_9236,N_9912);
nor UO_1349 (O_1349,N_9020,N_9917);
or UO_1350 (O_1350,N_9508,N_9992);
nor UO_1351 (O_1351,N_9422,N_9011);
and UO_1352 (O_1352,N_9393,N_9890);
or UO_1353 (O_1353,N_9709,N_9400);
or UO_1354 (O_1354,N_9106,N_9610);
nor UO_1355 (O_1355,N_9099,N_9370);
nand UO_1356 (O_1356,N_9583,N_9685);
and UO_1357 (O_1357,N_9209,N_9583);
nand UO_1358 (O_1358,N_9979,N_9511);
and UO_1359 (O_1359,N_9683,N_9448);
xnor UO_1360 (O_1360,N_9783,N_9096);
nor UO_1361 (O_1361,N_9412,N_9091);
nand UO_1362 (O_1362,N_9328,N_9161);
nor UO_1363 (O_1363,N_9003,N_9240);
nand UO_1364 (O_1364,N_9030,N_9906);
or UO_1365 (O_1365,N_9412,N_9591);
nor UO_1366 (O_1366,N_9077,N_9976);
or UO_1367 (O_1367,N_9164,N_9618);
nor UO_1368 (O_1368,N_9384,N_9323);
nor UO_1369 (O_1369,N_9588,N_9172);
and UO_1370 (O_1370,N_9165,N_9750);
and UO_1371 (O_1371,N_9856,N_9822);
or UO_1372 (O_1372,N_9026,N_9579);
or UO_1373 (O_1373,N_9043,N_9387);
or UO_1374 (O_1374,N_9124,N_9383);
nand UO_1375 (O_1375,N_9477,N_9533);
xnor UO_1376 (O_1376,N_9228,N_9697);
nor UO_1377 (O_1377,N_9791,N_9845);
and UO_1378 (O_1378,N_9228,N_9242);
nor UO_1379 (O_1379,N_9506,N_9487);
or UO_1380 (O_1380,N_9811,N_9194);
nand UO_1381 (O_1381,N_9412,N_9623);
nand UO_1382 (O_1382,N_9676,N_9928);
nor UO_1383 (O_1383,N_9036,N_9709);
xnor UO_1384 (O_1384,N_9284,N_9874);
nor UO_1385 (O_1385,N_9190,N_9110);
nor UO_1386 (O_1386,N_9264,N_9915);
or UO_1387 (O_1387,N_9123,N_9050);
xnor UO_1388 (O_1388,N_9820,N_9876);
and UO_1389 (O_1389,N_9061,N_9097);
nand UO_1390 (O_1390,N_9710,N_9970);
or UO_1391 (O_1391,N_9955,N_9947);
or UO_1392 (O_1392,N_9742,N_9933);
and UO_1393 (O_1393,N_9209,N_9337);
nor UO_1394 (O_1394,N_9702,N_9115);
nor UO_1395 (O_1395,N_9093,N_9416);
or UO_1396 (O_1396,N_9489,N_9335);
and UO_1397 (O_1397,N_9418,N_9742);
nand UO_1398 (O_1398,N_9654,N_9713);
xnor UO_1399 (O_1399,N_9434,N_9085);
or UO_1400 (O_1400,N_9287,N_9088);
xor UO_1401 (O_1401,N_9414,N_9706);
nand UO_1402 (O_1402,N_9406,N_9569);
or UO_1403 (O_1403,N_9550,N_9651);
or UO_1404 (O_1404,N_9478,N_9849);
and UO_1405 (O_1405,N_9174,N_9255);
nand UO_1406 (O_1406,N_9449,N_9370);
xor UO_1407 (O_1407,N_9662,N_9431);
and UO_1408 (O_1408,N_9847,N_9505);
nor UO_1409 (O_1409,N_9191,N_9543);
or UO_1410 (O_1410,N_9442,N_9766);
or UO_1411 (O_1411,N_9572,N_9419);
nor UO_1412 (O_1412,N_9445,N_9415);
and UO_1413 (O_1413,N_9035,N_9617);
nor UO_1414 (O_1414,N_9546,N_9522);
nand UO_1415 (O_1415,N_9479,N_9497);
nand UO_1416 (O_1416,N_9978,N_9399);
and UO_1417 (O_1417,N_9345,N_9004);
or UO_1418 (O_1418,N_9839,N_9513);
nor UO_1419 (O_1419,N_9821,N_9888);
or UO_1420 (O_1420,N_9266,N_9709);
nand UO_1421 (O_1421,N_9060,N_9423);
nand UO_1422 (O_1422,N_9425,N_9517);
or UO_1423 (O_1423,N_9996,N_9577);
or UO_1424 (O_1424,N_9041,N_9806);
or UO_1425 (O_1425,N_9746,N_9420);
nor UO_1426 (O_1426,N_9498,N_9122);
or UO_1427 (O_1427,N_9861,N_9521);
nor UO_1428 (O_1428,N_9399,N_9965);
xor UO_1429 (O_1429,N_9381,N_9403);
and UO_1430 (O_1430,N_9914,N_9442);
xor UO_1431 (O_1431,N_9935,N_9425);
or UO_1432 (O_1432,N_9144,N_9176);
and UO_1433 (O_1433,N_9875,N_9491);
or UO_1434 (O_1434,N_9908,N_9074);
and UO_1435 (O_1435,N_9360,N_9468);
nor UO_1436 (O_1436,N_9230,N_9454);
nor UO_1437 (O_1437,N_9399,N_9601);
nor UO_1438 (O_1438,N_9112,N_9781);
and UO_1439 (O_1439,N_9297,N_9382);
nor UO_1440 (O_1440,N_9081,N_9329);
and UO_1441 (O_1441,N_9839,N_9937);
or UO_1442 (O_1442,N_9755,N_9456);
nor UO_1443 (O_1443,N_9196,N_9493);
xor UO_1444 (O_1444,N_9788,N_9374);
xnor UO_1445 (O_1445,N_9954,N_9338);
xor UO_1446 (O_1446,N_9266,N_9245);
and UO_1447 (O_1447,N_9830,N_9327);
and UO_1448 (O_1448,N_9846,N_9463);
xnor UO_1449 (O_1449,N_9248,N_9079);
nor UO_1450 (O_1450,N_9068,N_9265);
and UO_1451 (O_1451,N_9413,N_9102);
or UO_1452 (O_1452,N_9234,N_9647);
nand UO_1453 (O_1453,N_9564,N_9620);
and UO_1454 (O_1454,N_9813,N_9799);
and UO_1455 (O_1455,N_9613,N_9104);
nand UO_1456 (O_1456,N_9863,N_9589);
or UO_1457 (O_1457,N_9869,N_9586);
or UO_1458 (O_1458,N_9467,N_9026);
or UO_1459 (O_1459,N_9184,N_9994);
nand UO_1460 (O_1460,N_9039,N_9994);
or UO_1461 (O_1461,N_9437,N_9456);
nand UO_1462 (O_1462,N_9913,N_9653);
or UO_1463 (O_1463,N_9047,N_9745);
xnor UO_1464 (O_1464,N_9985,N_9918);
or UO_1465 (O_1465,N_9625,N_9830);
nor UO_1466 (O_1466,N_9216,N_9778);
and UO_1467 (O_1467,N_9691,N_9937);
and UO_1468 (O_1468,N_9357,N_9157);
and UO_1469 (O_1469,N_9190,N_9947);
and UO_1470 (O_1470,N_9396,N_9227);
nor UO_1471 (O_1471,N_9712,N_9079);
nand UO_1472 (O_1472,N_9729,N_9832);
nor UO_1473 (O_1473,N_9597,N_9074);
nor UO_1474 (O_1474,N_9748,N_9047);
nor UO_1475 (O_1475,N_9985,N_9082);
or UO_1476 (O_1476,N_9288,N_9334);
xor UO_1477 (O_1477,N_9431,N_9354);
or UO_1478 (O_1478,N_9996,N_9792);
or UO_1479 (O_1479,N_9366,N_9992);
and UO_1480 (O_1480,N_9979,N_9628);
nand UO_1481 (O_1481,N_9116,N_9308);
or UO_1482 (O_1482,N_9637,N_9380);
nand UO_1483 (O_1483,N_9752,N_9207);
and UO_1484 (O_1484,N_9716,N_9373);
and UO_1485 (O_1485,N_9365,N_9186);
nand UO_1486 (O_1486,N_9251,N_9655);
or UO_1487 (O_1487,N_9932,N_9636);
and UO_1488 (O_1488,N_9645,N_9247);
nand UO_1489 (O_1489,N_9037,N_9269);
nor UO_1490 (O_1490,N_9258,N_9903);
and UO_1491 (O_1491,N_9537,N_9411);
nor UO_1492 (O_1492,N_9182,N_9342);
and UO_1493 (O_1493,N_9385,N_9424);
nor UO_1494 (O_1494,N_9833,N_9703);
nor UO_1495 (O_1495,N_9177,N_9547);
nand UO_1496 (O_1496,N_9782,N_9374);
and UO_1497 (O_1497,N_9476,N_9024);
and UO_1498 (O_1498,N_9173,N_9552);
nor UO_1499 (O_1499,N_9107,N_9098);
endmodule