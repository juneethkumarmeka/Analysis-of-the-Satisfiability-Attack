module basic_1500_15000_2000_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_777,In_1315);
and U1 (N_1,In_659,In_1107);
or U2 (N_2,In_1351,In_503);
or U3 (N_3,In_842,In_125);
or U4 (N_4,In_471,In_89);
or U5 (N_5,In_276,In_1233);
nand U6 (N_6,In_315,In_778);
xnor U7 (N_7,In_197,In_1087);
or U8 (N_8,In_361,In_1289);
xnor U9 (N_9,In_1323,In_1177);
and U10 (N_10,In_1096,In_507);
xor U11 (N_11,In_456,In_453);
or U12 (N_12,In_769,In_615);
or U13 (N_13,In_1286,In_1260);
and U14 (N_14,In_1085,In_1368);
nand U15 (N_15,In_1420,In_852);
xor U16 (N_16,In_535,In_1275);
and U17 (N_17,In_31,In_1019);
and U18 (N_18,In_10,In_933);
nor U19 (N_19,In_727,In_1415);
or U20 (N_20,In_173,In_674);
nand U21 (N_21,In_1156,In_1431);
xnor U22 (N_22,In_825,In_1179);
or U23 (N_23,In_520,In_1261);
xor U24 (N_24,In_848,In_735);
xor U25 (N_25,In_1367,In_1201);
nor U26 (N_26,In_90,In_128);
nand U27 (N_27,In_1349,In_1290);
nand U28 (N_28,In_969,In_865);
nand U29 (N_29,In_839,In_1317);
xor U30 (N_30,In_499,In_355);
or U31 (N_31,In_1460,In_1330);
or U32 (N_32,In_892,In_338);
or U33 (N_33,In_360,In_310);
xor U34 (N_34,In_857,In_1126);
xnor U35 (N_35,In_475,In_1336);
xnor U36 (N_36,In_981,In_140);
and U37 (N_37,In_193,In_34);
and U38 (N_38,In_849,In_352);
nor U39 (N_39,In_190,In_318);
nand U40 (N_40,In_1099,In_1429);
xnor U41 (N_41,In_78,In_1326);
and U42 (N_42,In_1377,In_1157);
xor U43 (N_43,In_677,In_689);
nand U44 (N_44,In_783,In_18);
or U45 (N_45,In_1333,In_448);
nand U46 (N_46,In_1239,In_1237);
nor U47 (N_47,In_867,In_108);
nor U48 (N_48,In_163,In_28);
nand U49 (N_49,In_80,In_288);
nor U50 (N_50,In_142,In_915);
or U51 (N_51,In_544,In_962);
xnor U52 (N_52,In_1144,In_1218);
nor U53 (N_53,In_122,In_881);
nor U54 (N_54,In_464,In_566);
and U55 (N_55,In_372,In_472);
nor U56 (N_56,In_1325,In_1443);
xor U57 (N_57,In_1070,In_397);
nand U58 (N_58,In_785,In_562);
and U59 (N_59,In_802,In_212);
or U60 (N_60,In_1297,In_1258);
nand U61 (N_61,In_1303,In_353);
nand U62 (N_62,In_730,In_781);
or U63 (N_63,In_421,In_557);
and U64 (N_64,In_174,In_648);
xor U65 (N_65,In_183,In_661);
nand U66 (N_66,In_1259,In_223);
and U67 (N_67,In_687,In_329);
or U68 (N_68,In_401,In_905);
or U69 (N_69,In_607,In_949);
nor U70 (N_70,In_1145,In_652);
nor U71 (N_71,In_886,In_920);
nand U72 (N_72,In_683,In_556);
and U73 (N_73,In_35,In_1244);
and U74 (N_74,In_1418,In_1127);
nor U75 (N_75,In_866,In_328);
xnor U76 (N_76,In_1441,In_637);
nor U77 (N_77,In_171,In_653);
or U78 (N_78,In_793,In_1396);
or U79 (N_79,In_337,In_40);
nor U80 (N_80,In_253,In_216);
and U81 (N_81,In_1301,In_470);
or U82 (N_82,In_1210,In_257);
xnor U83 (N_83,In_1473,In_658);
nor U84 (N_84,In_927,In_1133);
xor U85 (N_85,In_895,In_1158);
xnor U86 (N_86,In_1161,In_761);
and U87 (N_87,In_316,In_359);
nand U88 (N_88,In_1089,In_1120);
nand U89 (N_89,In_113,In_1498);
and U90 (N_90,In_750,In_1007);
nor U91 (N_91,In_756,In_53);
nor U92 (N_92,In_259,In_342);
and U93 (N_93,In_935,In_1168);
or U94 (N_94,In_970,In_725);
and U95 (N_95,In_221,In_875);
nand U96 (N_96,In_411,In_1449);
nand U97 (N_97,In_1219,In_1043);
xor U98 (N_98,In_1190,In_581);
nor U99 (N_99,In_244,In_670);
and U100 (N_100,In_322,In_1474);
nor U101 (N_101,In_1294,In_226);
nand U102 (N_102,In_700,In_107);
or U103 (N_103,In_691,In_344);
nand U104 (N_104,In_672,In_151);
or U105 (N_105,In_1214,In_968);
nor U106 (N_106,In_195,In_1054);
or U107 (N_107,In_1184,In_994);
nor U108 (N_108,In_790,In_1348);
xor U109 (N_109,In_26,In_801);
nor U110 (N_110,In_747,In_1083);
xor U111 (N_111,In_2,In_178);
or U112 (N_112,In_204,In_1495);
and U113 (N_113,In_512,In_440);
nor U114 (N_114,In_1124,In_1472);
and U115 (N_115,In_297,In_371);
nand U116 (N_116,In_1012,In_1018);
or U117 (N_117,In_1309,In_1139);
or U118 (N_118,In_1065,In_367);
or U119 (N_119,In_519,In_874);
or U120 (N_120,In_462,In_410);
nor U121 (N_121,In_719,In_1427);
xor U122 (N_122,In_907,In_1355);
nand U123 (N_123,In_686,In_926);
nand U124 (N_124,In_1140,In_709);
xor U125 (N_125,In_388,In_1162);
nor U126 (N_126,In_1378,In_600);
nor U127 (N_127,In_1409,In_294);
or U128 (N_128,In_1395,In_1366);
nand U129 (N_129,In_991,In_161);
nor U130 (N_130,In_243,In_59);
xnor U131 (N_131,In_1117,In_693);
nor U132 (N_132,In_1468,In_1393);
nand U133 (N_133,In_638,In_270);
nor U134 (N_134,In_1492,In_1082);
xor U135 (N_135,In_1350,In_1483);
or U136 (N_136,In_491,In_831);
and U137 (N_137,In_433,In_385);
nor U138 (N_138,In_249,In_1115);
nor U139 (N_139,In_16,In_647);
nand U140 (N_140,In_43,In_1224);
and U141 (N_141,In_856,In_83);
and U142 (N_142,In_746,In_127);
or U143 (N_143,In_1255,In_889);
and U144 (N_144,In_1052,In_1481);
or U145 (N_145,In_1142,In_714);
nor U146 (N_146,In_664,In_639);
nand U147 (N_147,In_1277,In_41);
or U148 (N_148,In_304,In_534);
or U149 (N_149,In_1006,In_551);
nor U150 (N_150,In_711,In_224);
nand U151 (N_151,In_135,In_285);
and U152 (N_152,In_4,In_1375);
xor U153 (N_153,In_597,In_1181);
and U154 (N_154,In_954,In_573);
or U155 (N_155,In_992,In_893);
and U156 (N_156,In_541,In_989);
or U157 (N_157,In_1002,In_1112);
nand U158 (N_158,In_1146,In_309);
and U159 (N_159,In_215,In_540);
nand U160 (N_160,In_816,In_1320);
or U161 (N_161,In_586,In_8);
nor U162 (N_162,In_37,In_738);
or U163 (N_163,In_1167,In_906);
nor U164 (N_164,In_811,In_1452);
and U165 (N_165,In_1391,In_770);
nor U166 (N_166,In_1362,In_998);
nor U167 (N_167,In_1359,In_1307);
xnor U168 (N_168,In_77,In_1364);
or U169 (N_169,In_1268,In_1094);
and U170 (N_170,In_1496,In_424);
nand U171 (N_171,In_722,In_1058);
and U172 (N_172,In_1357,In_91);
or U173 (N_173,In_1147,In_312);
or U174 (N_174,In_971,In_1376);
or U175 (N_175,In_1337,In_369);
nor U176 (N_176,In_104,In_763);
or U177 (N_177,In_326,In_1199);
nand U178 (N_178,In_744,In_986);
and U179 (N_179,In_1067,In_1050);
nor U180 (N_180,In_864,In_619);
nand U181 (N_181,In_1302,In_898);
nor U182 (N_182,In_692,In_1414);
or U183 (N_183,In_1225,In_589);
nand U184 (N_184,In_103,In_1417);
xnor U185 (N_185,In_914,In_751);
nand U186 (N_186,In_495,In_579);
nor U187 (N_187,In_251,In_948);
nand U188 (N_188,In_629,In_1152);
nor U189 (N_189,In_1432,In_912);
nor U190 (N_190,In_44,In_872);
nor U191 (N_191,In_828,In_655);
or U192 (N_192,In_443,In_73);
nand U193 (N_193,In_1159,In_596);
nand U194 (N_194,In_917,In_563);
xor U195 (N_195,In_167,In_281);
or U196 (N_196,In_479,In_218);
nand U197 (N_197,In_1344,In_513);
xnor U198 (N_198,In_736,In_68);
and U199 (N_199,In_694,In_696);
or U200 (N_200,In_1232,In_529);
and U201 (N_201,In_430,In_1068);
and U202 (N_202,In_227,In_960);
nand U203 (N_203,In_669,In_102);
nand U204 (N_204,In_530,In_524);
or U205 (N_205,In_965,In_1469);
xor U206 (N_206,In_1478,In_1457);
xor U207 (N_207,In_599,In_1392);
nand U208 (N_208,In_650,In_780);
nor U209 (N_209,In_308,In_584);
xnor U210 (N_210,In_796,In_1381);
nor U211 (N_211,In_1280,In_602);
nor U212 (N_212,In_331,In_273);
or U213 (N_213,In_121,In_200);
nand U214 (N_214,In_49,In_788);
or U215 (N_215,In_740,In_116);
or U216 (N_216,In_1245,In_1374);
nor U217 (N_217,In_545,In_964);
xor U218 (N_218,In_305,In_358);
nand U219 (N_219,In_22,In_1160);
xnor U220 (N_220,In_445,In_1461);
xor U221 (N_221,In_625,In_36);
xnor U222 (N_222,In_794,In_1170);
or U223 (N_223,In_585,In_765);
nor U224 (N_224,In_565,In_890);
or U225 (N_225,In_643,In_608);
and U226 (N_226,In_284,In_487);
nor U227 (N_227,In_984,In_48);
nor U228 (N_228,In_1300,In_29);
or U229 (N_229,In_767,In_274);
nand U230 (N_230,In_583,In_465);
nor U231 (N_231,In_1370,In_293);
nor U232 (N_232,In_668,In_903);
nor U233 (N_233,In_206,In_560);
or U234 (N_234,In_649,In_386);
nand U235 (N_235,In_87,In_766);
and U236 (N_236,In_247,In_690);
and U237 (N_237,In_396,In_612);
nor U238 (N_238,In_577,In_1234);
nand U239 (N_239,In_363,In_1151);
nand U240 (N_240,In_241,In_1251);
nor U241 (N_241,In_977,In_979);
or U242 (N_242,In_955,In_1192);
xor U243 (N_243,In_362,In_1078);
or U244 (N_244,In_821,In_675);
nor U245 (N_245,In_263,In_1235);
nand U246 (N_246,In_1137,In_518);
or U247 (N_247,In_716,In_9);
nor U248 (N_248,In_158,In_240);
and U249 (N_249,In_1476,In_921);
xor U250 (N_250,In_380,In_33);
or U251 (N_251,In_393,In_517);
and U252 (N_252,In_1397,In_208);
nor U253 (N_253,In_1121,In_1271);
nor U254 (N_254,In_282,In_737);
nand U255 (N_255,In_633,In_980);
nor U256 (N_256,In_729,In_1466);
xnor U257 (N_257,In_1205,In_883);
or U258 (N_258,In_1111,In_1073);
nor U259 (N_259,In_900,In_1130);
and U260 (N_260,In_804,In_1421);
and U261 (N_261,In_651,In_853);
and U262 (N_262,In_527,In_861);
or U263 (N_263,In_814,In_909);
and U264 (N_264,In_833,In_1113);
nand U265 (N_265,In_147,In_119);
xor U266 (N_266,In_1299,In_999);
or U267 (N_267,In_1278,In_705);
or U268 (N_268,In_306,In_138);
xnor U269 (N_269,In_1486,In_806);
or U270 (N_270,In_120,In_67);
nor U271 (N_271,In_1293,In_510);
or U272 (N_272,In_1484,In_454);
xor U273 (N_273,In_473,In_42);
nor U274 (N_274,In_1022,In_707);
nand U275 (N_275,In_975,In_296);
and U276 (N_276,In_822,In_478);
xnor U277 (N_277,In_868,In_459);
or U278 (N_278,In_569,In_888);
nand U279 (N_279,In_879,In_1343);
or U280 (N_280,In_1084,In_1281);
and U281 (N_281,In_194,In_922);
or U282 (N_282,In_1338,In_972);
and U283 (N_283,In_548,In_232);
nand U284 (N_284,In_1231,In_759);
nand U285 (N_285,In_1213,In_1455);
nor U286 (N_286,In_325,In_1487);
and U287 (N_287,In_1428,In_1352);
and U288 (N_288,In_1382,In_112);
xnor U289 (N_289,In_745,In_1056);
nand U290 (N_290,In_51,In_1091);
and U291 (N_291,In_1141,In_100);
or U292 (N_292,In_724,In_869);
nor U293 (N_293,In_712,In_787);
and U294 (N_294,In_290,In_115);
nor U295 (N_295,In_911,In_749);
or U296 (N_296,In_95,In_758);
and U297 (N_297,In_713,In_1077);
and U298 (N_298,In_1358,In_1437);
and U299 (N_299,In_514,In_15);
xor U300 (N_300,In_1185,In_663);
nand U301 (N_301,In_1222,In_30);
nor U302 (N_302,In_1240,N_184);
or U303 (N_303,In_63,In_606);
nand U304 (N_304,N_133,In_1456);
or U305 (N_305,N_15,In_1027);
or U306 (N_306,In_434,N_235);
or U307 (N_307,In_307,In_98);
nand U308 (N_308,In_165,In_610);
nand U309 (N_309,In_137,In_1438);
or U310 (N_310,N_24,N_260);
or U311 (N_311,In_460,In_400);
or U312 (N_312,N_23,In_203);
or U313 (N_313,In_379,In_54);
or U314 (N_314,In_1497,In_628);
xor U315 (N_315,N_61,N_78);
and U316 (N_316,N_95,In_644);
xor U317 (N_317,In_85,In_365);
or U318 (N_318,In_374,In_1230);
nor U319 (N_319,In_841,In_343);
nand U320 (N_320,In_133,In_109);
and U321 (N_321,In_748,N_220);
or U322 (N_322,In_1227,In_1206);
nor U323 (N_323,In_149,N_251);
nor U324 (N_324,N_7,In_809);
nand U325 (N_325,In_1308,N_156);
or U326 (N_326,In_1257,N_17);
and U327 (N_327,In_576,In_1204);
nor U328 (N_328,In_81,In_1175);
nand U329 (N_329,In_407,In_908);
xor U330 (N_330,In_418,In_645);
or U331 (N_331,In_139,In_1413);
xnor U332 (N_332,In_1405,N_12);
or U333 (N_333,In_1114,N_232);
xor U334 (N_334,In_330,In_941);
xor U335 (N_335,In_721,N_10);
nand U336 (N_336,In_860,N_102);
nor U337 (N_337,In_1017,In_680);
or U338 (N_338,In_1459,In_236);
and U339 (N_339,In_86,N_25);
or U340 (N_340,In_345,In_1369);
nor U341 (N_341,In_1086,In_1129);
xnor U342 (N_342,In_1105,In_673);
or U343 (N_343,N_225,N_192);
nor U344 (N_344,In_214,In_1493);
nor U345 (N_345,In_1211,N_41);
nand U346 (N_346,In_71,In_202);
or U347 (N_347,In_0,In_1384);
xnor U348 (N_348,In_1020,In_982);
nand U349 (N_349,In_947,In_952);
nand U350 (N_350,In_899,In_419);
nor U351 (N_351,In_1329,N_190);
nor U352 (N_352,In_1347,In_1403);
nand U353 (N_353,In_1412,In_429);
and U354 (N_354,In_118,In_452);
nor U355 (N_355,In_1475,In_377);
nand U356 (N_356,N_155,In_490);
or U357 (N_357,N_66,In_800);
xnor U358 (N_358,In_395,N_65);
or U359 (N_359,In_536,N_214);
xor U360 (N_360,In_191,In_1470);
and U361 (N_361,In_646,In_538);
nand U362 (N_362,N_195,In_997);
xor U363 (N_363,In_552,In_1064);
and U364 (N_364,N_106,In_772);
or U365 (N_365,In_829,N_80);
or U366 (N_366,N_236,In_186);
nand U367 (N_367,In_258,In_558);
or U368 (N_368,N_230,N_108);
nand U369 (N_369,In_1042,In_605);
xnor U370 (N_370,In_1295,In_717);
xnor U371 (N_371,In_792,In_771);
nor U372 (N_372,In_1200,In_522);
or U373 (N_373,N_216,In_1328);
or U374 (N_374,N_196,In_500);
xor U375 (N_375,N_27,In_1061);
xnor U376 (N_376,N_29,N_53);
and U377 (N_377,In_84,In_1266);
or U378 (N_378,In_1274,N_60);
xnor U379 (N_379,In_1051,In_1186);
and U380 (N_380,In_162,In_1223);
or U381 (N_381,In_409,In_1093);
nand U382 (N_382,In_1216,N_204);
or U383 (N_383,In_805,In_498);
and U384 (N_384,In_595,In_145);
or U385 (N_385,In_1090,N_50);
nor U386 (N_386,N_54,In_489);
nor U387 (N_387,In_726,In_1136);
xnor U388 (N_388,In_988,In_335);
xnor U389 (N_389,In_376,In_580);
xor U390 (N_390,In_32,In_1040);
nor U391 (N_391,N_152,N_209);
and U392 (N_392,N_285,In_446);
nand U393 (N_393,In_1331,In_61);
nand U394 (N_394,In_1062,In_414);
nor U395 (N_395,In_1116,N_186);
nor U396 (N_396,In_254,N_5);
nor U397 (N_397,In_635,N_271);
and U398 (N_398,In_930,In_931);
nand U399 (N_399,In_803,In_1276);
nor U400 (N_400,N_163,In_832);
nand U401 (N_401,In_444,N_74);
or U402 (N_402,In_242,In_511);
nand U403 (N_403,N_39,In_292);
xor U404 (N_404,N_292,In_1189);
or U405 (N_405,In_23,In_1169);
and U406 (N_406,In_169,In_603);
or U407 (N_407,In_936,In_111);
nand U408 (N_408,In_564,In_1026);
xnor U409 (N_409,In_413,In_1041);
or U410 (N_410,In_373,In_447);
xor U411 (N_411,In_590,In_1436);
or U412 (N_412,N_121,In_148);
xnor U413 (N_413,In_1380,In_568);
nand U414 (N_414,In_928,In_555);
or U415 (N_415,N_168,In_734);
xor U416 (N_416,In_1106,In_268);
and U417 (N_417,N_208,In_1118);
or U418 (N_418,In_143,N_185);
nor U419 (N_419,In_1310,In_614);
nor U420 (N_420,In_134,In_426);
or U421 (N_421,In_389,In_463);
xnor U422 (N_422,In_1171,In_1148);
nor U423 (N_423,In_438,In_1265);
nand U424 (N_424,In_618,In_1306);
nand U425 (N_425,In_1379,In_46);
nor U426 (N_426,In_817,In_1182);
nor U427 (N_427,In_1226,N_188);
or U428 (N_428,In_1220,In_298);
xnor U429 (N_429,N_256,N_151);
xnor U430 (N_430,In_676,In_157);
or U431 (N_431,In_877,In_1322);
and U432 (N_432,In_532,In_350);
nor U433 (N_433,In_575,In_82);
xnor U434 (N_434,In_11,N_122);
and U435 (N_435,N_221,N_139);
nand U436 (N_436,In_1188,N_4);
xor U437 (N_437,In_1416,In_333);
nand U438 (N_438,In_485,In_117);
or U439 (N_439,N_176,In_731);
nand U440 (N_440,In_1311,In_482);
xor U441 (N_441,N_288,In_1372);
nand U442 (N_442,N_277,In_791);
xnor U443 (N_443,In_1425,In_1453);
or U444 (N_444,N_11,In_431);
nor U445 (N_445,In_1057,In_671);
and U446 (N_446,N_269,In_1433);
or U447 (N_447,N_147,In_876);
nand U448 (N_448,In_1408,In_559);
xor U449 (N_449,In_732,In_820);
or U450 (N_450,In_185,In_320);
nor U451 (N_451,In_578,In_1283);
and U452 (N_452,In_681,In_406);
nor U453 (N_453,In_1327,In_124);
and U454 (N_454,In_990,N_134);
and U455 (N_455,In_238,In_382);
and U456 (N_456,In_92,In_617);
xnor U457 (N_457,In_958,In_843);
and U458 (N_458,N_20,N_160);
and U459 (N_459,In_261,In_951);
and U460 (N_460,In_623,In_334);
nor U461 (N_461,In_1287,In_974);
xor U462 (N_462,In_812,In_136);
nor U463 (N_463,In_685,N_91);
and U464 (N_464,N_21,N_72);
and U465 (N_465,In_1176,In_913);
nor U466 (N_466,In_1149,In_815);
nand U467 (N_467,In_264,In_69);
or U468 (N_468,In_1150,In_141);
or U469 (N_469,In_93,N_104);
xor U470 (N_470,In_515,In_267);
or U471 (N_471,In_1047,In_1272);
nand U472 (N_472,In_231,In_188);
nor U473 (N_473,N_205,In_1217);
nand U474 (N_474,N_193,In_348);
nor U475 (N_475,In_1025,In_854);
or U476 (N_476,In_441,N_234);
xor U477 (N_477,N_46,In_542);
xor U478 (N_478,In_851,In_953);
or U479 (N_479,In_220,In_567);
and U480 (N_480,In_1060,In_1033);
nor U481 (N_481,In_657,In_837);
nand U482 (N_482,In_1447,In_347);
nand U483 (N_483,In_640,In_1402);
xor U484 (N_484,In_1030,In_873);
nor U485 (N_485,N_92,In_789);
xor U486 (N_486,In_70,In_1263);
nand U487 (N_487,N_242,N_244);
nor U488 (N_488,N_42,In_753);
or U489 (N_489,In_1228,In_1029);
nand U490 (N_490,In_237,In_266);
or U491 (N_491,N_237,In_1053);
xnor U492 (N_492,In_381,In_764);
and U493 (N_493,In_782,In_255);
nor U494 (N_494,In_1045,N_161);
nand U495 (N_495,In_1010,In_1003);
and U496 (N_496,In_182,In_1097);
and U497 (N_497,In_179,In_632);
nor U498 (N_498,In_235,In_642);
or U499 (N_499,In_497,In_1296);
nor U500 (N_500,N_117,In_1236);
nand U501 (N_501,N_127,N_13);
and U502 (N_502,In_408,In_13);
xnor U503 (N_503,In_354,N_58);
or U504 (N_504,In_64,N_274);
nor U505 (N_505,In_1491,In_423);
and U506 (N_506,In_47,In_1122);
xnor U507 (N_507,In_880,In_144);
nor U508 (N_508,N_142,In_546);
or U509 (N_509,In_1482,In_1305);
nand U510 (N_510,In_1499,N_68);
or U511 (N_511,In_272,In_682);
or U512 (N_512,N_206,In_435);
xor U513 (N_513,In_1389,N_84);
xor U514 (N_514,In_349,In_1342);
or U515 (N_515,In_336,In_1442);
or U516 (N_516,In_688,In_375);
nand U517 (N_517,In_225,In_878);
nor U518 (N_518,In_295,In_1319);
xor U519 (N_519,In_74,In_1490);
or U520 (N_520,N_90,N_181);
xnor U521 (N_521,N_76,In_52);
and U522 (N_522,In_1477,In_768);
nand U523 (N_523,In_356,In_269);
xor U524 (N_524,N_241,In_1464);
nand U525 (N_525,N_197,In_469);
or U526 (N_526,N_71,N_137);
nor U527 (N_527,In_1288,In_256);
nand U528 (N_528,In_1373,N_296);
nand U529 (N_529,In_904,In_718);
or U530 (N_530,In_383,In_1267);
or U531 (N_531,In_1180,In_474);
xor U532 (N_532,N_231,N_298);
nor U533 (N_533,In_553,In_1195);
and U534 (N_534,In_547,N_62);
nand U535 (N_535,In_170,In_205);
and U536 (N_536,In_428,In_757);
xnor U537 (N_537,In_286,In_65);
xnor U538 (N_538,In_291,In_684);
xor U539 (N_539,In_187,In_715);
and U540 (N_540,N_33,N_273);
nor U541 (N_541,In_416,In_624);
and U542 (N_542,N_140,In_175);
or U543 (N_543,In_808,In_834);
nand U544 (N_544,In_1203,In_1254);
nand U545 (N_545,N_154,N_99);
and U546 (N_546,In_62,In_1356);
nor U547 (N_547,In_1422,In_289);
and U548 (N_548,In_384,In_887);
xor U549 (N_549,In_234,N_6);
or U550 (N_550,In_1318,In_180);
or U551 (N_551,In_287,In_1172);
xnor U552 (N_552,In_846,In_160);
or U553 (N_553,In_679,N_259);
xnor U554 (N_554,In_591,In_896);
nor U555 (N_555,N_279,In_213);
and U556 (N_556,In_660,In_1187);
and U557 (N_557,In_403,In_415);
or U558 (N_558,In_976,In_483);
nor U559 (N_559,In_959,In_902);
nand U560 (N_560,In_1066,In_492);
and U561 (N_561,In_311,In_502);
nand U562 (N_562,In_1371,In_1059);
and U563 (N_563,In_493,In_101);
or U564 (N_564,In_1092,In_1080);
nand U565 (N_565,N_22,In_897);
nor U566 (N_566,In_508,In_6);
nand U567 (N_567,N_100,In_146);
nor U568 (N_568,In_937,In_387);
nor U569 (N_569,In_1075,In_351);
xor U570 (N_570,In_1411,In_477);
nor U571 (N_571,In_1419,In_1451);
nand U572 (N_572,In_466,In_1131);
xor U573 (N_573,In_1119,N_229);
xnor U574 (N_574,In_1346,In_1314);
nand U575 (N_575,In_1284,N_83);
nor U576 (N_576,N_247,In_250);
nand U577 (N_577,N_144,In_1044);
nand U578 (N_578,In_942,In_774);
xnor U579 (N_579,In_245,In_827);
nand U580 (N_580,In_570,In_863);
xor U581 (N_581,In_1016,In_1174);
nand U582 (N_582,N_253,In_594);
xor U583 (N_583,In_1049,In_1354);
and U584 (N_584,N_162,N_243);
and U585 (N_585,In_799,N_217);
xor U586 (N_586,In_38,In_96);
nor U587 (N_587,In_950,N_110);
and U588 (N_588,N_170,N_120);
xor U589 (N_589,In_303,N_276);
nor U590 (N_590,In_1081,In_1153);
or U591 (N_591,In_1247,In_754);
or U592 (N_592,N_43,N_126);
xnor U593 (N_593,In_1385,In_1039);
xnor U594 (N_594,In_755,In_929);
nor U595 (N_595,In_467,N_112);
nor U596 (N_596,In_1011,N_40);
or U597 (N_597,In_1390,N_19);
and U598 (N_598,N_30,In_1383);
or U599 (N_599,In_966,In_978);
and U600 (N_600,In_278,N_512);
nor U601 (N_601,N_18,N_410);
nand U602 (N_602,N_215,In_105);
nand U603 (N_603,N_339,In_1335);
or U604 (N_604,N_352,In_332);
nand U605 (N_605,N_383,In_1212);
and U606 (N_606,N_596,In_995);
or U607 (N_607,N_581,N_498);
and U608 (N_608,N_320,In_1243);
and U609 (N_609,N_57,N_447);
nor U610 (N_610,In_932,In_210);
and U611 (N_611,N_562,In_72);
nand U612 (N_612,In_417,In_1109);
nor U613 (N_613,In_230,N_385);
or U614 (N_614,N_541,In_1173);
or U615 (N_615,N_573,N_489);
nand U616 (N_616,N_200,N_371);
xor U617 (N_617,N_449,N_218);
or U618 (N_618,N_89,In_1386);
or U619 (N_619,N_429,In_1454);
nor U620 (N_620,In_1467,N_557);
or U621 (N_621,N_389,N_522);
and U622 (N_622,In_129,N_566);
or U623 (N_623,N_294,In_1423);
and U624 (N_624,In_1069,In_1363);
or U625 (N_625,In_302,N_36);
and U626 (N_626,N_169,N_480);
or U627 (N_627,N_345,N_159);
and U628 (N_628,N_378,N_331);
and U629 (N_629,N_212,In_1229);
xor U630 (N_630,N_107,In_587);
or U631 (N_631,N_337,In_934);
and U632 (N_632,In_1248,N_474);
nor U633 (N_633,In_699,N_0);
nor U634 (N_634,In_901,N_299);
nor U635 (N_635,In_1191,In_1291);
or U636 (N_636,In_12,N_426);
xnor U637 (N_637,In_910,N_481);
xnor U638 (N_638,N_403,N_384);
nand U639 (N_639,N_487,In_1196);
xnor U640 (N_640,N_490,In_17);
nor U641 (N_641,N_388,In_192);
or U642 (N_642,N_550,In_1448);
nand U643 (N_643,N_433,N_419);
and U644 (N_644,N_310,In_420);
nor U645 (N_645,In_321,In_58);
and U646 (N_646,N_521,In_341);
or U647 (N_647,N_213,In_252);
nor U648 (N_648,N_338,N_262);
nand U649 (N_649,In_963,In_1100);
xnor U650 (N_650,In_775,In_56);
or U651 (N_651,In_1183,N_402);
and U652 (N_652,In_301,In_506);
xor U653 (N_653,N_219,N_48);
nor U654 (N_654,In_626,N_308);
xnor U655 (N_655,In_702,N_495);
nor U656 (N_656,In_509,In_706);
nor U657 (N_657,N_435,In_1340);
nand U658 (N_658,In_1132,In_1292);
or U659 (N_659,In_1208,N_471);
nand U660 (N_660,In_539,In_75);
and U661 (N_661,In_698,In_176);
nor U662 (N_662,In_1298,In_439);
nor U663 (N_663,N_129,In_1324);
nor U664 (N_664,N_572,N_406);
and U665 (N_665,N_393,In_938);
or U666 (N_666,In_993,In_24);
nand U667 (N_667,In_1446,N_281);
nor U668 (N_668,In_704,N_94);
xnor U669 (N_669,In_425,In_760);
nor U670 (N_670,In_1128,In_956);
xor U671 (N_671,N_451,In_1103);
and U672 (N_672,N_85,In_1238);
xnor U673 (N_673,N_556,N_202);
and U674 (N_674,N_228,N_407);
nand U675 (N_675,N_64,In_181);
nor U676 (N_676,N_575,N_366);
nor U677 (N_677,N_325,N_398);
and U678 (N_678,In_1135,N_355);
or U679 (N_679,In_1063,In_476);
nor U680 (N_680,In_1055,N_536);
nand U681 (N_681,In_229,In_1098);
nor U682 (N_682,N_254,N_98);
nand U683 (N_683,In_925,N_179);
or U684 (N_684,In_521,N_413);
or U685 (N_685,N_199,In_1462);
and U686 (N_686,In_943,N_263);
nor U687 (N_687,In_45,In_1138);
xor U688 (N_688,N_382,In_1404);
xor U689 (N_689,N_317,In_1285);
and U690 (N_690,In_1479,In_1071);
or U691 (N_691,In_378,N_96);
xnor U692 (N_692,In_432,N_145);
nor U693 (N_693,In_275,In_620);
or U694 (N_694,N_315,In_773);
and U695 (N_695,N_466,In_21);
or U696 (N_696,In_1341,N_509);
nor U697 (N_697,N_238,In_449);
nor U698 (N_698,N_286,N_559);
nor U699 (N_699,In_1256,N_82);
nor U700 (N_700,N_322,In_391);
nand U701 (N_701,N_397,N_529);
or U702 (N_702,N_307,In_1032);
nor U703 (N_703,N_484,N_390);
xor U704 (N_704,In_168,N_539);
and U705 (N_705,In_1038,N_118);
nor U706 (N_706,In_209,N_290);
nor U707 (N_707,In_1028,In_1110);
or U708 (N_708,N_386,In_279);
nand U709 (N_709,In_1108,In_1163);
nand U710 (N_710,N_592,In_436);
nand U711 (N_711,N_555,In_177);
nor U712 (N_712,N_75,N_38);
xor U713 (N_713,In_458,N_207);
nor U714 (N_714,N_128,In_1072);
nand U715 (N_715,In_189,In_708);
nor U716 (N_716,N_63,N_347);
xnor U717 (N_717,N_488,N_577);
nand U718 (N_718,N_125,In_1102);
and U719 (N_719,N_565,N_376);
nand U720 (N_720,In_1361,N_93);
or U721 (N_721,In_370,N_172);
xnor U722 (N_722,N_587,In_1009);
and U723 (N_723,N_153,N_59);
and U724 (N_724,N_305,In_19);
or U725 (N_725,N_2,In_1445);
and U726 (N_726,In_1035,N_37);
nor U727 (N_727,N_324,N_270);
nand U728 (N_728,N_157,N_578);
or U729 (N_729,In_1178,N_264);
nand U730 (N_730,In_1485,N_440);
nand U731 (N_731,N_227,In_246);
and U732 (N_732,N_593,N_545);
and U733 (N_733,N_396,In_1036);
xor U734 (N_734,N_450,In_50);
or U735 (N_735,N_551,N_86);
nand U736 (N_736,N_114,N_586);
nand U737 (N_737,In_627,In_262);
and U738 (N_738,In_1440,N_493);
nor U739 (N_739,N_143,In_703);
nor U740 (N_740,In_1242,N_470);
nor U741 (N_741,N_417,N_252);
or U742 (N_742,In_1365,In_1154);
xnor U743 (N_743,N_375,In_528);
or U744 (N_744,N_165,In_422);
nor U745 (N_745,In_450,In_826);
nand U746 (N_746,In_402,In_1321);
nand U747 (N_747,In_505,N_547);
xnor U748 (N_748,In_940,In_1031);
and U749 (N_749,In_219,N_569);
nand U750 (N_750,In_813,N_377);
nor U751 (N_751,N_524,N_588);
nor U752 (N_752,N_56,In_55);
or U753 (N_753,N_295,N_424);
or U754 (N_754,N_591,N_67);
and U755 (N_755,N_462,N_585);
nor U756 (N_756,In_723,In_884);
nand U757 (N_757,N_544,In_366);
nor U758 (N_758,N_239,N_138);
nand U759 (N_759,N_367,In_823);
nand U760 (N_760,In_368,In_919);
nor U761 (N_761,N_554,N_431);
xnor U762 (N_762,In_1480,N_394);
or U763 (N_763,In_480,N_479);
xor U764 (N_764,N_261,In_807);
or U765 (N_765,In_437,N_226);
nand U766 (N_766,In_131,In_1401);
or U767 (N_767,In_894,In_847);
or U768 (N_768,N_284,In_1304);
or U769 (N_769,In_340,In_1123);
xnor U770 (N_770,In_207,In_1450);
xor U771 (N_771,N_415,In_1005);
and U772 (N_772,In_1165,N_428);
and U773 (N_773,N_416,N_579);
xor U774 (N_774,In_1262,In_840);
and U775 (N_775,In_1394,In_1194);
or U776 (N_776,In_891,N_458);
nand U777 (N_777,In_442,N_459);
nand U778 (N_778,In_836,In_1000);
xnor U779 (N_779,In_1246,N_330);
xnor U780 (N_780,In_1209,In_198);
nor U781 (N_781,N_457,N_28);
or U782 (N_782,In_741,In_451);
xnor U783 (N_783,In_516,N_87);
or U784 (N_784,N_571,In_1104);
nand U785 (N_785,In_123,N_594);
and U786 (N_786,In_601,In_14);
nand U787 (N_787,N_548,N_446);
and U788 (N_788,In_390,In_1353);
nand U789 (N_789,N_327,In_488);
xnor U790 (N_790,N_8,In_248);
nand U791 (N_791,In_845,N_527);
nand U792 (N_792,In_957,N_420);
nand U793 (N_793,In_79,N_411);
or U794 (N_794,N_583,N_278);
xnor U795 (N_795,N_513,N_370);
and U796 (N_796,N_131,In_611);
or U797 (N_797,N_344,N_359);
nand U798 (N_798,In_150,In_742);
nor U799 (N_799,In_277,N_434);
or U800 (N_800,N_364,In_739);
and U801 (N_801,N_265,N_341);
nand U802 (N_802,N_174,N_353);
nor U803 (N_803,N_334,N_405);
and U804 (N_804,In_1021,In_622);
nor U805 (N_805,In_549,In_265);
xor U806 (N_806,N_267,N_499);
xnor U807 (N_807,N_520,N_14);
xnor U808 (N_808,In_57,In_870);
nor U809 (N_809,In_233,N_201);
xor U810 (N_810,In_1004,N_531);
xor U811 (N_811,N_472,N_70);
xor U812 (N_812,N_477,N_525);
or U813 (N_813,N_283,In_616);
or U814 (N_814,N_31,N_350);
and U815 (N_815,In_5,N_590);
and U816 (N_816,N_47,N_537);
nor U817 (N_817,N_368,In_153);
nor U818 (N_818,N_52,In_1134);
xnor U819 (N_819,In_1241,N_148);
nand U820 (N_820,N_469,N_306);
and U821 (N_821,N_356,N_304);
and U822 (N_822,In_1046,In_339);
xnor U823 (N_823,N_182,In_399);
nand U824 (N_824,N_348,In_1279);
nand U825 (N_825,In_531,N_570);
nand U826 (N_826,In_1074,N_507);
and U827 (N_827,In_923,N_515);
and U828 (N_828,In_945,In_60);
xnor U829 (N_829,In_1037,N_198);
nor U830 (N_830,In_324,In_300);
xor U831 (N_831,N_523,N_343);
and U832 (N_832,N_248,In_697);
nor U833 (N_833,N_475,In_525);
or U834 (N_834,In_1270,N_69);
nand U835 (N_835,In_27,N_503);
or U836 (N_836,N_399,N_282);
and U837 (N_837,N_316,In_39);
or U838 (N_838,In_398,In_228);
or U839 (N_839,In_468,In_987);
and U840 (N_840,N_369,In_710);
xnor U841 (N_841,In_795,In_1444);
nor U842 (N_842,In_571,N_346);
nor U843 (N_843,N_275,N_135);
nand U844 (N_844,N_483,N_506);
or U845 (N_845,N_476,N_3);
or U846 (N_846,In_604,In_239);
nand U847 (N_847,In_114,In_1332);
or U848 (N_848,In_967,In_427);
nor U849 (N_849,In_1197,N_448);
nand U850 (N_850,N_223,In_662);
nand U851 (N_851,In_1125,In_172);
or U852 (N_852,N_211,In_1489);
nor U853 (N_853,In_504,N_560);
nor U854 (N_854,N_576,N_311);
and U855 (N_855,In_631,N_105);
nor U856 (N_856,In_217,N_518);
xor U857 (N_857,In_996,In_533);
nor U858 (N_858,In_1269,In_665);
nor U859 (N_859,N_599,N_467);
nand U860 (N_860,N_444,In_1095);
nor U861 (N_861,N_191,In_88);
and U862 (N_862,N_597,N_77);
xnor U863 (N_863,N_441,N_508);
or U864 (N_864,In_786,In_314);
nor U865 (N_865,In_543,N_32);
nor U866 (N_866,In_404,N_132);
xor U867 (N_867,N_319,In_76);
and U868 (N_868,N_297,N_561);
nand U869 (N_869,In_1387,In_537);
nor U870 (N_870,N_329,In_1465);
nand U871 (N_871,In_1166,In_486);
nand U872 (N_872,In_973,N_210);
and U873 (N_873,In_762,N_26);
and U874 (N_874,In_1471,In_392);
xnor U875 (N_875,N_540,In_1249);
nand U876 (N_876,N_412,N_414);
nor U877 (N_877,In_574,In_810);
and U878 (N_878,In_593,N_425);
xnor U879 (N_879,N_233,N_9);
or U880 (N_880,N_314,In_1434);
xor U881 (N_881,N_421,In_94);
xnor U882 (N_882,N_504,N_460);
nand U883 (N_883,N_580,In_1076);
or U884 (N_884,N_222,N_497);
nand U885 (N_885,N_123,N_392);
and U886 (N_886,N_249,N_543);
xor U887 (N_887,N_49,N_465);
nor U888 (N_888,N_568,N_113);
or U889 (N_889,In_983,In_1252);
or U890 (N_890,In_66,N_564);
or U891 (N_891,N_486,N_354);
nand U892 (N_892,In_1,N_34);
nand U893 (N_893,In_184,In_752);
xnor U894 (N_894,N_173,N_35);
nand U895 (N_895,N_340,N_500);
nand U896 (N_896,N_391,N_177);
or U897 (N_897,In_1388,In_156);
and U898 (N_898,In_728,In_634);
and U899 (N_899,In_1048,In_1207);
and U900 (N_900,N_654,In_271);
nor U901 (N_901,N_641,N_656);
or U902 (N_902,In_641,N_784);
nand U903 (N_903,In_1312,N_817);
nand U904 (N_904,N_764,In_1198);
xor U905 (N_905,N_603,N_582);
xnor U906 (N_906,N_806,N_792);
and U907 (N_907,N_146,N_695);
or U908 (N_908,N_240,In_882);
and U909 (N_909,N_250,N_627);
xor U910 (N_910,In_598,N_430);
xor U911 (N_911,N_778,N_595);
xnor U912 (N_912,N_834,N_395);
nand U913 (N_913,N_268,N_404);
xor U914 (N_914,N_838,In_1014);
or U915 (N_915,N_718,N_762);
and U916 (N_916,N_141,N_625);
nand U917 (N_917,In_327,N_187);
xnor U918 (N_918,N_609,N_829);
nor U919 (N_919,In_784,N_532);
and U920 (N_920,N_701,N_516);
xnor U921 (N_921,N_822,N_584);
or U922 (N_922,N_700,In_201);
nor U923 (N_923,N_867,N_485);
nand U924 (N_924,N_633,N_837);
or U925 (N_925,N_845,N_705);
xor U926 (N_926,N_719,N_683);
nand U927 (N_927,N_671,N_801);
xor U928 (N_928,N_149,N_864);
and U929 (N_929,N_749,N_883);
or U930 (N_930,In_1430,In_1024);
xnor U931 (N_931,N_178,N_589);
nand U932 (N_932,N_715,N_688);
xnor U933 (N_933,N_797,N_635);
or U934 (N_934,In_1250,In_592);
nand U935 (N_935,In_733,N_534);
nor U936 (N_936,In_152,N_567);
nor U937 (N_937,N_847,In_199);
and U938 (N_938,N_678,N_739);
and U939 (N_939,N_620,N_381);
xnor U940 (N_940,In_818,In_346);
xor U941 (N_941,N_628,N_362);
nor U942 (N_942,In_885,N_681);
and U943 (N_943,N_626,In_97);
or U944 (N_944,N_839,N_731);
nand U945 (N_945,N_850,N_763);
and U946 (N_946,N_728,N_863);
nor U947 (N_947,N_538,N_614);
xor U948 (N_948,N_245,In_106);
nor U949 (N_949,N_546,In_196);
and U950 (N_950,N_736,N_755);
nand U951 (N_951,N_783,N_703);
and U952 (N_952,N_750,N_618);
or U953 (N_953,In_1400,N_716);
or U954 (N_954,In_126,N_437);
xor U955 (N_955,N_709,N_840);
or U956 (N_956,N_781,N_194);
nand U957 (N_957,N_667,N_598);
or U958 (N_958,N_861,N_166);
nor U959 (N_959,N_427,N_707);
and U960 (N_960,N_613,N_768);
nor U961 (N_961,N_349,N_807);
nand U962 (N_962,In_283,N_103);
nand U963 (N_963,N_636,N_663);
xnor U964 (N_964,N_738,N_732);
nor U965 (N_965,N_835,N_335);
or U966 (N_966,In_871,N_640);
nand U967 (N_967,In_1143,N_757);
or U968 (N_968,In_155,N_436);
xnor U969 (N_969,N_824,N_798);
nor U970 (N_970,In_862,N_789);
xor U971 (N_971,N_727,N_786);
nand U972 (N_972,N_841,N_702);
nor U973 (N_973,N_312,N_492);
nand U974 (N_974,In_695,In_654);
and U975 (N_975,N_836,In_211);
nand U976 (N_976,In_779,In_260);
nand U977 (N_977,In_319,N_675);
and U978 (N_978,N_409,N_891);
nand U979 (N_979,In_918,N_44);
xnor U980 (N_980,N_203,N_810);
xnor U981 (N_981,N_878,N_119);
nor U982 (N_982,N_258,N_300);
nand U983 (N_983,N_687,N_638);
or U984 (N_984,In_501,N_699);
and U985 (N_985,N_690,N_623);
nor U986 (N_986,In_99,N_765);
xor U987 (N_987,In_130,N_16);
and U988 (N_988,N_860,N_189);
xnor U989 (N_989,N_720,N_51);
xor U990 (N_990,N_610,N_766);
or U991 (N_991,N_788,N_514);
nand U992 (N_992,N_88,N_183);
nand U993 (N_993,N_442,N_857);
nand U994 (N_994,N_790,N_624);
nor U995 (N_995,N_361,In_481);
and U996 (N_996,In_916,In_412);
nand U997 (N_997,N_893,In_550);
nor U998 (N_998,N_898,N_747);
xnor U999 (N_999,In_132,N_713);
xor U1000 (N_1000,N_723,N_109);
or U1001 (N_1001,In_985,N_502);
nor U1002 (N_1002,N_528,N_124);
and U1003 (N_1003,N_97,N_832);
xor U1004 (N_1004,N_722,N_814);
xor U1005 (N_1005,N_323,N_879);
nand U1006 (N_1006,N_771,In_961);
or U1007 (N_1007,N_775,N_712);
xnor U1008 (N_1008,N_733,N_272);
xor U1009 (N_1009,In_609,In_850);
or U1010 (N_1010,N_328,N_443);
nand U1011 (N_1011,N_735,N_884);
nand U1012 (N_1012,N_363,N_679);
xor U1013 (N_1013,In_1008,N_849);
nand U1014 (N_1014,In_494,N_740);
nor U1015 (N_1015,N_744,N_647);
nor U1016 (N_1016,In_323,N_453);
xnor U1017 (N_1017,N_111,In_1494);
nand U1018 (N_1018,N_828,N_869);
nand U1019 (N_1019,In_364,N_795);
xnor U1020 (N_1020,In_110,N_130);
xnor U1021 (N_1021,N_655,In_666);
nor U1022 (N_1022,N_608,N_530);
nand U1023 (N_1023,N_351,N_676);
and U1024 (N_1024,N_606,In_838);
nor U1025 (N_1025,In_1215,N_800);
and U1026 (N_1026,N_666,N_650);
nor U1027 (N_1027,N_365,N_380);
and U1028 (N_1028,N_805,N_897);
xor U1029 (N_1029,N_820,In_1001);
xor U1030 (N_1030,N_890,In_523);
nor U1031 (N_1031,N_372,N_680);
nand U1032 (N_1032,N_721,In_621);
xnor U1033 (N_1033,N_646,N_756);
xnor U1034 (N_1034,N_802,N_164);
nor U1035 (N_1035,In_1313,N_1);
xnor U1036 (N_1036,N_856,N_400);
nor U1037 (N_1037,N_604,N_379);
nor U1038 (N_1038,N_882,N_692);
xnor U1039 (N_1039,N_895,N_754);
nand U1040 (N_1040,In_944,N_478);
or U1041 (N_1041,N_704,N_611);
or U1042 (N_1042,In_720,In_701);
xnor U1043 (N_1043,N_387,N_813);
xnor U1044 (N_1044,N_794,N_892);
xnor U1045 (N_1045,In_572,In_1282);
nor U1046 (N_1046,N_658,N_651);
and U1047 (N_1047,N_664,In_776);
nor U1048 (N_1048,In_484,N_896);
or U1049 (N_1049,N_357,In_317);
nand U1050 (N_1050,N_616,In_1406);
and U1051 (N_1051,In_824,In_1088);
or U1052 (N_1052,N_136,N_843);
or U1053 (N_1053,N_742,N_491);
or U1054 (N_1054,N_708,In_946);
or U1055 (N_1055,N_714,In_1407);
and U1056 (N_1056,N_336,N_770);
or U1057 (N_1057,N_621,N_619);
or U1058 (N_1058,N_662,In_313);
nand U1059 (N_1059,N_830,In_1426);
nand U1060 (N_1060,N_661,N_266);
nor U1061 (N_1061,N_482,In_299);
nand U1062 (N_1062,N_865,N_574);
nor U1063 (N_1063,N_734,N_438);
or U1064 (N_1064,In_1410,N_684);
or U1065 (N_1065,N_808,In_461);
nor U1066 (N_1066,In_582,In_858);
xnor U1067 (N_1067,In_394,N_876);
nor U1068 (N_1068,N_558,In_405);
nand U1069 (N_1069,N_649,N_842);
or U1070 (N_1070,In_561,N_871);
xor U1071 (N_1071,In_588,N_852);
or U1072 (N_1072,N_677,N_673);
nand U1073 (N_1073,In_357,N_823);
and U1074 (N_1074,N_774,N_746);
nor U1075 (N_1075,N_793,N_669);
or U1076 (N_1076,In_855,N_706);
and U1077 (N_1077,N_710,N_759);
xnor U1078 (N_1078,N_657,N_542);
and U1079 (N_1079,N_686,N_158);
nand U1080 (N_1080,In_1264,N_748);
and U1081 (N_1081,N_445,In_222);
and U1082 (N_1082,In_1023,In_455);
nor U1083 (N_1083,In_636,N_885);
and U1084 (N_1084,N_854,In_159);
nand U1085 (N_1085,In_1013,N_615);
nor U1086 (N_1086,In_830,N_461);
or U1087 (N_1087,In_1101,N_873);
and U1088 (N_1088,In_1079,N_870);
or U1089 (N_1089,N_517,In_1034);
and U1090 (N_1090,N_553,In_613);
nand U1091 (N_1091,N_725,N_639);
or U1092 (N_1092,N_332,N_894);
xor U1093 (N_1093,N_672,In_1273);
xor U1094 (N_1094,N_552,N_293);
nand U1095 (N_1095,N_693,In_656);
nor U1096 (N_1096,N_776,N_729);
or U1097 (N_1097,N_605,N_607);
and U1098 (N_1098,N_401,N_496);
nand U1099 (N_1099,N_318,N_321);
xnor U1100 (N_1100,N_642,N_785);
and U1101 (N_1101,N_745,N_629);
and U1102 (N_1102,N_289,N_665);
or U1103 (N_1103,N_510,In_924);
or U1104 (N_1104,In_630,N_886);
nor U1105 (N_1105,N_224,N_511);
or U1106 (N_1106,N_180,N_150);
xnor U1107 (N_1107,N_333,N_408);
nand U1108 (N_1108,N_81,N_769);
nor U1109 (N_1109,N_772,N_862);
xor U1110 (N_1110,N_780,N_811);
xor U1111 (N_1111,N_115,N_833);
xor U1112 (N_1112,In_859,N_812);
nand U1113 (N_1113,N_549,N_612);
nand U1114 (N_1114,N_859,N_696);
and U1115 (N_1115,N_652,N_779);
nor U1116 (N_1116,N_79,In_526);
or U1117 (N_1117,N_45,In_1399);
nor U1118 (N_1118,N_670,N_563);
and U1119 (N_1119,N_851,In_1398);
and U1120 (N_1120,N_535,N_287);
and U1121 (N_1121,N_473,N_101);
or U1122 (N_1122,N_533,N_777);
and U1123 (N_1123,N_825,N_455);
xnor U1124 (N_1124,N_358,N_726);
and U1125 (N_1125,In_1424,N_758);
xnor U1126 (N_1126,N_55,N_602);
nor U1127 (N_1127,In_3,In_1435);
nor U1128 (N_1128,N_831,N_804);
nor U1129 (N_1129,N_631,N_432);
or U1130 (N_1130,In_798,N_724);
xnor U1131 (N_1131,N_373,N_648);
and U1132 (N_1132,N_601,N_257);
and U1133 (N_1133,N_753,In_1345);
xnor U1134 (N_1134,N_456,In_25);
nand U1135 (N_1135,N_175,In_1439);
and U1136 (N_1136,N_116,N_760);
or U1137 (N_1137,N_877,N_819);
or U1138 (N_1138,In_1360,N_303);
and U1139 (N_1139,N_313,In_797);
or U1140 (N_1140,In_1193,N_698);
nand U1141 (N_1141,In_166,In_1463);
nand U1142 (N_1142,N_809,N_691);
nor U1143 (N_1143,N_875,N_682);
and U1144 (N_1144,N_791,In_496);
or U1145 (N_1145,N_171,N_787);
xor U1146 (N_1146,N_632,N_660);
nand U1147 (N_1147,In_7,N_643);
xor U1148 (N_1148,In_1155,In_164);
nor U1149 (N_1149,N_844,N_803);
xnor U1150 (N_1150,N_302,N_752);
nor U1151 (N_1151,N_741,N_888);
and U1152 (N_1152,N_246,N_796);
nand U1153 (N_1153,N_653,N_422);
xnor U1154 (N_1154,N_846,N_622);
or U1155 (N_1155,N_848,N_881);
nand U1156 (N_1156,N_617,N_855);
or U1157 (N_1157,In_835,In_1253);
and U1158 (N_1158,In_1164,In_280);
or U1159 (N_1159,N_342,N_767);
nand U1160 (N_1160,N_659,In_1015);
and U1161 (N_1161,In_678,N_866);
xor U1162 (N_1162,N_526,N_309);
xor U1163 (N_1163,N_464,N_600);
xor U1164 (N_1164,In_819,N_880);
or U1165 (N_1165,N_668,N_637);
nor U1166 (N_1166,N_899,N_685);
and U1167 (N_1167,N_326,N_674);
nand U1168 (N_1168,N_374,N_730);
nand U1169 (N_1169,N_645,N_782);
or U1170 (N_1170,N_821,N_717);
nand U1171 (N_1171,N_255,N_454);
and U1172 (N_1172,N_853,In_1202);
and U1173 (N_1173,N_418,N_423);
or U1174 (N_1174,N_773,In_844);
nand U1175 (N_1175,N_816,N_463);
xor U1176 (N_1176,In_939,In_20);
nand U1177 (N_1177,N_291,In_154);
xnor U1178 (N_1178,N_874,N_494);
or U1179 (N_1179,In_743,N_858);
and U1180 (N_1180,N_439,N_452);
nand U1181 (N_1181,N_889,N_872);
xnor U1182 (N_1182,N_167,N_360);
nand U1183 (N_1183,N_301,In_1458);
and U1184 (N_1184,N_519,N_689);
nand U1185 (N_1185,In_667,In_457);
xor U1186 (N_1186,N_644,N_694);
xnor U1187 (N_1187,In_1334,N_697);
nand U1188 (N_1188,N_826,N_799);
xnor U1189 (N_1189,N_751,N_818);
or U1190 (N_1190,N_737,In_1316);
nand U1191 (N_1191,N_280,In_1488);
nand U1192 (N_1192,In_1339,N_501);
xor U1193 (N_1193,N_634,N_887);
nand U1194 (N_1194,N_827,N_73);
and U1195 (N_1195,N_505,In_1221);
or U1196 (N_1196,N_761,N_868);
xnor U1197 (N_1197,N_630,N_815);
xor U1198 (N_1198,N_743,N_711);
nor U1199 (N_1199,In_554,N_468);
nor U1200 (N_1200,N_1098,N_901);
nand U1201 (N_1201,N_1026,N_986);
and U1202 (N_1202,N_977,N_919);
nand U1203 (N_1203,N_924,N_973);
xor U1204 (N_1204,N_972,N_988);
xor U1205 (N_1205,N_949,N_1024);
xor U1206 (N_1206,N_1015,N_942);
nand U1207 (N_1207,N_948,N_938);
or U1208 (N_1208,N_1171,N_1181);
nand U1209 (N_1209,N_1004,N_1187);
nor U1210 (N_1210,N_1000,N_960);
xor U1211 (N_1211,N_1137,N_1174);
nand U1212 (N_1212,N_1168,N_1061);
xor U1213 (N_1213,N_1057,N_931);
or U1214 (N_1214,N_1089,N_1052);
nand U1215 (N_1215,N_1065,N_962);
or U1216 (N_1216,N_922,N_914);
nor U1217 (N_1217,N_1009,N_990);
or U1218 (N_1218,N_917,N_1092);
xnor U1219 (N_1219,N_936,N_1049);
xnor U1220 (N_1220,N_1097,N_979);
or U1221 (N_1221,N_1178,N_980);
xnor U1222 (N_1222,N_1063,N_1161);
or U1223 (N_1223,N_991,N_1190);
nor U1224 (N_1224,N_964,N_900);
xnor U1225 (N_1225,N_1184,N_928);
xor U1226 (N_1226,N_933,N_1058);
nor U1227 (N_1227,N_910,N_1101);
and U1228 (N_1228,N_995,N_1122);
xor U1229 (N_1229,N_1016,N_1060);
nand U1230 (N_1230,N_1199,N_981);
and U1231 (N_1231,N_1055,N_1121);
or U1232 (N_1232,N_957,N_968);
nand U1233 (N_1233,N_1076,N_955);
and U1234 (N_1234,N_1054,N_1160);
nor U1235 (N_1235,N_999,N_918);
xnor U1236 (N_1236,N_1093,N_956);
nand U1237 (N_1237,N_932,N_1164);
nor U1238 (N_1238,N_1045,N_1118);
nor U1239 (N_1239,N_1188,N_934);
nor U1240 (N_1240,N_1166,N_1038);
or U1241 (N_1241,N_1050,N_1152);
and U1242 (N_1242,N_1147,N_1078);
and U1243 (N_1243,N_961,N_1149);
nand U1244 (N_1244,N_1180,N_969);
or U1245 (N_1245,N_1081,N_915);
or U1246 (N_1246,N_1145,N_1017);
nand U1247 (N_1247,N_1023,N_1048);
nor U1248 (N_1248,N_950,N_902);
xnor U1249 (N_1249,N_1080,N_1069);
nand U1250 (N_1250,N_1044,N_1102);
xnor U1251 (N_1251,N_920,N_1019);
nand U1252 (N_1252,N_907,N_1127);
xor U1253 (N_1253,N_1109,N_1028);
nor U1254 (N_1254,N_1036,N_1194);
and U1255 (N_1255,N_952,N_913);
or U1256 (N_1256,N_1096,N_1157);
nor U1257 (N_1257,N_1172,N_1099);
nor U1258 (N_1258,N_1010,N_1070);
nor U1259 (N_1259,N_1128,N_1001);
nor U1260 (N_1260,N_1129,N_1020);
nand U1261 (N_1261,N_1091,N_1189);
nand U1262 (N_1262,N_1022,N_1130);
nor U1263 (N_1263,N_1170,N_1186);
or U1264 (N_1264,N_1124,N_1126);
or U1265 (N_1265,N_997,N_1154);
and U1266 (N_1266,N_905,N_1179);
xnor U1267 (N_1267,N_1095,N_1140);
nor U1268 (N_1268,N_1008,N_1197);
and U1269 (N_1269,N_1047,N_1046);
or U1270 (N_1270,N_1011,N_1173);
nor U1271 (N_1271,N_1159,N_1162);
nor U1272 (N_1272,N_1033,N_1111);
and U1273 (N_1273,N_1191,N_966);
and U1274 (N_1274,N_939,N_937);
or U1275 (N_1275,N_1002,N_1059);
nand U1276 (N_1276,N_1086,N_1125);
nor U1277 (N_1277,N_994,N_1071);
and U1278 (N_1278,N_1037,N_1082);
nand U1279 (N_1279,N_1083,N_1087);
xor U1280 (N_1280,N_1151,N_978);
nor U1281 (N_1281,N_998,N_1135);
nor U1282 (N_1282,N_1163,N_941);
xor U1283 (N_1283,N_983,N_1195);
and U1284 (N_1284,N_954,N_953);
xnor U1285 (N_1285,N_1088,N_911);
xnor U1286 (N_1286,N_1156,N_1074);
nand U1287 (N_1287,N_944,N_1039);
nor U1288 (N_1288,N_1169,N_1075);
xnor U1289 (N_1289,N_1192,N_929);
nand U1290 (N_1290,N_1040,N_1107);
nand U1291 (N_1291,N_1072,N_1114);
xnor U1292 (N_1292,N_1133,N_951);
or U1293 (N_1293,N_1103,N_1073);
nand U1294 (N_1294,N_1123,N_1013);
or U1295 (N_1295,N_1112,N_1176);
nand U1296 (N_1296,N_993,N_1029);
nand U1297 (N_1297,N_1113,N_1077);
nor U1298 (N_1298,N_1079,N_1014);
xnor U1299 (N_1299,N_945,N_1108);
or U1300 (N_1300,N_1120,N_1084);
xor U1301 (N_1301,N_1155,N_1090);
and U1302 (N_1302,N_1064,N_1132);
nor U1303 (N_1303,N_1018,N_967);
and U1304 (N_1304,N_1056,N_1175);
and U1305 (N_1305,N_923,N_1148);
nand U1306 (N_1306,N_909,N_1167);
nand U1307 (N_1307,N_1177,N_1143);
nand U1308 (N_1308,N_1138,N_1003);
nand U1309 (N_1309,N_1025,N_1035);
nor U1310 (N_1310,N_1100,N_989);
nor U1311 (N_1311,N_903,N_1031);
or U1312 (N_1312,N_921,N_912);
nor U1313 (N_1313,N_996,N_1150);
xnor U1314 (N_1314,N_965,N_1005);
nor U1315 (N_1315,N_984,N_1182);
nor U1316 (N_1316,N_1034,N_1116);
nand U1317 (N_1317,N_1062,N_1153);
and U1318 (N_1318,N_1067,N_987);
xnor U1319 (N_1319,N_916,N_985);
xor U1320 (N_1320,N_970,N_943);
and U1321 (N_1321,N_1027,N_940);
and U1322 (N_1322,N_1146,N_1198);
and U1323 (N_1323,N_1142,N_1021);
or U1324 (N_1324,N_1139,N_974);
nand U1325 (N_1325,N_1006,N_904);
and U1326 (N_1326,N_1032,N_1012);
nor U1327 (N_1327,N_1165,N_1158);
or U1328 (N_1328,N_1104,N_1053);
nor U1329 (N_1329,N_958,N_930);
nand U1330 (N_1330,N_1051,N_1041);
nor U1331 (N_1331,N_908,N_1136);
nand U1332 (N_1332,N_1144,N_976);
or U1333 (N_1333,N_906,N_992);
nor U1334 (N_1334,N_1042,N_1106);
or U1335 (N_1335,N_1105,N_926);
nor U1336 (N_1336,N_1119,N_1085);
and U1337 (N_1337,N_1068,N_1066);
nor U1338 (N_1338,N_1141,N_975);
nor U1339 (N_1339,N_1043,N_982);
xor U1340 (N_1340,N_971,N_1196);
and U1341 (N_1341,N_963,N_947);
or U1342 (N_1342,N_1117,N_925);
nor U1343 (N_1343,N_1183,N_1193);
or U1344 (N_1344,N_1110,N_1115);
and U1345 (N_1345,N_1007,N_935);
nand U1346 (N_1346,N_946,N_1094);
nor U1347 (N_1347,N_1030,N_959);
or U1348 (N_1348,N_1134,N_1131);
xor U1349 (N_1349,N_927,N_1185);
nor U1350 (N_1350,N_1072,N_922);
nor U1351 (N_1351,N_1197,N_1172);
xor U1352 (N_1352,N_972,N_994);
nor U1353 (N_1353,N_1060,N_903);
or U1354 (N_1354,N_1043,N_1105);
nand U1355 (N_1355,N_937,N_999);
or U1356 (N_1356,N_1065,N_928);
or U1357 (N_1357,N_965,N_1135);
nand U1358 (N_1358,N_1191,N_967);
nor U1359 (N_1359,N_1107,N_994);
and U1360 (N_1360,N_927,N_976);
xnor U1361 (N_1361,N_988,N_1194);
or U1362 (N_1362,N_923,N_906);
nor U1363 (N_1363,N_990,N_1115);
nand U1364 (N_1364,N_1129,N_928);
nand U1365 (N_1365,N_926,N_1198);
xnor U1366 (N_1366,N_972,N_1100);
and U1367 (N_1367,N_1191,N_1111);
xnor U1368 (N_1368,N_1037,N_991);
or U1369 (N_1369,N_990,N_909);
nor U1370 (N_1370,N_1164,N_923);
and U1371 (N_1371,N_915,N_1096);
and U1372 (N_1372,N_935,N_1080);
or U1373 (N_1373,N_1170,N_950);
xnor U1374 (N_1374,N_1023,N_1015);
or U1375 (N_1375,N_942,N_904);
and U1376 (N_1376,N_1027,N_976);
nand U1377 (N_1377,N_1105,N_1131);
nor U1378 (N_1378,N_1145,N_1140);
or U1379 (N_1379,N_1162,N_1037);
xnor U1380 (N_1380,N_1009,N_1183);
or U1381 (N_1381,N_1022,N_974);
xnor U1382 (N_1382,N_955,N_1174);
xnor U1383 (N_1383,N_923,N_1018);
nor U1384 (N_1384,N_952,N_984);
nor U1385 (N_1385,N_1148,N_980);
nand U1386 (N_1386,N_1026,N_962);
or U1387 (N_1387,N_1187,N_918);
and U1388 (N_1388,N_1058,N_1106);
or U1389 (N_1389,N_970,N_1168);
and U1390 (N_1390,N_949,N_910);
nand U1391 (N_1391,N_1017,N_1125);
xnor U1392 (N_1392,N_1015,N_1003);
nand U1393 (N_1393,N_1021,N_949);
or U1394 (N_1394,N_1162,N_922);
or U1395 (N_1395,N_970,N_1014);
and U1396 (N_1396,N_1172,N_992);
or U1397 (N_1397,N_1005,N_1038);
nor U1398 (N_1398,N_1062,N_986);
xnor U1399 (N_1399,N_1035,N_1108);
xnor U1400 (N_1400,N_1025,N_902);
nor U1401 (N_1401,N_1082,N_1032);
nor U1402 (N_1402,N_1091,N_992);
nor U1403 (N_1403,N_998,N_1122);
xnor U1404 (N_1404,N_1008,N_1037);
and U1405 (N_1405,N_997,N_1065);
or U1406 (N_1406,N_913,N_1133);
xor U1407 (N_1407,N_932,N_1159);
nand U1408 (N_1408,N_932,N_1175);
nand U1409 (N_1409,N_1123,N_950);
nand U1410 (N_1410,N_1068,N_1105);
and U1411 (N_1411,N_1157,N_1070);
nand U1412 (N_1412,N_1185,N_1123);
nor U1413 (N_1413,N_1008,N_1108);
nor U1414 (N_1414,N_1102,N_1160);
xor U1415 (N_1415,N_1077,N_1105);
xor U1416 (N_1416,N_1048,N_925);
nor U1417 (N_1417,N_908,N_1077);
nand U1418 (N_1418,N_924,N_1034);
nor U1419 (N_1419,N_1115,N_1081);
xnor U1420 (N_1420,N_1190,N_1102);
nand U1421 (N_1421,N_900,N_966);
or U1422 (N_1422,N_1123,N_1120);
and U1423 (N_1423,N_1145,N_973);
nand U1424 (N_1424,N_1107,N_902);
nor U1425 (N_1425,N_993,N_1039);
and U1426 (N_1426,N_938,N_1071);
or U1427 (N_1427,N_1174,N_1199);
nand U1428 (N_1428,N_1103,N_1083);
xor U1429 (N_1429,N_902,N_1018);
or U1430 (N_1430,N_952,N_901);
nor U1431 (N_1431,N_929,N_1030);
or U1432 (N_1432,N_928,N_992);
and U1433 (N_1433,N_1094,N_1099);
and U1434 (N_1434,N_1048,N_1009);
or U1435 (N_1435,N_981,N_1166);
nor U1436 (N_1436,N_966,N_1174);
and U1437 (N_1437,N_917,N_1143);
or U1438 (N_1438,N_1019,N_1013);
nand U1439 (N_1439,N_1193,N_912);
or U1440 (N_1440,N_982,N_1092);
xnor U1441 (N_1441,N_1027,N_999);
and U1442 (N_1442,N_1144,N_930);
and U1443 (N_1443,N_1072,N_1066);
and U1444 (N_1444,N_1022,N_1048);
and U1445 (N_1445,N_1025,N_1028);
nor U1446 (N_1446,N_1032,N_1063);
or U1447 (N_1447,N_907,N_920);
or U1448 (N_1448,N_1083,N_966);
nor U1449 (N_1449,N_1016,N_952);
nor U1450 (N_1450,N_929,N_1069);
or U1451 (N_1451,N_913,N_992);
or U1452 (N_1452,N_1050,N_915);
and U1453 (N_1453,N_1139,N_1128);
and U1454 (N_1454,N_1009,N_1095);
xor U1455 (N_1455,N_1110,N_921);
nor U1456 (N_1456,N_1190,N_959);
xnor U1457 (N_1457,N_971,N_1016);
or U1458 (N_1458,N_923,N_1054);
nor U1459 (N_1459,N_947,N_950);
nor U1460 (N_1460,N_1063,N_965);
nand U1461 (N_1461,N_1191,N_1053);
nor U1462 (N_1462,N_1064,N_932);
xnor U1463 (N_1463,N_1006,N_999);
and U1464 (N_1464,N_1110,N_1059);
nor U1465 (N_1465,N_930,N_1068);
nor U1466 (N_1466,N_1109,N_1197);
or U1467 (N_1467,N_1179,N_1118);
xor U1468 (N_1468,N_947,N_1128);
or U1469 (N_1469,N_948,N_1055);
nor U1470 (N_1470,N_920,N_947);
xnor U1471 (N_1471,N_901,N_1099);
and U1472 (N_1472,N_1058,N_1182);
nor U1473 (N_1473,N_1043,N_1024);
and U1474 (N_1474,N_973,N_1020);
or U1475 (N_1475,N_929,N_1120);
nand U1476 (N_1476,N_1145,N_1171);
nor U1477 (N_1477,N_1185,N_964);
nand U1478 (N_1478,N_943,N_1114);
nor U1479 (N_1479,N_915,N_1173);
nand U1480 (N_1480,N_1175,N_1183);
xnor U1481 (N_1481,N_914,N_1087);
nor U1482 (N_1482,N_1032,N_997);
nand U1483 (N_1483,N_1170,N_1158);
or U1484 (N_1484,N_919,N_967);
nor U1485 (N_1485,N_1135,N_1133);
xor U1486 (N_1486,N_998,N_1048);
nor U1487 (N_1487,N_1095,N_907);
nand U1488 (N_1488,N_1156,N_1126);
nor U1489 (N_1489,N_1019,N_1003);
and U1490 (N_1490,N_919,N_1120);
nor U1491 (N_1491,N_972,N_1056);
xnor U1492 (N_1492,N_1054,N_1196);
nor U1493 (N_1493,N_968,N_1134);
and U1494 (N_1494,N_977,N_1139);
nand U1495 (N_1495,N_1028,N_975);
xnor U1496 (N_1496,N_1042,N_996);
nor U1497 (N_1497,N_1136,N_1140);
xor U1498 (N_1498,N_951,N_1151);
and U1499 (N_1499,N_932,N_907);
nand U1500 (N_1500,N_1207,N_1331);
and U1501 (N_1501,N_1368,N_1301);
or U1502 (N_1502,N_1235,N_1415);
nor U1503 (N_1503,N_1426,N_1459);
nor U1504 (N_1504,N_1396,N_1239);
and U1505 (N_1505,N_1366,N_1454);
nand U1506 (N_1506,N_1431,N_1326);
nor U1507 (N_1507,N_1261,N_1482);
nand U1508 (N_1508,N_1441,N_1248);
xor U1509 (N_1509,N_1494,N_1412);
nor U1510 (N_1510,N_1478,N_1462);
or U1511 (N_1511,N_1325,N_1357);
xor U1512 (N_1512,N_1234,N_1211);
nor U1513 (N_1513,N_1479,N_1440);
or U1514 (N_1514,N_1379,N_1255);
and U1515 (N_1515,N_1270,N_1318);
nor U1516 (N_1516,N_1260,N_1215);
xor U1517 (N_1517,N_1269,N_1477);
or U1518 (N_1518,N_1423,N_1250);
or U1519 (N_1519,N_1443,N_1252);
xor U1520 (N_1520,N_1303,N_1485);
nand U1521 (N_1521,N_1306,N_1391);
nand U1522 (N_1522,N_1382,N_1469);
and U1523 (N_1523,N_1259,N_1218);
nand U1524 (N_1524,N_1253,N_1434);
nor U1525 (N_1525,N_1344,N_1458);
or U1526 (N_1526,N_1292,N_1319);
xnor U1527 (N_1527,N_1332,N_1435);
xor U1528 (N_1528,N_1275,N_1204);
nor U1529 (N_1529,N_1402,N_1237);
xnor U1530 (N_1530,N_1463,N_1293);
nor U1531 (N_1531,N_1413,N_1465);
xnor U1532 (N_1532,N_1442,N_1499);
nand U1533 (N_1533,N_1311,N_1496);
or U1534 (N_1534,N_1475,N_1315);
and U1535 (N_1535,N_1381,N_1279);
and U1536 (N_1536,N_1480,N_1405);
nand U1537 (N_1537,N_1324,N_1380);
or U1538 (N_1538,N_1450,N_1421);
nand U1539 (N_1539,N_1305,N_1358);
or U1540 (N_1540,N_1445,N_1340);
nor U1541 (N_1541,N_1376,N_1350);
nor U1542 (N_1542,N_1457,N_1466);
xnor U1543 (N_1543,N_1205,N_1460);
and U1544 (N_1544,N_1386,N_1302);
xnor U1545 (N_1545,N_1409,N_1287);
and U1546 (N_1546,N_1476,N_1369);
and U1547 (N_1547,N_1309,N_1233);
nand U1548 (N_1548,N_1456,N_1313);
xor U1549 (N_1549,N_1359,N_1438);
nor U1550 (N_1550,N_1263,N_1256);
xnor U1551 (N_1551,N_1401,N_1323);
xnor U1552 (N_1552,N_1246,N_1224);
nor U1553 (N_1553,N_1300,N_1492);
or U1554 (N_1554,N_1419,N_1467);
nand U1555 (N_1555,N_1371,N_1484);
and U1556 (N_1556,N_1243,N_1449);
or U1557 (N_1557,N_1493,N_1210);
nor U1558 (N_1558,N_1343,N_1422);
nand U1559 (N_1559,N_1404,N_1247);
nor U1560 (N_1560,N_1451,N_1372);
or U1561 (N_1561,N_1498,N_1427);
or U1562 (N_1562,N_1251,N_1214);
and U1563 (N_1563,N_1348,N_1294);
nand U1564 (N_1564,N_1437,N_1221);
or U1565 (N_1565,N_1228,N_1274);
nor U1566 (N_1566,N_1406,N_1212);
nand U1567 (N_1567,N_1220,N_1314);
or U1568 (N_1568,N_1238,N_1276);
nor U1569 (N_1569,N_1489,N_1297);
nand U1570 (N_1570,N_1241,N_1227);
or U1571 (N_1571,N_1452,N_1461);
xnor U1572 (N_1572,N_1266,N_1487);
or U1573 (N_1573,N_1341,N_1429);
and U1574 (N_1574,N_1353,N_1361);
xor U1575 (N_1575,N_1201,N_1219);
and U1576 (N_1576,N_1362,N_1295);
or U1577 (N_1577,N_1455,N_1225);
nand U1578 (N_1578,N_1417,N_1439);
nor U1579 (N_1579,N_1351,N_1310);
and U1580 (N_1580,N_1268,N_1448);
xor U1581 (N_1581,N_1283,N_1328);
xnor U1582 (N_1582,N_1453,N_1290);
xnor U1583 (N_1583,N_1394,N_1335);
nand U1584 (N_1584,N_1262,N_1345);
nand U1585 (N_1585,N_1392,N_1307);
and U1586 (N_1586,N_1285,N_1231);
xor U1587 (N_1587,N_1329,N_1216);
and U1588 (N_1588,N_1308,N_1399);
and U1589 (N_1589,N_1444,N_1245);
and U1590 (N_1590,N_1375,N_1286);
or U1591 (N_1591,N_1258,N_1471);
or U1592 (N_1592,N_1390,N_1490);
nor U1593 (N_1593,N_1349,N_1223);
and U1594 (N_1594,N_1240,N_1356);
nand U1595 (N_1595,N_1430,N_1271);
nor U1596 (N_1596,N_1355,N_1424);
or U1597 (N_1597,N_1472,N_1398);
nor U1598 (N_1598,N_1208,N_1254);
nor U1599 (N_1599,N_1363,N_1447);
and U1600 (N_1600,N_1229,N_1374);
nand U1601 (N_1601,N_1364,N_1433);
xnor U1602 (N_1602,N_1410,N_1277);
or U1603 (N_1603,N_1473,N_1354);
xor U1604 (N_1604,N_1385,N_1408);
nor U1605 (N_1605,N_1436,N_1342);
nor U1606 (N_1606,N_1428,N_1336);
xnor U1607 (N_1607,N_1296,N_1464);
and U1608 (N_1608,N_1373,N_1418);
or U1609 (N_1609,N_1497,N_1333);
xnor U1610 (N_1610,N_1367,N_1388);
and U1611 (N_1611,N_1378,N_1304);
or U1612 (N_1612,N_1339,N_1491);
or U1613 (N_1613,N_1312,N_1317);
xnor U1614 (N_1614,N_1299,N_1327);
and U1615 (N_1615,N_1416,N_1316);
or U1616 (N_1616,N_1347,N_1232);
and U1617 (N_1617,N_1384,N_1206);
and U1618 (N_1618,N_1244,N_1273);
xor U1619 (N_1619,N_1346,N_1264);
xnor U1620 (N_1620,N_1414,N_1202);
or U1621 (N_1621,N_1281,N_1334);
nand U1622 (N_1622,N_1383,N_1200);
or U1623 (N_1623,N_1322,N_1257);
nand U1624 (N_1624,N_1289,N_1272);
or U1625 (N_1625,N_1395,N_1265);
or U1626 (N_1626,N_1403,N_1468);
or U1627 (N_1627,N_1470,N_1242);
nand U1628 (N_1628,N_1360,N_1446);
nor U1629 (N_1629,N_1222,N_1213);
and U1630 (N_1630,N_1203,N_1236);
nand U1631 (N_1631,N_1209,N_1411);
or U1632 (N_1632,N_1280,N_1284);
xnor U1633 (N_1633,N_1320,N_1337);
xnor U1634 (N_1634,N_1267,N_1249);
xnor U1635 (N_1635,N_1338,N_1278);
or U1636 (N_1636,N_1226,N_1377);
nor U1637 (N_1637,N_1365,N_1425);
and U1638 (N_1638,N_1330,N_1420);
nor U1639 (N_1639,N_1481,N_1389);
xor U1640 (N_1640,N_1488,N_1387);
and U1641 (N_1641,N_1486,N_1291);
xnor U1642 (N_1642,N_1298,N_1400);
nor U1643 (N_1643,N_1288,N_1474);
or U1644 (N_1644,N_1483,N_1495);
or U1645 (N_1645,N_1282,N_1407);
xnor U1646 (N_1646,N_1352,N_1230);
nor U1647 (N_1647,N_1393,N_1370);
nor U1648 (N_1648,N_1432,N_1217);
xnor U1649 (N_1649,N_1321,N_1397);
xor U1650 (N_1650,N_1244,N_1298);
and U1651 (N_1651,N_1389,N_1282);
xnor U1652 (N_1652,N_1242,N_1386);
and U1653 (N_1653,N_1228,N_1276);
and U1654 (N_1654,N_1321,N_1204);
xnor U1655 (N_1655,N_1365,N_1318);
or U1656 (N_1656,N_1207,N_1405);
and U1657 (N_1657,N_1445,N_1416);
and U1658 (N_1658,N_1277,N_1268);
or U1659 (N_1659,N_1219,N_1225);
xnor U1660 (N_1660,N_1497,N_1408);
xnor U1661 (N_1661,N_1296,N_1387);
or U1662 (N_1662,N_1308,N_1220);
nor U1663 (N_1663,N_1484,N_1335);
nor U1664 (N_1664,N_1313,N_1202);
or U1665 (N_1665,N_1466,N_1336);
and U1666 (N_1666,N_1495,N_1300);
or U1667 (N_1667,N_1480,N_1489);
or U1668 (N_1668,N_1339,N_1348);
and U1669 (N_1669,N_1329,N_1315);
or U1670 (N_1670,N_1451,N_1473);
xnor U1671 (N_1671,N_1208,N_1226);
nand U1672 (N_1672,N_1265,N_1259);
nor U1673 (N_1673,N_1413,N_1341);
xnor U1674 (N_1674,N_1335,N_1220);
xnor U1675 (N_1675,N_1213,N_1492);
nand U1676 (N_1676,N_1260,N_1406);
and U1677 (N_1677,N_1327,N_1464);
xnor U1678 (N_1678,N_1330,N_1492);
nand U1679 (N_1679,N_1236,N_1371);
xor U1680 (N_1680,N_1327,N_1417);
nand U1681 (N_1681,N_1229,N_1235);
and U1682 (N_1682,N_1262,N_1289);
and U1683 (N_1683,N_1326,N_1271);
nand U1684 (N_1684,N_1348,N_1247);
and U1685 (N_1685,N_1473,N_1327);
xnor U1686 (N_1686,N_1463,N_1425);
and U1687 (N_1687,N_1225,N_1272);
nand U1688 (N_1688,N_1249,N_1403);
xor U1689 (N_1689,N_1200,N_1206);
and U1690 (N_1690,N_1261,N_1393);
nor U1691 (N_1691,N_1218,N_1240);
nor U1692 (N_1692,N_1478,N_1473);
or U1693 (N_1693,N_1242,N_1373);
or U1694 (N_1694,N_1205,N_1226);
and U1695 (N_1695,N_1342,N_1330);
nand U1696 (N_1696,N_1343,N_1277);
nand U1697 (N_1697,N_1233,N_1319);
or U1698 (N_1698,N_1463,N_1287);
and U1699 (N_1699,N_1409,N_1487);
xor U1700 (N_1700,N_1429,N_1496);
xnor U1701 (N_1701,N_1387,N_1294);
and U1702 (N_1702,N_1302,N_1467);
or U1703 (N_1703,N_1343,N_1374);
and U1704 (N_1704,N_1499,N_1371);
and U1705 (N_1705,N_1294,N_1449);
nand U1706 (N_1706,N_1468,N_1431);
xor U1707 (N_1707,N_1384,N_1368);
or U1708 (N_1708,N_1335,N_1204);
and U1709 (N_1709,N_1274,N_1395);
or U1710 (N_1710,N_1494,N_1308);
and U1711 (N_1711,N_1393,N_1330);
xnor U1712 (N_1712,N_1242,N_1253);
and U1713 (N_1713,N_1338,N_1335);
and U1714 (N_1714,N_1460,N_1438);
nand U1715 (N_1715,N_1355,N_1365);
and U1716 (N_1716,N_1397,N_1334);
nand U1717 (N_1717,N_1252,N_1476);
and U1718 (N_1718,N_1334,N_1277);
nor U1719 (N_1719,N_1464,N_1417);
nor U1720 (N_1720,N_1297,N_1426);
nand U1721 (N_1721,N_1317,N_1347);
xor U1722 (N_1722,N_1485,N_1451);
nor U1723 (N_1723,N_1219,N_1388);
and U1724 (N_1724,N_1263,N_1408);
nand U1725 (N_1725,N_1246,N_1223);
nand U1726 (N_1726,N_1253,N_1453);
xnor U1727 (N_1727,N_1239,N_1498);
and U1728 (N_1728,N_1320,N_1298);
xor U1729 (N_1729,N_1319,N_1439);
nand U1730 (N_1730,N_1235,N_1342);
xnor U1731 (N_1731,N_1260,N_1310);
nor U1732 (N_1732,N_1298,N_1227);
nand U1733 (N_1733,N_1303,N_1468);
nand U1734 (N_1734,N_1365,N_1286);
or U1735 (N_1735,N_1266,N_1373);
and U1736 (N_1736,N_1381,N_1219);
xor U1737 (N_1737,N_1255,N_1309);
or U1738 (N_1738,N_1443,N_1303);
xor U1739 (N_1739,N_1388,N_1364);
and U1740 (N_1740,N_1219,N_1394);
xnor U1741 (N_1741,N_1357,N_1300);
or U1742 (N_1742,N_1207,N_1385);
or U1743 (N_1743,N_1370,N_1205);
nor U1744 (N_1744,N_1372,N_1298);
nand U1745 (N_1745,N_1205,N_1473);
xor U1746 (N_1746,N_1243,N_1223);
xnor U1747 (N_1747,N_1293,N_1333);
and U1748 (N_1748,N_1374,N_1288);
or U1749 (N_1749,N_1317,N_1429);
nor U1750 (N_1750,N_1452,N_1251);
or U1751 (N_1751,N_1254,N_1412);
or U1752 (N_1752,N_1447,N_1401);
nor U1753 (N_1753,N_1256,N_1473);
or U1754 (N_1754,N_1431,N_1456);
nor U1755 (N_1755,N_1320,N_1465);
and U1756 (N_1756,N_1319,N_1446);
nor U1757 (N_1757,N_1256,N_1395);
nand U1758 (N_1758,N_1451,N_1336);
nor U1759 (N_1759,N_1433,N_1269);
and U1760 (N_1760,N_1404,N_1430);
xnor U1761 (N_1761,N_1326,N_1439);
and U1762 (N_1762,N_1406,N_1417);
and U1763 (N_1763,N_1266,N_1349);
nor U1764 (N_1764,N_1310,N_1469);
xnor U1765 (N_1765,N_1374,N_1221);
nor U1766 (N_1766,N_1251,N_1474);
and U1767 (N_1767,N_1260,N_1255);
or U1768 (N_1768,N_1281,N_1263);
or U1769 (N_1769,N_1396,N_1473);
or U1770 (N_1770,N_1431,N_1297);
nand U1771 (N_1771,N_1351,N_1336);
xor U1772 (N_1772,N_1347,N_1250);
xor U1773 (N_1773,N_1383,N_1217);
nand U1774 (N_1774,N_1484,N_1416);
nor U1775 (N_1775,N_1371,N_1349);
xor U1776 (N_1776,N_1444,N_1496);
and U1777 (N_1777,N_1463,N_1222);
xnor U1778 (N_1778,N_1382,N_1454);
xor U1779 (N_1779,N_1266,N_1375);
nor U1780 (N_1780,N_1387,N_1215);
nand U1781 (N_1781,N_1367,N_1305);
and U1782 (N_1782,N_1455,N_1391);
nand U1783 (N_1783,N_1364,N_1322);
nor U1784 (N_1784,N_1245,N_1379);
nor U1785 (N_1785,N_1344,N_1473);
nand U1786 (N_1786,N_1353,N_1448);
or U1787 (N_1787,N_1430,N_1388);
or U1788 (N_1788,N_1338,N_1442);
nor U1789 (N_1789,N_1466,N_1352);
or U1790 (N_1790,N_1233,N_1406);
and U1791 (N_1791,N_1455,N_1245);
nor U1792 (N_1792,N_1393,N_1433);
and U1793 (N_1793,N_1411,N_1210);
nor U1794 (N_1794,N_1359,N_1320);
nand U1795 (N_1795,N_1378,N_1412);
nor U1796 (N_1796,N_1381,N_1252);
or U1797 (N_1797,N_1277,N_1204);
nand U1798 (N_1798,N_1351,N_1340);
or U1799 (N_1799,N_1385,N_1233);
nor U1800 (N_1800,N_1607,N_1794);
xnor U1801 (N_1801,N_1687,N_1769);
xnor U1802 (N_1802,N_1770,N_1563);
nand U1803 (N_1803,N_1795,N_1616);
xnor U1804 (N_1804,N_1638,N_1599);
and U1805 (N_1805,N_1705,N_1504);
and U1806 (N_1806,N_1623,N_1682);
nand U1807 (N_1807,N_1503,N_1606);
nor U1808 (N_1808,N_1571,N_1768);
nor U1809 (N_1809,N_1653,N_1772);
nor U1810 (N_1810,N_1570,N_1520);
xnor U1811 (N_1811,N_1610,N_1539);
xor U1812 (N_1812,N_1509,N_1629);
nand U1813 (N_1813,N_1760,N_1654);
nand U1814 (N_1814,N_1630,N_1625);
or U1815 (N_1815,N_1685,N_1664);
and U1816 (N_1816,N_1510,N_1666);
or U1817 (N_1817,N_1578,N_1559);
nor U1818 (N_1818,N_1688,N_1678);
and U1819 (N_1819,N_1528,N_1542);
or U1820 (N_1820,N_1798,N_1581);
nor U1821 (N_1821,N_1576,N_1555);
xnor U1822 (N_1822,N_1675,N_1604);
and U1823 (N_1823,N_1518,N_1639);
nor U1824 (N_1824,N_1649,N_1776);
nor U1825 (N_1825,N_1501,N_1573);
and U1826 (N_1826,N_1697,N_1751);
nor U1827 (N_1827,N_1673,N_1535);
or U1828 (N_1828,N_1667,N_1575);
and U1829 (N_1829,N_1620,N_1763);
nor U1830 (N_1830,N_1766,N_1741);
xnor U1831 (N_1831,N_1712,N_1618);
xnor U1832 (N_1832,N_1747,N_1686);
nor U1833 (N_1833,N_1611,N_1782);
nor U1834 (N_1834,N_1758,N_1695);
and U1835 (N_1835,N_1786,N_1718);
and U1836 (N_1836,N_1566,N_1700);
xor U1837 (N_1837,N_1554,N_1734);
and U1838 (N_1838,N_1561,N_1597);
xor U1839 (N_1839,N_1680,N_1586);
and U1840 (N_1840,N_1543,N_1600);
nand U1841 (N_1841,N_1753,N_1544);
nand U1842 (N_1842,N_1784,N_1761);
or U1843 (N_1843,N_1722,N_1515);
nor U1844 (N_1844,N_1721,N_1635);
xnor U1845 (N_1845,N_1689,N_1529);
nor U1846 (N_1846,N_1752,N_1565);
nand U1847 (N_1847,N_1725,N_1694);
nand U1848 (N_1848,N_1548,N_1762);
and U1849 (N_1849,N_1550,N_1779);
or U1850 (N_1850,N_1632,N_1726);
and U1851 (N_1851,N_1661,N_1790);
nor U1852 (N_1852,N_1523,N_1711);
nor U1853 (N_1853,N_1531,N_1552);
or U1854 (N_1854,N_1742,N_1693);
nand U1855 (N_1855,N_1538,N_1647);
nand U1856 (N_1856,N_1502,N_1643);
xor U1857 (N_1857,N_1709,N_1743);
nor U1858 (N_1858,N_1698,N_1557);
nand U1859 (N_1859,N_1677,N_1720);
xnor U1860 (N_1860,N_1792,N_1773);
and U1861 (N_1861,N_1797,N_1780);
or U1862 (N_1862,N_1546,N_1777);
or U1863 (N_1863,N_1793,N_1671);
or U1864 (N_1864,N_1642,N_1602);
nor U1865 (N_1865,N_1572,N_1737);
and U1866 (N_1866,N_1749,N_1641);
or U1867 (N_1867,N_1651,N_1748);
and U1868 (N_1868,N_1615,N_1534);
xnor U1869 (N_1869,N_1624,N_1696);
nor U1870 (N_1870,N_1704,N_1580);
nor U1871 (N_1871,N_1530,N_1622);
or U1872 (N_1872,N_1701,N_1540);
or U1873 (N_1873,N_1662,N_1567);
xnor U1874 (N_1874,N_1676,N_1799);
and U1875 (N_1875,N_1719,N_1739);
and U1876 (N_1876,N_1755,N_1791);
nand U1877 (N_1877,N_1582,N_1738);
nor U1878 (N_1878,N_1516,N_1603);
xor U1879 (N_1879,N_1584,N_1583);
xor U1880 (N_1880,N_1723,N_1590);
or U1881 (N_1881,N_1560,N_1558);
nor U1882 (N_1882,N_1706,N_1591);
nor U1883 (N_1883,N_1507,N_1536);
nand U1884 (N_1884,N_1553,N_1512);
or U1885 (N_1885,N_1506,N_1759);
and U1886 (N_1886,N_1577,N_1729);
nand U1887 (N_1887,N_1733,N_1521);
and U1888 (N_1888,N_1505,N_1633);
nand U1889 (N_1889,N_1674,N_1598);
xnor U1890 (N_1890,N_1796,N_1594);
or U1891 (N_1891,N_1650,N_1707);
and U1892 (N_1892,N_1774,N_1670);
and U1893 (N_1893,N_1541,N_1735);
nand U1894 (N_1894,N_1728,N_1549);
or U1895 (N_1895,N_1640,N_1508);
nor U1896 (N_1896,N_1778,N_1621);
nand U1897 (N_1897,N_1568,N_1692);
nor U1898 (N_1898,N_1595,N_1781);
xor U1899 (N_1899,N_1659,N_1646);
and U1900 (N_1900,N_1765,N_1787);
nand U1901 (N_1901,N_1665,N_1519);
nand U1902 (N_1902,N_1522,N_1757);
nor U1903 (N_1903,N_1613,N_1783);
nand U1904 (N_1904,N_1690,N_1703);
nor U1905 (N_1905,N_1652,N_1710);
nand U1906 (N_1906,N_1744,N_1589);
and U1907 (N_1907,N_1672,N_1525);
xnor U1908 (N_1908,N_1785,N_1513);
nor U1909 (N_1909,N_1526,N_1663);
xor U1910 (N_1910,N_1545,N_1699);
or U1911 (N_1911,N_1619,N_1569);
nand U1912 (N_1912,N_1756,N_1631);
and U1913 (N_1913,N_1724,N_1562);
xor U1914 (N_1914,N_1681,N_1617);
nand U1915 (N_1915,N_1551,N_1679);
nor U1916 (N_1916,N_1746,N_1547);
and U1917 (N_1917,N_1736,N_1740);
or U1918 (N_1918,N_1533,N_1585);
nand U1919 (N_1919,N_1669,N_1636);
nor U1920 (N_1920,N_1702,N_1648);
xor U1921 (N_1921,N_1532,N_1609);
or U1922 (N_1922,N_1574,N_1750);
xnor U1923 (N_1923,N_1788,N_1655);
nand U1924 (N_1924,N_1668,N_1658);
or U1925 (N_1925,N_1691,N_1731);
nand U1926 (N_1926,N_1601,N_1716);
nor U1927 (N_1927,N_1564,N_1517);
nor U1928 (N_1928,N_1714,N_1789);
or U1929 (N_1929,N_1634,N_1645);
and U1930 (N_1930,N_1713,N_1596);
nand U1931 (N_1931,N_1579,N_1657);
nor U1932 (N_1932,N_1592,N_1684);
xor U1933 (N_1933,N_1527,N_1605);
xnor U1934 (N_1934,N_1745,N_1514);
or U1935 (N_1935,N_1587,N_1732);
nand U1936 (N_1936,N_1608,N_1644);
or U1937 (N_1937,N_1771,N_1754);
or U1938 (N_1938,N_1727,N_1637);
nor U1939 (N_1939,N_1717,N_1524);
nand U1940 (N_1940,N_1730,N_1593);
xnor U1941 (N_1941,N_1660,N_1556);
nor U1942 (N_1942,N_1626,N_1500);
xor U1943 (N_1943,N_1656,N_1767);
nor U1944 (N_1944,N_1764,N_1511);
nand U1945 (N_1945,N_1627,N_1775);
xnor U1946 (N_1946,N_1537,N_1683);
and U1947 (N_1947,N_1588,N_1628);
nor U1948 (N_1948,N_1612,N_1715);
nand U1949 (N_1949,N_1708,N_1614);
nor U1950 (N_1950,N_1768,N_1747);
or U1951 (N_1951,N_1647,N_1586);
nor U1952 (N_1952,N_1602,N_1623);
nor U1953 (N_1953,N_1566,N_1734);
nand U1954 (N_1954,N_1586,N_1600);
nor U1955 (N_1955,N_1741,N_1714);
xor U1956 (N_1956,N_1737,N_1516);
nor U1957 (N_1957,N_1640,N_1765);
or U1958 (N_1958,N_1762,N_1566);
or U1959 (N_1959,N_1506,N_1653);
nand U1960 (N_1960,N_1764,N_1701);
or U1961 (N_1961,N_1635,N_1777);
and U1962 (N_1962,N_1644,N_1661);
nor U1963 (N_1963,N_1727,N_1768);
nand U1964 (N_1964,N_1780,N_1676);
nor U1965 (N_1965,N_1730,N_1567);
or U1966 (N_1966,N_1627,N_1770);
and U1967 (N_1967,N_1644,N_1797);
xnor U1968 (N_1968,N_1729,N_1734);
nand U1969 (N_1969,N_1546,N_1623);
or U1970 (N_1970,N_1623,N_1663);
or U1971 (N_1971,N_1667,N_1624);
and U1972 (N_1972,N_1604,N_1729);
nand U1973 (N_1973,N_1540,N_1768);
and U1974 (N_1974,N_1721,N_1707);
or U1975 (N_1975,N_1585,N_1502);
nand U1976 (N_1976,N_1647,N_1548);
nor U1977 (N_1977,N_1606,N_1698);
xnor U1978 (N_1978,N_1551,N_1666);
or U1979 (N_1979,N_1699,N_1509);
or U1980 (N_1980,N_1650,N_1779);
nor U1981 (N_1981,N_1756,N_1512);
or U1982 (N_1982,N_1702,N_1518);
xnor U1983 (N_1983,N_1538,N_1509);
xor U1984 (N_1984,N_1696,N_1582);
xor U1985 (N_1985,N_1742,N_1600);
nand U1986 (N_1986,N_1531,N_1795);
and U1987 (N_1987,N_1662,N_1523);
nand U1988 (N_1988,N_1662,N_1514);
or U1989 (N_1989,N_1597,N_1675);
nor U1990 (N_1990,N_1567,N_1559);
or U1991 (N_1991,N_1519,N_1635);
nor U1992 (N_1992,N_1600,N_1566);
nand U1993 (N_1993,N_1666,N_1583);
nand U1994 (N_1994,N_1715,N_1704);
nor U1995 (N_1995,N_1737,N_1547);
and U1996 (N_1996,N_1527,N_1603);
and U1997 (N_1997,N_1763,N_1726);
and U1998 (N_1998,N_1616,N_1703);
nand U1999 (N_1999,N_1562,N_1504);
or U2000 (N_2000,N_1539,N_1758);
and U2001 (N_2001,N_1717,N_1669);
nor U2002 (N_2002,N_1640,N_1686);
nand U2003 (N_2003,N_1770,N_1737);
xor U2004 (N_2004,N_1627,N_1596);
nor U2005 (N_2005,N_1716,N_1541);
and U2006 (N_2006,N_1629,N_1575);
nor U2007 (N_2007,N_1649,N_1555);
or U2008 (N_2008,N_1602,N_1505);
nor U2009 (N_2009,N_1630,N_1687);
or U2010 (N_2010,N_1759,N_1572);
xor U2011 (N_2011,N_1678,N_1779);
or U2012 (N_2012,N_1545,N_1593);
nor U2013 (N_2013,N_1627,N_1657);
or U2014 (N_2014,N_1583,N_1509);
or U2015 (N_2015,N_1536,N_1609);
nand U2016 (N_2016,N_1651,N_1798);
nand U2017 (N_2017,N_1576,N_1727);
nor U2018 (N_2018,N_1725,N_1708);
xor U2019 (N_2019,N_1594,N_1652);
nand U2020 (N_2020,N_1623,N_1592);
nand U2021 (N_2021,N_1565,N_1660);
xor U2022 (N_2022,N_1657,N_1753);
or U2023 (N_2023,N_1727,N_1742);
nand U2024 (N_2024,N_1511,N_1651);
and U2025 (N_2025,N_1769,N_1614);
or U2026 (N_2026,N_1782,N_1724);
nand U2027 (N_2027,N_1587,N_1540);
nand U2028 (N_2028,N_1756,N_1548);
nand U2029 (N_2029,N_1744,N_1576);
xor U2030 (N_2030,N_1588,N_1795);
or U2031 (N_2031,N_1672,N_1615);
nand U2032 (N_2032,N_1706,N_1662);
and U2033 (N_2033,N_1635,N_1580);
nor U2034 (N_2034,N_1625,N_1799);
and U2035 (N_2035,N_1732,N_1754);
nor U2036 (N_2036,N_1708,N_1662);
nand U2037 (N_2037,N_1758,N_1626);
and U2038 (N_2038,N_1637,N_1513);
or U2039 (N_2039,N_1709,N_1650);
or U2040 (N_2040,N_1583,N_1773);
or U2041 (N_2041,N_1526,N_1508);
and U2042 (N_2042,N_1562,N_1755);
nor U2043 (N_2043,N_1738,N_1642);
nand U2044 (N_2044,N_1674,N_1517);
nor U2045 (N_2045,N_1792,N_1515);
or U2046 (N_2046,N_1611,N_1771);
nor U2047 (N_2047,N_1763,N_1581);
nand U2048 (N_2048,N_1779,N_1581);
nor U2049 (N_2049,N_1575,N_1541);
and U2050 (N_2050,N_1591,N_1791);
xnor U2051 (N_2051,N_1539,N_1770);
nor U2052 (N_2052,N_1737,N_1553);
nand U2053 (N_2053,N_1792,N_1536);
or U2054 (N_2054,N_1735,N_1781);
nor U2055 (N_2055,N_1688,N_1684);
xnor U2056 (N_2056,N_1646,N_1738);
xor U2057 (N_2057,N_1539,N_1561);
or U2058 (N_2058,N_1661,N_1747);
xor U2059 (N_2059,N_1798,N_1712);
or U2060 (N_2060,N_1784,N_1529);
and U2061 (N_2061,N_1725,N_1686);
nor U2062 (N_2062,N_1688,N_1529);
xor U2063 (N_2063,N_1676,N_1683);
nor U2064 (N_2064,N_1790,N_1684);
and U2065 (N_2065,N_1596,N_1520);
nand U2066 (N_2066,N_1634,N_1642);
and U2067 (N_2067,N_1579,N_1510);
xor U2068 (N_2068,N_1571,N_1548);
or U2069 (N_2069,N_1668,N_1681);
nor U2070 (N_2070,N_1668,N_1787);
xnor U2071 (N_2071,N_1682,N_1586);
or U2072 (N_2072,N_1778,N_1723);
nor U2073 (N_2073,N_1792,N_1753);
and U2074 (N_2074,N_1617,N_1638);
xnor U2075 (N_2075,N_1514,N_1597);
nor U2076 (N_2076,N_1784,N_1562);
nor U2077 (N_2077,N_1525,N_1517);
xnor U2078 (N_2078,N_1706,N_1765);
or U2079 (N_2079,N_1799,N_1744);
xnor U2080 (N_2080,N_1750,N_1731);
xnor U2081 (N_2081,N_1585,N_1598);
and U2082 (N_2082,N_1785,N_1742);
and U2083 (N_2083,N_1533,N_1719);
and U2084 (N_2084,N_1526,N_1748);
nand U2085 (N_2085,N_1775,N_1535);
and U2086 (N_2086,N_1790,N_1698);
nor U2087 (N_2087,N_1527,N_1622);
xnor U2088 (N_2088,N_1565,N_1767);
and U2089 (N_2089,N_1635,N_1641);
or U2090 (N_2090,N_1582,N_1508);
and U2091 (N_2091,N_1576,N_1782);
xor U2092 (N_2092,N_1555,N_1776);
xnor U2093 (N_2093,N_1682,N_1772);
xnor U2094 (N_2094,N_1721,N_1527);
xor U2095 (N_2095,N_1567,N_1725);
nand U2096 (N_2096,N_1769,N_1701);
nand U2097 (N_2097,N_1528,N_1772);
xor U2098 (N_2098,N_1620,N_1616);
xor U2099 (N_2099,N_1618,N_1673);
xnor U2100 (N_2100,N_1889,N_1909);
and U2101 (N_2101,N_1928,N_2052);
nor U2102 (N_2102,N_2033,N_1978);
nand U2103 (N_2103,N_2086,N_1929);
nor U2104 (N_2104,N_1869,N_2001);
nand U2105 (N_2105,N_1985,N_2094);
nor U2106 (N_2106,N_1936,N_1916);
xnor U2107 (N_2107,N_1847,N_2020);
or U2108 (N_2108,N_1894,N_1850);
and U2109 (N_2109,N_1980,N_2006);
xnor U2110 (N_2110,N_2024,N_1812);
and U2111 (N_2111,N_1808,N_1924);
xnor U2112 (N_2112,N_1870,N_1991);
nor U2113 (N_2113,N_1998,N_2064);
xor U2114 (N_2114,N_1961,N_2012);
nor U2115 (N_2115,N_2059,N_2055);
xor U2116 (N_2116,N_2084,N_1873);
or U2117 (N_2117,N_2078,N_2021);
nor U2118 (N_2118,N_1811,N_1988);
and U2119 (N_2119,N_1885,N_1835);
or U2120 (N_2120,N_1856,N_2060);
xor U2121 (N_2121,N_2007,N_1815);
and U2122 (N_2122,N_1953,N_1992);
or U2123 (N_2123,N_2058,N_1891);
xnor U2124 (N_2124,N_2071,N_1802);
nor U2125 (N_2125,N_2005,N_1933);
and U2126 (N_2126,N_1945,N_1838);
nand U2127 (N_2127,N_1878,N_1901);
or U2128 (N_2128,N_1841,N_1881);
xnor U2129 (N_2129,N_2062,N_1923);
xor U2130 (N_2130,N_1912,N_1834);
and U2131 (N_2131,N_2053,N_1984);
and U2132 (N_2132,N_1962,N_1903);
nand U2133 (N_2133,N_2054,N_2010);
or U2134 (N_2134,N_2034,N_1810);
or U2135 (N_2135,N_2087,N_1860);
nand U2136 (N_2136,N_1824,N_1946);
nand U2137 (N_2137,N_1877,N_1906);
and U2138 (N_2138,N_2030,N_2045);
nand U2139 (N_2139,N_1966,N_1858);
nand U2140 (N_2140,N_1803,N_2063);
xor U2141 (N_2141,N_1976,N_2080);
nand U2142 (N_2142,N_2017,N_1979);
and U2143 (N_2143,N_1943,N_1995);
and U2144 (N_2144,N_1967,N_1816);
xnor U2145 (N_2145,N_1819,N_1944);
and U2146 (N_2146,N_2038,N_1855);
nand U2147 (N_2147,N_1987,N_2066);
and U2148 (N_2148,N_1868,N_1994);
nor U2149 (N_2149,N_2013,N_2073);
and U2150 (N_2150,N_1921,N_2061);
nand U2151 (N_2151,N_2029,N_1817);
and U2152 (N_2152,N_2070,N_2077);
xor U2153 (N_2153,N_1892,N_1820);
and U2154 (N_2154,N_1954,N_1968);
nor U2155 (N_2155,N_2085,N_1874);
or U2156 (N_2156,N_1920,N_2009);
and U2157 (N_2157,N_1938,N_2072);
xor U2158 (N_2158,N_2015,N_2003);
and U2159 (N_2159,N_1910,N_1843);
xnor U2160 (N_2160,N_1872,N_1829);
xor U2161 (N_2161,N_2044,N_1848);
or U2162 (N_2162,N_2076,N_1989);
xor U2163 (N_2163,N_2023,N_1934);
nor U2164 (N_2164,N_1864,N_1899);
or U2165 (N_2165,N_1958,N_1908);
nor U2166 (N_2166,N_1852,N_2074);
nor U2167 (N_2167,N_2093,N_2041);
nor U2168 (N_2168,N_1975,N_1837);
nand U2169 (N_2169,N_1917,N_1836);
and U2170 (N_2170,N_1982,N_2043);
nand U2171 (N_2171,N_1922,N_1828);
xor U2172 (N_2172,N_2097,N_1830);
xnor U2173 (N_2173,N_1871,N_1857);
nor U2174 (N_2174,N_1840,N_1949);
or U2175 (N_2175,N_1902,N_2048);
nor U2176 (N_2176,N_2089,N_1950);
nand U2177 (N_2177,N_1986,N_1801);
and U2178 (N_2178,N_1983,N_1895);
and U2179 (N_2179,N_1931,N_1963);
and U2180 (N_2180,N_1970,N_2018);
or U2181 (N_2181,N_1955,N_2090);
and U2182 (N_2182,N_1971,N_1940);
nor U2183 (N_2183,N_1935,N_1926);
and U2184 (N_2184,N_1886,N_1867);
xnor U2185 (N_2185,N_2008,N_1806);
and U2186 (N_2186,N_1911,N_2004);
and U2187 (N_2187,N_2081,N_1900);
nor U2188 (N_2188,N_1800,N_1904);
xnor U2189 (N_2189,N_1898,N_1959);
or U2190 (N_2190,N_1876,N_1964);
nor U2191 (N_2191,N_1947,N_1839);
nor U2192 (N_2192,N_1844,N_1996);
or U2193 (N_2193,N_2047,N_1833);
or U2194 (N_2194,N_2057,N_1880);
nor U2195 (N_2195,N_1939,N_2011);
xnor U2196 (N_2196,N_2056,N_1969);
and U2197 (N_2197,N_1842,N_1927);
and U2198 (N_2198,N_1853,N_1814);
and U2199 (N_2199,N_1951,N_2031);
nand U2200 (N_2200,N_2095,N_1809);
nor U2201 (N_2201,N_1818,N_1914);
nor U2202 (N_2202,N_2092,N_1849);
nor U2203 (N_2203,N_2096,N_1879);
or U2204 (N_2204,N_1804,N_2027);
or U2205 (N_2205,N_2067,N_1960);
nor U2206 (N_2206,N_1866,N_1977);
nor U2207 (N_2207,N_2025,N_1981);
nor U2208 (N_2208,N_1974,N_1854);
xor U2209 (N_2209,N_2091,N_2022);
nand U2210 (N_2210,N_1965,N_1863);
xnor U2211 (N_2211,N_1957,N_1883);
nand U2212 (N_2212,N_1807,N_2028);
nor U2213 (N_2213,N_1915,N_1846);
xor U2214 (N_2214,N_1887,N_2046);
or U2215 (N_2215,N_1941,N_1862);
or U2216 (N_2216,N_1937,N_1999);
xnor U2217 (N_2217,N_1942,N_2019);
or U2218 (N_2218,N_1825,N_1925);
and U2219 (N_2219,N_1956,N_1859);
xor U2220 (N_2220,N_2099,N_2002);
xor U2221 (N_2221,N_1888,N_2037);
nand U2222 (N_2222,N_1907,N_1821);
xnor U2223 (N_2223,N_1919,N_1827);
nor U2224 (N_2224,N_2036,N_1932);
nor U2225 (N_2225,N_1948,N_1952);
nand U2226 (N_2226,N_1831,N_2088);
nor U2227 (N_2227,N_2079,N_1845);
and U2228 (N_2228,N_2039,N_1823);
nor U2229 (N_2229,N_1832,N_2051);
nand U2230 (N_2230,N_1905,N_1972);
and U2231 (N_2231,N_1897,N_2065);
or U2232 (N_2232,N_1813,N_2068);
nor U2233 (N_2233,N_1875,N_1882);
nor U2234 (N_2234,N_1884,N_1826);
or U2235 (N_2235,N_2069,N_2050);
nand U2236 (N_2236,N_1890,N_1851);
or U2237 (N_2237,N_1896,N_1865);
and U2238 (N_2238,N_1913,N_2032);
nor U2239 (N_2239,N_2098,N_1990);
or U2240 (N_2240,N_2075,N_2035);
nand U2241 (N_2241,N_2082,N_1861);
or U2242 (N_2242,N_2040,N_2016);
nand U2243 (N_2243,N_1993,N_2083);
xnor U2244 (N_2244,N_1930,N_2000);
or U2245 (N_2245,N_1822,N_1973);
nand U2246 (N_2246,N_1918,N_2049);
nand U2247 (N_2247,N_2042,N_2026);
nor U2248 (N_2248,N_1805,N_1997);
or U2249 (N_2249,N_2014,N_1893);
or U2250 (N_2250,N_2001,N_1891);
xor U2251 (N_2251,N_2089,N_1807);
nand U2252 (N_2252,N_2003,N_1838);
or U2253 (N_2253,N_1831,N_1913);
xor U2254 (N_2254,N_1953,N_1864);
nor U2255 (N_2255,N_1949,N_1897);
nor U2256 (N_2256,N_1981,N_1895);
or U2257 (N_2257,N_2069,N_2071);
xnor U2258 (N_2258,N_1984,N_1990);
nand U2259 (N_2259,N_1943,N_2094);
xnor U2260 (N_2260,N_2062,N_2020);
nand U2261 (N_2261,N_2096,N_1922);
and U2262 (N_2262,N_1949,N_1908);
and U2263 (N_2263,N_1879,N_1921);
nor U2264 (N_2264,N_2083,N_1997);
nand U2265 (N_2265,N_1985,N_2070);
nand U2266 (N_2266,N_1819,N_1893);
nor U2267 (N_2267,N_1817,N_1993);
or U2268 (N_2268,N_2099,N_2066);
nor U2269 (N_2269,N_2065,N_1835);
nand U2270 (N_2270,N_1931,N_2046);
nor U2271 (N_2271,N_1900,N_2027);
nor U2272 (N_2272,N_1911,N_1946);
or U2273 (N_2273,N_2045,N_2046);
and U2274 (N_2274,N_2076,N_1814);
nand U2275 (N_2275,N_2058,N_1854);
or U2276 (N_2276,N_1804,N_2075);
or U2277 (N_2277,N_1905,N_1826);
and U2278 (N_2278,N_1808,N_1946);
xor U2279 (N_2279,N_2014,N_1831);
xnor U2280 (N_2280,N_1929,N_2003);
nor U2281 (N_2281,N_1940,N_1804);
and U2282 (N_2282,N_1816,N_1835);
nand U2283 (N_2283,N_2043,N_1924);
nand U2284 (N_2284,N_1828,N_1992);
nand U2285 (N_2285,N_1991,N_2067);
or U2286 (N_2286,N_1994,N_2050);
xor U2287 (N_2287,N_1911,N_1881);
and U2288 (N_2288,N_2095,N_1819);
nor U2289 (N_2289,N_1853,N_1864);
or U2290 (N_2290,N_1977,N_1975);
and U2291 (N_2291,N_2018,N_1996);
nand U2292 (N_2292,N_2058,N_1905);
nand U2293 (N_2293,N_1950,N_1973);
or U2294 (N_2294,N_1953,N_1930);
xnor U2295 (N_2295,N_1977,N_1875);
xor U2296 (N_2296,N_1868,N_2085);
nor U2297 (N_2297,N_1853,N_1909);
nand U2298 (N_2298,N_1977,N_2022);
xnor U2299 (N_2299,N_1991,N_2023);
or U2300 (N_2300,N_1851,N_1857);
nand U2301 (N_2301,N_1894,N_2085);
or U2302 (N_2302,N_1886,N_1900);
nand U2303 (N_2303,N_1907,N_1959);
and U2304 (N_2304,N_2027,N_2071);
or U2305 (N_2305,N_1809,N_1928);
and U2306 (N_2306,N_1806,N_1985);
nand U2307 (N_2307,N_1882,N_2076);
or U2308 (N_2308,N_1994,N_2006);
xnor U2309 (N_2309,N_1872,N_1939);
xnor U2310 (N_2310,N_1826,N_1827);
nand U2311 (N_2311,N_2061,N_1979);
nor U2312 (N_2312,N_1980,N_2005);
and U2313 (N_2313,N_1964,N_1883);
or U2314 (N_2314,N_1842,N_1921);
xnor U2315 (N_2315,N_1802,N_2038);
xor U2316 (N_2316,N_1822,N_1949);
xnor U2317 (N_2317,N_1925,N_2077);
or U2318 (N_2318,N_2033,N_2060);
and U2319 (N_2319,N_1868,N_2094);
or U2320 (N_2320,N_2087,N_1829);
or U2321 (N_2321,N_1967,N_1968);
or U2322 (N_2322,N_1863,N_2030);
and U2323 (N_2323,N_2011,N_1981);
and U2324 (N_2324,N_2022,N_1911);
and U2325 (N_2325,N_2070,N_1979);
nor U2326 (N_2326,N_2045,N_2001);
nand U2327 (N_2327,N_1828,N_1968);
xnor U2328 (N_2328,N_1862,N_1840);
nand U2329 (N_2329,N_1886,N_2025);
or U2330 (N_2330,N_1928,N_2088);
nor U2331 (N_2331,N_1958,N_1842);
nand U2332 (N_2332,N_1948,N_2047);
xnor U2333 (N_2333,N_1956,N_1888);
and U2334 (N_2334,N_2030,N_1982);
nor U2335 (N_2335,N_2053,N_1950);
xnor U2336 (N_2336,N_1961,N_1954);
nand U2337 (N_2337,N_1974,N_1901);
or U2338 (N_2338,N_1847,N_1860);
nand U2339 (N_2339,N_2026,N_1974);
and U2340 (N_2340,N_1895,N_1810);
xor U2341 (N_2341,N_1855,N_1941);
nor U2342 (N_2342,N_1864,N_1849);
nand U2343 (N_2343,N_1896,N_1804);
xnor U2344 (N_2344,N_2003,N_1966);
xnor U2345 (N_2345,N_1809,N_2093);
nor U2346 (N_2346,N_2062,N_2048);
xor U2347 (N_2347,N_1819,N_1882);
nand U2348 (N_2348,N_1903,N_1899);
and U2349 (N_2349,N_1975,N_1931);
or U2350 (N_2350,N_1946,N_2018);
and U2351 (N_2351,N_1877,N_1847);
xor U2352 (N_2352,N_2053,N_1933);
nor U2353 (N_2353,N_1923,N_2024);
nand U2354 (N_2354,N_1883,N_2090);
nand U2355 (N_2355,N_1990,N_1826);
or U2356 (N_2356,N_2037,N_2077);
nand U2357 (N_2357,N_1925,N_1818);
xor U2358 (N_2358,N_2067,N_2027);
xnor U2359 (N_2359,N_1890,N_1812);
nor U2360 (N_2360,N_2091,N_1954);
xnor U2361 (N_2361,N_1947,N_1896);
or U2362 (N_2362,N_2081,N_2073);
nand U2363 (N_2363,N_1802,N_1921);
nor U2364 (N_2364,N_2058,N_2036);
and U2365 (N_2365,N_1829,N_1970);
nor U2366 (N_2366,N_1986,N_2000);
or U2367 (N_2367,N_1924,N_1865);
nor U2368 (N_2368,N_1996,N_2025);
xor U2369 (N_2369,N_1912,N_2041);
nor U2370 (N_2370,N_1878,N_2058);
or U2371 (N_2371,N_1999,N_1843);
and U2372 (N_2372,N_1883,N_1976);
nor U2373 (N_2373,N_1923,N_1881);
nor U2374 (N_2374,N_1978,N_1862);
or U2375 (N_2375,N_1893,N_1874);
xnor U2376 (N_2376,N_1911,N_2016);
xnor U2377 (N_2377,N_1834,N_1931);
and U2378 (N_2378,N_1955,N_1910);
or U2379 (N_2379,N_1880,N_1851);
or U2380 (N_2380,N_2006,N_1947);
nand U2381 (N_2381,N_1910,N_1993);
or U2382 (N_2382,N_1914,N_2046);
nor U2383 (N_2383,N_1912,N_1890);
nor U2384 (N_2384,N_1898,N_1919);
and U2385 (N_2385,N_2022,N_1923);
xnor U2386 (N_2386,N_2047,N_2022);
xnor U2387 (N_2387,N_1831,N_1888);
nor U2388 (N_2388,N_2037,N_2007);
and U2389 (N_2389,N_1829,N_1817);
xnor U2390 (N_2390,N_1809,N_2052);
xnor U2391 (N_2391,N_2065,N_1888);
nor U2392 (N_2392,N_2006,N_1915);
nor U2393 (N_2393,N_2020,N_2044);
nand U2394 (N_2394,N_1929,N_2082);
xnor U2395 (N_2395,N_1865,N_2014);
or U2396 (N_2396,N_1991,N_1815);
nand U2397 (N_2397,N_2026,N_2034);
nand U2398 (N_2398,N_1995,N_1986);
xnor U2399 (N_2399,N_1964,N_1839);
nand U2400 (N_2400,N_2288,N_2351);
nand U2401 (N_2401,N_2386,N_2119);
nand U2402 (N_2402,N_2310,N_2175);
and U2403 (N_2403,N_2194,N_2138);
or U2404 (N_2404,N_2127,N_2329);
and U2405 (N_2405,N_2352,N_2214);
or U2406 (N_2406,N_2221,N_2371);
nor U2407 (N_2407,N_2174,N_2297);
nand U2408 (N_2408,N_2286,N_2301);
or U2409 (N_2409,N_2195,N_2375);
xor U2410 (N_2410,N_2167,N_2392);
xor U2411 (N_2411,N_2285,N_2284);
nor U2412 (N_2412,N_2249,N_2384);
and U2413 (N_2413,N_2134,N_2341);
and U2414 (N_2414,N_2343,N_2205);
nand U2415 (N_2415,N_2391,N_2115);
nand U2416 (N_2416,N_2185,N_2325);
xor U2417 (N_2417,N_2118,N_2184);
xor U2418 (N_2418,N_2238,N_2208);
nor U2419 (N_2419,N_2355,N_2105);
nor U2420 (N_2420,N_2299,N_2233);
nor U2421 (N_2421,N_2120,N_2260);
xor U2422 (N_2422,N_2101,N_2168);
or U2423 (N_2423,N_2227,N_2287);
nand U2424 (N_2424,N_2157,N_2378);
xor U2425 (N_2425,N_2346,N_2109);
or U2426 (N_2426,N_2222,N_2318);
nand U2427 (N_2427,N_2296,N_2149);
nand U2428 (N_2428,N_2158,N_2156);
nand U2429 (N_2429,N_2394,N_2182);
or U2430 (N_2430,N_2348,N_2376);
or U2431 (N_2431,N_2212,N_2294);
or U2432 (N_2432,N_2103,N_2319);
nor U2433 (N_2433,N_2316,N_2326);
nor U2434 (N_2434,N_2183,N_2271);
xor U2435 (N_2435,N_2177,N_2148);
nor U2436 (N_2436,N_2322,N_2209);
and U2437 (N_2437,N_2180,N_2330);
and U2438 (N_2438,N_2229,N_2144);
or U2439 (N_2439,N_2372,N_2360);
nor U2440 (N_2440,N_2151,N_2226);
xnor U2441 (N_2441,N_2273,N_2317);
or U2442 (N_2442,N_2276,N_2283);
or U2443 (N_2443,N_2201,N_2303);
xor U2444 (N_2444,N_2161,N_2267);
nand U2445 (N_2445,N_2363,N_2154);
and U2446 (N_2446,N_2126,N_2274);
or U2447 (N_2447,N_2112,N_2170);
xor U2448 (N_2448,N_2110,N_2121);
and U2449 (N_2449,N_2179,N_2186);
nor U2450 (N_2450,N_2137,N_2150);
and U2451 (N_2451,N_2388,N_2128);
nand U2452 (N_2452,N_2390,N_2256);
nand U2453 (N_2453,N_2277,N_2198);
xnor U2454 (N_2454,N_2344,N_2236);
xor U2455 (N_2455,N_2328,N_2162);
xor U2456 (N_2456,N_2262,N_2106);
and U2457 (N_2457,N_2247,N_2298);
nand U2458 (N_2458,N_2171,N_2333);
nor U2459 (N_2459,N_2327,N_2129);
nand U2460 (N_2460,N_2231,N_2114);
nand U2461 (N_2461,N_2200,N_2189);
or U2462 (N_2462,N_2241,N_2377);
nor U2463 (N_2463,N_2315,N_2323);
or U2464 (N_2464,N_2374,N_2246);
nor U2465 (N_2465,N_2237,N_2136);
xnor U2466 (N_2466,N_2362,N_2204);
nand U2467 (N_2467,N_2396,N_2337);
xnor U2468 (N_2468,N_2387,N_2336);
and U2469 (N_2469,N_2385,N_2311);
or U2470 (N_2470,N_2359,N_2218);
nand U2471 (N_2471,N_2223,N_2232);
nand U2472 (N_2472,N_2193,N_2141);
or U2473 (N_2473,N_2219,N_2293);
nor U2474 (N_2474,N_2117,N_2187);
xnor U2475 (N_2475,N_2111,N_2133);
nand U2476 (N_2476,N_2230,N_2353);
and U2477 (N_2477,N_2313,N_2216);
xnor U2478 (N_2478,N_2291,N_2248);
xor U2479 (N_2479,N_2305,N_2347);
and U2480 (N_2480,N_2381,N_2124);
or U2481 (N_2481,N_2269,N_2272);
and U2482 (N_2482,N_2373,N_2142);
xor U2483 (N_2483,N_2196,N_2250);
or U2484 (N_2484,N_2321,N_2253);
or U2485 (N_2485,N_2261,N_2320);
nor U2486 (N_2486,N_2116,N_2102);
nor U2487 (N_2487,N_2251,N_2395);
nor U2488 (N_2488,N_2345,N_2181);
nor U2489 (N_2489,N_2255,N_2113);
or U2490 (N_2490,N_2278,N_2338);
nand U2491 (N_2491,N_2289,N_2135);
xnor U2492 (N_2492,N_2398,N_2140);
nor U2493 (N_2493,N_2191,N_2324);
and U2494 (N_2494,N_2339,N_2202);
and U2495 (N_2495,N_2139,N_2163);
and U2496 (N_2496,N_2302,N_2397);
or U2497 (N_2497,N_2370,N_2122);
nand U2498 (N_2498,N_2350,N_2281);
and U2499 (N_2499,N_2306,N_2169);
nor U2500 (N_2500,N_2280,N_2234);
and U2501 (N_2501,N_2257,N_2143);
nor U2502 (N_2502,N_2357,N_2153);
xor U2503 (N_2503,N_2146,N_2178);
and U2504 (N_2504,N_2107,N_2332);
nor U2505 (N_2505,N_2308,N_2279);
nor U2506 (N_2506,N_2243,N_2244);
xnor U2507 (N_2507,N_2266,N_2399);
or U2508 (N_2508,N_2217,N_2354);
xor U2509 (N_2509,N_2123,N_2155);
nor U2510 (N_2510,N_2188,N_2206);
nand U2511 (N_2511,N_2264,N_2309);
xnor U2512 (N_2512,N_2259,N_2225);
nand U2513 (N_2513,N_2252,N_2240);
and U2514 (N_2514,N_2164,N_2331);
and U2515 (N_2515,N_2125,N_2145);
nand U2516 (N_2516,N_2369,N_2270);
xnor U2517 (N_2517,N_2295,N_2176);
xor U2518 (N_2518,N_2265,N_2300);
nor U2519 (N_2519,N_2361,N_2379);
nand U2520 (N_2520,N_2131,N_2173);
nand U2521 (N_2521,N_2132,N_2211);
nand U2522 (N_2522,N_2356,N_2393);
or U2523 (N_2523,N_2389,N_2340);
or U2524 (N_2524,N_2349,N_2235);
and U2525 (N_2525,N_2258,N_2160);
or U2526 (N_2526,N_2380,N_2314);
nor U2527 (N_2527,N_2292,N_2197);
and U2528 (N_2528,N_2282,N_2165);
or U2529 (N_2529,N_2335,N_2224);
nor U2530 (N_2530,N_2213,N_2290);
nand U2531 (N_2531,N_2242,N_2108);
nor U2532 (N_2532,N_2220,N_2239);
and U2533 (N_2533,N_2228,N_2130);
or U2534 (N_2534,N_2342,N_2268);
and U2535 (N_2535,N_2192,N_2312);
nand U2536 (N_2536,N_2245,N_2334);
xnor U2537 (N_2537,N_2304,N_2364);
nor U2538 (N_2538,N_2383,N_2166);
or U2539 (N_2539,N_2263,N_2203);
xnor U2540 (N_2540,N_2199,N_2207);
nor U2541 (N_2541,N_2368,N_2152);
nor U2542 (N_2542,N_2210,N_2159);
nand U2543 (N_2543,N_2367,N_2365);
nand U2544 (N_2544,N_2100,N_2215);
xor U2545 (N_2545,N_2172,N_2366);
nor U2546 (N_2546,N_2275,N_2254);
nor U2547 (N_2547,N_2190,N_2382);
or U2548 (N_2548,N_2307,N_2104);
nand U2549 (N_2549,N_2358,N_2147);
nor U2550 (N_2550,N_2383,N_2136);
nor U2551 (N_2551,N_2133,N_2238);
and U2552 (N_2552,N_2294,N_2398);
and U2553 (N_2553,N_2221,N_2363);
xor U2554 (N_2554,N_2113,N_2117);
or U2555 (N_2555,N_2244,N_2151);
nand U2556 (N_2556,N_2185,N_2178);
or U2557 (N_2557,N_2311,N_2376);
nand U2558 (N_2558,N_2179,N_2299);
xnor U2559 (N_2559,N_2314,N_2254);
nand U2560 (N_2560,N_2276,N_2217);
or U2561 (N_2561,N_2124,N_2302);
and U2562 (N_2562,N_2349,N_2366);
nand U2563 (N_2563,N_2226,N_2391);
xor U2564 (N_2564,N_2109,N_2262);
nor U2565 (N_2565,N_2246,N_2373);
or U2566 (N_2566,N_2249,N_2191);
nand U2567 (N_2567,N_2271,N_2374);
nand U2568 (N_2568,N_2310,N_2301);
and U2569 (N_2569,N_2229,N_2246);
and U2570 (N_2570,N_2156,N_2213);
nor U2571 (N_2571,N_2299,N_2304);
nand U2572 (N_2572,N_2346,N_2100);
xnor U2573 (N_2573,N_2122,N_2339);
or U2574 (N_2574,N_2319,N_2142);
and U2575 (N_2575,N_2125,N_2128);
and U2576 (N_2576,N_2191,N_2360);
and U2577 (N_2577,N_2255,N_2389);
or U2578 (N_2578,N_2277,N_2203);
and U2579 (N_2579,N_2351,N_2103);
and U2580 (N_2580,N_2263,N_2348);
nand U2581 (N_2581,N_2388,N_2281);
or U2582 (N_2582,N_2125,N_2299);
nor U2583 (N_2583,N_2253,N_2328);
nand U2584 (N_2584,N_2145,N_2253);
nand U2585 (N_2585,N_2310,N_2116);
and U2586 (N_2586,N_2281,N_2376);
xnor U2587 (N_2587,N_2290,N_2141);
nand U2588 (N_2588,N_2158,N_2251);
nor U2589 (N_2589,N_2275,N_2112);
xnor U2590 (N_2590,N_2288,N_2246);
and U2591 (N_2591,N_2252,N_2155);
and U2592 (N_2592,N_2120,N_2189);
or U2593 (N_2593,N_2382,N_2377);
and U2594 (N_2594,N_2265,N_2220);
or U2595 (N_2595,N_2254,N_2382);
nor U2596 (N_2596,N_2205,N_2290);
and U2597 (N_2597,N_2293,N_2246);
nor U2598 (N_2598,N_2340,N_2213);
xnor U2599 (N_2599,N_2352,N_2170);
and U2600 (N_2600,N_2229,N_2274);
nor U2601 (N_2601,N_2253,N_2139);
nand U2602 (N_2602,N_2281,N_2317);
and U2603 (N_2603,N_2355,N_2214);
xor U2604 (N_2604,N_2238,N_2103);
nand U2605 (N_2605,N_2186,N_2352);
nor U2606 (N_2606,N_2312,N_2266);
and U2607 (N_2607,N_2207,N_2188);
xnor U2608 (N_2608,N_2306,N_2118);
nand U2609 (N_2609,N_2297,N_2393);
nor U2610 (N_2610,N_2244,N_2358);
or U2611 (N_2611,N_2190,N_2176);
and U2612 (N_2612,N_2205,N_2207);
nor U2613 (N_2613,N_2100,N_2388);
nand U2614 (N_2614,N_2228,N_2119);
nand U2615 (N_2615,N_2288,N_2326);
xnor U2616 (N_2616,N_2300,N_2120);
xnor U2617 (N_2617,N_2121,N_2308);
nor U2618 (N_2618,N_2373,N_2169);
nor U2619 (N_2619,N_2101,N_2249);
nor U2620 (N_2620,N_2267,N_2142);
nand U2621 (N_2621,N_2239,N_2232);
nand U2622 (N_2622,N_2228,N_2304);
or U2623 (N_2623,N_2247,N_2325);
or U2624 (N_2624,N_2332,N_2331);
and U2625 (N_2625,N_2392,N_2244);
nor U2626 (N_2626,N_2315,N_2120);
nor U2627 (N_2627,N_2301,N_2129);
nand U2628 (N_2628,N_2388,N_2215);
nor U2629 (N_2629,N_2228,N_2292);
nor U2630 (N_2630,N_2216,N_2201);
and U2631 (N_2631,N_2155,N_2151);
nor U2632 (N_2632,N_2306,N_2275);
or U2633 (N_2633,N_2374,N_2367);
or U2634 (N_2634,N_2389,N_2214);
xnor U2635 (N_2635,N_2305,N_2241);
nor U2636 (N_2636,N_2214,N_2378);
and U2637 (N_2637,N_2216,N_2271);
or U2638 (N_2638,N_2175,N_2160);
xor U2639 (N_2639,N_2224,N_2160);
or U2640 (N_2640,N_2213,N_2286);
and U2641 (N_2641,N_2205,N_2187);
and U2642 (N_2642,N_2221,N_2117);
and U2643 (N_2643,N_2145,N_2116);
or U2644 (N_2644,N_2231,N_2189);
xnor U2645 (N_2645,N_2221,N_2227);
xor U2646 (N_2646,N_2292,N_2101);
xor U2647 (N_2647,N_2301,N_2163);
nand U2648 (N_2648,N_2103,N_2216);
and U2649 (N_2649,N_2292,N_2104);
xnor U2650 (N_2650,N_2253,N_2213);
or U2651 (N_2651,N_2196,N_2237);
nor U2652 (N_2652,N_2386,N_2248);
or U2653 (N_2653,N_2259,N_2135);
and U2654 (N_2654,N_2382,N_2126);
or U2655 (N_2655,N_2119,N_2118);
xor U2656 (N_2656,N_2248,N_2297);
and U2657 (N_2657,N_2154,N_2150);
or U2658 (N_2658,N_2299,N_2277);
nand U2659 (N_2659,N_2385,N_2330);
nand U2660 (N_2660,N_2209,N_2297);
nor U2661 (N_2661,N_2260,N_2237);
or U2662 (N_2662,N_2327,N_2126);
or U2663 (N_2663,N_2159,N_2125);
or U2664 (N_2664,N_2386,N_2154);
or U2665 (N_2665,N_2133,N_2124);
or U2666 (N_2666,N_2297,N_2344);
nor U2667 (N_2667,N_2111,N_2184);
xor U2668 (N_2668,N_2325,N_2341);
nor U2669 (N_2669,N_2303,N_2210);
or U2670 (N_2670,N_2319,N_2338);
xnor U2671 (N_2671,N_2262,N_2149);
nand U2672 (N_2672,N_2396,N_2345);
or U2673 (N_2673,N_2294,N_2251);
and U2674 (N_2674,N_2226,N_2207);
xnor U2675 (N_2675,N_2391,N_2247);
or U2676 (N_2676,N_2241,N_2162);
and U2677 (N_2677,N_2284,N_2212);
nor U2678 (N_2678,N_2356,N_2303);
xor U2679 (N_2679,N_2269,N_2302);
nor U2680 (N_2680,N_2178,N_2124);
nand U2681 (N_2681,N_2332,N_2115);
nor U2682 (N_2682,N_2383,N_2125);
nand U2683 (N_2683,N_2112,N_2221);
xnor U2684 (N_2684,N_2153,N_2318);
and U2685 (N_2685,N_2300,N_2262);
and U2686 (N_2686,N_2315,N_2247);
nor U2687 (N_2687,N_2175,N_2297);
and U2688 (N_2688,N_2250,N_2386);
xor U2689 (N_2689,N_2328,N_2222);
nor U2690 (N_2690,N_2217,N_2308);
nor U2691 (N_2691,N_2102,N_2223);
nand U2692 (N_2692,N_2107,N_2348);
nor U2693 (N_2693,N_2335,N_2312);
xnor U2694 (N_2694,N_2205,N_2359);
xor U2695 (N_2695,N_2325,N_2182);
nand U2696 (N_2696,N_2301,N_2177);
and U2697 (N_2697,N_2209,N_2240);
or U2698 (N_2698,N_2279,N_2351);
nand U2699 (N_2699,N_2254,N_2133);
and U2700 (N_2700,N_2441,N_2623);
and U2701 (N_2701,N_2548,N_2587);
or U2702 (N_2702,N_2619,N_2620);
nor U2703 (N_2703,N_2459,N_2417);
or U2704 (N_2704,N_2500,N_2425);
nand U2705 (N_2705,N_2685,N_2554);
xor U2706 (N_2706,N_2515,N_2527);
nor U2707 (N_2707,N_2535,N_2525);
nor U2708 (N_2708,N_2482,N_2485);
nor U2709 (N_2709,N_2547,N_2690);
nand U2710 (N_2710,N_2454,N_2456);
or U2711 (N_2711,N_2446,N_2696);
xnor U2712 (N_2712,N_2511,N_2656);
and U2713 (N_2713,N_2664,N_2444);
nor U2714 (N_2714,N_2610,N_2418);
or U2715 (N_2715,N_2676,N_2595);
nand U2716 (N_2716,N_2533,N_2571);
and U2717 (N_2717,N_2488,N_2671);
or U2718 (N_2718,N_2529,N_2594);
or U2719 (N_2719,N_2470,N_2497);
or U2720 (N_2720,N_2622,N_2627);
or U2721 (N_2721,N_2419,N_2407);
or U2722 (N_2722,N_2439,N_2581);
nand U2723 (N_2723,N_2659,N_2504);
nor U2724 (N_2724,N_2578,N_2647);
nor U2725 (N_2725,N_2411,N_2635);
and U2726 (N_2726,N_2568,N_2556);
xnor U2727 (N_2727,N_2637,N_2626);
xnor U2728 (N_2728,N_2450,N_2674);
xor U2729 (N_2729,N_2406,N_2606);
xnor U2730 (N_2730,N_2557,N_2592);
and U2731 (N_2731,N_2435,N_2599);
and U2732 (N_2732,N_2634,N_2508);
or U2733 (N_2733,N_2445,N_2546);
nand U2734 (N_2734,N_2426,N_2458);
nor U2735 (N_2735,N_2440,N_2496);
nor U2736 (N_2736,N_2624,N_2538);
xor U2737 (N_2737,N_2513,N_2648);
xnor U2738 (N_2738,N_2598,N_2400);
nand U2739 (N_2739,N_2693,N_2494);
xnor U2740 (N_2740,N_2506,N_2583);
and U2741 (N_2741,N_2603,N_2574);
xor U2742 (N_2742,N_2668,N_2545);
nand U2743 (N_2743,N_2638,N_2608);
xor U2744 (N_2744,N_2537,N_2499);
nor U2745 (N_2745,N_2694,N_2692);
nand U2746 (N_2746,N_2457,N_2570);
xor U2747 (N_2747,N_2605,N_2510);
xor U2748 (N_2748,N_2474,N_2478);
xnor U2749 (N_2749,N_2484,N_2699);
or U2750 (N_2750,N_2616,N_2649);
nand U2751 (N_2751,N_2401,N_2489);
or U2752 (N_2752,N_2507,N_2531);
nand U2753 (N_2753,N_2675,N_2415);
nor U2754 (N_2754,N_2580,N_2480);
nand U2755 (N_2755,N_2503,N_2673);
nor U2756 (N_2756,N_2536,N_2633);
and U2757 (N_2757,N_2405,N_2629);
nor U2758 (N_2758,N_2588,N_2621);
or U2759 (N_2759,N_2644,N_2697);
nor U2760 (N_2760,N_2591,N_2684);
nand U2761 (N_2761,N_2609,N_2490);
nand U2762 (N_2762,N_2514,N_2472);
or U2763 (N_2763,N_2639,N_2560);
and U2764 (N_2764,N_2698,N_2462);
nand U2765 (N_2765,N_2534,N_2522);
and U2766 (N_2766,N_2453,N_2584);
nor U2767 (N_2767,N_2561,N_2614);
or U2768 (N_2768,N_2573,N_2617);
or U2769 (N_2769,N_2409,N_2577);
nand U2770 (N_2770,N_2495,N_2452);
and U2771 (N_2771,N_2688,N_2670);
or U2772 (N_2772,N_2467,N_2640);
or U2773 (N_2773,N_2564,N_2681);
or U2774 (N_2774,N_2569,N_2597);
nor U2775 (N_2775,N_2483,N_2553);
xor U2776 (N_2776,N_2412,N_2442);
or U2777 (N_2777,N_2526,N_2516);
and U2778 (N_2778,N_2505,N_2416);
xor U2779 (N_2779,N_2589,N_2437);
xor U2780 (N_2780,N_2487,N_2660);
and U2781 (N_2781,N_2424,N_2555);
xnor U2782 (N_2782,N_2543,N_2582);
nand U2783 (N_2783,N_2651,N_2601);
and U2784 (N_2784,N_2475,N_2461);
xnor U2785 (N_2785,N_2563,N_2524);
nor U2786 (N_2786,N_2566,N_2408);
nand U2787 (N_2787,N_2695,N_2518);
and U2788 (N_2788,N_2691,N_2476);
nand U2789 (N_2789,N_2469,N_2559);
or U2790 (N_2790,N_2471,N_2652);
or U2791 (N_2791,N_2679,N_2544);
nand U2792 (N_2792,N_2451,N_2613);
and U2793 (N_2793,N_2443,N_2641);
nand U2794 (N_2794,N_2414,N_2687);
or U2795 (N_2795,N_2643,N_2429);
xor U2796 (N_2796,N_2666,N_2632);
nor U2797 (N_2797,N_2539,N_2686);
and U2798 (N_2798,N_2593,N_2665);
xor U2799 (N_2799,N_2575,N_2654);
xnor U2800 (N_2800,N_2541,N_2572);
nor U2801 (N_2801,N_2473,N_2630);
or U2802 (N_2802,N_2540,N_2607);
and U2803 (N_2803,N_2512,N_2662);
nand U2804 (N_2804,N_2628,N_2523);
xor U2805 (N_2805,N_2669,N_2567);
or U2806 (N_2806,N_2667,N_2492);
xnor U2807 (N_2807,N_2600,N_2672);
and U2808 (N_2808,N_2436,N_2430);
xor U2809 (N_2809,N_2466,N_2528);
or U2810 (N_2810,N_2658,N_2447);
nand U2811 (N_2811,N_2428,N_2427);
nor U2812 (N_2812,N_2530,N_2565);
and U2813 (N_2813,N_2479,N_2657);
or U2814 (N_2814,N_2460,N_2455);
nand U2815 (N_2815,N_2551,N_2502);
or U2816 (N_2816,N_2596,N_2642);
and U2817 (N_2817,N_2618,N_2420);
and U2818 (N_2818,N_2585,N_2604);
xor U2819 (N_2819,N_2402,N_2520);
or U2820 (N_2820,N_2602,N_2653);
nand U2821 (N_2821,N_2631,N_2493);
nand U2822 (N_2822,N_2678,N_2612);
nand U2823 (N_2823,N_2663,N_2491);
nand U2824 (N_2824,N_2465,N_2615);
or U2825 (N_2825,N_2677,N_2661);
xnor U2826 (N_2826,N_2410,N_2517);
nor U2827 (N_2827,N_2645,N_2433);
nor U2828 (N_2828,N_2421,N_2432);
xor U2829 (N_2829,N_2636,N_2519);
nand U2830 (N_2830,N_2403,N_2650);
nand U2831 (N_2831,N_2683,N_2552);
xor U2832 (N_2832,N_2404,N_2434);
nand U2833 (N_2833,N_2611,N_2501);
and U2834 (N_2834,N_2431,N_2413);
nand U2835 (N_2835,N_2549,N_2463);
or U2836 (N_2836,N_2477,N_2422);
nor U2837 (N_2837,N_2486,N_2655);
or U2838 (N_2838,N_2448,N_2646);
xor U2839 (N_2839,N_2550,N_2586);
or U2840 (N_2840,N_2579,N_2562);
nor U2841 (N_2841,N_2590,N_2498);
and U2842 (N_2842,N_2558,N_2532);
nand U2843 (N_2843,N_2509,N_2682);
xnor U2844 (N_2844,N_2438,N_2576);
and U2845 (N_2845,N_2464,N_2468);
and U2846 (N_2846,N_2542,N_2680);
nor U2847 (N_2847,N_2449,N_2625);
xnor U2848 (N_2848,N_2481,N_2521);
xor U2849 (N_2849,N_2423,N_2689);
xnor U2850 (N_2850,N_2675,N_2577);
or U2851 (N_2851,N_2563,N_2571);
and U2852 (N_2852,N_2443,N_2465);
or U2853 (N_2853,N_2600,N_2632);
xnor U2854 (N_2854,N_2490,N_2678);
xnor U2855 (N_2855,N_2446,N_2623);
and U2856 (N_2856,N_2667,N_2516);
and U2857 (N_2857,N_2635,N_2453);
nand U2858 (N_2858,N_2507,N_2529);
nand U2859 (N_2859,N_2669,N_2481);
xnor U2860 (N_2860,N_2626,N_2458);
or U2861 (N_2861,N_2536,N_2435);
nand U2862 (N_2862,N_2651,N_2421);
nand U2863 (N_2863,N_2527,N_2599);
nor U2864 (N_2864,N_2514,N_2530);
and U2865 (N_2865,N_2576,N_2644);
or U2866 (N_2866,N_2425,N_2593);
or U2867 (N_2867,N_2451,N_2685);
nor U2868 (N_2868,N_2540,N_2465);
and U2869 (N_2869,N_2414,N_2452);
or U2870 (N_2870,N_2454,N_2581);
or U2871 (N_2871,N_2514,N_2582);
xor U2872 (N_2872,N_2537,N_2578);
nor U2873 (N_2873,N_2683,N_2589);
nor U2874 (N_2874,N_2520,N_2468);
nor U2875 (N_2875,N_2591,N_2465);
nor U2876 (N_2876,N_2629,N_2404);
xnor U2877 (N_2877,N_2563,N_2676);
or U2878 (N_2878,N_2494,N_2430);
nand U2879 (N_2879,N_2546,N_2578);
xnor U2880 (N_2880,N_2426,N_2606);
or U2881 (N_2881,N_2534,N_2584);
and U2882 (N_2882,N_2620,N_2502);
and U2883 (N_2883,N_2436,N_2463);
nor U2884 (N_2884,N_2616,N_2607);
nor U2885 (N_2885,N_2412,N_2504);
xor U2886 (N_2886,N_2431,N_2443);
xnor U2887 (N_2887,N_2449,N_2566);
or U2888 (N_2888,N_2600,N_2660);
nor U2889 (N_2889,N_2698,N_2548);
nor U2890 (N_2890,N_2603,N_2468);
nor U2891 (N_2891,N_2479,N_2594);
or U2892 (N_2892,N_2509,N_2401);
or U2893 (N_2893,N_2626,N_2634);
and U2894 (N_2894,N_2541,N_2638);
xnor U2895 (N_2895,N_2409,N_2464);
nand U2896 (N_2896,N_2472,N_2674);
and U2897 (N_2897,N_2580,N_2526);
nor U2898 (N_2898,N_2583,N_2648);
and U2899 (N_2899,N_2641,N_2562);
and U2900 (N_2900,N_2561,N_2410);
nand U2901 (N_2901,N_2423,N_2581);
and U2902 (N_2902,N_2497,N_2410);
and U2903 (N_2903,N_2482,N_2569);
xnor U2904 (N_2904,N_2613,N_2632);
and U2905 (N_2905,N_2436,N_2478);
and U2906 (N_2906,N_2685,N_2448);
nand U2907 (N_2907,N_2404,N_2549);
or U2908 (N_2908,N_2581,N_2526);
xnor U2909 (N_2909,N_2455,N_2534);
and U2910 (N_2910,N_2552,N_2439);
and U2911 (N_2911,N_2508,N_2431);
nand U2912 (N_2912,N_2550,N_2589);
or U2913 (N_2913,N_2575,N_2587);
nor U2914 (N_2914,N_2624,N_2663);
xnor U2915 (N_2915,N_2686,N_2676);
or U2916 (N_2916,N_2639,N_2503);
nor U2917 (N_2917,N_2528,N_2559);
xor U2918 (N_2918,N_2643,N_2630);
or U2919 (N_2919,N_2430,N_2605);
and U2920 (N_2920,N_2452,N_2694);
or U2921 (N_2921,N_2404,N_2662);
nor U2922 (N_2922,N_2588,N_2454);
xor U2923 (N_2923,N_2421,N_2552);
or U2924 (N_2924,N_2457,N_2462);
xnor U2925 (N_2925,N_2637,N_2527);
xor U2926 (N_2926,N_2620,N_2669);
nand U2927 (N_2927,N_2575,N_2474);
nor U2928 (N_2928,N_2520,N_2646);
and U2929 (N_2929,N_2614,N_2644);
nand U2930 (N_2930,N_2685,N_2498);
nor U2931 (N_2931,N_2635,N_2586);
xor U2932 (N_2932,N_2461,N_2449);
or U2933 (N_2933,N_2442,N_2402);
nand U2934 (N_2934,N_2402,N_2679);
or U2935 (N_2935,N_2537,N_2614);
or U2936 (N_2936,N_2664,N_2662);
xor U2937 (N_2937,N_2478,N_2443);
and U2938 (N_2938,N_2578,N_2406);
nand U2939 (N_2939,N_2664,N_2555);
nand U2940 (N_2940,N_2501,N_2492);
or U2941 (N_2941,N_2432,N_2516);
or U2942 (N_2942,N_2513,N_2653);
and U2943 (N_2943,N_2417,N_2457);
or U2944 (N_2944,N_2642,N_2612);
or U2945 (N_2945,N_2580,N_2623);
or U2946 (N_2946,N_2516,N_2498);
nand U2947 (N_2947,N_2645,N_2554);
or U2948 (N_2948,N_2697,N_2674);
or U2949 (N_2949,N_2408,N_2684);
and U2950 (N_2950,N_2479,N_2542);
or U2951 (N_2951,N_2460,N_2667);
or U2952 (N_2952,N_2554,N_2684);
or U2953 (N_2953,N_2553,N_2601);
and U2954 (N_2954,N_2586,N_2656);
nor U2955 (N_2955,N_2465,N_2427);
and U2956 (N_2956,N_2528,N_2409);
xor U2957 (N_2957,N_2539,N_2417);
nand U2958 (N_2958,N_2694,N_2676);
or U2959 (N_2959,N_2522,N_2626);
nor U2960 (N_2960,N_2438,N_2402);
xnor U2961 (N_2961,N_2502,N_2489);
nand U2962 (N_2962,N_2582,N_2404);
or U2963 (N_2963,N_2598,N_2682);
or U2964 (N_2964,N_2433,N_2466);
or U2965 (N_2965,N_2541,N_2592);
nand U2966 (N_2966,N_2670,N_2470);
and U2967 (N_2967,N_2605,N_2693);
nor U2968 (N_2968,N_2614,N_2475);
nor U2969 (N_2969,N_2652,N_2583);
or U2970 (N_2970,N_2553,N_2685);
or U2971 (N_2971,N_2411,N_2668);
nor U2972 (N_2972,N_2480,N_2640);
xor U2973 (N_2973,N_2476,N_2619);
xnor U2974 (N_2974,N_2639,N_2576);
nor U2975 (N_2975,N_2564,N_2574);
or U2976 (N_2976,N_2686,N_2690);
or U2977 (N_2977,N_2575,N_2588);
nand U2978 (N_2978,N_2608,N_2685);
nand U2979 (N_2979,N_2576,N_2582);
and U2980 (N_2980,N_2538,N_2622);
nand U2981 (N_2981,N_2668,N_2454);
and U2982 (N_2982,N_2617,N_2412);
nand U2983 (N_2983,N_2580,N_2683);
and U2984 (N_2984,N_2510,N_2453);
and U2985 (N_2985,N_2670,N_2481);
and U2986 (N_2986,N_2514,N_2466);
nand U2987 (N_2987,N_2480,N_2538);
or U2988 (N_2988,N_2614,N_2699);
nor U2989 (N_2989,N_2689,N_2520);
nor U2990 (N_2990,N_2588,N_2633);
and U2991 (N_2991,N_2612,N_2558);
and U2992 (N_2992,N_2418,N_2565);
nand U2993 (N_2993,N_2633,N_2433);
or U2994 (N_2994,N_2686,N_2457);
xor U2995 (N_2995,N_2530,N_2577);
nor U2996 (N_2996,N_2593,N_2522);
nor U2997 (N_2997,N_2546,N_2463);
nor U2998 (N_2998,N_2483,N_2423);
nor U2999 (N_2999,N_2430,N_2440);
nand U3000 (N_3000,N_2846,N_2777);
xor U3001 (N_3001,N_2880,N_2864);
or U3002 (N_3002,N_2878,N_2989);
nand U3003 (N_3003,N_2859,N_2705);
or U3004 (N_3004,N_2908,N_2960);
nand U3005 (N_3005,N_2722,N_2941);
xor U3006 (N_3006,N_2885,N_2884);
or U3007 (N_3007,N_2958,N_2854);
or U3008 (N_3008,N_2714,N_2966);
nor U3009 (N_3009,N_2724,N_2856);
nand U3010 (N_3010,N_2766,N_2788);
nand U3011 (N_3011,N_2725,N_2794);
nand U3012 (N_3012,N_2991,N_2821);
nand U3013 (N_3013,N_2817,N_2959);
xnor U3014 (N_3014,N_2848,N_2986);
and U3015 (N_3015,N_2801,N_2944);
nand U3016 (N_3016,N_2963,N_2962);
and U3017 (N_3017,N_2978,N_2759);
or U3018 (N_3018,N_2950,N_2793);
nor U3019 (N_3019,N_2851,N_2935);
xnor U3020 (N_3020,N_2765,N_2713);
nand U3021 (N_3021,N_2955,N_2928);
and U3022 (N_3022,N_2778,N_2707);
nor U3023 (N_3023,N_2740,N_2737);
xnor U3024 (N_3024,N_2853,N_2905);
and U3025 (N_3025,N_2761,N_2728);
nand U3026 (N_3026,N_2816,N_2920);
nand U3027 (N_3027,N_2805,N_2804);
xor U3028 (N_3028,N_2889,N_2918);
or U3029 (N_3029,N_2755,N_2814);
and U3030 (N_3030,N_2719,N_2985);
or U3031 (N_3031,N_2729,N_2818);
and U3032 (N_3032,N_2731,N_2974);
and U3033 (N_3033,N_2822,N_2927);
and U3034 (N_3034,N_2969,N_2939);
nor U3035 (N_3035,N_2909,N_2971);
xor U3036 (N_3036,N_2833,N_2942);
and U3037 (N_3037,N_2844,N_2839);
nor U3038 (N_3038,N_2704,N_2973);
and U3039 (N_3039,N_2734,N_2826);
nor U3040 (N_3040,N_2977,N_2715);
nor U3041 (N_3041,N_2862,N_2925);
nor U3042 (N_3042,N_2911,N_2983);
or U3043 (N_3043,N_2745,N_2797);
xor U3044 (N_3044,N_2947,N_2741);
nand U3045 (N_3045,N_2926,N_2799);
xor U3046 (N_3046,N_2965,N_2748);
xor U3047 (N_3047,N_2872,N_2727);
nand U3048 (N_3048,N_2735,N_2783);
nand U3049 (N_3049,N_2775,N_2840);
or U3050 (N_3050,N_2823,N_2994);
xor U3051 (N_3051,N_2847,N_2943);
or U3052 (N_3052,N_2838,N_2903);
xor U3053 (N_3053,N_2866,N_2841);
nand U3054 (N_3054,N_2824,N_2855);
xnor U3055 (N_3055,N_2896,N_2800);
nor U3056 (N_3056,N_2954,N_2786);
nand U3057 (N_3057,N_2747,N_2998);
or U3058 (N_3058,N_2730,N_2875);
nand U3059 (N_3059,N_2850,N_2753);
or U3060 (N_3060,N_2931,N_2791);
xnor U3061 (N_3061,N_2767,N_2837);
and U3062 (N_3062,N_2913,N_2723);
or U3063 (N_3063,N_2970,N_2988);
nor U3064 (N_3064,N_2716,N_2764);
xnor U3065 (N_3065,N_2802,N_2710);
or U3066 (N_3066,N_2781,N_2882);
nand U3067 (N_3067,N_2999,N_2789);
nand U3068 (N_3068,N_2803,N_2987);
and U3069 (N_3069,N_2934,N_2938);
or U3070 (N_3070,N_2770,N_2795);
and U3071 (N_3071,N_2711,N_2899);
and U3072 (N_3072,N_2744,N_2709);
nor U3073 (N_3073,N_2964,N_2924);
and U3074 (N_3074,N_2733,N_2750);
nor U3075 (N_3075,N_2769,N_2852);
nand U3076 (N_3076,N_2790,N_2886);
xnor U3077 (N_3077,N_2807,N_2949);
or U3078 (N_3078,N_2742,N_2910);
nand U3079 (N_3079,N_2961,N_2873);
or U3080 (N_3080,N_2808,N_2749);
or U3081 (N_3081,N_2771,N_2849);
or U3082 (N_3082,N_2825,N_2888);
nand U3083 (N_3083,N_2945,N_2923);
or U3084 (N_3084,N_2835,N_2891);
or U3085 (N_3085,N_2979,N_2809);
and U3086 (N_3086,N_2787,N_2813);
or U3087 (N_3087,N_2860,N_2952);
xnor U3088 (N_3088,N_2901,N_2915);
nand U3089 (N_3089,N_2746,N_2967);
and U3090 (N_3090,N_2917,N_2871);
nor U3091 (N_3091,N_2904,N_2890);
or U3092 (N_3092,N_2976,N_2701);
xor U3093 (N_3093,N_2990,N_2812);
or U3094 (N_3094,N_2776,N_2946);
nor U3095 (N_3095,N_2914,N_2900);
nor U3096 (N_3096,N_2857,N_2831);
or U3097 (N_3097,N_2932,N_2758);
xnor U3098 (N_3098,N_2876,N_2907);
nand U3099 (N_3099,N_2912,N_2726);
nand U3100 (N_3100,N_2754,N_2868);
and U3101 (N_3101,N_2763,N_2992);
and U3102 (N_3102,N_2982,N_2736);
or U3103 (N_3103,N_2780,N_2836);
or U3104 (N_3104,N_2951,N_2757);
nand U3105 (N_3105,N_2739,N_2832);
or U3106 (N_3106,N_2702,N_2718);
nor U3107 (N_3107,N_2732,N_2865);
and U3108 (N_3108,N_2842,N_2993);
or U3109 (N_3109,N_2929,N_2883);
nor U3110 (N_3110,N_2751,N_2861);
nor U3111 (N_3111,N_2972,N_2706);
or U3112 (N_3112,N_2922,N_2898);
nand U3113 (N_3113,N_2933,N_2829);
xor U3114 (N_3114,N_2984,N_2957);
and U3115 (N_3115,N_2717,N_2708);
and U3116 (N_3116,N_2834,N_2811);
xnor U3117 (N_3117,N_2877,N_2981);
or U3118 (N_3118,N_2863,N_2936);
xnor U3119 (N_3119,N_2806,N_2956);
xnor U3120 (N_3120,N_2784,N_2738);
nor U3121 (N_3121,N_2997,N_2874);
and U3122 (N_3122,N_2980,N_2895);
nor U3123 (N_3123,N_2869,N_2870);
or U3124 (N_3124,N_2995,N_2768);
nor U3125 (N_3125,N_2700,N_2828);
nand U3126 (N_3126,N_2703,N_2940);
or U3127 (N_3127,N_2712,N_2975);
and U3128 (N_3128,N_2892,N_2782);
nor U3129 (N_3129,N_2830,N_2792);
nor U3130 (N_3130,N_2760,N_2820);
and U3131 (N_3131,N_2919,N_2815);
or U3132 (N_3132,N_2774,N_2721);
nor U3133 (N_3133,N_2879,N_2720);
xor U3134 (N_3134,N_2843,N_2858);
nand U3135 (N_3135,N_2894,N_2897);
xnor U3136 (N_3136,N_2881,N_2827);
and U3137 (N_3137,N_2968,N_2906);
nor U3138 (N_3138,N_2798,N_2937);
nand U3139 (N_3139,N_2772,N_2867);
nor U3140 (N_3140,N_2762,N_2743);
nand U3141 (N_3141,N_2902,N_2893);
nor U3142 (N_3142,N_2752,N_2930);
and U3143 (N_3143,N_2756,N_2810);
and U3144 (N_3144,N_2996,N_2921);
and U3145 (N_3145,N_2819,N_2953);
nand U3146 (N_3146,N_2948,N_2916);
xnor U3147 (N_3147,N_2773,N_2845);
and U3148 (N_3148,N_2779,N_2887);
or U3149 (N_3149,N_2785,N_2796);
xor U3150 (N_3150,N_2797,N_2717);
nor U3151 (N_3151,N_2885,N_2896);
xor U3152 (N_3152,N_2737,N_2857);
xor U3153 (N_3153,N_2770,N_2766);
nor U3154 (N_3154,N_2718,N_2839);
xnor U3155 (N_3155,N_2765,N_2839);
and U3156 (N_3156,N_2914,N_2733);
or U3157 (N_3157,N_2997,N_2790);
or U3158 (N_3158,N_2941,N_2758);
or U3159 (N_3159,N_2889,N_2995);
xnor U3160 (N_3160,N_2949,N_2937);
or U3161 (N_3161,N_2953,N_2756);
or U3162 (N_3162,N_2924,N_2910);
nor U3163 (N_3163,N_2860,N_2967);
nor U3164 (N_3164,N_2956,N_2785);
or U3165 (N_3165,N_2933,N_2739);
and U3166 (N_3166,N_2855,N_2801);
and U3167 (N_3167,N_2946,N_2829);
nand U3168 (N_3168,N_2722,N_2752);
nor U3169 (N_3169,N_2989,N_2974);
nor U3170 (N_3170,N_2981,N_2829);
nor U3171 (N_3171,N_2705,N_2901);
and U3172 (N_3172,N_2770,N_2978);
xnor U3173 (N_3173,N_2763,N_2768);
nand U3174 (N_3174,N_2739,N_2702);
or U3175 (N_3175,N_2739,N_2734);
nor U3176 (N_3176,N_2941,N_2761);
or U3177 (N_3177,N_2716,N_2941);
nand U3178 (N_3178,N_2746,N_2827);
and U3179 (N_3179,N_2865,N_2959);
nor U3180 (N_3180,N_2705,N_2841);
nand U3181 (N_3181,N_2917,N_2704);
nor U3182 (N_3182,N_2757,N_2761);
or U3183 (N_3183,N_2754,N_2914);
and U3184 (N_3184,N_2975,N_2959);
or U3185 (N_3185,N_2996,N_2711);
or U3186 (N_3186,N_2952,N_2992);
nor U3187 (N_3187,N_2740,N_2739);
nand U3188 (N_3188,N_2772,N_2973);
nand U3189 (N_3189,N_2868,N_2894);
xor U3190 (N_3190,N_2967,N_2951);
and U3191 (N_3191,N_2747,N_2969);
and U3192 (N_3192,N_2762,N_2948);
xnor U3193 (N_3193,N_2847,N_2981);
or U3194 (N_3194,N_2848,N_2921);
and U3195 (N_3195,N_2956,N_2706);
or U3196 (N_3196,N_2832,N_2763);
or U3197 (N_3197,N_2773,N_2808);
xor U3198 (N_3198,N_2959,N_2931);
xnor U3199 (N_3199,N_2878,N_2891);
or U3200 (N_3200,N_2848,N_2879);
or U3201 (N_3201,N_2889,N_2983);
or U3202 (N_3202,N_2863,N_2934);
nand U3203 (N_3203,N_2765,N_2853);
or U3204 (N_3204,N_2830,N_2849);
xnor U3205 (N_3205,N_2758,N_2715);
or U3206 (N_3206,N_2723,N_2865);
xor U3207 (N_3207,N_2830,N_2890);
nor U3208 (N_3208,N_2966,N_2882);
nor U3209 (N_3209,N_2707,N_2903);
or U3210 (N_3210,N_2746,N_2892);
nand U3211 (N_3211,N_2990,N_2999);
nand U3212 (N_3212,N_2941,N_2995);
nor U3213 (N_3213,N_2877,N_2870);
nand U3214 (N_3214,N_2836,N_2843);
xor U3215 (N_3215,N_2832,N_2700);
nand U3216 (N_3216,N_2940,N_2717);
or U3217 (N_3217,N_2719,N_2727);
nor U3218 (N_3218,N_2986,N_2972);
nor U3219 (N_3219,N_2703,N_2828);
xnor U3220 (N_3220,N_2874,N_2969);
nor U3221 (N_3221,N_2952,N_2916);
nand U3222 (N_3222,N_2929,N_2822);
xor U3223 (N_3223,N_2856,N_2903);
nor U3224 (N_3224,N_2710,N_2789);
nand U3225 (N_3225,N_2900,N_2967);
xnor U3226 (N_3226,N_2971,N_2945);
nor U3227 (N_3227,N_2740,N_2843);
and U3228 (N_3228,N_2869,N_2971);
and U3229 (N_3229,N_2941,N_2756);
nor U3230 (N_3230,N_2700,N_2934);
nand U3231 (N_3231,N_2919,N_2914);
nor U3232 (N_3232,N_2986,N_2825);
nand U3233 (N_3233,N_2868,N_2865);
nor U3234 (N_3234,N_2972,N_2878);
and U3235 (N_3235,N_2930,N_2736);
xor U3236 (N_3236,N_2770,N_2726);
xor U3237 (N_3237,N_2898,N_2823);
or U3238 (N_3238,N_2909,N_2868);
or U3239 (N_3239,N_2975,N_2921);
xor U3240 (N_3240,N_2848,N_2906);
and U3241 (N_3241,N_2708,N_2770);
xnor U3242 (N_3242,N_2867,N_2887);
xor U3243 (N_3243,N_2882,N_2962);
and U3244 (N_3244,N_2872,N_2770);
xor U3245 (N_3245,N_2854,N_2793);
nor U3246 (N_3246,N_2868,N_2983);
nor U3247 (N_3247,N_2785,N_2906);
nand U3248 (N_3248,N_2993,N_2838);
or U3249 (N_3249,N_2721,N_2897);
nor U3250 (N_3250,N_2818,N_2710);
xnor U3251 (N_3251,N_2942,N_2795);
nor U3252 (N_3252,N_2779,N_2910);
xnor U3253 (N_3253,N_2807,N_2795);
or U3254 (N_3254,N_2990,N_2768);
and U3255 (N_3255,N_2797,N_2781);
or U3256 (N_3256,N_2908,N_2953);
nand U3257 (N_3257,N_2825,N_2865);
or U3258 (N_3258,N_2718,N_2833);
nand U3259 (N_3259,N_2805,N_2807);
or U3260 (N_3260,N_2933,N_2735);
and U3261 (N_3261,N_2796,N_2827);
nand U3262 (N_3262,N_2746,N_2824);
nand U3263 (N_3263,N_2781,N_2870);
nor U3264 (N_3264,N_2797,N_2863);
and U3265 (N_3265,N_2875,N_2972);
and U3266 (N_3266,N_2850,N_2960);
xor U3267 (N_3267,N_2782,N_2952);
nor U3268 (N_3268,N_2923,N_2912);
or U3269 (N_3269,N_2892,N_2903);
and U3270 (N_3270,N_2760,N_2982);
or U3271 (N_3271,N_2789,N_2706);
and U3272 (N_3272,N_2773,N_2822);
and U3273 (N_3273,N_2842,N_2848);
nand U3274 (N_3274,N_2930,N_2952);
nor U3275 (N_3275,N_2946,N_2791);
and U3276 (N_3276,N_2993,N_2854);
nand U3277 (N_3277,N_2873,N_2985);
xnor U3278 (N_3278,N_2887,N_2740);
xor U3279 (N_3279,N_2804,N_2942);
or U3280 (N_3280,N_2988,N_2926);
xnor U3281 (N_3281,N_2886,N_2918);
and U3282 (N_3282,N_2851,N_2747);
nor U3283 (N_3283,N_2841,N_2900);
xor U3284 (N_3284,N_2721,N_2817);
and U3285 (N_3285,N_2756,N_2760);
nand U3286 (N_3286,N_2739,N_2859);
nand U3287 (N_3287,N_2793,N_2795);
nand U3288 (N_3288,N_2893,N_2959);
xor U3289 (N_3289,N_2857,N_2920);
or U3290 (N_3290,N_2972,N_2954);
and U3291 (N_3291,N_2767,N_2981);
nor U3292 (N_3292,N_2956,N_2918);
or U3293 (N_3293,N_2711,N_2737);
nor U3294 (N_3294,N_2973,N_2792);
or U3295 (N_3295,N_2751,N_2758);
nand U3296 (N_3296,N_2830,N_2713);
nor U3297 (N_3297,N_2859,N_2720);
nor U3298 (N_3298,N_2885,N_2879);
and U3299 (N_3299,N_2835,N_2865);
or U3300 (N_3300,N_3200,N_3139);
nor U3301 (N_3301,N_3185,N_3075);
and U3302 (N_3302,N_3280,N_3134);
and U3303 (N_3303,N_3003,N_3255);
and U3304 (N_3304,N_3293,N_3024);
nor U3305 (N_3305,N_3167,N_3298);
or U3306 (N_3306,N_3269,N_3160);
or U3307 (N_3307,N_3154,N_3274);
and U3308 (N_3308,N_3251,N_3135);
and U3309 (N_3309,N_3085,N_3203);
or U3310 (N_3310,N_3172,N_3074);
nor U3311 (N_3311,N_3210,N_3041);
nand U3312 (N_3312,N_3263,N_3292);
and U3313 (N_3313,N_3052,N_3032);
nor U3314 (N_3314,N_3209,N_3174);
or U3315 (N_3315,N_3063,N_3213);
xor U3316 (N_3316,N_3267,N_3219);
or U3317 (N_3317,N_3101,N_3230);
and U3318 (N_3318,N_3073,N_3038);
nor U3319 (N_3319,N_3168,N_3001);
xnor U3320 (N_3320,N_3206,N_3272);
nand U3321 (N_3321,N_3067,N_3049);
nand U3322 (N_3322,N_3009,N_3090);
and U3323 (N_3323,N_3146,N_3109);
and U3324 (N_3324,N_3247,N_3008);
or U3325 (N_3325,N_3045,N_3201);
or U3326 (N_3326,N_3130,N_3002);
or U3327 (N_3327,N_3028,N_3264);
and U3328 (N_3328,N_3088,N_3114);
and U3329 (N_3329,N_3241,N_3012);
or U3330 (N_3330,N_3187,N_3061);
nor U3331 (N_3331,N_3016,N_3112);
nand U3332 (N_3332,N_3020,N_3047);
or U3333 (N_3333,N_3176,N_3126);
nor U3334 (N_3334,N_3148,N_3031);
nand U3335 (N_3335,N_3068,N_3297);
xor U3336 (N_3336,N_3093,N_3216);
and U3337 (N_3337,N_3244,N_3190);
and U3338 (N_3338,N_3159,N_3042);
and U3339 (N_3339,N_3055,N_3158);
and U3340 (N_3340,N_3277,N_3260);
or U3341 (N_3341,N_3107,N_3117);
nand U3342 (N_3342,N_3243,N_3278);
or U3343 (N_3343,N_3091,N_3248);
xnor U3344 (N_3344,N_3223,N_3258);
and U3345 (N_3345,N_3207,N_3137);
xor U3346 (N_3346,N_3053,N_3170);
xnor U3347 (N_3347,N_3100,N_3026);
nand U3348 (N_3348,N_3034,N_3262);
nor U3349 (N_3349,N_3083,N_3150);
xnor U3350 (N_3350,N_3268,N_3182);
nor U3351 (N_3351,N_3145,N_3071);
nor U3352 (N_3352,N_3197,N_3108);
nand U3353 (N_3353,N_3023,N_3022);
xor U3354 (N_3354,N_3081,N_3196);
xor U3355 (N_3355,N_3084,N_3129);
nor U3356 (N_3356,N_3184,N_3044);
xor U3357 (N_3357,N_3133,N_3218);
xor U3358 (N_3358,N_3070,N_3141);
xnor U3359 (N_3359,N_3040,N_3180);
nor U3360 (N_3360,N_3005,N_3198);
or U3361 (N_3361,N_3118,N_3163);
or U3362 (N_3362,N_3221,N_3286);
xnor U3363 (N_3363,N_3127,N_3078);
and U3364 (N_3364,N_3236,N_3122);
or U3365 (N_3365,N_3238,N_3110);
and U3366 (N_3366,N_3030,N_3065);
and U3367 (N_3367,N_3037,N_3283);
or U3368 (N_3368,N_3069,N_3120);
nand U3369 (N_3369,N_3270,N_3102);
and U3370 (N_3370,N_3115,N_3025);
or U3371 (N_3371,N_3036,N_3017);
and U3372 (N_3372,N_3193,N_3128);
nand U3373 (N_3373,N_3010,N_3169);
xnor U3374 (N_3374,N_3189,N_3132);
and U3375 (N_3375,N_3291,N_3076);
xnor U3376 (N_3376,N_3224,N_3246);
nor U3377 (N_3377,N_3296,N_3097);
and U3378 (N_3378,N_3089,N_3029);
xor U3379 (N_3379,N_3153,N_3188);
nand U3380 (N_3380,N_3059,N_3181);
nand U3381 (N_3381,N_3051,N_3217);
xnor U3382 (N_3382,N_3048,N_3199);
nor U3383 (N_3383,N_3254,N_3057);
or U3384 (N_3384,N_3046,N_3062);
and U3385 (N_3385,N_3099,N_3152);
or U3386 (N_3386,N_3166,N_3098);
or U3387 (N_3387,N_3155,N_3231);
and U3388 (N_3388,N_3156,N_3281);
xor U3389 (N_3389,N_3054,N_3094);
or U3390 (N_3390,N_3289,N_3228);
nor U3391 (N_3391,N_3173,N_3004);
nand U3392 (N_3392,N_3215,N_3104);
and U3393 (N_3393,N_3257,N_3271);
nand U3394 (N_3394,N_3125,N_3131);
and U3395 (N_3395,N_3205,N_3233);
and U3396 (N_3396,N_3266,N_3095);
nor U3397 (N_3397,N_3252,N_3214);
and U3398 (N_3398,N_3232,N_3211);
nor U3399 (N_3399,N_3013,N_3276);
or U3400 (N_3400,N_3006,N_3178);
nand U3401 (N_3401,N_3007,N_3242);
nor U3402 (N_3402,N_3039,N_3119);
and U3403 (N_3403,N_3240,N_3014);
or U3404 (N_3404,N_3227,N_3287);
nor U3405 (N_3405,N_3082,N_3234);
or U3406 (N_3406,N_3229,N_3275);
nand U3407 (N_3407,N_3080,N_3195);
xnor U3408 (N_3408,N_3225,N_3050);
nand U3409 (N_3409,N_3140,N_3259);
nand U3410 (N_3410,N_3290,N_3285);
or U3411 (N_3411,N_3179,N_3124);
xnor U3412 (N_3412,N_3245,N_3256);
xor U3413 (N_3413,N_3011,N_3273);
or U3414 (N_3414,N_3033,N_3019);
nor U3415 (N_3415,N_3186,N_3027);
and U3416 (N_3416,N_3092,N_3250);
or U3417 (N_3417,N_3237,N_3220);
or U3418 (N_3418,N_3018,N_3202);
or U3419 (N_3419,N_3123,N_3157);
or U3420 (N_3420,N_3015,N_3239);
and U3421 (N_3421,N_3058,N_3235);
nor U3422 (N_3422,N_3106,N_3295);
and U3423 (N_3423,N_3294,N_3149);
nand U3424 (N_3424,N_3208,N_3087);
xnor U3425 (N_3425,N_3265,N_3035);
xnor U3426 (N_3426,N_3226,N_3105);
nand U3427 (N_3427,N_3175,N_3177);
and U3428 (N_3428,N_3165,N_3253);
xor U3429 (N_3429,N_3204,N_3111);
xor U3430 (N_3430,N_3079,N_3144);
or U3431 (N_3431,N_3161,N_3192);
and U3432 (N_3432,N_3261,N_3113);
nand U3433 (N_3433,N_3249,N_3086);
nor U3434 (N_3434,N_3212,N_3072);
nand U3435 (N_3435,N_3096,N_3056);
or U3436 (N_3436,N_3162,N_3043);
and U3437 (N_3437,N_3060,N_3151);
xor U3438 (N_3438,N_3143,N_3066);
nor U3439 (N_3439,N_3136,N_3279);
or U3440 (N_3440,N_3121,N_3299);
xor U3441 (N_3441,N_3138,N_3077);
nor U3442 (N_3442,N_3000,N_3194);
nor U3443 (N_3443,N_3147,N_3171);
and U3444 (N_3444,N_3284,N_3064);
nand U3445 (N_3445,N_3142,N_3222);
or U3446 (N_3446,N_3191,N_3116);
and U3447 (N_3447,N_3103,N_3021);
or U3448 (N_3448,N_3288,N_3282);
and U3449 (N_3449,N_3164,N_3183);
nand U3450 (N_3450,N_3027,N_3283);
or U3451 (N_3451,N_3171,N_3127);
xnor U3452 (N_3452,N_3284,N_3086);
nor U3453 (N_3453,N_3289,N_3206);
nand U3454 (N_3454,N_3094,N_3128);
nor U3455 (N_3455,N_3210,N_3183);
and U3456 (N_3456,N_3221,N_3186);
nand U3457 (N_3457,N_3053,N_3073);
nor U3458 (N_3458,N_3111,N_3029);
nor U3459 (N_3459,N_3268,N_3261);
or U3460 (N_3460,N_3049,N_3230);
nor U3461 (N_3461,N_3171,N_3043);
and U3462 (N_3462,N_3174,N_3289);
xor U3463 (N_3463,N_3283,N_3288);
nor U3464 (N_3464,N_3068,N_3221);
nor U3465 (N_3465,N_3207,N_3279);
and U3466 (N_3466,N_3273,N_3294);
xnor U3467 (N_3467,N_3283,N_3150);
xor U3468 (N_3468,N_3212,N_3046);
nand U3469 (N_3469,N_3022,N_3008);
or U3470 (N_3470,N_3196,N_3129);
and U3471 (N_3471,N_3038,N_3230);
nand U3472 (N_3472,N_3112,N_3248);
xnor U3473 (N_3473,N_3114,N_3242);
nand U3474 (N_3474,N_3241,N_3082);
or U3475 (N_3475,N_3020,N_3072);
xnor U3476 (N_3476,N_3172,N_3072);
and U3477 (N_3477,N_3103,N_3202);
and U3478 (N_3478,N_3031,N_3164);
nor U3479 (N_3479,N_3227,N_3058);
or U3480 (N_3480,N_3028,N_3198);
nand U3481 (N_3481,N_3287,N_3117);
and U3482 (N_3482,N_3201,N_3016);
and U3483 (N_3483,N_3084,N_3288);
and U3484 (N_3484,N_3099,N_3151);
nor U3485 (N_3485,N_3235,N_3190);
nor U3486 (N_3486,N_3252,N_3044);
nand U3487 (N_3487,N_3184,N_3283);
or U3488 (N_3488,N_3267,N_3167);
nor U3489 (N_3489,N_3225,N_3270);
nand U3490 (N_3490,N_3258,N_3040);
or U3491 (N_3491,N_3136,N_3173);
nor U3492 (N_3492,N_3267,N_3041);
xnor U3493 (N_3493,N_3123,N_3011);
or U3494 (N_3494,N_3143,N_3031);
xor U3495 (N_3495,N_3088,N_3110);
xnor U3496 (N_3496,N_3069,N_3010);
xnor U3497 (N_3497,N_3076,N_3253);
or U3498 (N_3498,N_3148,N_3160);
xor U3499 (N_3499,N_3279,N_3209);
xor U3500 (N_3500,N_3149,N_3096);
xnor U3501 (N_3501,N_3142,N_3111);
nand U3502 (N_3502,N_3251,N_3182);
xor U3503 (N_3503,N_3041,N_3000);
nor U3504 (N_3504,N_3147,N_3225);
and U3505 (N_3505,N_3252,N_3212);
nand U3506 (N_3506,N_3004,N_3128);
and U3507 (N_3507,N_3080,N_3116);
nor U3508 (N_3508,N_3084,N_3095);
and U3509 (N_3509,N_3258,N_3029);
nor U3510 (N_3510,N_3037,N_3094);
nor U3511 (N_3511,N_3171,N_3254);
nor U3512 (N_3512,N_3269,N_3277);
or U3513 (N_3513,N_3060,N_3184);
nor U3514 (N_3514,N_3071,N_3149);
or U3515 (N_3515,N_3275,N_3270);
nand U3516 (N_3516,N_3086,N_3220);
and U3517 (N_3517,N_3246,N_3101);
and U3518 (N_3518,N_3267,N_3116);
and U3519 (N_3519,N_3078,N_3233);
xnor U3520 (N_3520,N_3242,N_3071);
nand U3521 (N_3521,N_3035,N_3049);
xor U3522 (N_3522,N_3145,N_3136);
or U3523 (N_3523,N_3285,N_3108);
and U3524 (N_3524,N_3166,N_3277);
and U3525 (N_3525,N_3026,N_3189);
or U3526 (N_3526,N_3010,N_3018);
xor U3527 (N_3527,N_3230,N_3072);
nor U3528 (N_3528,N_3189,N_3109);
nand U3529 (N_3529,N_3065,N_3251);
xor U3530 (N_3530,N_3002,N_3053);
nor U3531 (N_3531,N_3151,N_3219);
nor U3532 (N_3532,N_3181,N_3058);
or U3533 (N_3533,N_3111,N_3152);
nand U3534 (N_3534,N_3139,N_3295);
xnor U3535 (N_3535,N_3255,N_3062);
or U3536 (N_3536,N_3226,N_3229);
xor U3537 (N_3537,N_3021,N_3185);
and U3538 (N_3538,N_3078,N_3237);
nand U3539 (N_3539,N_3225,N_3072);
xor U3540 (N_3540,N_3164,N_3253);
nand U3541 (N_3541,N_3075,N_3121);
or U3542 (N_3542,N_3090,N_3219);
nand U3543 (N_3543,N_3287,N_3190);
or U3544 (N_3544,N_3161,N_3186);
and U3545 (N_3545,N_3256,N_3263);
xnor U3546 (N_3546,N_3214,N_3181);
xnor U3547 (N_3547,N_3294,N_3102);
xnor U3548 (N_3548,N_3150,N_3203);
nor U3549 (N_3549,N_3211,N_3118);
nor U3550 (N_3550,N_3185,N_3032);
or U3551 (N_3551,N_3282,N_3270);
or U3552 (N_3552,N_3274,N_3047);
and U3553 (N_3553,N_3029,N_3247);
nand U3554 (N_3554,N_3108,N_3039);
and U3555 (N_3555,N_3218,N_3060);
and U3556 (N_3556,N_3221,N_3100);
xor U3557 (N_3557,N_3109,N_3285);
or U3558 (N_3558,N_3087,N_3049);
nand U3559 (N_3559,N_3196,N_3013);
nand U3560 (N_3560,N_3012,N_3292);
and U3561 (N_3561,N_3109,N_3098);
nand U3562 (N_3562,N_3227,N_3216);
or U3563 (N_3563,N_3106,N_3130);
nor U3564 (N_3564,N_3256,N_3042);
or U3565 (N_3565,N_3212,N_3026);
nor U3566 (N_3566,N_3153,N_3287);
nor U3567 (N_3567,N_3162,N_3087);
and U3568 (N_3568,N_3184,N_3073);
nor U3569 (N_3569,N_3017,N_3146);
and U3570 (N_3570,N_3172,N_3222);
nand U3571 (N_3571,N_3156,N_3290);
xnor U3572 (N_3572,N_3002,N_3045);
nor U3573 (N_3573,N_3079,N_3021);
nor U3574 (N_3574,N_3190,N_3018);
nand U3575 (N_3575,N_3061,N_3021);
nand U3576 (N_3576,N_3230,N_3214);
nor U3577 (N_3577,N_3299,N_3123);
nand U3578 (N_3578,N_3121,N_3066);
or U3579 (N_3579,N_3153,N_3020);
nand U3580 (N_3580,N_3070,N_3119);
and U3581 (N_3581,N_3058,N_3082);
or U3582 (N_3582,N_3103,N_3162);
and U3583 (N_3583,N_3092,N_3009);
nand U3584 (N_3584,N_3045,N_3145);
nor U3585 (N_3585,N_3173,N_3121);
and U3586 (N_3586,N_3040,N_3210);
xor U3587 (N_3587,N_3085,N_3023);
or U3588 (N_3588,N_3110,N_3112);
or U3589 (N_3589,N_3253,N_3213);
xor U3590 (N_3590,N_3039,N_3217);
xnor U3591 (N_3591,N_3280,N_3020);
and U3592 (N_3592,N_3144,N_3261);
xnor U3593 (N_3593,N_3145,N_3030);
nor U3594 (N_3594,N_3194,N_3185);
xnor U3595 (N_3595,N_3169,N_3131);
and U3596 (N_3596,N_3271,N_3102);
xnor U3597 (N_3597,N_3183,N_3013);
nand U3598 (N_3598,N_3078,N_3251);
or U3599 (N_3599,N_3036,N_3262);
nand U3600 (N_3600,N_3339,N_3559);
nand U3601 (N_3601,N_3372,N_3389);
nor U3602 (N_3602,N_3452,N_3497);
xnor U3603 (N_3603,N_3532,N_3522);
nand U3604 (N_3604,N_3549,N_3370);
and U3605 (N_3605,N_3561,N_3552);
nor U3606 (N_3606,N_3328,N_3547);
xor U3607 (N_3607,N_3446,N_3430);
nor U3608 (N_3608,N_3373,N_3584);
or U3609 (N_3609,N_3346,N_3324);
and U3610 (N_3610,N_3479,N_3423);
or U3611 (N_3611,N_3553,N_3465);
and U3612 (N_3612,N_3411,N_3344);
xor U3613 (N_3613,N_3428,N_3431);
and U3614 (N_3614,N_3494,N_3413);
or U3615 (N_3615,N_3379,N_3540);
or U3616 (N_3616,N_3571,N_3354);
and U3617 (N_3617,N_3315,N_3459);
or U3618 (N_3618,N_3486,N_3516);
or U3619 (N_3619,N_3581,N_3517);
and U3620 (N_3620,N_3595,N_3352);
nor U3621 (N_3621,N_3322,N_3503);
nand U3622 (N_3622,N_3310,N_3577);
and U3623 (N_3623,N_3371,N_3330);
nor U3624 (N_3624,N_3392,N_3468);
nand U3625 (N_3625,N_3591,N_3480);
nand U3626 (N_3626,N_3323,N_3524);
nand U3627 (N_3627,N_3526,N_3519);
and U3628 (N_3628,N_3491,N_3560);
or U3629 (N_3629,N_3576,N_3362);
or U3630 (N_3630,N_3343,N_3566);
or U3631 (N_3631,N_3306,N_3331);
nor U3632 (N_3632,N_3574,N_3329);
or U3633 (N_3633,N_3320,N_3550);
xor U3634 (N_3634,N_3409,N_3510);
nand U3635 (N_3635,N_3400,N_3347);
nor U3636 (N_3636,N_3304,N_3425);
nand U3637 (N_3637,N_3590,N_3583);
or U3638 (N_3638,N_3495,N_3449);
and U3639 (N_3639,N_3327,N_3496);
xnor U3640 (N_3640,N_3504,N_3333);
or U3641 (N_3641,N_3565,N_3312);
nor U3642 (N_3642,N_3437,N_3335);
nor U3643 (N_3643,N_3393,N_3403);
and U3644 (N_3644,N_3377,N_3490);
nor U3645 (N_3645,N_3300,N_3415);
nand U3646 (N_3646,N_3453,N_3585);
xnor U3647 (N_3647,N_3388,N_3301);
nand U3648 (N_3648,N_3457,N_3309);
nand U3649 (N_3649,N_3515,N_3391);
nor U3650 (N_3650,N_3355,N_3447);
nand U3651 (N_3651,N_3511,N_3325);
xor U3652 (N_3652,N_3341,N_3387);
nand U3653 (N_3653,N_3404,N_3464);
and U3654 (N_3654,N_3375,N_3338);
nor U3655 (N_3655,N_3458,N_3448);
nor U3656 (N_3656,N_3402,N_3365);
xnor U3657 (N_3657,N_3502,N_3390);
nand U3658 (N_3658,N_3472,N_3498);
or U3659 (N_3659,N_3462,N_3407);
xnor U3660 (N_3660,N_3442,N_3311);
or U3661 (N_3661,N_3363,N_3523);
nand U3662 (N_3662,N_3481,N_3454);
nor U3663 (N_3663,N_3527,N_3358);
nor U3664 (N_3664,N_3434,N_3353);
nor U3665 (N_3665,N_3420,N_3531);
nor U3666 (N_3666,N_3412,N_3460);
and U3667 (N_3667,N_3509,N_3314);
and U3668 (N_3668,N_3345,N_3483);
xor U3669 (N_3669,N_3334,N_3360);
and U3670 (N_3670,N_3512,N_3493);
and U3671 (N_3671,N_3432,N_3520);
xor U3672 (N_3672,N_3303,N_3421);
nor U3673 (N_3673,N_3544,N_3445);
nand U3674 (N_3674,N_3426,N_3588);
and U3675 (N_3675,N_3507,N_3348);
and U3676 (N_3676,N_3364,N_3416);
or U3677 (N_3677,N_3485,N_3313);
or U3678 (N_3678,N_3418,N_3538);
and U3679 (N_3679,N_3535,N_3518);
nor U3680 (N_3680,N_3349,N_3429);
and U3681 (N_3681,N_3487,N_3533);
nand U3682 (N_3682,N_3476,N_3427);
nor U3683 (N_3683,N_3405,N_3378);
and U3684 (N_3684,N_3546,N_3580);
or U3685 (N_3685,N_3489,N_3541);
nor U3686 (N_3686,N_3380,N_3488);
or U3687 (N_3687,N_3382,N_3567);
nand U3688 (N_3688,N_3451,N_3302);
nand U3689 (N_3689,N_3351,N_3384);
xnor U3690 (N_3690,N_3564,N_3484);
and U3691 (N_3691,N_3573,N_3381);
and U3692 (N_3692,N_3383,N_3319);
xor U3693 (N_3693,N_3529,N_3555);
nor U3694 (N_3694,N_3492,N_3593);
and U3695 (N_3695,N_3477,N_3395);
nand U3696 (N_3696,N_3435,N_3357);
nor U3697 (N_3697,N_3367,N_3337);
nor U3698 (N_3698,N_3436,N_3368);
or U3699 (N_3699,N_3386,N_3443);
nor U3700 (N_3700,N_3394,N_3305);
nand U3701 (N_3701,N_3525,N_3568);
nor U3702 (N_3702,N_3414,N_3422);
or U3703 (N_3703,N_3586,N_3599);
or U3704 (N_3704,N_3545,N_3572);
nand U3705 (N_3705,N_3398,N_3543);
or U3706 (N_3706,N_3506,N_3563);
or U3707 (N_3707,N_3321,N_3417);
nand U3708 (N_3708,N_3500,N_3406);
xnor U3709 (N_3709,N_3359,N_3508);
nand U3710 (N_3710,N_3408,N_3350);
xnor U3711 (N_3711,N_3557,N_3579);
and U3712 (N_3712,N_3307,N_3410);
or U3713 (N_3713,N_3318,N_3356);
nor U3714 (N_3714,N_3475,N_3528);
nand U3715 (N_3715,N_3374,N_3340);
xor U3716 (N_3716,N_3505,N_3551);
or U3717 (N_3717,N_3463,N_3433);
xnor U3718 (N_3718,N_3332,N_3537);
and U3719 (N_3719,N_3558,N_3562);
and U3720 (N_3720,N_3548,N_3385);
or U3721 (N_3721,N_3441,N_3456);
or U3722 (N_3722,N_3466,N_3569);
and U3723 (N_3723,N_3419,N_3575);
nand U3724 (N_3724,N_3317,N_3424);
nor U3725 (N_3725,N_3440,N_3396);
and U3726 (N_3726,N_3482,N_3342);
and U3727 (N_3727,N_3397,N_3450);
nand U3728 (N_3728,N_3594,N_3534);
and U3729 (N_3729,N_3514,N_3539);
and U3730 (N_3730,N_3474,N_3542);
nand U3731 (N_3731,N_3467,N_3316);
xnor U3732 (N_3732,N_3439,N_3455);
and U3733 (N_3733,N_3473,N_3471);
nor U3734 (N_3734,N_3596,N_3530);
nand U3735 (N_3735,N_3308,N_3578);
xnor U3736 (N_3736,N_3336,N_3587);
and U3737 (N_3737,N_3478,N_3589);
nor U3738 (N_3738,N_3366,N_3470);
and U3739 (N_3739,N_3399,N_3461);
xor U3740 (N_3740,N_3361,N_3582);
or U3741 (N_3741,N_3536,N_3592);
nand U3742 (N_3742,N_3376,N_3554);
xor U3743 (N_3743,N_3570,N_3444);
xor U3744 (N_3744,N_3369,N_3556);
or U3745 (N_3745,N_3469,N_3521);
xnor U3746 (N_3746,N_3513,N_3438);
or U3747 (N_3747,N_3326,N_3499);
and U3748 (N_3748,N_3597,N_3501);
nor U3749 (N_3749,N_3401,N_3598);
and U3750 (N_3750,N_3300,N_3587);
and U3751 (N_3751,N_3307,N_3300);
and U3752 (N_3752,N_3465,N_3586);
nor U3753 (N_3753,N_3344,N_3503);
or U3754 (N_3754,N_3392,N_3346);
nand U3755 (N_3755,N_3400,N_3324);
and U3756 (N_3756,N_3565,N_3442);
xnor U3757 (N_3757,N_3570,N_3384);
nand U3758 (N_3758,N_3440,N_3531);
nand U3759 (N_3759,N_3545,N_3341);
xnor U3760 (N_3760,N_3551,N_3336);
and U3761 (N_3761,N_3390,N_3486);
or U3762 (N_3762,N_3462,N_3532);
or U3763 (N_3763,N_3574,N_3475);
nor U3764 (N_3764,N_3554,N_3560);
and U3765 (N_3765,N_3431,N_3450);
or U3766 (N_3766,N_3450,N_3555);
nand U3767 (N_3767,N_3350,N_3558);
nor U3768 (N_3768,N_3380,N_3334);
xnor U3769 (N_3769,N_3454,N_3393);
nand U3770 (N_3770,N_3303,N_3389);
and U3771 (N_3771,N_3395,N_3535);
xor U3772 (N_3772,N_3354,N_3472);
xnor U3773 (N_3773,N_3384,N_3305);
and U3774 (N_3774,N_3525,N_3588);
or U3775 (N_3775,N_3401,N_3544);
nor U3776 (N_3776,N_3535,N_3456);
or U3777 (N_3777,N_3308,N_3304);
nand U3778 (N_3778,N_3327,N_3462);
nand U3779 (N_3779,N_3440,N_3318);
and U3780 (N_3780,N_3570,N_3303);
xor U3781 (N_3781,N_3307,N_3509);
and U3782 (N_3782,N_3411,N_3546);
and U3783 (N_3783,N_3555,N_3383);
and U3784 (N_3784,N_3536,N_3302);
or U3785 (N_3785,N_3373,N_3451);
xor U3786 (N_3786,N_3480,N_3477);
nor U3787 (N_3787,N_3596,N_3533);
xor U3788 (N_3788,N_3337,N_3424);
and U3789 (N_3789,N_3407,N_3488);
nand U3790 (N_3790,N_3359,N_3589);
xnor U3791 (N_3791,N_3388,N_3310);
xnor U3792 (N_3792,N_3597,N_3506);
nor U3793 (N_3793,N_3495,N_3574);
xnor U3794 (N_3794,N_3472,N_3336);
or U3795 (N_3795,N_3544,N_3475);
nand U3796 (N_3796,N_3360,N_3321);
and U3797 (N_3797,N_3336,N_3554);
nor U3798 (N_3798,N_3420,N_3515);
and U3799 (N_3799,N_3514,N_3366);
and U3800 (N_3800,N_3367,N_3366);
nor U3801 (N_3801,N_3449,N_3373);
nor U3802 (N_3802,N_3518,N_3348);
nand U3803 (N_3803,N_3583,N_3584);
nand U3804 (N_3804,N_3564,N_3346);
nor U3805 (N_3805,N_3539,N_3374);
and U3806 (N_3806,N_3318,N_3497);
or U3807 (N_3807,N_3361,N_3463);
and U3808 (N_3808,N_3462,N_3451);
and U3809 (N_3809,N_3487,N_3420);
xnor U3810 (N_3810,N_3418,N_3320);
nand U3811 (N_3811,N_3374,N_3587);
and U3812 (N_3812,N_3316,N_3433);
and U3813 (N_3813,N_3583,N_3471);
or U3814 (N_3814,N_3399,N_3540);
nor U3815 (N_3815,N_3364,N_3301);
xor U3816 (N_3816,N_3354,N_3466);
and U3817 (N_3817,N_3547,N_3511);
xnor U3818 (N_3818,N_3408,N_3485);
nand U3819 (N_3819,N_3424,N_3591);
and U3820 (N_3820,N_3323,N_3392);
or U3821 (N_3821,N_3561,N_3365);
nand U3822 (N_3822,N_3468,N_3576);
and U3823 (N_3823,N_3528,N_3364);
nor U3824 (N_3824,N_3323,N_3463);
xor U3825 (N_3825,N_3542,N_3490);
or U3826 (N_3826,N_3463,N_3362);
or U3827 (N_3827,N_3413,N_3329);
nand U3828 (N_3828,N_3466,N_3572);
or U3829 (N_3829,N_3379,N_3440);
nand U3830 (N_3830,N_3322,N_3349);
xor U3831 (N_3831,N_3389,N_3411);
xor U3832 (N_3832,N_3341,N_3563);
or U3833 (N_3833,N_3528,N_3418);
and U3834 (N_3834,N_3463,N_3375);
and U3835 (N_3835,N_3499,N_3480);
xnor U3836 (N_3836,N_3564,N_3523);
and U3837 (N_3837,N_3556,N_3399);
or U3838 (N_3838,N_3411,N_3578);
or U3839 (N_3839,N_3442,N_3384);
nor U3840 (N_3840,N_3381,N_3375);
and U3841 (N_3841,N_3500,N_3314);
or U3842 (N_3842,N_3316,N_3379);
xnor U3843 (N_3843,N_3485,N_3376);
or U3844 (N_3844,N_3525,N_3427);
and U3845 (N_3845,N_3574,N_3448);
and U3846 (N_3846,N_3305,N_3457);
xnor U3847 (N_3847,N_3340,N_3442);
nand U3848 (N_3848,N_3392,N_3345);
nor U3849 (N_3849,N_3598,N_3443);
and U3850 (N_3850,N_3423,N_3321);
and U3851 (N_3851,N_3317,N_3407);
or U3852 (N_3852,N_3383,N_3317);
or U3853 (N_3853,N_3417,N_3594);
or U3854 (N_3854,N_3310,N_3484);
xnor U3855 (N_3855,N_3536,N_3501);
nor U3856 (N_3856,N_3478,N_3305);
xor U3857 (N_3857,N_3373,N_3500);
xnor U3858 (N_3858,N_3342,N_3436);
xor U3859 (N_3859,N_3419,N_3514);
and U3860 (N_3860,N_3552,N_3382);
and U3861 (N_3861,N_3570,N_3544);
or U3862 (N_3862,N_3598,N_3575);
nor U3863 (N_3863,N_3422,N_3541);
xnor U3864 (N_3864,N_3454,N_3582);
or U3865 (N_3865,N_3543,N_3304);
and U3866 (N_3866,N_3578,N_3429);
or U3867 (N_3867,N_3440,N_3316);
xnor U3868 (N_3868,N_3590,N_3587);
and U3869 (N_3869,N_3321,N_3554);
nor U3870 (N_3870,N_3339,N_3412);
or U3871 (N_3871,N_3345,N_3384);
or U3872 (N_3872,N_3450,N_3599);
xor U3873 (N_3873,N_3458,N_3472);
nand U3874 (N_3874,N_3452,N_3374);
or U3875 (N_3875,N_3471,N_3362);
xnor U3876 (N_3876,N_3523,N_3356);
nor U3877 (N_3877,N_3501,N_3322);
nand U3878 (N_3878,N_3475,N_3505);
nand U3879 (N_3879,N_3388,N_3326);
or U3880 (N_3880,N_3550,N_3371);
nor U3881 (N_3881,N_3526,N_3482);
and U3882 (N_3882,N_3431,N_3553);
and U3883 (N_3883,N_3542,N_3401);
or U3884 (N_3884,N_3467,N_3461);
or U3885 (N_3885,N_3584,N_3485);
or U3886 (N_3886,N_3388,N_3596);
nand U3887 (N_3887,N_3553,N_3504);
or U3888 (N_3888,N_3417,N_3514);
nand U3889 (N_3889,N_3494,N_3300);
xor U3890 (N_3890,N_3574,N_3490);
and U3891 (N_3891,N_3528,N_3371);
or U3892 (N_3892,N_3430,N_3589);
or U3893 (N_3893,N_3342,N_3388);
nand U3894 (N_3894,N_3550,N_3402);
xnor U3895 (N_3895,N_3492,N_3552);
xnor U3896 (N_3896,N_3520,N_3554);
nor U3897 (N_3897,N_3388,N_3469);
xor U3898 (N_3898,N_3359,N_3326);
nand U3899 (N_3899,N_3509,N_3500);
xor U3900 (N_3900,N_3650,N_3798);
and U3901 (N_3901,N_3723,N_3787);
nand U3902 (N_3902,N_3858,N_3608);
or U3903 (N_3903,N_3744,N_3857);
xor U3904 (N_3904,N_3852,N_3739);
and U3905 (N_3905,N_3878,N_3618);
and U3906 (N_3906,N_3621,N_3745);
nor U3907 (N_3907,N_3772,N_3773);
or U3908 (N_3908,N_3642,N_3888);
or U3909 (N_3909,N_3721,N_3889);
nand U3910 (N_3910,N_3755,N_3818);
xor U3911 (N_3911,N_3761,N_3716);
nand U3912 (N_3912,N_3705,N_3623);
nand U3913 (N_3913,N_3733,N_3769);
or U3914 (N_3914,N_3704,N_3720);
nand U3915 (N_3915,N_3838,N_3826);
nor U3916 (N_3916,N_3861,N_3811);
xor U3917 (N_3917,N_3795,N_3614);
or U3918 (N_3918,N_3688,N_3833);
or U3919 (N_3919,N_3625,N_3758);
xnor U3920 (N_3920,N_3805,N_3725);
and U3921 (N_3921,N_3699,N_3813);
xnor U3922 (N_3922,N_3868,N_3724);
xor U3923 (N_3923,N_3710,N_3830);
nand U3924 (N_3924,N_3604,N_3763);
nor U3925 (N_3925,N_3771,N_3749);
xor U3926 (N_3926,N_3702,N_3680);
nand U3927 (N_3927,N_3631,N_3675);
or U3928 (N_3928,N_3844,N_3767);
and U3929 (N_3929,N_3689,N_3788);
nor U3930 (N_3930,N_3896,N_3753);
nand U3931 (N_3931,N_3863,N_3692);
and U3932 (N_3932,N_3867,N_3655);
xnor U3933 (N_3933,N_3683,N_3869);
nor U3934 (N_3934,N_3780,N_3803);
or U3935 (N_3935,N_3652,N_3762);
xor U3936 (N_3936,N_3827,N_3862);
xor U3937 (N_3937,N_3777,N_3801);
nand U3938 (N_3938,N_3624,N_3898);
nor U3939 (N_3939,N_3842,N_3690);
xor U3940 (N_3940,N_3809,N_3885);
and U3941 (N_3941,N_3620,N_3600);
or U3942 (N_3942,N_3845,N_3674);
nor U3943 (N_3943,N_3843,N_3782);
nor U3944 (N_3944,N_3866,N_3684);
and U3945 (N_3945,N_3816,N_3626);
nand U3946 (N_3946,N_3606,N_3848);
nand U3947 (N_3947,N_3627,N_3828);
or U3948 (N_3948,N_3815,N_3776);
nand U3949 (N_3949,N_3884,N_3865);
xor U3950 (N_3950,N_3644,N_3778);
nand U3951 (N_3951,N_3685,N_3601);
nor U3952 (N_3952,N_3647,N_3797);
or U3953 (N_3953,N_3832,N_3645);
and U3954 (N_3954,N_3874,N_3810);
xnor U3955 (N_3955,N_3817,N_3636);
xor U3956 (N_3956,N_3668,N_3659);
nor U3957 (N_3957,N_3876,N_3808);
nor U3958 (N_3958,N_3719,N_3611);
nor U3959 (N_3959,N_3728,N_3766);
nand U3960 (N_3960,N_3839,N_3836);
nor U3961 (N_3961,N_3617,N_3629);
nand U3962 (N_3962,N_3887,N_3882);
or U3963 (N_3963,N_3717,N_3691);
nor U3964 (N_3964,N_3612,N_3737);
xnor U3965 (N_3965,N_3754,N_3694);
xor U3966 (N_3966,N_3605,N_3660);
nor U3967 (N_3967,N_3651,N_3802);
xor U3968 (N_3968,N_3610,N_3697);
nand U3969 (N_3969,N_3854,N_3709);
and U3970 (N_3970,N_3841,N_3784);
and U3971 (N_3971,N_3678,N_3873);
nor U3972 (N_3972,N_3708,N_3757);
nand U3973 (N_3973,N_3639,N_3853);
xor U3974 (N_3974,N_3894,N_3768);
or U3975 (N_3975,N_3892,N_3875);
nor U3976 (N_3976,N_3791,N_3883);
nor U3977 (N_3977,N_3738,N_3796);
or U3978 (N_3978,N_3880,N_3657);
xnor U3979 (N_3979,N_3695,N_3871);
nand U3980 (N_3980,N_3664,N_3877);
and U3981 (N_3981,N_3609,N_3829);
and U3982 (N_3982,N_3872,N_3638);
nand U3983 (N_3983,N_3712,N_3756);
xnor U3984 (N_3984,N_3670,N_3646);
xnor U3985 (N_3985,N_3822,N_3648);
nand U3986 (N_3986,N_3726,N_3669);
xnor U3987 (N_3987,N_3732,N_3673);
xnor U3988 (N_3988,N_3825,N_3814);
xor U3989 (N_3989,N_3835,N_3748);
nand U3990 (N_3990,N_3603,N_3682);
nand U3991 (N_3991,N_3775,N_3635);
and U3992 (N_3992,N_3654,N_3734);
nor U3993 (N_3993,N_3794,N_3790);
nand U3994 (N_3994,N_3886,N_3718);
and U3995 (N_3995,N_3715,N_3711);
nor U3996 (N_3996,N_3633,N_3849);
nand U3997 (N_3997,N_3831,N_3607);
and U3998 (N_3998,N_3698,N_3851);
or U3999 (N_3999,N_3740,N_3731);
or U4000 (N_4000,N_3703,N_3727);
nand U4001 (N_4001,N_3779,N_3759);
xor U4002 (N_4002,N_3730,N_3671);
xnor U4003 (N_4003,N_3895,N_3837);
xnor U4004 (N_4004,N_3634,N_3856);
nor U4005 (N_4005,N_3806,N_3824);
and U4006 (N_4006,N_3879,N_3804);
or U4007 (N_4007,N_3774,N_3765);
or U4008 (N_4008,N_3742,N_3860);
or U4009 (N_4009,N_3707,N_3665);
xnor U4010 (N_4010,N_3679,N_3864);
or U4011 (N_4011,N_3820,N_3736);
or U4012 (N_4012,N_3750,N_3653);
or U4013 (N_4013,N_3812,N_3819);
or U4014 (N_4014,N_3602,N_3619);
xor U4015 (N_4015,N_3722,N_3677);
nand U4016 (N_4016,N_3799,N_3643);
nor U4017 (N_4017,N_3785,N_3800);
nor U4018 (N_4018,N_3899,N_3713);
nand U4019 (N_4019,N_3667,N_3847);
or U4020 (N_4020,N_3821,N_3890);
nand U4021 (N_4021,N_3700,N_3741);
or U4022 (N_4022,N_3714,N_3628);
nand U4023 (N_4023,N_3613,N_3686);
or U4024 (N_4024,N_3662,N_3792);
and U4025 (N_4025,N_3630,N_3615);
or U4026 (N_4026,N_3786,N_3747);
nor U4027 (N_4027,N_3893,N_3656);
or U4028 (N_4028,N_3770,N_3746);
xor U4029 (N_4029,N_3706,N_3632);
nand U4030 (N_4030,N_3793,N_3676);
nand U4031 (N_4031,N_3696,N_3640);
xnor U4032 (N_4032,N_3840,N_3616);
nand U4033 (N_4033,N_3687,N_3823);
xor U4034 (N_4034,N_3752,N_3649);
xnor U4035 (N_4035,N_3751,N_3870);
xnor U4036 (N_4036,N_3672,N_3760);
and U4037 (N_4037,N_3681,N_3855);
and U4038 (N_4038,N_3658,N_3789);
xnor U4039 (N_4039,N_3897,N_3743);
nand U4040 (N_4040,N_3783,N_3859);
or U4041 (N_4041,N_3661,N_3701);
nor U4042 (N_4042,N_3846,N_3881);
or U4043 (N_4043,N_3622,N_3637);
nand U4044 (N_4044,N_3834,N_3807);
nor U4045 (N_4045,N_3729,N_3693);
or U4046 (N_4046,N_3641,N_3891);
xor U4047 (N_4047,N_3663,N_3735);
nand U4048 (N_4048,N_3666,N_3764);
xnor U4049 (N_4049,N_3850,N_3781);
nand U4050 (N_4050,N_3885,N_3840);
and U4051 (N_4051,N_3690,N_3837);
nor U4052 (N_4052,N_3869,N_3815);
and U4053 (N_4053,N_3620,N_3681);
nor U4054 (N_4054,N_3726,N_3635);
xor U4055 (N_4055,N_3894,N_3864);
nor U4056 (N_4056,N_3897,N_3733);
and U4057 (N_4057,N_3816,N_3717);
nor U4058 (N_4058,N_3723,N_3834);
xor U4059 (N_4059,N_3794,N_3884);
nor U4060 (N_4060,N_3748,N_3750);
nand U4061 (N_4061,N_3881,N_3869);
or U4062 (N_4062,N_3810,N_3665);
nor U4063 (N_4063,N_3819,N_3813);
or U4064 (N_4064,N_3728,N_3761);
nand U4065 (N_4065,N_3714,N_3755);
nor U4066 (N_4066,N_3769,N_3862);
or U4067 (N_4067,N_3758,N_3708);
nand U4068 (N_4068,N_3881,N_3873);
xor U4069 (N_4069,N_3627,N_3746);
or U4070 (N_4070,N_3833,N_3704);
and U4071 (N_4071,N_3842,N_3887);
nor U4072 (N_4072,N_3676,N_3736);
and U4073 (N_4073,N_3886,N_3863);
xnor U4074 (N_4074,N_3712,N_3883);
or U4075 (N_4075,N_3646,N_3610);
and U4076 (N_4076,N_3747,N_3691);
and U4077 (N_4077,N_3723,N_3785);
and U4078 (N_4078,N_3858,N_3829);
xnor U4079 (N_4079,N_3870,N_3775);
nand U4080 (N_4080,N_3791,N_3613);
xnor U4081 (N_4081,N_3695,N_3658);
nor U4082 (N_4082,N_3675,N_3822);
or U4083 (N_4083,N_3783,N_3786);
or U4084 (N_4084,N_3886,N_3741);
and U4085 (N_4085,N_3604,N_3813);
nor U4086 (N_4086,N_3815,N_3714);
nor U4087 (N_4087,N_3712,N_3784);
nand U4088 (N_4088,N_3619,N_3622);
nand U4089 (N_4089,N_3888,N_3871);
nand U4090 (N_4090,N_3622,N_3835);
nand U4091 (N_4091,N_3646,N_3621);
nor U4092 (N_4092,N_3721,N_3604);
xor U4093 (N_4093,N_3703,N_3685);
xor U4094 (N_4094,N_3624,N_3699);
nand U4095 (N_4095,N_3632,N_3875);
and U4096 (N_4096,N_3628,N_3715);
and U4097 (N_4097,N_3899,N_3806);
xor U4098 (N_4098,N_3780,N_3664);
or U4099 (N_4099,N_3697,N_3846);
and U4100 (N_4100,N_3801,N_3871);
nand U4101 (N_4101,N_3760,N_3870);
nor U4102 (N_4102,N_3856,N_3675);
xor U4103 (N_4103,N_3852,N_3825);
nor U4104 (N_4104,N_3705,N_3600);
nand U4105 (N_4105,N_3676,N_3773);
nand U4106 (N_4106,N_3821,N_3664);
or U4107 (N_4107,N_3849,N_3832);
or U4108 (N_4108,N_3778,N_3663);
nor U4109 (N_4109,N_3822,N_3715);
and U4110 (N_4110,N_3895,N_3827);
nor U4111 (N_4111,N_3604,N_3713);
nand U4112 (N_4112,N_3761,N_3738);
xnor U4113 (N_4113,N_3617,N_3662);
nor U4114 (N_4114,N_3615,N_3890);
nand U4115 (N_4115,N_3640,N_3869);
nand U4116 (N_4116,N_3621,N_3812);
or U4117 (N_4117,N_3663,N_3690);
and U4118 (N_4118,N_3771,N_3871);
and U4119 (N_4119,N_3814,N_3746);
and U4120 (N_4120,N_3686,N_3701);
and U4121 (N_4121,N_3740,N_3774);
xnor U4122 (N_4122,N_3813,N_3791);
or U4123 (N_4123,N_3887,N_3719);
and U4124 (N_4124,N_3659,N_3812);
or U4125 (N_4125,N_3742,N_3780);
nor U4126 (N_4126,N_3609,N_3806);
and U4127 (N_4127,N_3840,N_3631);
nor U4128 (N_4128,N_3754,N_3791);
xor U4129 (N_4129,N_3676,N_3696);
and U4130 (N_4130,N_3887,N_3881);
or U4131 (N_4131,N_3779,N_3787);
and U4132 (N_4132,N_3659,N_3736);
nand U4133 (N_4133,N_3761,N_3890);
and U4134 (N_4134,N_3636,N_3757);
nand U4135 (N_4135,N_3657,N_3640);
nand U4136 (N_4136,N_3898,N_3710);
and U4137 (N_4137,N_3719,N_3737);
nor U4138 (N_4138,N_3884,N_3737);
or U4139 (N_4139,N_3730,N_3850);
nand U4140 (N_4140,N_3729,N_3715);
nor U4141 (N_4141,N_3636,N_3659);
xnor U4142 (N_4142,N_3771,N_3716);
and U4143 (N_4143,N_3622,N_3828);
or U4144 (N_4144,N_3840,N_3625);
xor U4145 (N_4145,N_3785,N_3612);
or U4146 (N_4146,N_3874,N_3702);
nand U4147 (N_4147,N_3708,N_3848);
nor U4148 (N_4148,N_3617,N_3893);
nor U4149 (N_4149,N_3806,N_3603);
and U4150 (N_4150,N_3699,N_3785);
nor U4151 (N_4151,N_3878,N_3667);
nand U4152 (N_4152,N_3815,N_3861);
and U4153 (N_4153,N_3762,N_3721);
xor U4154 (N_4154,N_3652,N_3824);
and U4155 (N_4155,N_3835,N_3644);
nand U4156 (N_4156,N_3820,N_3840);
xnor U4157 (N_4157,N_3717,N_3685);
nand U4158 (N_4158,N_3760,N_3605);
nor U4159 (N_4159,N_3652,N_3849);
or U4160 (N_4160,N_3805,N_3728);
xnor U4161 (N_4161,N_3846,N_3691);
xor U4162 (N_4162,N_3764,N_3830);
or U4163 (N_4163,N_3831,N_3624);
and U4164 (N_4164,N_3633,N_3812);
nor U4165 (N_4165,N_3828,N_3709);
nand U4166 (N_4166,N_3723,N_3745);
nand U4167 (N_4167,N_3766,N_3794);
nand U4168 (N_4168,N_3762,N_3675);
or U4169 (N_4169,N_3723,N_3891);
nand U4170 (N_4170,N_3724,N_3715);
or U4171 (N_4171,N_3872,N_3850);
nand U4172 (N_4172,N_3730,N_3748);
or U4173 (N_4173,N_3817,N_3887);
nand U4174 (N_4174,N_3699,N_3700);
or U4175 (N_4175,N_3893,N_3687);
and U4176 (N_4176,N_3618,N_3755);
or U4177 (N_4177,N_3731,N_3693);
xnor U4178 (N_4178,N_3624,N_3709);
nand U4179 (N_4179,N_3640,N_3639);
nand U4180 (N_4180,N_3887,N_3814);
xor U4181 (N_4181,N_3634,N_3718);
nand U4182 (N_4182,N_3681,N_3835);
nand U4183 (N_4183,N_3890,N_3893);
xor U4184 (N_4184,N_3838,N_3699);
nand U4185 (N_4185,N_3849,N_3778);
nor U4186 (N_4186,N_3827,N_3838);
xnor U4187 (N_4187,N_3712,N_3789);
or U4188 (N_4188,N_3684,N_3638);
xnor U4189 (N_4189,N_3751,N_3806);
nand U4190 (N_4190,N_3711,N_3785);
or U4191 (N_4191,N_3760,N_3888);
nand U4192 (N_4192,N_3830,N_3658);
xnor U4193 (N_4193,N_3649,N_3792);
nor U4194 (N_4194,N_3875,N_3729);
or U4195 (N_4195,N_3704,N_3621);
and U4196 (N_4196,N_3805,N_3851);
xor U4197 (N_4197,N_3668,N_3827);
nand U4198 (N_4198,N_3885,N_3671);
and U4199 (N_4199,N_3741,N_3815);
nand U4200 (N_4200,N_4114,N_4146);
and U4201 (N_4201,N_4019,N_3992);
xor U4202 (N_4202,N_4142,N_3996);
nand U4203 (N_4203,N_4123,N_4075);
and U4204 (N_4204,N_4120,N_4002);
nor U4205 (N_4205,N_4101,N_3990);
xnor U4206 (N_4206,N_4148,N_3911);
nor U4207 (N_4207,N_4097,N_3970);
nand U4208 (N_4208,N_4087,N_4004);
nor U4209 (N_4209,N_4069,N_3901);
nor U4210 (N_4210,N_4168,N_4041);
and U4211 (N_4211,N_4195,N_4180);
or U4212 (N_4212,N_4115,N_4045);
nand U4213 (N_4213,N_4196,N_3931);
nor U4214 (N_4214,N_4086,N_3977);
nor U4215 (N_4215,N_3966,N_3985);
or U4216 (N_4216,N_3935,N_4162);
xor U4217 (N_4217,N_4178,N_4031);
or U4218 (N_4218,N_3971,N_3917);
xor U4219 (N_4219,N_4159,N_4014);
xnor U4220 (N_4220,N_4003,N_4105);
xor U4221 (N_4221,N_4192,N_4116);
or U4222 (N_4222,N_4053,N_3995);
and U4223 (N_4223,N_4155,N_4052);
nand U4224 (N_4224,N_4156,N_4108);
and U4225 (N_4225,N_4026,N_3941);
xnor U4226 (N_4226,N_4141,N_4076);
nor U4227 (N_4227,N_3979,N_4030);
nand U4228 (N_4228,N_3900,N_3948);
and U4229 (N_4229,N_3957,N_3950);
or U4230 (N_4230,N_4175,N_4079);
xnor U4231 (N_4231,N_3905,N_4193);
and U4232 (N_4232,N_4138,N_4092);
and U4233 (N_4233,N_4073,N_3997);
or U4234 (N_4234,N_4006,N_4048);
nor U4235 (N_4235,N_3933,N_3936);
nor U4236 (N_4236,N_3923,N_4085);
xnor U4237 (N_4237,N_4157,N_4022);
nor U4238 (N_4238,N_4181,N_4100);
or U4239 (N_4239,N_3910,N_4040);
nor U4240 (N_4240,N_4043,N_4152);
xnor U4241 (N_4241,N_4096,N_3953);
xnor U4242 (N_4242,N_4128,N_4130);
nor U4243 (N_4243,N_4169,N_4182);
nand U4244 (N_4244,N_4125,N_3945);
and U4245 (N_4245,N_4074,N_4027);
xnor U4246 (N_4246,N_4067,N_4140);
nand U4247 (N_4247,N_3903,N_4112);
nand U4248 (N_4248,N_3959,N_4005);
xnor U4249 (N_4249,N_3969,N_3934);
nand U4250 (N_4250,N_4088,N_3943);
or U4251 (N_4251,N_4176,N_3989);
or U4252 (N_4252,N_3968,N_4197);
or U4253 (N_4253,N_4017,N_4143);
nand U4254 (N_4254,N_4185,N_3922);
and U4255 (N_4255,N_3956,N_4190);
nor U4256 (N_4256,N_4135,N_3906);
and U4257 (N_4257,N_4084,N_4110);
xnor U4258 (N_4258,N_4124,N_4150);
xnor U4259 (N_4259,N_4051,N_4117);
and U4260 (N_4260,N_4012,N_3920);
or U4261 (N_4261,N_4153,N_4059);
nand U4262 (N_4262,N_3904,N_4072);
or U4263 (N_4263,N_4145,N_4177);
nor U4264 (N_4264,N_3926,N_3967);
nand U4265 (N_4265,N_4095,N_4165);
or U4266 (N_4266,N_3998,N_4009);
or U4267 (N_4267,N_4093,N_4136);
nand U4268 (N_4268,N_3980,N_4071);
nor U4269 (N_4269,N_4010,N_4047);
or U4270 (N_4270,N_4164,N_3958);
xor U4271 (N_4271,N_4050,N_4122);
xnor U4272 (N_4272,N_4023,N_3938);
and U4273 (N_4273,N_3973,N_4166);
nor U4274 (N_4274,N_4194,N_4104);
nand U4275 (N_4275,N_3984,N_4144);
or U4276 (N_4276,N_4066,N_3913);
nor U4277 (N_4277,N_4151,N_4083);
xor U4278 (N_4278,N_3949,N_4107);
xnor U4279 (N_4279,N_4060,N_4080);
and U4280 (N_4280,N_3991,N_4139);
nor U4281 (N_4281,N_4063,N_4163);
xor U4282 (N_4282,N_3932,N_4106);
or U4283 (N_4283,N_4111,N_3919);
nand U4284 (N_4284,N_4013,N_4029);
nand U4285 (N_4285,N_3981,N_4173);
xnor U4286 (N_4286,N_4154,N_4158);
nand U4287 (N_4287,N_3975,N_4054);
or U4288 (N_4288,N_4077,N_3921);
xor U4289 (N_4289,N_3915,N_3940);
xor U4290 (N_4290,N_4046,N_4131);
nor U4291 (N_4291,N_4068,N_4134);
or U4292 (N_4292,N_4149,N_4109);
or U4293 (N_4293,N_4036,N_4078);
nand U4294 (N_4294,N_3982,N_4191);
xor U4295 (N_4295,N_3965,N_4170);
or U4296 (N_4296,N_4121,N_3929);
nor U4297 (N_4297,N_4189,N_3952);
nand U4298 (N_4298,N_3947,N_4113);
nor U4299 (N_4299,N_4147,N_3994);
nor U4300 (N_4300,N_3962,N_4021);
or U4301 (N_4301,N_3978,N_4184);
nand U4302 (N_4302,N_3964,N_4160);
and U4303 (N_4303,N_4055,N_4000);
nor U4304 (N_4304,N_4016,N_4133);
or U4305 (N_4305,N_4061,N_4082);
and U4306 (N_4306,N_4118,N_3944);
nor U4307 (N_4307,N_4057,N_3927);
nor U4308 (N_4308,N_3908,N_3916);
nand U4309 (N_4309,N_4044,N_3983);
or U4310 (N_4310,N_4042,N_4167);
nor U4311 (N_4311,N_3955,N_4037);
or U4312 (N_4312,N_4119,N_4102);
and U4313 (N_4313,N_3960,N_3914);
or U4314 (N_4314,N_4174,N_3902);
and U4315 (N_4315,N_4161,N_4094);
xnor U4316 (N_4316,N_3918,N_4001);
nand U4317 (N_4317,N_4187,N_4033);
and U4318 (N_4318,N_4015,N_4081);
nor U4319 (N_4319,N_4098,N_3928);
and U4320 (N_4320,N_4198,N_4132);
nor U4321 (N_4321,N_3987,N_4039);
or U4322 (N_4322,N_4199,N_4056);
or U4323 (N_4323,N_4058,N_3912);
nor U4324 (N_4324,N_3999,N_4018);
xnor U4325 (N_4325,N_3963,N_4090);
nor U4326 (N_4326,N_3986,N_4011);
xor U4327 (N_4327,N_3954,N_3976);
or U4328 (N_4328,N_4129,N_4183);
or U4329 (N_4329,N_3946,N_4137);
nor U4330 (N_4330,N_4008,N_4091);
or U4331 (N_4331,N_4049,N_4028);
nor U4332 (N_4332,N_3937,N_4032);
nor U4333 (N_4333,N_4064,N_3930);
and U4334 (N_4334,N_4035,N_4186);
nor U4335 (N_4335,N_4065,N_3942);
xnor U4336 (N_4336,N_4062,N_3909);
xor U4337 (N_4337,N_4179,N_4127);
xnor U4338 (N_4338,N_3951,N_3907);
xor U4339 (N_4339,N_3925,N_4089);
nand U4340 (N_4340,N_3961,N_3988);
and U4341 (N_4341,N_3939,N_4024);
and U4342 (N_4342,N_3924,N_4007);
and U4343 (N_4343,N_4025,N_4099);
nand U4344 (N_4344,N_3993,N_4034);
or U4345 (N_4345,N_4103,N_3972);
xor U4346 (N_4346,N_3974,N_4188);
and U4347 (N_4347,N_4171,N_4172);
and U4348 (N_4348,N_4020,N_4038);
nor U4349 (N_4349,N_4126,N_4070);
nand U4350 (N_4350,N_4107,N_4056);
nor U4351 (N_4351,N_4013,N_3985);
xnor U4352 (N_4352,N_4074,N_3982);
or U4353 (N_4353,N_4092,N_4067);
and U4354 (N_4354,N_3995,N_3976);
nand U4355 (N_4355,N_4171,N_4117);
nor U4356 (N_4356,N_4086,N_4029);
nor U4357 (N_4357,N_4080,N_3989);
xnor U4358 (N_4358,N_3971,N_4035);
xnor U4359 (N_4359,N_3912,N_3911);
and U4360 (N_4360,N_3960,N_3910);
and U4361 (N_4361,N_4155,N_4056);
nor U4362 (N_4362,N_4189,N_4180);
or U4363 (N_4363,N_4127,N_3946);
nor U4364 (N_4364,N_4109,N_3995);
nand U4365 (N_4365,N_3919,N_4103);
or U4366 (N_4366,N_3961,N_4052);
and U4367 (N_4367,N_3915,N_4150);
xnor U4368 (N_4368,N_3916,N_3920);
nand U4369 (N_4369,N_3930,N_4029);
xnor U4370 (N_4370,N_3964,N_4137);
or U4371 (N_4371,N_4140,N_4059);
nor U4372 (N_4372,N_4174,N_4053);
or U4373 (N_4373,N_4134,N_3944);
or U4374 (N_4374,N_3943,N_4055);
nand U4375 (N_4375,N_3965,N_3920);
nand U4376 (N_4376,N_4043,N_4101);
xor U4377 (N_4377,N_4183,N_4098);
and U4378 (N_4378,N_4182,N_4149);
xor U4379 (N_4379,N_4055,N_3979);
and U4380 (N_4380,N_3917,N_3927);
xnor U4381 (N_4381,N_3927,N_4005);
or U4382 (N_4382,N_3924,N_3917);
xor U4383 (N_4383,N_4052,N_4024);
nor U4384 (N_4384,N_4133,N_3990);
nor U4385 (N_4385,N_4017,N_4146);
nor U4386 (N_4386,N_4180,N_4013);
nand U4387 (N_4387,N_3990,N_3983);
nor U4388 (N_4388,N_4173,N_4134);
xor U4389 (N_4389,N_4072,N_4006);
nand U4390 (N_4390,N_4015,N_3994);
nand U4391 (N_4391,N_4099,N_3923);
and U4392 (N_4392,N_3978,N_4032);
nand U4393 (N_4393,N_3908,N_4005);
nor U4394 (N_4394,N_4198,N_4163);
nand U4395 (N_4395,N_3960,N_4013);
or U4396 (N_4396,N_4047,N_4046);
xnor U4397 (N_4397,N_4193,N_4028);
or U4398 (N_4398,N_4165,N_3933);
or U4399 (N_4399,N_4067,N_3960);
xnor U4400 (N_4400,N_4115,N_4030);
xnor U4401 (N_4401,N_4131,N_4019);
nand U4402 (N_4402,N_3928,N_3961);
and U4403 (N_4403,N_4014,N_3917);
nand U4404 (N_4404,N_3904,N_4108);
or U4405 (N_4405,N_4121,N_4181);
and U4406 (N_4406,N_4055,N_4163);
xor U4407 (N_4407,N_3999,N_3939);
and U4408 (N_4408,N_3927,N_3932);
xnor U4409 (N_4409,N_4104,N_3946);
or U4410 (N_4410,N_4030,N_4182);
xnor U4411 (N_4411,N_4148,N_4090);
or U4412 (N_4412,N_3970,N_3987);
nand U4413 (N_4413,N_4147,N_3961);
nand U4414 (N_4414,N_4111,N_3981);
and U4415 (N_4415,N_4000,N_4001);
or U4416 (N_4416,N_3974,N_4117);
or U4417 (N_4417,N_4190,N_4133);
nor U4418 (N_4418,N_4007,N_3985);
xnor U4419 (N_4419,N_4036,N_4007);
and U4420 (N_4420,N_4105,N_4122);
nor U4421 (N_4421,N_4124,N_4009);
nand U4422 (N_4422,N_3999,N_4068);
nor U4423 (N_4423,N_3988,N_3913);
nand U4424 (N_4424,N_4100,N_4179);
xor U4425 (N_4425,N_4108,N_4127);
and U4426 (N_4426,N_4077,N_3947);
and U4427 (N_4427,N_4143,N_3984);
nor U4428 (N_4428,N_4153,N_4169);
xor U4429 (N_4429,N_4081,N_4162);
nor U4430 (N_4430,N_3922,N_4162);
and U4431 (N_4431,N_4162,N_4018);
nand U4432 (N_4432,N_4137,N_4006);
nand U4433 (N_4433,N_4019,N_4030);
nor U4434 (N_4434,N_4067,N_4136);
or U4435 (N_4435,N_4027,N_3991);
nor U4436 (N_4436,N_3900,N_3952);
or U4437 (N_4437,N_3976,N_4182);
and U4438 (N_4438,N_3974,N_3926);
nor U4439 (N_4439,N_4003,N_4123);
nand U4440 (N_4440,N_3948,N_3922);
nand U4441 (N_4441,N_4001,N_4017);
and U4442 (N_4442,N_3972,N_4028);
xor U4443 (N_4443,N_4126,N_4069);
nor U4444 (N_4444,N_4095,N_4082);
nand U4445 (N_4445,N_3999,N_3912);
nand U4446 (N_4446,N_3933,N_3970);
xnor U4447 (N_4447,N_4198,N_3924);
or U4448 (N_4448,N_4119,N_4133);
nand U4449 (N_4449,N_4017,N_4187);
or U4450 (N_4450,N_4188,N_3951);
or U4451 (N_4451,N_3992,N_3953);
nand U4452 (N_4452,N_4165,N_4041);
or U4453 (N_4453,N_4049,N_3973);
and U4454 (N_4454,N_4028,N_4190);
or U4455 (N_4455,N_4100,N_4048);
xor U4456 (N_4456,N_3959,N_3969);
nor U4457 (N_4457,N_3961,N_3913);
nor U4458 (N_4458,N_4013,N_3984);
or U4459 (N_4459,N_3927,N_4163);
nor U4460 (N_4460,N_3925,N_4054);
nand U4461 (N_4461,N_4086,N_3989);
nor U4462 (N_4462,N_4198,N_3914);
nor U4463 (N_4463,N_4093,N_4028);
or U4464 (N_4464,N_4027,N_3957);
nor U4465 (N_4465,N_4184,N_4026);
nand U4466 (N_4466,N_3977,N_4116);
and U4467 (N_4467,N_3989,N_3971);
xnor U4468 (N_4468,N_4176,N_4198);
and U4469 (N_4469,N_4016,N_4118);
nand U4470 (N_4470,N_4187,N_3938);
or U4471 (N_4471,N_4150,N_4189);
nand U4472 (N_4472,N_3942,N_4068);
nand U4473 (N_4473,N_4004,N_4166);
nor U4474 (N_4474,N_4018,N_3970);
xor U4475 (N_4475,N_4125,N_4136);
xnor U4476 (N_4476,N_4150,N_4157);
xnor U4477 (N_4477,N_4171,N_4102);
and U4478 (N_4478,N_3972,N_3940);
xor U4479 (N_4479,N_3912,N_4175);
and U4480 (N_4480,N_4116,N_3940);
or U4481 (N_4481,N_4148,N_4103);
and U4482 (N_4482,N_4039,N_4103);
xnor U4483 (N_4483,N_4139,N_3953);
and U4484 (N_4484,N_4062,N_3987);
xor U4485 (N_4485,N_4127,N_4060);
or U4486 (N_4486,N_4089,N_4067);
nand U4487 (N_4487,N_4067,N_4169);
nor U4488 (N_4488,N_4070,N_4051);
and U4489 (N_4489,N_4070,N_4035);
xor U4490 (N_4490,N_4058,N_4035);
nor U4491 (N_4491,N_3994,N_4003);
nand U4492 (N_4492,N_4151,N_4060);
or U4493 (N_4493,N_3974,N_4020);
nand U4494 (N_4494,N_3974,N_3967);
nor U4495 (N_4495,N_3940,N_4034);
nor U4496 (N_4496,N_4059,N_3984);
or U4497 (N_4497,N_3965,N_4035);
nand U4498 (N_4498,N_4021,N_4107);
nand U4499 (N_4499,N_3972,N_3956);
nand U4500 (N_4500,N_4354,N_4405);
and U4501 (N_4501,N_4301,N_4280);
xnor U4502 (N_4502,N_4262,N_4315);
and U4503 (N_4503,N_4383,N_4219);
nand U4504 (N_4504,N_4366,N_4493);
xor U4505 (N_4505,N_4424,N_4390);
or U4506 (N_4506,N_4455,N_4420);
nor U4507 (N_4507,N_4391,N_4297);
nor U4508 (N_4508,N_4249,N_4233);
or U4509 (N_4509,N_4256,N_4258);
and U4510 (N_4510,N_4477,N_4369);
nand U4511 (N_4511,N_4353,N_4328);
and U4512 (N_4512,N_4430,N_4260);
nor U4513 (N_4513,N_4373,N_4403);
nand U4514 (N_4514,N_4423,N_4488);
and U4515 (N_4515,N_4441,N_4209);
nor U4516 (N_4516,N_4302,N_4474);
nor U4517 (N_4517,N_4339,N_4463);
xor U4518 (N_4518,N_4214,N_4313);
and U4519 (N_4519,N_4446,N_4444);
and U4520 (N_4520,N_4412,N_4485);
nand U4521 (N_4521,N_4284,N_4386);
xnor U4522 (N_4522,N_4375,N_4295);
and U4523 (N_4523,N_4498,N_4257);
nor U4524 (N_4524,N_4343,N_4232);
or U4525 (N_4525,N_4201,N_4407);
nand U4526 (N_4526,N_4345,N_4250);
nor U4527 (N_4527,N_4346,N_4290);
nand U4528 (N_4528,N_4235,N_4389);
nand U4529 (N_4529,N_4228,N_4494);
nor U4530 (N_4530,N_4229,N_4350);
and U4531 (N_4531,N_4453,N_4406);
and U4532 (N_4532,N_4274,N_4293);
xor U4533 (N_4533,N_4422,N_4259);
nand U4534 (N_4534,N_4234,N_4336);
and U4535 (N_4535,N_4253,N_4267);
xor U4536 (N_4536,N_4247,N_4427);
or U4537 (N_4537,N_4499,N_4223);
xnor U4538 (N_4538,N_4211,N_4400);
and U4539 (N_4539,N_4401,N_4478);
nand U4540 (N_4540,N_4337,N_4252);
xnor U4541 (N_4541,N_4268,N_4319);
nand U4542 (N_4542,N_4460,N_4398);
xnor U4543 (N_4543,N_4299,N_4322);
xnor U4544 (N_4544,N_4464,N_4459);
nand U4545 (N_4545,N_4410,N_4226);
nand U4546 (N_4546,N_4497,N_4372);
nand U4547 (N_4547,N_4426,N_4241);
nor U4548 (N_4548,N_4487,N_4292);
xnor U4549 (N_4549,N_4324,N_4320);
nand U4550 (N_4550,N_4447,N_4205);
or U4551 (N_4551,N_4334,N_4273);
nor U4552 (N_4552,N_4458,N_4291);
nand U4553 (N_4553,N_4392,N_4456);
or U4554 (N_4554,N_4222,N_4445);
nand U4555 (N_4555,N_4462,N_4311);
nand U4556 (N_4556,N_4448,N_4342);
nor U4557 (N_4557,N_4344,N_4415);
nand U4558 (N_4558,N_4206,N_4432);
nand U4559 (N_4559,N_4425,N_4321);
xor U4560 (N_4560,N_4307,N_4409);
and U4561 (N_4561,N_4326,N_4246);
nor U4562 (N_4562,N_4495,N_4238);
or U4563 (N_4563,N_4378,N_4368);
nor U4564 (N_4564,N_4340,N_4467);
nand U4565 (N_4565,N_4387,N_4379);
or U4566 (N_4566,N_4385,N_4479);
nor U4567 (N_4567,N_4363,N_4442);
nor U4568 (N_4568,N_4288,N_4461);
xnor U4569 (N_4569,N_4347,N_4490);
nor U4570 (N_4570,N_4207,N_4298);
and U4571 (N_4571,N_4281,N_4335);
xor U4572 (N_4572,N_4255,N_4397);
xnor U4573 (N_4573,N_4382,N_4395);
nor U4574 (N_4574,N_4220,N_4491);
xor U4575 (N_4575,N_4483,N_4312);
and U4576 (N_4576,N_4470,N_4367);
nor U4577 (N_4577,N_4231,N_4359);
and U4578 (N_4578,N_4221,N_4381);
nor U4579 (N_4579,N_4351,N_4314);
xor U4580 (N_4580,N_4362,N_4454);
and U4581 (N_4581,N_4417,N_4263);
and U4582 (N_4582,N_4254,N_4300);
or U4583 (N_4583,N_4308,N_4449);
and U4584 (N_4584,N_4333,N_4468);
and U4585 (N_4585,N_4419,N_4393);
or U4586 (N_4586,N_4275,N_4356);
and U4587 (N_4587,N_4279,N_4271);
nand U4588 (N_4588,N_4438,N_4332);
or U4589 (N_4589,N_4489,N_4416);
and U4590 (N_4590,N_4473,N_4411);
and U4591 (N_4591,N_4245,N_4304);
nor U4592 (N_4592,N_4421,N_4305);
xor U4593 (N_4593,N_4331,N_4352);
nand U4594 (N_4594,N_4278,N_4481);
and U4595 (N_4595,N_4436,N_4208);
nor U4596 (N_4596,N_4451,N_4466);
xnor U4597 (N_4597,N_4428,N_4360);
and U4598 (N_4598,N_4418,N_4434);
nand U4599 (N_4599,N_4227,N_4212);
nor U4600 (N_4600,N_4429,N_4371);
xnor U4601 (N_4601,N_4361,N_4244);
or U4602 (N_4602,N_4402,N_4435);
or U4603 (N_4603,N_4303,N_4408);
and U4604 (N_4604,N_4325,N_4437);
nor U4605 (N_4605,N_4443,N_4277);
xor U4606 (N_4606,N_4388,N_4457);
or U4607 (N_4607,N_4215,N_4380);
or U4608 (N_4608,N_4203,N_4480);
nand U4609 (N_4609,N_4218,N_4204);
nor U4610 (N_4610,N_4341,N_4309);
and U4611 (N_4611,N_4266,N_4296);
nand U4612 (N_4612,N_4225,N_4394);
xor U4613 (N_4613,N_4202,N_4374);
and U4614 (N_4614,N_4283,N_4475);
and U4615 (N_4615,N_4348,N_4240);
nand U4616 (N_4616,N_4377,N_4465);
nor U4617 (N_4617,N_4413,N_4349);
or U4618 (N_4618,N_4327,N_4294);
nor U4619 (N_4619,N_4399,N_4492);
and U4620 (N_4620,N_4310,N_4264);
and U4621 (N_4621,N_4431,N_4482);
and U4622 (N_4622,N_4289,N_4216);
or U4623 (N_4623,N_4265,N_4338);
nand U4624 (N_4624,N_4414,N_4439);
nand U4625 (N_4625,N_4318,N_4472);
and U4626 (N_4626,N_4239,N_4236);
nor U4627 (N_4627,N_4306,N_4476);
xor U4628 (N_4628,N_4276,N_4316);
or U4629 (N_4629,N_4237,N_4323);
nand U4630 (N_4630,N_4486,N_4358);
xor U4631 (N_4631,N_4242,N_4248);
nand U4632 (N_4632,N_4217,N_4450);
nor U4633 (N_4633,N_4452,N_4329);
and U4634 (N_4634,N_4404,N_4210);
nor U4635 (N_4635,N_4370,N_4224);
or U4636 (N_4636,N_4286,N_4484);
nand U4637 (N_4637,N_4269,N_4317);
nor U4638 (N_4638,N_4365,N_4469);
nor U4639 (N_4639,N_4330,N_4496);
or U4640 (N_4640,N_4251,N_4261);
and U4641 (N_4641,N_4396,N_4384);
nand U4642 (N_4642,N_4376,N_4433);
nor U4643 (N_4643,N_4272,N_4230);
xnor U4644 (N_4644,N_4200,N_4285);
nand U4645 (N_4645,N_4471,N_4364);
xnor U4646 (N_4646,N_4357,N_4355);
or U4647 (N_4647,N_4243,N_4440);
xnor U4648 (N_4648,N_4287,N_4213);
nor U4649 (N_4649,N_4282,N_4270);
or U4650 (N_4650,N_4405,N_4276);
or U4651 (N_4651,N_4224,N_4219);
nand U4652 (N_4652,N_4357,N_4410);
nor U4653 (N_4653,N_4466,N_4342);
and U4654 (N_4654,N_4223,N_4262);
xnor U4655 (N_4655,N_4279,N_4379);
or U4656 (N_4656,N_4468,N_4341);
or U4657 (N_4657,N_4362,N_4476);
and U4658 (N_4658,N_4212,N_4451);
nand U4659 (N_4659,N_4319,N_4340);
or U4660 (N_4660,N_4487,N_4351);
xnor U4661 (N_4661,N_4376,N_4370);
xnor U4662 (N_4662,N_4245,N_4482);
and U4663 (N_4663,N_4256,N_4293);
and U4664 (N_4664,N_4442,N_4274);
xnor U4665 (N_4665,N_4261,N_4207);
nor U4666 (N_4666,N_4375,N_4423);
or U4667 (N_4667,N_4490,N_4222);
and U4668 (N_4668,N_4244,N_4353);
and U4669 (N_4669,N_4217,N_4323);
xor U4670 (N_4670,N_4222,N_4362);
xor U4671 (N_4671,N_4484,N_4338);
nor U4672 (N_4672,N_4276,N_4437);
or U4673 (N_4673,N_4204,N_4333);
nor U4674 (N_4674,N_4393,N_4340);
xor U4675 (N_4675,N_4294,N_4376);
xor U4676 (N_4676,N_4454,N_4482);
and U4677 (N_4677,N_4372,N_4486);
and U4678 (N_4678,N_4280,N_4442);
xnor U4679 (N_4679,N_4314,N_4237);
or U4680 (N_4680,N_4256,N_4389);
nor U4681 (N_4681,N_4329,N_4244);
or U4682 (N_4682,N_4485,N_4495);
nor U4683 (N_4683,N_4416,N_4398);
nor U4684 (N_4684,N_4258,N_4224);
and U4685 (N_4685,N_4231,N_4324);
or U4686 (N_4686,N_4298,N_4380);
or U4687 (N_4687,N_4433,N_4367);
nor U4688 (N_4688,N_4415,N_4283);
nand U4689 (N_4689,N_4443,N_4432);
nand U4690 (N_4690,N_4492,N_4344);
or U4691 (N_4691,N_4449,N_4368);
or U4692 (N_4692,N_4491,N_4225);
xor U4693 (N_4693,N_4321,N_4298);
and U4694 (N_4694,N_4346,N_4279);
nor U4695 (N_4695,N_4417,N_4396);
xor U4696 (N_4696,N_4343,N_4393);
xor U4697 (N_4697,N_4327,N_4311);
nor U4698 (N_4698,N_4343,N_4249);
nand U4699 (N_4699,N_4309,N_4306);
nor U4700 (N_4700,N_4453,N_4412);
xor U4701 (N_4701,N_4271,N_4343);
nand U4702 (N_4702,N_4458,N_4334);
and U4703 (N_4703,N_4495,N_4399);
nor U4704 (N_4704,N_4223,N_4234);
and U4705 (N_4705,N_4275,N_4311);
xnor U4706 (N_4706,N_4308,N_4286);
xnor U4707 (N_4707,N_4330,N_4349);
and U4708 (N_4708,N_4449,N_4354);
nand U4709 (N_4709,N_4367,N_4318);
and U4710 (N_4710,N_4282,N_4398);
and U4711 (N_4711,N_4416,N_4316);
and U4712 (N_4712,N_4203,N_4448);
and U4713 (N_4713,N_4384,N_4375);
or U4714 (N_4714,N_4258,N_4414);
nand U4715 (N_4715,N_4275,N_4236);
or U4716 (N_4716,N_4290,N_4415);
or U4717 (N_4717,N_4355,N_4390);
xnor U4718 (N_4718,N_4394,N_4327);
and U4719 (N_4719,N_4250,N_4322);
xnor U4720 (N_4720,N_4495,N_4328);
or U4721 (N_4721,N_4248,N_4404);
nand U4722 (N_4722,N_4228,N_4200);
xnor U4723 (N_4723,N_4473,N_4330);
xor U4724 (N_4724,N_4477,N_4482);
nand U4725 (N_4725,N_4281,N_4457);
xnor U4726 (N_4726,N_4360,N_4215);
nor U4727 (N_4727,N_4396,N_4241);
or U4728 (N_4728,N_4433,N_4246);
nand U4729 (N_4729,N_4482,N_4219);
xor U4730 (N_4730,N_4449,N_4320);
nor U4731 (N_4731,N_4252,N_4278);
nand U4732 (N_4732,N_4220,N_4375);
nand U4733 (N_4733,N_4450,N_4251);
nor U4734 (N_4734,N_4429,N_4288);
and U4735 (N_4735,N_4461,N_4470);
nor U4736 (N_4736,N_4358,N_4302);
nor U4737 (N_4737,N_4441,N_4387);
or U4738 (N_4738,N_4282,N_4297);
and U4739 (N_4739,N_4271,N_4412);
or U4740 (N_4740,N_4380,N_4286);
nand U4741 (N_4741,N_4262,N_4260);
xor U4742 (N_4742,N_4479,N_4493);
nand U4743 (N_4743,N_4478,N_4347);
and U4744 (N_4744,N_4453,N_4341);
nor U4745 (N_4745,N_4313,N_4304);
nand U4746 (N_4746,N_4200,N_4478);
or U4747 (N_4747,N_4248,N_4438);
nand U4748 (N_4748,N_4272,N_4469);
xnor U4749 (N_4749,N_4365,N_4463);
or U4750 (N_4750,N_4282,N_4471);
or U4751 (N_4751,N_4439,N_4478);
and U4752 (N_4752,N_4240,N_4252);
and U4753 (N_4753,N_4480,N_4243);
and U4754 (N_4754,N_4368,N_4442);
or U4755 (N_4755,N_4360,N_4252);
xnor U4756 (N_4756,N_4423,N_4403);
nand U4757 (N_4757,N_4499,N_4414);
xor U4758 (N_4758,N_4348,N_4353);
nand U4759 (N_4759,N_4205,N_4280);
or U4760 (N_4760,N_4385,N_4298);
nor U4761 (N_4761,N_4398,N_4437);
nand U4762 (N_4762,N_4328,N_4479);
or U4763 (N_4763,N_4309,N_4464);
nor U4764 (N_4764,N_4430,N_4205);
or U4765 (N_4765,N_4359,N_4426);
nand U4766 (N_4766,N_4427,N_4399);
nor U4767 (N_4767,N_4249,N_4413);
and U4768 (N_4768,N_4211,N_4495);
and U4769 (N_4769,N_4391,N_4265);
nor U4770 (N_4770,N_4313,N_4372);
nor U4771 (N_4771,N_4340,N_4430);
xnor U4772 (N_4772,N_4265,N_4475);
nor U4773 (N_4773,N_4368,N_4284);
and U4774 (N_4774,N_4453,N_4392);
xnor U4775 (N_4775,N_4368,N_4295);
and U4776 (N_4776,N_4219,N_4377);
and U4777 (N_4777,N_4257,N_4440);
or U4778 (N_4778,N_4346,N_4204);
and U4779 (N_4779,N_4287,N_4328);
nand U4780 (N_4780,N_4317,N_4251);
and U4781 (N_4781,N_4361,N_4212);
nor U4782 (N_4782,N_4312,N_4437);
xnor U4783 (N_4783,N_4492,N_4393);
xnor U4784 (N_4784,N_4332,N_4313);
nor U4785 (N_4785,N_4438,N_4278);
or U4786 (N_4786,N_4262,N_4372);
xnor U4787 (N_4787,N_4468,N_4235);
nor U4788 (N_4788,N_4330,N_4484);
nor U4789 (N_4789,N_4396,N_4434);
nand U4790 (N_4790,N_4358,N_4217);
nand U4791 (N_4791,N_4221,N_4238);
nor U4792 (N_4792,N_4266,N_4433);
xnor U4793 (N_4793,N_4329,N_4428);
or U4794 (N_4794,N_4293,N_4318);
nor U4795 (N_4795,N_4400,N_4268);
xor U4796 (N_4796,N_4302,N_4355);
or U4797 (N_4797,N_4453,N_4214);
xor U4798 (N_4798,N_4370,N_4225);
xnor U4799 (N_4799,N_4481,N_4382);
xor U4800 (N_4800,N_4589,N_4565);
xor U4801 (N_4801,N_4675,N_4531);
nor U4802 (N_4802,N_4791,N_4528);
nand U4803 (N_4803,N_4797,N_4525);
nor U4804 (N_4804,N_4511,N_4640);
nor U4805 (N_4805,N_4600,N_4731);
nor U4806 (N_4806,N_4611,N_4766);
and U4807 (N_4807,N_4720,N_4738);
nand U4808 (N_4808,N_4631,N_4752);
nor U4809 (N_4809,N_4756,N_4561);
nor U4810 (N_4810,N_4614,N_4655);
and U4811 (N_4811,N_4653,N_4771);
or U4812 (N_4812,N_4633,N_4693);
or U4813 (N_4813,N_4566,N_4699);
or U4814 (N_4814,N_4586,N_4728);
and U4815 (N_4815,N_4568,N_4734);
and U4816 (N_4816,N_4799,N_4585);
nand U4817 (N_4817,N_4588,N_4639);
nand U4818 (N_4818,N_4500,N_4740);
xnor U4819 (N_4819,N_4700,N_4770);
and U4820 (N_4820,N_4562,N_4609);
xnor U4821 (N_4821,N_4613,N_4570);
or U4822 (N_4822,N_4524,N_4748);
or U4823 (N_4823,N_4519,N_4713);
or U4824 (N_4824,N_4768,N_4571);
xor U4825 (N_4825,N_4597,N_4607);
or U4826 (N_4826,N_4628,N_4627);
xnor U4827 (N_4827,N_4711,N_4648);
nor U4828 (N_4828,N_4735,N_4520);
xnor U4829 (N_4829,N_4694,N_4754);
nand U4830 (N_4830,N_4643,N_4721);
and U4831 (N_4831,N_4666,N_4564);
nand U4832 (N_4832,N_4642,N_4764);
xnor U4833 (N_4833,N_4676,N_4767);
nand U4834 (N_4834,N_4579,N_4783);
nand U4835 (N_4835,N_4606,N_4557);
nand U4836 (N_4836,N_4618,N_4595);
and U4837 (N_4837,N_4681,N_4707);
or U4838 (N_4838,N_4773,N_4533);
nor U4839 (N_4839,N_4708,N_4513);
and U4840 (N_4840,N_4719,N_4775);
or U4841 (N_4841,N_4795,N_4651);
nor U4842 (N_4842,N_4736,N_4677);
nand U4843 (N_4843,N_4506,N_4745);
or U4844 (N_4844,N_4584,N_4776);
nor U4845 (N_4845,N_4787,N_4619);
nand U4846 (N_4846,N_4554,N_4674);
xor U4847 (N_4847,N_4501,N_4730);
and U4848 (N_4848,N_4701,N_4503);
or U4849 (N_4849,N_4656,N_4502);
xnor U4850 (N_4850,N_4781,N_4757);
and U4851 (N_4851,N_4690,N_4784);
and U4852 (N_4852,N_4567,N_4749);
nor U4853 (N_4853,N_4669,N_4542);
and U4854 (N_4854,N_4536,N_4665);
xor U4855 (N_4855,N_4794,N_4788);
nor U4856 (N_4856,N_4569,N_4539);
nand U4857 (N_4857,N_4516,N_4594);
nor U4858 (N_4858,N_4723,N_4729);
nor U4859 (N_4859,N_4644,N_4543);
nor U4860 (N_4860,N_4509,N_4761);
nand U4861 (N_4861,N_4538,N_4685);
and U4862 (N_4862,N_4626,N_4512);
xor U4863 (N_4863,N_4551,N_4632);
and U4864 (N_4864,N_4591,N_4650);
or U4865 (N_4865,N_4762,N_4544);
nor U4866 (N_4866,N_4532,N_4673);
nor U4867 (N_4867,N_4523,N_4630);
nand U4868 (N_4868,N_4652,N_4535);
nand U4869 (N_4869,N_4744,N_4504);
nand U4870 (N_4870,N_4641,N_4581);
nor U4871 (N_4871,N_4601,N_4548);
nand U4872 (N_4872,N_4592,N_4629);
nor U4873 (N_4873,N_4559,N_4649);
nor U4874 (N_4874,N_4507,N_4605);
nand U4875 (N_4875,N_4555,N_4578);
or U4876 (N_4876,N_4662,N_4737);
or U4877 (N_4877,N_4508,N_4540);
or U4878 (N_4878,N_4654,N_4657);
xnor U4879 (N_4879,N_4560,N_4610);
nor U4880 (N_4880,N_4722,N_4704);
or U4881 (N_4881,N_4697,N_4705);
nand U4882 (N_4882,N_4663,N_4637);
xor U4883 (N_4883,N_4634,N_4715);
xor U4884 (N_4884,N_4658,N_4537);
nor U4885 (N_4885,N_4659,N_4716);
xor U4886 (N_4886,N_4798,N_4772);
xnor U4887 (N_4887,N_4689,N_4750);
nand U4888 (N_4888,N_4563,N_4726);
and U4889 (N_4889,N_4647,N_4598);
nand U4890 (N_4890,N_4518,N_4514);
or U4891 (N_4891,N_4746,N_4688);
xor U4892 (N_4892,N_4696,N_4671);
and U4893 (N_4893,N_4620,N_4703);
or U4894 (N_4894,N_4769,N_4617);
xnor U4895 (N_4895,N_4616,N_4576);
or U4896 (N_4896,N_4751,N_4515);
nor U4897 (N_4897,N_4583,N_4683);
xor U4898 (N_4898,N_4777,N_4765);
nand U4899 (N_4899,N_4505,N_4792);
nor U4900 (N_4900,N_4733,N_4552);
or U4901 (N_4901,N_4779,N_4623);
xnor U4902 (N_4902,N_4574,N_4739);
and U4903 (N_4903,N_4702,N_4624);
or U4904 (N_4904,N_4695,N_4760);
and U4905 (N_4905,N_4789,N_4575);
nand U4906 (N_4906,N_4692,N_4712);
and U4907 (N_4907,N_4796,N_4686);
or U4908 (N_4908,N_4558,N_4573);
nand U4909 (N_4909,N_4763,N_4774);
or U4910 (N_4910,N_4710,N_4755);
nand U4911 (N_4911,N_4793,N_4778);
and U4912 (N_4912,N_4638,N_4680);
nor U4913 (N_4913,N_4660,N_4621);
nor U4914 (N_4914,N_4672,N_4526);
nor U4915 (N_4915,N_4608,N_4661);
nand U4916 (N_4916,N_4667,N_4615);
nor U4917 (N_4917,N_4790,N_4596);
xor U4918 (N_4918,N_4580,N_4590);
nor U4919 (N_4919,N_4530,N_4550);
or U4920 (N_4920,N_4599,N_4521);
xor U4921 (N_4921,N_4517,N_4541);
nor U4922 (N_4922,N_4725,N_4529);
and U4923 (N_4923,N_4684,N_4759);
nand U4924 (N_4924,N_4742,N_4545);
xnor U4925 (N_4925,N_4678,N_4646);
xor U4926 (N_4926,N_4727,N_4709);
and U4927 (N_4927,N_4572,N_4682);
or U4928 (N_4928,N_4602,N_4603);
or U4929 (N_4929,N_4743,N_4679);
and U4930 (N_4930,N_4753,N_4758);
or U4931 (N_4931,N_4625,N_4717);
nand U4932 (N_4932,N_4556,N_4547);
nor U4933 (N_4933,N_4741,N_4622);
or U4934 (N_4934,N_4612,N_4786);
xor U4935 (N_4935,N_4645,N_4732);
or U4936 (N_4936,N_4582,N_4691);
nor U4937 (N_4937,N_4534,N_4698);
xnor U4938 (N_4938,N_4718,N_4549);
nand U4939 (N_4939,N_4636,N_4747);
or U4940 (N_4940,N_4782,N_4780);
nor U4941 (N_4941,N_4668,N_4664);
nand U4942 (N_4942,N_4577,N_4553);
xnor U4943 (N_4943,N_4635,N_4546);
nand U4944 (N_4944,N_4785,N_4670);
and U4945 (N_4945,N_4687,N_4604);
nand U4946 (N_4946,N_4510,N_4714);
xnor U4947 (N_4947,N_4527,N_4706);
and U4948 (N_4948,N_4522,N_4724);
and U4949 (N_4949,N_4587,N_4593);
xnor U4950 (N_4950,N_4525,N_4731);
xor U4951 (N_4951,N_4535,N_4633);
xor U4952 (N_4952,N_4782,N_4695);
or U4953 (N_4953,N_4635,N_4524);
or U4954 (N_4954,N_4640,N_4671);
nor U4955 (N_4955,N_4643,N_4504);
nor U4956 (N_4956,N_4551,N_4644);
nand U4957 (N_4957,N_4791,N_4609);
nor U4958 (N_4958,N_4568,N_4732);
or U4959 (N_4959,N_4692,N_4639);
nor U4960 (N_4960,N_4668,N_4710);
nand U4961 (N_4961,N_4644,N_4793);
or U4962 (N_4962,N_4644,N_4668);
or U4963 (N_4963,N_4521,N_4727);
xnor U4964 (N_4964,N_4691,N_4515);
or U4965 (N_4965,N_4561,N_4713);
xor U4966 (N_4966,N_4768,N_4589);
nand U4967 (N_4967,N_4596,N_4728);
and U4968 (N_4968,N_4680,N_4797);
xor U4969 (N_4969,N_4615,N_4735);
nor U4970 (N_4970,N_4677,N_4759);
and U4971 (N_4971,N_4779,N_4603);
or U4972 (N_4972,N_4763,N_4620);
and U4973 (N_4973,N_4607,N_4751);
xor U4974 (N_4974,N_4621,N_4506);
nand U4975 (N_4975,N_4534,N_4528);
or U4976 (N_4976,N_4777,N_4670);
or U4977 (N_4977,N_4765,N_4569);
and U4978 (N_4978,N_4618,N_4787);
and U4979 (N_4979,N_4727,N_4665);
nor U4980 (N_4980,N_4766,N_4781);
and U4981 (N_4981,N_4767,N_4567);
and U4982 (N_4982,N_4609,N_4569);
xor U4983 (N_4983,N_4737,N_4773);
xor U4984 (N_4984,N_4673,N_4500);
nor U4985 (N_4985,N_4504,N_4593);
or U4986 (N_4986,N_4609,N_4728);
nor U4987 (N_4987,N_4798,N_4500);
or U4988 (N_4988,N_4620,N_4584);
xor U4989 (N_4989,N_4512,N_4665);
or U4990 (N_4990,N_4647,N_4570);
nor U4991 (N_4991,N_4614,N_4575);
nor U4992 (N_4992,N_4527,N_4707);
xnor U4993 (N_4993,N_4738,N_4751);
nand U4994 (N_4994,N_4785,N_4763);
nor U4995 (N_4995,N_4630,N_4758);
or U4996 (N_4996,N_4674,N_4503);
nand U4997 (N_4997,N_4503,N_4583);
nor U4998 (N_4998,N_4675,N_4766);
or U4999 (N_4999,N_4609,N_4701);
and U5000 (N_5000,N_4770,N_4763);
or U5001 (N_5001,N_4506,N_4655);
xor U5002 (N_5002,N_4601,N_4709);
nand U5003 (N_5003,N_4766,N_4719);
or U5004 (N_5004,N_4630,N_4671);
nand U5005 (N_5005,N_4788,N_4527);
or U5006 (N_5006,N_4698,N_4671);
nand U5007 (N_5007,N_4730,N_4774);
and U5008 (N_5008,N_4557,N_4795);
xnor U5009 (N_5009,N_4543,N_4765);
xor U5010 (N_5010,N_4548,N_4779);
nand U5011 (N_5011,N_4722,N_4577);
nand U5012 (N_5012,N_4529,N_4581);
nor U5013 (N_5013,N_4513,N_4525);
xnor U5014 (N_5014,N_4651,N_4792);
nand U5015 (N_5015,N_4661,N_4634);
or U5016 (N_5016,N_4768,N_4502);
nand U5017 (N_5017,N_4524,N_4736);
and U5018 (N_5018,N_4599,N_4733);
nand U5019 (N_5019,N_4785,N_4575);
or U5020 (N_5020,N_4554,N_4787);
or U5021 (N_5021,N_4773,N_4525);
or U5022 (N_5022,N_4698,N_4584);
and U5023 (N_5023,N_4544,N_4642);
or U5024 (N_5024,N_4595,N_4508);
xnor U5025 (N_5025,N_4550,N_4628);
or U5026 (N_5026,N_4687,N_4511);
nor U5027 (N_5027,N_4610,N_4633);
xnor U5028 (N_5028,N_4652,N_4538);
nand U5029 (N_5029,N_4650,N_4630);
or U5030 (N_5030,N_4550,N_4566);
nor U5031 (N_5031,N_4541,N_4682);
nand U5032 (N_5032,N_4767,N_4659);
xnor U5033 (N_5033,N_4614,N_4579);
nand U5034 (N_5034,N_4569,N_4671);
and U5035 (N_5035,N_4560,N_4683);
nor U5036 (N_5036,N_4700,N_4615);
nor U5037 (N_5037,N_4748,N_4695);
or U5038 (N_5038,N_4545,N_4752);
xnor U5039 (N_5039,N_4751,N_4567);
and U5040 (N_5040,N_4757,N_4696);
xor U5041 (N_5041,N_4648,N_4721);
nor U5042 (N_5042,N_4759,N_4505);
xnor U5043 (N_5043,N_4675,N_4653);
nor U5044 (N_5044,N_4597,N_4779);
and U5045 (N_5045,N_4603,N_4505);
or U5046 (N_5046,N_4624,N_4742);
nor U5047 (N_5047,N_4757,N_4635);
and U5048 (N_5048,N_4753,N_4576);
xor U5049 (N_5049,N_4522,N_4520);
or U5050 (N_5050,N_4692,N_4659);
xnor U5051 (N_5051,N_4557,N_4631);
nor U5052 (N_5052,N_4692,N_4697);
nor U5053 (N_5053,N_4778,N_4780);
xor U5054 (N_5054,N_4736,N_4564);
and U5055 (N_5055,N_4645,N_4614);
and U5056 (N_5056,N_4657,N_4796);
nor U5057 (N_5057,N_4565,N_4765);
or U5058 (N_5058,N_4651,N_4774);
xor U5059 (N_5059,N_4525,N_4648);
xor U5060 (N_5060,N_4714,N_4501);
nor U5061 (N_5061,N_4715,N_4513);
nand U5062 (N_5062,N_4772,N_4641);
and U5063 (N_5063,N_4604,N_4770);
xnor U5064 (N_5064,N_4594,N_4521);
nor U5065 (N_5065,N_4621,N_4728);
xnor U5066 (N_5066,N_4640,N_4601);
and U5067 (N_5067,N_4590,N_4793);
nand U5068 (N_5068,N_4631,N_4518);
or U5069 (N_5069,N_4720,N_4517);
xor U5070 (N_5070,N_4602,N_4599);
or U5071 (N_5071,N_4705,N_4600);
nor U5072 (N_5072,N_4794,N_4656);
nand U5073 (N_5073,N_4593,N_4631);
and U5074 (N_5074,N_4555,N_4648);
nand U5075 (N_5075,N_4689,N_4720);
or U5076 (N_5076,N_4692,N_4778);
nor U5077 (N_5077,N_4744,N_4558);
and U5078 (N_5078,N_4581,N_4652);
nand U5079 (N_5079,N_4588,N_4575);
nor U5080 (N_5080,N_4673,N_4501);
nand U5081 (N_5081,N_4533,N_4718);
xor U5082 (N_5082,N_4708,N_4709);
xor U5083 (N_5083,N_4792,N_4767);
and U5084 (N_5084,N_4592,N_4603);
nor U5085 (N_5085,N_4569,N_4512);
and U5086 (N_5086,N_4614,N_4708);
or U5087 (N_5087,N_4647,N_4710);
nand U5088 (N_5088,N_4733,N_4590);
or U5089 (N_5089,N_4759,N_4716);
nand U5090 (N_5090,N_4506,N_4567);
nor U5091 (N_5091,N_4787,N_4561);
nor U5092 (N_5092,N_4678,N_4703);
xor U5093 (N_5093,N_4723,N_4536);
xnor U5094 (N_5094,N_4522,N_4551);
or U5095 (N_5095,N_4714,N_4742);
or U5096 (N_5096,N_4768,N_4746);
nand U5097 (N_5097,N_4587,N_4571);
and U5098 (N_5098,N_4633,N_4525);
or U5099 (N_5099,N_4615,N_4740);
xnor U5100 (N_5100,N_5087,N_5070);
or U5101 (N_5101,N_4834,N_4815);
and U5102 (N_5102,N_4879,N_4968);
and U5103 (N_5103,N_4803,N_4985);
nand U5104 (N_5104,N_5044,N_5084);
xor U5105 (N_5105,N_5075,N_4813);
nand U5106 (N_5106,N_4853,N_5045);
nand U5107 (N_5107,N_4911,N_4923);
and U5108 (N_5108,N_5007,N_4971);
xnor U5109 (N_5109,N_4938,N_4890);
nor U5110 (N_5110,N_4842,N_5065);
or U5111 (N_5111,N_4986,N_5052);
xor U5112 (N_5112,N_5018,N_4989);
xor U5113 (N_5113,N_4870,N_5085);
or U5114 (N_5114,N_5020,N_4949);
nand U5115 (N_5115,N_5046,N_4980);
xor U5116 (N_5116,N_5004,N_5005);
or U5117 (N_5117,N_4983,N_5032);
and U5118 (N_5118,N_4955,N_4916);
nor U5119 (N_5119,N_5014,N_4977);
or U5120 (N_5120,N_4832,N_4881);
nand U5121 (N_5121,N_4909,N_5013);
or U5122 (N_5122,N_4958,N_5074);
xnor U5123 (N_5123,N_4867,N_4818);
xnor U5124 (N_5124,N_4892,N_5025);
xnor U5125 (N_5125,N_5029,N_4970);
nand U5126 (N_5126,N_5080,N_4947);
nand U5127 (N_5127,N_4952,N_4910);
or U5128 (N_5128,N_4921,N_4844);
nor U5129 (N_5129,N_4954,N_5028);
or U5130 (N_5130,N_5050,N_4998);
nor U5131 (N_5131,N_5094,N_5095);
xnor U5132 (N_5132,N_4975,N_4808);
xnor U5133 (N_5133,N_5092,N_4886);
nor U5134 (N_5134,N_5097,N_4988);
nand U5135 (N_5135,N_4894,N_4807);
xnor U5136 (N_5136,N_5015,N_4864);
and U5137 (N_5137,N_4876,N_5069);
nor U5138 (N_5138,N_4825,N_4840);
nor U5139 (N_5139,N_4976,N_5000);
xor U5140 (N_5140,N_4805,N_4929);
xnor U5141 (N_5141,N_4979,N_5063);
and U5142 (N_5142,N_4974,N_4869);
or U5143 (N_5143,N_5035,N_4816);
nor U5144 (N_5144,N_4888,N_4871);
nor U5145 (N_5145,N_4927,N_4908);
and U5146 (N_5146,N_5039,N_5057);
xnor U5147 (N_5147,N_4982,N_5072);
nand U5148 (N_5148,N_5034,N_5026);
and U5149 (N_5149,N_4981,N_5043);
nor U5150 (N_5150,N_5086,N_4969);
nand U5151 (N_5151,N_5068,N_4914);
and U5152 (N_5152,N_4994,N_4862);
or U5153 (N_5153,N_4882,N_5099);
or U5154 (N_5154,N_4852,N_4854);
nand U5155 (N_5155,N_4802,N_4812);
xnor U5156 (N_5156,N_5091,N_5067);
xor U5157 (N_5157,N_4851,N_4865);
nor U5158 (N_5158,N_4933,N_5036);
or U5159 (N_5159,N_4861,N_5071);
or U5160 (N_5160,N_4904,N_4942);
and U5161 (N_5161,N_5049,N_5061);
nor U5162 (N_5162,N_5081,N_4822);
xor U5163 (N_5163,N_4884,N_4868);
or U5164 (N_5164,N_4887,N_4996);
xor U5165 (N_5165,N_5027,N_4841);
nand U5166 (N_5166,N_4936,N_4823);
nand U5167 (N_5167,N_4992,N_4846);
or U5168 (N_5168,N_4913,N_4827);
and U5169 (N_5169,N_4866,N_5064);
and U5170 (N_5170,N_4801,N_5019);
and U5171 (N_5171,N_4848,N_5022);
or U5172 (N_5172,N_4880,N_4814);
or U5173 (N_5173,N_4895,N_5006);
or U5174 (N_5174,N_5073,N_4900);
nor U5175 (N_5175,N_4837,N_4993);
nor U5176 (N_5176,N_4984,N_5066);
and U5177 (N_5177,N_4961,N_4875);
or U5178 (N_5178,N_4917,N_5078);
or U5179 (N_5179,N_5079,N_4883);
xnor U5180 (N_5180,N_4847,N_4964);
xor U5181 (N_5181,N_4906,N_5089);
or U5182 (N_5182,N_4850,N_4943);
or U5183 (N_5183,N_4941,N_5033);
xnor U5184 (N_5184,N_4944,N_5010);
or U5185 (N_5185,N_4838,N_4946);
and U5186 (N_5186,N_4856,N_5047);
nand U5187 (N_5187,N_4824,N_4963);
xor U5188 (N_5188,N_4907,N_4819);
xnor U5189 (N_5189,N_4912,N_4836);
or U5190 (N_5190,N_5060,N_5055);
nor U5191 (N_5191,N_5053,N_4903);
xor U5192 (N_5192,N_5051,N_4967);
or U5193 (N_5193,N_5076,N_4962);
and U5194 (N_5194,N_4897,N_4831);
nand U5195 (N_5195,N_4873,N_5042);
nor U5196 (N_5196,N_5062,N_4804);
nand U5197 (N_5197,N_4925,N_4945);
and U5198 (N_5198,N_4920,N_4811);
or U5199 (N_5199,N_5016,N_4972);
nor U5200 (N_5200,N_4830,N_4889);
or U5201 (N_5201,N_4990,N_4833);
nor U5202 (N_5202,N_4826,N_5096);
and U5203 (N_5203,N_4839,N_5056);
xor U5204 (N_5204,N_5054,N_4924);
or U5205 (N_5205,N_4935,N_5083);
nand U5206 (N_5206,N_4934,N_4800);
or U5207 (N_5207,N_5003,N_5040);
and U5208 (N_5208,N_4960,N_5038);
nand U5209 (N_5209,N_4820,N_4821);
xnor U5210 (N_5210,N_5002,N_5001);
nand U5211 (N_5211,N_4806,N_4902);
or U5212 (N_5212,N_4966,N_5077);
xor U5213 (N_5213,N_4940,N_4973);
nand U5214 (N_5214,N_4872,N_4891);
and U5215 (N_5215,N_5008,N_4950);
xnor U5216 (N_5216,N_4857,N_4898);
xor U5217 (N_5217,N_5082,N_4863);
nand U5218 (N_5218,N_4931,N_4835);
or U5219 (N_5219,N_4987,N_4959);
nand U5220 (N_5220,N_4928,N_4858);
and U5221 (N_5221,N_4896,N_4995);
xor U5222 (N_5222,N_4951,N_4926);
nand U5223 (N_5223,N_4978,N_4965);
and U5224 (N_5224,N_4937,N_5017);
and U5225 (N_5225,N_4893,N_5058);
or U5226 (N_5226,N_5009,N_4809);
xnor U5227 (N_5227,N_4918,N_4919);
nor U5228 (N_5228,N_4953,N_5037);
or U5229 (N_5229,N_4874,N_4999);
nand U5230 (N_5230,N_5023,N_4860);
or U5231 (N_5231,N_4991,N_4997);
or U5232 (N_5232,N_4817,N_5024);
or U5233 (N_5233,N_5059,N_4878);
or U5234 (N_5234,N_4810,N_5041);
nand U5235 (N_5235,N_4957,N_5098);
nor U5236 (N_5236,N_4915,N_4849);
nand U5237 (N_5237,N_4939,N_5090);
and U5238 (N_5238,N_4843,N_4901);
xor U5239 (N_5239,N_4877,N_4922);
and U5240 (N_5240,N_5011,N_5031);
and U5241 (N_5241,N_4845,N_4855);
xnor U5242 (N_5242,N_5088,N_4885);
xor U5243 (N_5243,N_4930,N_4828);
nor U5244 (N_5244,N_5030,N_5048);
nor U5245 (N_5245,N_4829,N_5021);
or U5246 (N_5246,N_5093,N_4956);
nand U5247 (N_5247,N_4859,N_5012);
or U5248 (N_5248,N_4948,N_4932);
xor U5249 (N_5249,N_4899,N_4905);
xor U5250 (N_5250,N_4836,N_4831);
and U5251 (N_5251,N_5023,N_4979);
xnor U5252 (N_5252,N_4970,N_5095);
or U5253 (N_5253,N_4985,N_4952);
nand U5254 (N_5254,N_4966,N_4937);
nor U5255 (N_5255,N_5074,N_4968);
or U5256 (N_5256,N_4984,N_5062);
or U5257 (N_5257,N_4976,N_5007);
nand U5258 (N_5258,N_4898,N_4815);
xnor U5259 (N_5259,N_4832,N_5054);
and U5260 (N_5260,N_5051,N_4926);
or U5261 (N_5261,N_4898,N_4924);
xnor U5262 (N_5262,N_4969,N_4864);
nor U5263 (N_5263,N_4896,N_5030);
xor U5264 (N_5264,N_4946,N_4935);
nand U5265 (N_5265,N_4935,N_4806);
and U5266 (N_5266,N_5061,N_4978);
or U5267 (N_5267,N_5036,N_4935);
xnor U5268 (N_5268,N_4989,N_5089);
nand U5269 (N_5269,N_4805,N_4853);
or U5270 (N_5270,N_4868,N_5097);
nor U5271 (N_5271,N_4846,N_5062);
nand U5272 (N_5272,N_4941,N_4825);
xnor U5273 (N_5273,N_4846,N_5074);
and U5274 (N_5274,N_4894,N_5002);
nand U5275 (N_5275,N_4810,N_5022);
nor U5276 (N_5276,N_4950,N_5072);
or U5277 (N_5277,N_4995,N_5042);
and U5278 (N_5278,N_5087,N_4993);
and U5279 (N_5279,N_4830,N_4811);
nand U5280 (N_5280,N_4929,N_5028);
and U5281 (N_5281,N_4826,N_5037);
or U5282 (N_5282,N_4890,N_4915);
nand U5283 (N_5283,N_5018,N_4952);
xnor U5284 (N_5284,N_4834,N_5066);
nand U5285 (N_5285,N_4907,N_5039);
and U5286 (N_5286,N_5011,N_4877);
nand U5287 (N_5287,N_4945,N_5099);
xor U5288 (N_5288,N_4997,N_5084);
xnor U5289 (N_5289,N_5008,N_4906);
xor U5290 (N_5290,N_4883,N_5000);
xor U5291 (N_5291,N_4875,N_4803);
nand U5292 (N_5292,N_4968,N_4908);
nor U5293 (N_5293,N_5026,N_5062);
and U5294 (N_5294,N_4840,N_4847);
nor U5295 (N_5295,N_4815,N_5016);
or U5296 (N_5296,N_5020,N_5097);
and U5297 (N_5297,N_5003,N_4856);
or U5298 (N_5298,N_4973,N_5018);
and U5299 (N_5299,N_5059,N_4924);
and U5300 (N_5300,N_5011,N_4802);
or U5301 (N_5301,N_5073,N_5031);
nand U5302 (N_5302,N_5010,N_4885);
and U5303 (N_5303,N_4920,N_4871);
and U5304 (N_5304,N_4821,N_5053);
nand U5305 (N_5305,N_5094,N_5025);
and U5306 (N_5306,N_4874,N_4819);
xor U5307 (N_5307,N_4968,N_4994);
nor U5308 (N_5308,N_4921,N_4887);
nor U5309 (N_5309,N_4937,N_4877);
and U5310 (N_5310,N_5085,N_5032);
and U5311 (N_5311,N_5074,N_4857);
or U5312 (N_5312,N_4991,N_5072);
xor U5313 (N_5313,N_4998,N_5034);
or U5314 (N_5314,N_4809,N_4986);
nand U5315 (N_5315,N_4843,N_4857);
xnor U5316 (N_5316,N_4857,N_5012);
xor U5317 (N_5317,N_4992,N_5047);
or U5318 (N_5318,N_4876,N_4820);
and U5319 (N_5319,N_4962,N_4947);
nand U5320 (N_5320,N_5019,N_4854);
or U5321 (N_5321,N_4995,N_4945);
nand U5322 (N_5322,N_4914,N_4893);
xor U5323 (N_5323,N_5017,N_4959);
xnor U5324 (N_5324,N_4896,N_5026);
nand U5325 (N_5325,N_4801,N_4939);
nor U5326 (N_5326,N_5047,N_4924);
xor U5327 (N_5327,N_4983,N_4804);
nand U5328 (N_5328,N_4977,N_4900);
xnor U5329 (N_5329,N_4862,N_4878);
xnor U5330 (N_5330,N_4980,N_4807);
and U5331 (N_5331,N_4970,N_4993);
or U5332 (N_5332,N_4808,N_4985);
xnor U5333 (N_5333,N_5052,N_4940);
xnor U5334 (N_5334,N_4992,N_4832);
nor U5335 (N_5335,N_5004,N_4886);
and U5336 (N_5336,N_5063,N_4959);
nor U5337 (N_5337,N_4858,N_4924);
nor U5338 (N_5338,N_4990,N_4993);
or U5339 (N_5339,N_4995,N_4852);
nand U5340 (N_5340,N_4800,N_4962);
nand U5341 (N_5341,N_5047,N_5056);
xnor U5342 (N_5342,N_5012,N_5038);
nand U5343 (N_5343,N_5027,N_4930);
or U5344 (N_5344,N_4943,N_4891);
nand U5345 (N_5345,N_5008,N_5062);
nand U5346 (N_5346,N_5064,N_4977);
nor U5347 (N_5347,N_4834,N_4893);
or U5348 (N_5348,N_5050,N_4852);
nand U5349 (N_5349,N_5075,N_4867);
and U5350 (N_5350,N_5078,N_4860);
and U5351 (N_5351,N_4858,N_5037);
or U5352 (N_5352,N_5062,N_5033);
nand U5353 (N_5353,N_5034,N_4829);
or U5354 (N_5354,N_4905,N_4911);
nand U5355 (N_5355,N_5063,N_5087);
xor U5356 (N_5356,N_4918,N_5057);
nor U5357 (N_5357,N_4903,N_4999);
xor U5358 (N_5358,N_4899,N_4810);
or U5359 (N_5359,N_4802,N_4843);
or U5360 (N_5360,N_4845,N_4899);
xnor U5361 (N_5361,N_4850,N_4963);
or U5362 (N_5362,N_4919,N_4897);
nor U5363 (N_5363,N_4912,N_4926);
and U5364 (N_5364,N_5026,N_5010);
or U5365 (N_5365,N_5005,N_4945);
and U5366 (N_5366,N_4926,N_4996);
nand U5367 (N_5367,N_5096,N_4939);
nor U5368 (N_5368,N_4946,N_4933);
nor U5369 (N_5369,N_4931,N_4914);
and U5370 (N_5370,N_4818,N_4851);
and U5371 (N_5371,N_4944,N_5093);
and U5372 (N_5372,N_4833,N_4980);
and U5373 (N_5373,N_4988,N_4991);
and U5374 (N_5374,N_4995,N_5027);
and U5375 (N_5375,N_4942,N_4826);
nor U5376 (N_5376,N_4812,N_5059);
nand U5377 (N_5377,N_4923,N_5027);
and U5378 (N_5378,N_5014,N_4881);
xor U5379 (N_5379,N_4993,N_4828);
nor U5380 (N_5380,N_5092,N_5027);
xor U5381 (N_5381,N_4986,N_4827);
and U5382 (N_5382,N_5028,N_4953);
and U5383 (N_5383,N_5047,N_4900);
nor U5384 (N_5384,N_4832,N_4802);
nor U5385 (N_5385,N_4905,N_5032);
xor U5386 (N_5386,N_4932,N_4985);
nand U5387 (N_5387,N_4983,N_4965);
nor U5388 (N_5388,N_5086,N_4980);
nand U5389 (N_5389,N_4967,N_5006);
and U5390 (N_5390,N_4989,N_4859);
xnor U5391 (N_5391,N_4963,N_5004);
nor U5392 (N_5392,N_4937,N_5089);
xor U5393 (N_5393,N_4964,N_4808);
xor U5394 (N_5394,N_4864,N_4918);
xnor U5395 (N_5395,N_4886,N_4979);
and U5396 (N_5396,N_4931,N_4858);
and U5397 (N_5397,N_4859,N_5052);
xor U5398 (N_5398,N_5030,N_5047);
nor U5399 (N_5399,N_5054,N_4814);
xor U5400 (N_5400,N_5293,N_5285);
xnor U5401 (N_5401,N_5296,N_5182);
and U5402 (N_5402,N_5349,N_5327);
and U5403 (N_5403,N_5108,N_5256);
nor U5404 (N_5404,N_5211,N_5368);
nor U5405 (N_5405,N_5346,N_5394);
and U5406 (N_5406,N_5353,N_5376);
and U5407 (N_5407,N_5388,N_5371);
nand U5408 (N_5408,N_5221,N_5151);
nand U5409 (N_5409,N_5345,N_5137);
xnor U5410 (N_5410,N_5259,N_5319);
xnor U5411 (N_5411,N_5266,N_5145);
nand U5412 (N_5412,N_5250,N_5275);
xnor U5413 (N_5413,N_5372,N_5387);
and U5414 (N_5414,N_5391,N_5135);
nand U5415 (N_5415,N_5210,N_5140);
or U5416 (N_5416,N_5286,N_5240);
nor U5417 (N_5417,N_5272,N_5236);
xor U5418 (N_5418,N_5225,N_5183);
and U5419 (N_5419,N_5141,N_5320);
nor U5420 (N_5420,N_5191,N_5248);
nand U5421 (N_5421,N_5213,N_5118);
nand U5422 (N_5422,N_5334,N_5273);
and U5423 (N_5423,N_5129,N_5392);
xnor U5424 (N_5424,N_5157,N_5138);
and U5425 (N_5425,N_5350,N_5134);
or U5426 (N_5426,N_5190,N_5264);
xor U5427 (N_5427,N_5339,N_5174);
nor U5428 (N_5428,N_5245,N_5276);
and U5429 (N_5429,N_5215,N_5127);
or U5430 (N_5430,N_5364,N_5224);
xnor U5431 (N_5431,N_5366,N_5363);
or U5432 (N_5432,N_5374,N_5323);
nor U5433 (N_5433,N_5341,N_5208);
or U5434 (N_5434,N_5336,N_5186);
nor U5435 (N_5435,N_5283,N_5395);
nor U5436 (N_5436,N_5219,N_5197);
and U5437 (N_5437,N_5367,N_5315);
xnor U5438 (N_5438,N_5230,N_5185);
or U5439 (N_5439,N_5280,N_5270);
or U5440 (N_5440,N_5359,N_5122);
nor U5441 (N_5441,N_5389,N_5322);
xor U5442 (N_5442,N_5311,N_5321);
and U5443 (N_5443,N_5305,N_5284);
or U5444 (N_5444,N_5123,N_5136);
and U5445 (N_5445,N_5288,N_5238);
nand U5446 (N_5446,N_5379,N_5111);
nor U5447 (N_5447,N_5132,N_5106);
and U5448 (N_5448,N_5113,N_5310);
nand U5449 (N_5449,N_5365,N_5326);
xnor U5450 (N_5450,N_5206,N_5335);
nand U5451 (N_5451,N_5243,N_5119);
or U5452 (N_5452,N_5244,N_5258);
or U5453 (N_5453,N_5271,N_5189);
nand U5454 (N_5454,N_5205,N_5329);
or U5455 (N_5455,N_5342,N_5172);
and U5456 (N_5456,N_5229,N_5308);
xnor U5457 (N_5457,N_5198,N_5165);
and U5458 (N_5458,N_5159,N_5324);
and U5459 (N_5459,N_5214,N_5262);
xor U5460 (N_5460,N_5253,N_5314);
nor U5461 (N_5461,N_5139,N_5318);
and U5462 (N_5462,N_5166,N_5169);
nand U5463 (N_5463,N_5378,N_5187);
xor U5464 (N_5464,N_5161,N_5354);
and U5465 (N_5465,N_5199,N_5375);
or U5466 (N_5466,N_5218,N_5149);
nand U5467 (N_5467,N_5178,N_5393);
nor U5468 (N_5468,N_5184,N_5261);
or U5469 (N_5469,N_5175,N_5179);
and U5470 (N_5470,N_5239,N_5386);
or U5471 (N_5471,N_5398,N_5176);
or U5472 (N_5472,N_5124,N_5207);
or U5473 (N_5473,N_5130,N_5163);
or U5474 (N_5474,N_5233,N_5188);
nor U5475 (N_5475,N_5360,N_5298);
and U5476 (N_5476,N_5370,N_5337);
and U5477 (N_5477,N_5316,N_5116);
xor U5478 (N_5478,N_5103,N_5300);
xnor U5479 (N_5479,N_5201,N_5126);
nor U5480 (N_5480,N_5268,N_5144);
xor U5481 (N_5481,N_5196,N_5200);
and U5482 (N_5482,N_5269,N_5193);
and U5483 (N_5483,N_5146,N_5102);
and U5484 (N_5484,N_5249,N_5397);
nand U5485 (N_5485,N_5352,N_5306);
xnor U5486 (N_5486,N_5382,N_5154);
nand U5487 (N_5487,N_5343,N_5112);
and U5488 (N_5488,N_5192,N_5168);
nor U5489 (N_5489,N_5101,N_5361);
nand U5490 (N_5490,N_5309,N_5209);
and U5491 (N_5491,N_5155,N_5384);
and U5492 (N_5492,N_5235,N_5357);
xor U5493 (N_5493,N_5216,N_5332);
or U5494 (N_5494,N_5143,N_5381);
and U5495 (N_5495,N_5373,N_5297);
or U5496 (N_5496,N_5173,N_5125);
xor U5497 (N_5497,N_5330,N_5226);
or U5498 (N_5498,N_5195,N_5340);
xnor U5499 (N_5499,N_5278,N_5115);
nand U5500 (N_5500,N_5220,N_5133);
nor U5501 (N_5501,N_5162,N_5260);
or U5502 (N_5502,N_5114,N_5294);
or U5503 (N_5503,N_5302,N_5351);
xnor U5504 (N_5504,N_5328,N_5194);
xor U5505 (N_5505,N_5348,N_5105);
or U5506 (N_5506,N_5158,N_5100);
xnor U5507 (N_5507,N_5160,N_5304);
nor U5508 (N_5508,N_5274,N_5222);
or U5509 (N_5509,N_5299,N_5291);
nor U5510 (N_5510,N_5355,N_5109);
or U5511 (N_5511,N_5257,N_5252);
nand U5512 (N_5512,N_5234,N_5292);
and U5513 (N_5513,N_5121,N_5228);
and U5514 (N_5514,N_5241,N_5251);
and U5515 (N_5515,N_5344,N_5212);
nor U5516 (N_5516,N_5362,N_5347);
and U5517 (N_5517,N_5148,N_5279);
nand U5518 (N_5518,N_5203,N_5377);
nand U5519 (N_5519,N_5290,N_5277);
nor U5520 (N_5520,N_5153,N_5295);
nand U5521 (N_5521,N_5313,N_5325);
xnor U5522 (N_5522,N_5254,N_5170);
nor U5523 (N_5523,N_5171,N_5242);
and U5524 (N_5524,N_5289,N_5117);
and U5525 (N_5525,N_5142,N_5110);
and U5526 (N_5526,N_5307,N_5303);
xor U5527 (N_5527,N_5331,N_5217);
nor U5528 (N_5528,N_5204,N_5177);
and U5529 (N_5529,N_5152,N_5399);
or U5530 (N_5530,N_5131,N_5167);
and U5531 (N_5531,N_5107,N_5232);
nand U5532 (N_5532,N_5263,N_5380);
and U5533 (N_5533,N_5223,N_5147);
and U5534 (N_5534,N_5317,N_5120);
and U5535 (N_5535,N_5267,N_5202);
nand U5536 (N_5536,N_5255,N_5265);
nand U5537 (N_5537,N_5180,N_5231);
and U5538 (N_5538,N_5227,N_5156);
xnor U5539 (N_5539,N_5104,N_5333);
xnor U5540 (N_5540,N_5150,N_5287);
xnor U5541 (N_5541,N_5312,N_5246);
nor U5542 (N_5542,N_5385,N_5369);
xnor U5543 (N_5543,N_5390,N_5237);
and U5544 (N_5544,N_5301,N_5181);
and U5545 (N_5545,N_5128,N_5164);
nor U5546 (N_5546,N_5383,N_5247);
and U5547 (N_5547,N_5396,N_5358);
nor U5548 (N_5548,N_5356,N_5281);
nand U5549 (N_5549,N_5282,N_5338);
nor U5550 (N_5550,N_5193,N_5247);
and U5551 (N_5551,N_5256,N_5189);
nor U5552 (N_5552,N_5124,N_5152);
and U5553 (N_5553,N_5207,N_5292);
nor U5554 (N_5554,N_5130,N_5182);
nor U5555 (N_5555,N_5234,N_5377);
nand U5556 (N_5556,N_5360,N_5340);
and U5557 (N_5557,N_5120,N_5333);
nand U5558 (N_5558,N_5219,N_5295);
or U5559 (N_5559,N_5321,N_5169);
xnor U5560 (N_5560,N_5258,N_5378);
or U5561 (N_5561,N_5240,N_5199);
xor U5562 (N_5562,N_5219,N_5280);
nor U5563 (N_5563,N_5156,N_5192);
xnor U5564 (N_5564,N_5101,N_5208);
nand U5565 (N_5565,N_5158,N_5221);
xor U5566 (N_5566,N_5379,N_5332);
or U5567 (N_5567,N_5243,N_5304);
or U5568 (N_5568,N_5187,N_5230);
nor U5569 (N_5569,N_5286,N_5199);
and U5570 (N_5570,N_5106,N_5281);
or U5571 (N_5571,N_5321,N_5385);
nor U5572 (N_5572,N_5134,N_5229);
nand U5573 (N_5573,N_5289,N_5364);
nor U5574 (N_5574,N_5143,N_5380);
nor U5575 (N_5575,N_5391,N_5264);
nor U5576 (N_5576,N_5243,N_5259);
xor U5577 (N_5577,N_5252,N_5170);
nand U5578 (N_5578,N_5366,N_5223);
or U5579 (N_5579,N_5128,N_5224);
xnor U5580 (N_5580,N_5240,N_5185);
nor U5581 (N_5581,N_5333,N_5166);
xnor U5582 (N_5582,N_5349,N_5291);
nand U5583 (N_5583,N_5101,N_5191);
and U5584 (N_5584,N_5117,N_5166);
or U5585 (N_5585,N_5321,N_5292);
and U5586 (N_5586,N_5130,N_5109);
nor U5587 (N_5587,N_5373,N_5202);
and U5588 (N_5588,N_5151,N_5233);
nor U5589 (N_5589,N_5277,N_5265);
or U5590 (N_5590,N_5167,N_5199);
xor U5591 (N_5591,N_5186,N_5343);
or U5592 (N_5592,N_5312,N_5134);
nand U5593 (N_5593,N_5162,N_5380);
nor U5594 (N_5594,N_5247,N_5350);
nand U5595 (N_5595,N_5385,N_5119);
or U5596 (N_5596,N_5312,N_5227);
and U5597 (N_5597,N_5130,N_5372);
or U5598 (N_5598,N_5146,N_5398);
nor U5599 (N_5599,N_5274,N_5205);
nor U5600 (N_5600,N_5326,N_5191);
and U5601 (N_5601,N_5396,N_5381);
nor U5602 (N_5602,N_5279,N_5340);
nand U5603 (N_5603,N_5156,N_5108);
or U5604 (N_5604,N_5302,N_5156);
nor U5605 (N_5605,N_5242,N_5153);
and U5606 (N_5606,N_5161,N_5148);
and U5607 (N_5607,N_5300,N_5280);
nand U5608 (N_5608,N_5215,N_5255);
nor U5609 (N_5609,N_5228,N_5143);
or U5610 (N_5610,N_5144,N_5389);
xnor U5611 (N_5611,N_5372,N_5115);
nor U5612 (N_5612,N_5272,N_5176);
xor U5613 (N_5613,N_5341,N_5353);
nor U5614 (N_5614,N_5319,N_5115);
nor U5615 (N_5615,N_5234,N_5347);
xor U5616 (N_5616,N_5359,N_5235);
nand U5617 (N_5617,N_5341,N_5121);
and U5618 (N_5618,N_5268,N_5137);
and U5619 (N_5619,N_5324,N_5288);
nand U5620 (N_5620,N_5338,N_5329);
nand U5621 (N_5621,N_5165,N_5327);
xor U5622 (N_5622,N_5190,N_5312);
xnor U5623 (N_5623,N_5334,N_5354);
or U5624 (N_5624,N_5311,N_5341);
nand U5625 (N_5625,N_5259,N_5125);
or U5626 (N_5626,N_5152,N_5278);
or U5627 (N_5627,N_5122,N_5211);
nor U5628 (N_5628,N_5292,N_5262);
xor U5629 (N_5629,N_5381,N_5252);
or U5630 (N_5630,N_5386,N_5122);
or U5631 (N_5631,N_5229,N_5322);
or U5632 (N_5632,N_5342,N_5260);
xnor U5633 (N_5633,N_5210,N_5371);
and U5634 (N_5634,N_5263,N_5124);
xnor U5635 (N_5635,N_5300,N_5218);
xnor U5636 (N_5636,N_5259,N_5232);
xor U5637 (N_5637,N_5198,N_5292);
nand U5638 (N_5638,N_5294,N_5372);
and U5639 (N_5639,N_5139,N_5229);
or U5640 (N_5640,N_5262,N_5192);
xor U5641 (N_5641,N_5223,N_5144);
nand U5642 (N_5642,N_5195,N_5238);
nor U5643 (N_5643,N_5295,N_5290);
nand U5644 (N_5644,N_5249,N_5372);
and U5645 (N_5645,N_5168,N_5170);
xor U5646 (N_5646,N_5385,N_5160);
nand U5647 (N_5647,N_5119,N_5334);
or U5648 (N_5648,N_5348,N_5350);
nor U5649 (N_5649,N_5353,N_5227);
or U5650 (N_5650,N_5181,N_5204);
xnor U5651 (N_5651,N_5246,N_5273);
or U5652 (N_5652,N_5249,N_5295);
or U5653 (N_5653,N_5200,N_5318);
and U5654 (N_5654,N_5117,N_5154);
and U5655 (N_5655,N_5175,N_5110);
xor U5656 (N_5656,N_5144,N_5122);
and U5657 (N_5657,N_5360,N_5199);
nand U5658 (N_5658,N_5271,N_5365);
or U5659 (N_5659,N_5106,N_5302);
xor U5660 (N_5660,N_5287,N_5358);
or U5661 (N_5661,N_5124,N_5223);
xor U5662 (N_5662,N_5377,N_5112);
nor U5663 (N_5663,N_5182,N_5100);
nor U5664 (N_5664,N_5197,N_5328);
and U5665 (N_5665,N_5108,N_5209);
or U5666 (N_5666,N_5229,N_5180);
or U5667 (N_5667,N_5208,N_5229);
and U5668 (N_5668,N_5138,N_5121);
or U5669 (N_5669,N_5165,N_5224);
xnor U5670 (N_5670,N_5389,N_5131);
xor U5671 (N_5671,N_5252,N_5309);
xor U5672 (N_5672,N_5325,N_5264);
nand U5673 (N_5673,N_5156,N_5288);
or U5674 (N_5674,N_5284,N_5237);
xor U5675 (N_5675,N_5316,N_5312);
and U5676 (N_5676,N_5147,N_5391);
nand U5677 (N_5677,N_5222,N_5297);
and U5678 (N_5678,N_5275,N_5194);
xor U5679 (N_5679,N_5167,N_5235);
nand U5680 (N_5680,N_5374,N_5152);
xor U5681 (N_5681,N_5128,N_5267);
or U5682 (N_5682,N_5138,N_5384);
nand U5683 (N_5683,N_5242,N_5234);
nand U5684 (N_5684,N_5296,N_5218);
xor U5685 (N_5685,N_5238,N_5292);
or U5686 (N_5686,N_5282,N_5350);
xor U5687 (N_5687,N_5135,N_5313);
or U5688 (N_5688,N_5390,N_5171);
nand U5689 (N_5689,N_5346,N_5173);
xnor U5690 (N_5690,N_5190,N_5160);
xor U5691 (N_5691,N_5208,N_5174);
nor U5692 (N_5692,N_5385,N_5224);
nor U5693 (N_5693,N_5278,N_5376);
or U5694 (N_5694,N_5378,N_5367);
or U5695 (N_5695,N_5113,N_5196);
and U5696 (N_5696,N_5250,N_5225);
and U5697 (N_5697,N_5112,N_5296);
nor U5698 (N_5698,N_5160,N_5248);
and U5699 (N_5699,N_5310,N_5254);
nand U5700 (N_5700,N_5417,N_5644);
and U5701 (N_5701,N_5668,N_5457);
nor U5702 (N_5702,N_5578,N_5497);
or U5703 (N_5703,N_5597,N_5520);
nand U5704 (N_5704,N_5553,N_5413);
or U5705 (N_5705,N_5483,N_5408);
nor U5706 (N_5706,N_5546,N_5521);
nor U5707 (N_5707,N_5515,N_5599);
xnor U5708 (N_5708,N_5551,N_5486);
xnor U5709 (N_5709,N_5509,N_5536);
nor U5710 (N_5710,N_5460,N_5428);
and U5711 (N_5711,N_5659,N_5463);
xnor U5712 (N_5712,N_5568,N_5580);
and U5713 (N_5713,N_5502,N_5446);
xor U5714 (N_5714,N_5518,N_5665);
nand U5715 (N_5715,N_5444,N_5441);
nand U5716 (N_5716,N_5697,N_5484);
nor U5717 (N_5717,N_5436,N_5654);
nand U5718 (N_5718,N_5699,N_5577);
nand U5719 (N_5719,N_5545,N_5439);
nor U5720 (N_5720,N_5588,N_5661);
nand U5721 (N_5721,N_5527,N_5636);
or U5722 (N_5722,N_5513,N_5523);
or U5723 (N_5723,N_5626,N_5566);
and U5724 (N_5724,N_5487,N_5564);
xor U5725 (N_5725,N_5603,N_5563);
nor U5726 (N_5726,N_5456,N_5503);
nand U5727 (N_5727,N_5669,N_5570);
and U5728 (N_5728,N_5627,N_5500);
and U5729 (N_5729,N_5405,N_5572);
xor U5730 (N_5730,N_5681,N_5574);
nor U5731 (N_5731,N_5511,N_5620);
and U5732 (N_5732,N_5586,N_5579);
and U5733 (N_5733,N_5475,N_5535);
nor U5734 (N_5734,N_5696,N_5554);
or U5735 (N_5735,N_5604,N_5429);
nand U5736 (N_5736,N_5512,N_5453);
nor U5737 (N_5737,N_5581,N_5465);
and U5738 (N_5738,N_5610,N_5506);
or U5739 (N_5739,N_5476,N_5671);
xnor U5740 (N_5740,N_5537,N_5492);
and U5741 (N_5741,N_5589,N_5473);
nor U5742 (N_5742,N_5414,N_5623);
or U5743 (N_5743,N_5534,N_5609);
xnor U5744 (N_5744,N_5698,N_5451);
nand U5745 (N_5745,N_5538,N_5662);
nand U5746 (N_5746,N_5496,N_5433);
xor U5747 (N_5747,N_5533,N_5448);
and U5748 (N_5748,N_5642,N_5504);
nand U5749 (N_5749,N_5479,N_5495);
nor U5750 (N_5750,N_5582,N_5647);
xor U5751 (N_5751,N_5440,N_5633);
or U5752 (N_5752,N_5641,N_5525);
nor U5753 (N_5753,N_5548,N_5555);
and U5754 (N_5754,N_5556,N_5587);
xor U5755 (N_5755,N_5438,N_5672);
xnor U5756 (N_5756,N_5423,N_5516);
or U5757 (N_5757,N_5605,N_5445);
xnor U5758 (N_5758,N_5685,N_5459);
xor U5759 (N_5759,N_5667,N_5424);
or U5760 (N_5760,N_5557,N_5474);
and U5761 (N_5761,N_5655,N_5666);
and U5762 (N_5762,N_5540,N_5422);
and U5763 (N_5763,N_5567,N_5634);
or U5764 (N_5764,N_5443,N_5591);
xor U5765 (N_5765,N_5645,N_5585);
xnor U5766 (N_5766,N_5539,N_5409);
xnor U5767 (N_5767,N_5675,N_5430);
or U5768 (N_5768,N_5420,N_5435);
or U5769 (N_5769,N_5528,N_5690);
nand U5770 (N_5770,N_5426,N_5462);
and U5771 (N_5771,N_5499,N_5652);
nor U5772 (N_5772,N_5571,N_5622);
xor U5773 (N_5773,N_5600,N_5411);
and U5774 (N_5774,N_5469,N_5449);
xnor U5775 (N_5775,N_5559,N_5421);
nor U5776 (N_5776,N_5592,N_5618);
and U5777 (N_5777,N_5526,N_5478);
or U5778 (N_5778,N_5573,N_5606);
nor U5779 (N_5779,N_5455,N_5544);
and U5780 (N_5780,N_5458,N_5507);
nor U5781 (N_5781,N_5517,N_5615);
nor U5782 (N_5782,N_5648,N_5454);
xor U5783 (N_5783,N_5619,N_5468);
nand U5784 (N_5784,N_5691,N_5638);
and U5785 (N_5785,N_5561,N_5470);
or U5786 (N_5786,N_5531,N_5562);
nand U5787 (N_5787,N_5416,N_5410);
or U5788 (N_5788,N_5480,N_5649);
or U5789 (N_5789,N_5432,N_5658);
nand U5790 (N_5790,N_5498,N_5575);
nor U5791 (N_5791,N_5508,N_5660);
nand U5792 (N_5792,N_5694,N_5437);
and U5793 (N_5793,N_5519,N_5447);
nand U5794 (N_5794,N_5631,N_5682);
xnor U5795 (N_5795,N_5481,N_5677);
and U5796 (N_5796,N_5558,N_5529);
xor U5797 (N_5797,N_5689,N_5621);
or U5798 (N_5798,N_5412,N_5630);
and U5799 (N_5799,N_5402,N_5673);
or U5800 (N_5800,N_5612,N_5679);
xor U5801 (N_5801,N_5400,N_5617);
and U5802 (N_5802,N_5530,N_5688);
nand U5803 (N_5803,N_5657,N_5493);
nor U5804 (N_5804,N_5595,N_5425);
xor U5805 (N_5805,N_5646,N_5549);
and U5806 (N_5806,N_5650,N_5532);
and U5807 (N_5807,N_5404,N_5543);
and U5808 (N_5808,N_5467,N_5635);
nor U5809 (N_5809,N_5602,N_5637);
or U5810 (N_5810,N_5678,N_5427);
and U5811 (N_5811,N_5663,N_5550);
nor U5812 (N_5812,N_5505,N_5401);
and U5813 (N_5813,N_5489,N_5692);
or U5814 (N_5814,N_5541,N_5524);
xor U5815 (N_5815,N_5431,N_5674);
nand U5816 (N_5816,N_5643,N_5596);
and U5817 (N_5817,N_5461,N_5434);
nand U5818 (N_5818,N_5683,N_5466);
and U5819 (N_5819,N_5452,N_5613);
and U5820 (N_5820,N_5485,N_5501);
nand U5821 (N_5821,N_5542,N_5607);
nor U5822 (N_5822,N_5639,N_5472);
nor U5823 (N_5823,N_5680,N_5418);
nand U5824 (N_5824,N_5695,N_5624);
nand U5825 (N_5825,N_5601,N_5583);
and U5826 (N_5826,N_5611,N_5614);
and U5827 (N_5827,N_5415,N_5514);
and U5828 (N_5828,N_5488,N_5593);
nor U5829 (N_5829,N_5464,N_5406);
nand U5830 (N_5830,N_5594,N_5584);
nand U5831 (N_5831,N_5552,N_5419);
xnor U5832 (N_5832,N_5576,N_5522);
and U5833 (N_5833,N_5664,N_5616);
and U5834 (N_5834,N_5450,N_5590);
and U5835 (N_5835,N_5670,N_5640);
xor U5836 (N_5836,N_5471,N_5653);
nor U5837 (N_5837,N_5684,N_5407);
and U5838 (N_5838,N_5560,N_5565);
and U5839 (N_5839,N_5629,N_5687);
nand U5840 (N_5840,N_5686,N_5632);
or U5841 (N_5841,N_5656,N_5598);
xor U5842 (N_5842,N_5490,N_5477);
or U5843 (N_5843,N_5510,N_5693);
or U5844 (N_5844,N_5651,N_5403);
and U5845 (N_5845,N_5494,N_5676);
nor U5846 (N_5846,N_5547,N_5491);
or U5847 (N_5847,N_5625,N_5608);
or U5848 (N_5848,N_5482,N_5569);
or U5849 (N_5849,N_5442,N_5628);
nand U5850 (N_5850,N_5568,N_5517);
nand U5851 (N_5851,N_5431,N_5570);
xor U5852 (N_5852,N_5467,N_5455);
or U5853 (N_5853,N_5597,N_5477);
nand U5854 (N_5854,N_5439,N_5429);
or U5855 (N_5855,N_5516,N_5513);
xnor U5856 (N_5856,N_5566,N_5508);
nand U5857 (N_5857,N_5462,N_5579);
and U5858 (N_5858,N_5542,N_5626);
or U5859 (N_5859,N_5553,N_5563);
or U5860 (N_5860,N_5428,N_5484);
or U5861 (N_5861,N_5656,N_5586);
xnor U5862 (N_5862,N_5591,N_5503);
nor U5863 (N_5863,N_5466,N_5591);
or U5864 (N_5864,N_5638,N_5635);
xor U5865 (N_5865,N_5679,N_5672);
and U5866 (N_5866,N_5445,N_5595);
xnor U5867 (N_5867,N_5445,N_5450);
nand U5868 (N_5868,N_5564,N_5523);
and U5869 (N_5869,N_5484,N_5457);
nor U5870 (N_5870,N_5676,N_5465);
nand U5871 (N_5871,N_5631,N_5400);
nor U5872 (N_5872,N_5438,N_5636);
nor U5873 (N_5873,N_5672,N_5625);
or U5874 (N_5874,N_5622,N_5582);
or U5875 (N_5875,N_5518,N_5607);
xor U5876 (N_5876,N_5609,N_5634);
nand U5877 (N_5877,N_5512,N_5500);
nand U5878 (N_5878,N_5595,N_5622);
nor U5879 (N_5879,N_5557,N_5625);
or U5880 (N_5880,N_5692,N_5440);
nand U5881 (N_5881,N_5523,N_5594);
and U5882 (N_5882,N_5412,N_5420);
and U5883 (N_5883,N_5631,N_5673);
nor U5884 (N_5884,N_5550,N_5464);
and U5885 (N_5885,N_5444,N_5523);
and U5886 (N_5886,N_5575,N_5640);
or U5887 (N_5887,N_5417,N_5567);
nor U5888 (N_5888,N_5589,N_5513);
or U5889 (N_5889,N_5545,N_5452);
and U5890 (N_5890,N_5563,N_5401);
and U5891 (N_5891,N_5560,N_5687);
nor U5892 (N_5892,N_5684,N_5641);
nor U5893 (N_5893,N_5592,N_5512);
and U5894 (N_5894,N_5603,N_5458);
and U5895 (N_5895,N_5517,N_5509);
xnor U5896 (N_5896,N_5468,N_5656);
nand U5897 (N_5897,N_5622,N_5664);
nand U5898 (N_5898,N_5643,N_5681);
nand U5899 (N_5899,N_5634,N_5664);
or U5900 (N_5900,N_5571,N_5510);
and U5901 (N_5901,N_5585,N_5456);
nand U5902 (N_5902,N_5593,N_5501);
xnor U5903 (N_5903,N_5455,N_5642);
nand U5904 (N_5904,N_5556,N_5675);
or U5905 (N_5905,N_5602,N_5434);
nand U5906 (N_5906,N_5608,N_5578);
nor U5907 (N_5907,N_5495,N_5695);
and U5908 (N_5908,N_5680,N_5582);
and U5909 (N_5909,N_5482,N_5529);
nand U5910 (N_5910,N_5451,N_5591);
nand U5911 (N_5911,N_5579,N_5426);
nand U5912 (N_5912,N_5627,N_5607);
nor U5913 (N_5913,N_5415,N_5609);
nand U5914 (N_5914,N_5641,N_5537);
xnor U5915 (N_5915,N_5466,N_5462);
and U5916 (N_5916,N_5545,N_5448);
nand U5917 (N_5917,N_5632,N_5677);
or U5918 (N_5918,N_5411,N_5509);
xnor U5919 (N_5919,N_5422,N_5616);
xnor U5920 (N_5920,N_5403,N_5446);
nand U5921 (N_5921,N_5440,N_5661);
xor U5922 (N_5922,N_5424,N_5695);
or U5923 (N_5923,N_5646,N_5612);
nand U5924 (N_5924,N_5526,N_5403);
nor U5925 (N_5925,N_5673,N_5633);
nor U5926 (N_5926,N_5579,N_5627);
xor U5927 (N_5927,N_5559,N_5598);
or U5928 (N_5928,N_5683,N_5644);
nand U5929 (N_5929,N_5616,N_5689);
xnor U5930 (N_5930,N_5504,N_5454);
and U5931 (N_5931,N_5522,N_5678);
or U5932 (N_5932,N_5591,N_5429);
xor U5933 (N_5933,N_5500,N_5624);
and U5934 (N_5934,N_5499,N_5416);
and U5935 (N_5935,N_5475,N_5623);
nor U5936 (N_5936,N_5661,N_5498);
xnor U5937 (N_5937,N_5647,N_5553);
or U5938 (N_5938,N_5425,N_5602);
xor U5939 (N_5939,N_5584,N_5549);
nand U5940 (N_5940,N_5405,N_5469);
or U5941 (N_5941,N_5437,N_5645);
and U5942 (N_5942,N_5513,N_5419);
or U5943 (N_5943,N_5615,N_5523);
or U5944 (N_5944,N_5684,N_5416);
nand U5945 (N_5945,N_5447,N_5520);
and U5946 (N_5946,N_5406,N_5504);
or U5947 (N_5947,N_5407,N_5629);
nor U5948 (N_5948,N_5542,N_5664);
or U5949 (N_5949,N_5423,N_5411);
and U5950 (N_5950,N_5557,N_5617);
or U5951 (N_5951,N_5486,N_5451);
xnor U5952 (N_5952,N_5696,N_5561);
nand U5953 (N_5953,N_5662,N_5499);
xnor U5954 (N_5954,N_5583,N_5509);
or U5955 (N_5955,N_5535,N_5522);
nor U5956 (N_5956,N_5486,N_5466);
xor U5957 (N_5957,N_5651,N_5486);
and U5958 (N_5958,N_5453,N_5440);
xor U5959 (N_5959,N_5645,N_5581);
and U5960 (N_5960,N_5496,N_5541);
xor U5961 (N_5961,N_5433,N_5645);
and U5962 (N_5962,N_5405,N_5644);
nor U5963 (N_5963,N_5409,N_5556);
xor U5964 (N_5964,N_5466,N_5611);
xnor U5965 (N_5965,N_5434,N_5453);
nor U5966 (N_5966,N_5548,N_5480);
or U5967 (N_5967,N_5416,N_5419);
nor U5968 (N_5968,N_5607,N_5610);
or U5969 (N_5969,N_5583,N_5671);
and U5970 (N_5970,N_5451,N_5466);
xor U5971 (N_5971,N_5596,N_5406);
nand U5972 (N_5972,N_5413,N_5560);
nand U5973 (N_5973,N_5601,N_5444);
nand U5974 (N_5974,N_5601,N_5572);
and U5975 (N_5975,N_5433,N_5536);
nor U5976 (N_5976,N_5402,N_5618);
nand U5977 (N_5977,N_5414,N_5619);
xor U5978 (N_5978,N_5576,N_5487);
nor U5979 (N_5979,N_5524,N_5434);
nand U5980 (N_5980,N_5654,N_5683);
nand U5981 (N_5981,N_5609,N_5541);
or U5982 (N_5982,N_5576,N_5506);
or U5983 (N_5983,N_5670,N_5563);
nand U5984 (N_5984,N_5449,N_5437);
or U5985 (N_5985,N_5684,N_5588);
nor U5986 (N_5986,N_5521,N_5421);
xnor U5987 (N_5987,N_5465,N_5423);
nor U5988 (N_5988,N_5602,N_5406);
nand U5989 (N_5989,N_5536,N_5605);
and U5990 (N_5990,N_5466,N_5672);
and U5991 (N_5991,N_5597,N_5641);
and U5992 (N_5992,N_5671,N_5529);
xor U5993 (N_5993,N_5425,N_5601);
or U5994 (N_5994,N_5437,N_5447);
nor U5995 (N_5995,N_5574,N_5653);
nor U5996 (N_5996,N_5474,N_5446);
xor U5997 (N_5997,N_5698,N_5633);
and U5998 (N_5998,N_5429,N_5609);
nand U5999 (N_5999,N_5584,N_5672);
or U6000 (N_6000,N_5900,N_5918);
nor U6001 (N_6001,N_5733,N_5819);
nand U6002 (N_6002,N_5894,N_5903);
nand U6003 (N_6003,N_5947,N_5969);
or U6004 (N_6004,N_5796,N_5888);
xnor U6005 (N_6005,N_5791,N_5716);
or U6006 (N_6006,N_5766,N_5990);
and U6007 (N_6007,N_5767,N_5868);
or U6008 (N_6008,N_5797,N_5778);
or U6009 (N_6009,N_5787,N_5745);
nor U6010 (N_6010,N_5963,N_5960);
and U6011 (N_6011,N_5723,N_5709);
and U6012 (N_6012,N_5758,N_5887);
nor U6013 (N_6013,N_5884,N_5744);
and U6014 (N_6014,N_5817,N_5964);
xor U6015 (N_6015,N_5989,N_5768);
nor U6016 (N_6016,N_5911,N_5818);
or U6017 (N_6017,N_5908,N_5852);
or U6018 (N_6018,N_5798,N_5851);
or U6019 (N_6019,N_5764,N_5961);
nor U6020 (N_6020,N_5899,N_5777);
xnor U6021 (N_6021,N_5831,N_5741);
xnor U6022 (N_6022,N_5898,N_5905);
nand U6023 (N_6023,N_5932,N_5742);
nor U6024 (N_6024,N_5855,N_5986);
or U6025 (N_6025,N_5984,N_5843);
xnor U6026 (N_6026,N_5750,N_5922);
xor U6027 (N_6027,N_5846,N_5902);
or U6028 (N_6028,N_5953,N_5861);
nor U6029 (N_6029,N_5925,N_5746);
or U6030 (N_6030,N_5949,N_5747);
or U6031 (N_6031,N_5774,N_5734);
xnor U6032 (N_6032,N_5789,N_5836);
and U6033 (N_6033,N_5776,N_5948);
nand U6034 (N_6034,N_5783,N_5815);
and U6035 (N_6035,N_5935,N_5939);
and U6036 (N_6036,N_5755,N_5965);
xor U6037 (N_6037,N_5972,N_5840);
or U6038 (N_6038,N_5916,N_5743);
nor U6039 (N_6039,N_5890,N_5950);
nand U6040 (N_6040,N_5822,N_5848);
nor U6041 (N_6041,N_5813,N_5700);
and U6042 (N_6042,N_5999,N_5865);
or U6043 (N_6043,N_5993,N_5904);
or U6044 (N_6044,N_5892,N_5837);
xnor U6045 (N_6045,N_5872,N_5717);
xor U6046 (N_6046,N_5863,N_5866);
xor U6047 (N_6047,N_5858,N_5748);
and U6048 (N_6048,N_5707,N_5856);
or U6049 (N_6049,N_5775,N_5944);
or U6050 (N_6050,N_5847,N_5886);
nor U6051 (N_6051,N_5977,N_5906);
xnor U6052 (N_6052,N_5940,N_5729);
nand U6053 (N_6053,N_5907,N_5930);
nor U6054 (N_6054,N_5967,N_5811);
nor U6055 (N_6055,N_5844,N_5761);
xnor U6056 (N_6056,N_5952,N_5980);
and U6057 (N_6057,N_5973,N_5945);
nor U6058 (N_6058,N_5955,N_5715);
nor U6059 (N_6059,N_5937,N_5749);
nand U6060 (N_6060,N_5941,N_5857);
xor U6061 (N_6061,N_5769,N_5954);
or U6062 (N_6062,N_5985,N_5735);
nand U6063 (N_6063,N_5800,N_5966);
nand U6064 (N_6064,N_5752,N_5701);
xor U6065 (N_6065,N_5860,N_5909);
nand U6066 (N_6066,N_5958,N_5728);
or U6067 (N_6067,N_5706,N_5859);
or U6068 (N_6068,N_5740,N_5738);
or U6069 (N_6069,N_5880,N_5825);
or U6070 (N_6070,N_5810,N_5779);
or U6071 (N_6071,N_5968,N_5996);
xor U6072 (N_6072,N_5792,N_5849);
xnor U6073 (N_6073,N_5875,N_5923);
nand U6074 (N_6074,N_5754,N_5942);
nand U6075 (N_6075,N_5995,N_5921);
xor U6076 (N_6076,N_5771,N_5917);
xnor U6077 (N_6077,N_5951,N_5959);
nand U6078 (N_6078,N_5871,N_5876);
or U6079 (N_6079,N_5893,N_5896);
xor U6080 (N_6080,N_5920,N_5946);
and U6081 (N_6081,N_5877,N_5897);
and U6082 (N_6082,N_5773,N_5814);
and U6083 (N_6083,N_5727,N_5801);
nand U6084 (N_6084,N_5895,N_5933);
nor U6085 (N_6085,N_5807,N_5998);
xor U6086 (N_6086,N_5915,N_5820);
nand U6087 (N_6087,N_5703,N_5957);
xnor U6088 (N_6088,N_5845,N_5806);
xor U6089 (N_6089,N_5794,N_5816);
xor U6090 (N_6090,N_5710,N_5850);
and U6091 (N_6091,N_5823,N_5883);
nand U6092 (N_6092,N_5912,N_5782);
and U6093 (N_6093,N_5714,N_5943);
and U6094 (N_6094,N_5987,N_5913);
xnor U6095 (N_6095,N_5736,N_5828);
xnor U6096 (N_6096,N_5838,N_5862);
or U6097 (N_6097,N_5757,N_5722);
and U6098 (N_6098,N_5759,N_5718);
nand U6099 (N_6099,N_5751,N_5803);
and U6100 (N_6100,N_5730,N_5982);
and U6101 (N_6101,N_5780,N_5867);
or U6102 (N_6102,N_5731,N_5981);
nand U6103 (N_6103,N_5802,N_5784);
and U6104 (N_6104,N_5914,N_5991);
xor U6105 (N_6105,N_5885,N_5756);
or U6106 (N_6106,N_5997,N_5970);
or U6107 (N_6107,N_5938,N_5910);
or U6108 (N_6108,N_5835,N_5962);
nor U6109 (N_6109,N_5889,N_5864);
nand U6110 (N_6110,N_5971,N_5719);
nor U6111 (N_6111,N_5869,N_5781);
xor U6112 (N_6112,N_5874,N_5702);
nor U6113 (N_6113,N_5826,N_5901);
nor U6114 (N_6114,N_5708,N_5732);
nand U6115 (N_6115,N_5809,N_5934);
or U6116 (N_6116,N_5878,N_5786);
and U6117 (N_6117,N_5931,N_5853);
or U6118 (N_6118,N_5790,N_5979);
nand U6119 (N_6119,N_5832,N_5808);
xor U6120 (N_6120,N_5927,N_5882);
nand U6121 (N_6121,N_5737,N_5704);
nor U6122 (N_6122,N_5926,N_5873);
or U6123 (N_6123,N_5721,N_5725);
or U6124 (N_6124,N_5919,N_5712);
and U6125 (N_6125,N_5770,N_5724);
nand U6126 (N_6126,N_5929,N_5924);
and U6127 (N_6127,N_5833,N_5726);
or U6128 (N_6128,N_5763,N_5928);
xor U6129 (N_6129,N_5974,N_5936);
or U6130 (N_6130,N_5983,N_5793);
nor U6131 (N_6131,N_5760,N_5834);
or U6132 (N_6132,N_5804,N_5891);
nand U6133 (N_6133,N_5720,N_5881);
xor U6134 (N_6134,N_5854,N_5799);
nand U6135 (N_6135,N_5879,N_5842);
or U6136 (N_6136,N_5795,N_5788);
nor U6137 (N_6137,N_5824,N_5765);
nor U6138 (N_6138,N_5713,N_5978);
nand U6139 (N_6139,N_5812,N_5994);
and U6140 (N_6140,N_5841,N_5821);
nor U6141 (N_6141,N_5976,N_5711);
nor U6142 (N_6142,N_5827,N_5772);
nor U6143 (N_6143,N_5956,N_5705);
or U6144 (N_6144,N_5785,N_5805);
and U6145 (N_6145,N_5839,N_5829);
nand U6146 (N_6146,N_5830,N_5988);
nand U6147 (N_6147,N_5975,N_5992);
nand U6148 (N_6148,N_5870,N_5762);
nand U6149 (N_6149,N_5753,N_5739);
xnor U6150 (N_6150,N_5923,N_5913);
and U6151 (N_6151,N_5753,N_5794);
or U6152 (N_6152,N_5929,N_5831);
and U6153 (N_6153,N_5823,N_5925);
nor U6154 (N_6154,N_5859,N_5813);
xnor U6155 (N_6155,N_5913,N_5944);
nand U6156 (N_6156,N_5947,N_5973);
or U6157 (N_6157,N_5928,N_5810);
or U6158 (N_6158,N_5749,N_5720);
nor U6159 (N_6159,N_5804,N_5726);
xor U6160 (N_6160,N_5867,N_5766);
nand U6161 (N_6161,N_5920,N_5840);
and U6162 (N_6162,N_5990,N_5779);
nor U6163 (N_6163,N_5986,N_5998);
xor U6164 (N_6164,N_5944,N_5703);
and U6165 (N_6165,N_5950,N_5861);
xor U6166 (N_6166,N_5876,N_5904);
nand U6167 (N_6167,N_5769,N_5908);
xor U6168 (N_6168,N_5717,N_5929);
xnor U6169 (N_6169,N_5727,N_5872);
nor U6170 (N_6170,N_5908,N_5731);
and U6171 (N_6171,N_5972,N_5987);
xnor U6172 (N_6172,N_5874,N_5934);
or U6173 (N_6173,N_5900,N_5952);
nor U6174 (N_6174,N_5700,N_5726);
and U6175 (N_6175,N_5756,N_5866);
nor U6176 (N_6176,N_5815,N_5934);
and U6177 (N_6177,N_5714,N_5919);
or U6178 (N_6178,N_5866,N_5914);
nand U6179 (N_6179,N_5743,N_5940);
xor U6180 (N_6180,N_5934,N_5966);
and U6181 (N_6181,N_5893,N_5901);
xor U6182 (N_6182,N_5767,N_5709);
nand U6183 (N_6183,N_5879,N_5886);
nor U6184 (N_6184,N_5858,N_5863);
and U6185 (N_6185,N_5980,N_5769);
nor U6186 (N_6186,N_5798,N_5818);
or U6187 (N_6187,N_5858,N_5725);
xor U6188 (N_6188,N_5951,N_5800);
or U6189 (N_6189,N_5901,N_5957);
and U6190 (N_6190,N_5778,N_5903);
and U6191 (N_6191,N_5991,N_5903);
nor U6192 (N_6192,N_5985,N_5770);
or U6193 (N_6193,N_5737,N_5904);
nand U6194 (N_6194,N_5701,N_5824);
nor U6195 (N_6195,N_5941,N_5865);
nor U6196 (N_6196,N_5896,N_5879);
nor U6197 (N_6197,N_5818,N_5969);
nand U6198 (N_6198,N_5922,N_5825);
and U6199 (N_6199,N_5866,N_5842);
nand U6200 (N_6200,N_5746,N_5871);
and U6201 (N_6201,N_5805,N_5743);
nor U6202 (N_6202,N_5801,N_5793);
nand U6203 (N_6203,N_5830,N_5877);
xnor U6204 (N_6204,N_5864,N_5727);
nand U6205 (N_6205,N_5850,N_5886);
or U6206 (N_6206,N_5913,N_5710);
xnor U6207 (N_6207,N_5913,N_5850);
nor U6208 (N_6208,N_5975,N_5951);
and U6209 (N_6209,N_5868,N_5798);
nor U6210 (N_6210,N_5981,N_5843);
and U6211 (N_6211,N_5702,N_5813);
nor U6212 (N_6212,N_5844,N_5936);
xnor U6213 (N_6213,N_5804,N_5958);
nor U6214 (N_6214,N_5877,N_5828);
nand U6215 (N_6215,N_5775,N_5926);
and U6216 (N_6216,N_5702,N_5806);
or U6217 (N_6217,N_5705,N_5788);
nor U6218 (N_6218,N_5880,N_5765);
or U6219 (N_6219,N_5876,N_5716);
nor U6220 (N_6220,N_5821,N_5743);
nand U6221 (N_6221,N_5907,N_5747);
xnor U6222 (N_6222,N_5760,N_5764);
nand U6223 (N_6223,N_5790,N_5756);
nor U6224 (N_6224,N_5865,N_5954);
and U6225 (N_6225,N_5829,N_5739);
and U6226 (N_6226,N_5976,N_5916);
or U6227 (N_6227,N_5955,N_5925);
nor U6228 (N_6228,N_5726,N_5959);
or U6229 (N_6229,N_5711,N_5848);
xnor U6230 (N_6230,N_5848,N_5749);
nor U6231 (N_6231,N_5748,N_5777);
nor U6232 (N_6232,N_5930,N_5775);
xor U6233 (N_6233,N_5919,N_5965);
and U6234 (N_6234,N_5794,N_5979);
nor U6235 (N_6235,N_5840,N_5789);
nor U6236 (N_6236,N_5792,N_5776);
nor U6237 (N_6237,N_5924,N_5981);
xnor U6238 (N_6238,N_5833,N_5832);
and U6239 (N_6239,N_5907,N_5870);
xnor U6240 (N_6240,N_5982,N_5921);
or U6241 (N_6241,N_5948,N_5887);
nor U6242 (N_6242,N_5852,N_5932);
and U6243 (N_6243,N_5925,N_5731);
or U6244 (N_6244,N_5751,N_5890);
xnor U6245 (N_6245,N_5787,N_5811);
nand U6246 (N_6246,N_5885,N_5803);
xnor U6247 (N_6247,N_5931,N_5942);
nor U6248 (N_6248,N_5782,N_5787);
xor U6249 (N_6249,N_5959,N_5714);
xor U6250 (N_6250,N_5724,N_5952);
and U6251 (N_6251,N_5783,N_5827);
nand U6252 (N_6252,N_5834,N_5982);
nand U6253 (N_6253,N_5875,N_5807);
nor U6254 (N_6254,N_5726,N_5975);
nor U6255 (N_6255,N_5709,N_5887);
nand U6256 (N_6256,N_5831,N_5774);
and U6257 (N_6257,N_5806,N_5999);
and U6258 (N_6258,N_5881,N_5716);
or U6259 (N_6259,N_5703,N_5732);
or U6260 (N_6260,N_5711,N_5859);
and U6261 (N_6261,N_5818,N_5714);
nor U6262 (N_6262,N_5812,N_5766);
and U6263 (N_6263,N_5988,N_5852);
or U6264 (N_6264,N_5805,N_5907);
nand U6265 (N_6265,N_5786,N_5796);
nand U6266 (N_6266,N_5794,N_5838);
xor U6267 (N_6267,N_5882,N_5792);
nor U6268 (N_6268,N_5974,N_5766);
nor U6269 (N_6269,N_5874,N_5706);
or U6270 (N_6270,N_5958,N_5873);
xor U6271 (N_6271,N_5903,N_5858);
nand U6272 (N_6272,N_5966,N_5962);
or U6273 (N_6273,N_5900,N_5916);
xnor U6274 (N_6274,N_5818,N_5762);
nor U6275 (N_6275,N_5736,N_5796);
and U6276 (N_6276,N_5980,N_5993);
xor U6277 (N_6277,N_5830,N_5891);
nor U6278 (N_6278,N_5936,N_5716);
nor U6279 (N_6279,N_5809,N_5816);
or U6280 (N_6280,N_5818,N_5722);
and U6281 (N_6281,N_5781,N_5926);
xnor U6282 (N_6282,N_5845,N_5814);
xnor U6283 (N_6283,N_5894,N_5925);
xor U6284 (N_6284,N_5931,N_5848);
nor U6285 (N_6285,N_5748,N_5962);
nand U6286 (N_6286,N_5953,N_5941);
and U6287 (N_6287,N_5921,N_5833);
xnor U6288 (N_6288,N_5854,N_5889);
nor U6289 (N_6289,N_5755,N_5963);
xor U6290 (N_6290,N_5865,N_5825);
and U6291 (N_6291,N_5843,N_5792);
or U6292 (N_6292,N_5975,N_5917);
and U6293 (N_6293,N_5702,N_5892);
or U6294 (N_6294,N_5859,N_5795);
nand U6295 (N_6295,N_5760,N_5772);
or U6296 (N_6296,N_5862,N_5876);
nand U6297 (N_6297,N_5913,N_5705);
xor U6298 (N_6298,N_5740,N_5812);
and U6299 (N_6299,N_5962,N_5994);
or U6300 (N_6300,N_6069,N_6295);
xnor U6301 (N_6301,N_6074,N_6128);
or U6302 (N_6302,N_6275,N_6123);
xor U6303 (N_6303,N_6286,N_6134);
xnor U6304 (N_6304,N_6282,N_6152);
xor U6305 (N_6305,N_6034,N_6096);
or U6306 (N_6306,N_6171,N_6233);
nand U6307 (N_6307,N_6142,N_6216);
nor U6308 (N_6308,N_6028,N_6006);
nor U6309 (N_6309,N_6158,N_6110);
and U6310 (N_6310,N_6146,N_6047);
nor U6311 (N_6311,N_6088,N_6291);
nand U6312 (N_6312,N_6108,N_6240);
xnor U6313 (N_6313,N_6126,N_6101);
xnor U6314 (N_6314,N_6266,N_6247);
nand U6315 (N_6315,N_6170,N_6092);
or U6316 (N_6316,N_6221,N_6269);
xnor U6317 (N_6317,N_6104,N_6009);
and U6318 (N_6318,N_6227,N_6018);
and U6319 (N_6319,N_6013,N_6271);
or U6320 (N_6320,N_6080,N_6037);
xnor U6321 (N_6321,N_6193,N_6173);
xnor U6322 (N_6322,N_6056,N_6292);
and U6323 (N_6323,N_6157,N_6039);
and U6324 (N_6324,N_6132,N_6007);
xnor U6325 (N_6325,N_6002,N_6082);
nand U6326 (N_6326,N_6273,N_6197);
xnor U6327 (N_6327,N_6035,N_6213);
xnor U6328 (N_6328,N_6281,N_6019);
xor U6329 (N_6329,N_6089,N_6033);
and U6330 (N_6330,N_6091,N_6042);
nor U6331 (N_6331,N_6192,N_6078);
or U6332 (N_6332,N_6057,N_6022);
or U6333 (N_6333,N_6177,N_6141);
nand U6334 (N_6334,N_6118,N_6212);
nor U6335 (N_6335,N_6188,N_6169);
or U6336 (N_6336,N_6280,N_6087);
or U6337 (N_6337,N_6184,N_6287);
nor U6338 (N_6338,N_6099,N_6285);
nand U6339 (N_6339,N_6217,N_6114);
or U6340 (N_6340,N_6129,N_6038);
nor U6341 (N_6341,N_6021,N_6116);
or U6342 (N_6342,N_6139,N_6249);
and U6343 (N_6343,N_6050,N_6257);
xnor U6344 (N_6344,N_6235,N_6147);
or U6345 (N_6345,N_6117,N_6119);
nor U6346 (N_6346,N_6219,N_6276);
nand U6347 (N_6347,N_6025,N_6063);
nor U6348 (N_6348,N_6224,N_6115);
or U6349 (N_6349,N_6155,N_6127);
and U6350 (N_6350,N_6262,N_6030);
or U6351 (N_6351,N_6229,N_6293);
xor U6352 (N_6352,N_6014,N_6026);
or U6353 (N_6353,N_6189,N_6070);
nor U6354 (N_6354,N_6068,N_6162);
nand U6355 (N_6355,N_6183,N_6136);
and U6356 (N_6356,N_6060,N_6267);
and U6357 (N_6357,N_6196,N_6097);
nor U6358 (N_6358,N_6225,N_6234);
and U6359 (N_6359,N_6090,N_6036);
nand U6360 (N_6360,N_6186,N_6256);
nor U6361 (N_6361,N_6251,N_6046);
nor U6362 (N_6362,N_6236,N_6071);
nor U6363 (N_6363,N_6043,N_6250);
and U6364 (N_6364,N_6232,N_6145);
nand U6365 (N_6365,N_6143,N_6049);
nand U6366 (N_6366,N_6121,N_6261);
nand U6367 (N_6367,N_6029,N_6270);
xor U6368 (N_6368,N_6079,N_6100);
nand U6369 (N_6369,N_6176,N_6207);
xnor U6370 (N_6370,N_6182,N_6067);
or U6371 (N_6371,N_6020,N_6202);
nor U6372 (N_6372,N_6253,N_6214);
xor U6373 (N_6373,N_6055,N_6248);
and U6374 (N_6374,N_6045,N_6187);
xnor U6375 (N_6375,N_6125,N_6059);
xor U6376 (N_6376,N_6200,N_6120);
nor U6377 (N_6377,N_6284,N_6168);
and U6378 (N_6378,N_6137,N_6166);
xor U6379 (N_6379,N_6296,N_6077);
nand U6380 (N_6380,N_6133,N_6246);
and U6381 (N_6381,N_6160,N_6244);
nand U6382 (N_6382,N_6237,N_6205);
nand U6383 (N_6383,N_6209,N_6113);
xor U6384 (N_6384,N_6084,N_6138);
xor U6385 (N_6385,N_6231,N_6159);
or U6386 (N_6386,N_6041,N_6010);
nor U6387 (N_6387,N_6172,N_6072);
xnor U6388 (N_6388,N_6061,N_6005);
or U6389 (N_6389,N_6000,N_6179);
nand U6390 (N_6390,N_6095,N_6174);
or U6391 (N_6391,N_6064,N_6112);
nor U6392 (N_6392,N_6075,N_6272);
nor U6393 (N_6393,N_6297,N_6201);
nor U6394 (N_6394,N_6245,N_6161);
xnor U6395 (N_6395,N_6102,N_6148);
xnor U6396 (N_6396,N_6238,N_6058);
nor U6397 (N_6397,N_6230,N_6109);
xnor U6398 (N_6398,N_6279,N_6040);
nand U6399 (N_6399,N_6210,N_6011);
xnor U6400 (N_6400,N_6124,N_6298);
and U6401 (N_6401,N_6065,N_6191);
nand U6402 (N_6402,N_6203,N_6190);
nand U6403 (N_6403,N_6204,N_6180);
nor U6404 (N_6404,N_6259,N_6228);
or U6405 (N_6405,N_6027,N_6194);
xor U6406 (N_6406,N_6178,N_6218);
nor U6407 (N_6407,N_6085,N_6274);
nor U6408 (N_6408,N_6066,N_6054);
nor U6409 (N_6409,N_6023,N_6220);
nand U6410 (N_6410,N_6151,N_6016);
xnor U6411 (N_6411,N_6242,N_6001);
nor U6412 (N_6412,N_6052,N_6111);
xor U6413 (N_6413,N_6283,N_6181);
or U6414 (N_6414,N_6198,N_6122);
and U6415 (N_6415,N_6167,N_6044);
nand U6416 (N_6416,N_6003,N_6098);
or U6417 (N_6417,N_6243,N_6239);
and U6418 (N_6418,N_6268,N_6226);
nor U6419 (N_6419,N_6015,N_6106);
nor U6420 (N_6420,N_6255,N_6153);
xor U6421 (N_6421,N_6083,N_6206);
nand U6422 (N_6422,N_6008,N_6131);
nand U6423 (N_6423,N_6017,N_6130);
or U6424 (N_6424,N_6144,N_6165);
or U6425 (N_6425,N_6032,N_6048);
or U6426 (N_6426,N_6222,N_6140);
nand U6427 (N_6427,N_6288,N_6199);
nand U6428 (N_6428,N_6223,N_6149);
or U6429 (N_6429,N_6024,N_6093);
nor U6430 (N_6430,N_6241,N_6062);
nand U6431 (N_6431,N_6081,N_6278);
xnor U6432 (N_6432,N_6105,N_6277);
and U6433 (N_6433,N_6107,N_6175);
or U6434 (N_6434,N_6185,N_6086);
and U6435 (N_6435,N_6150,N_6299);
and U6436 (N_6436,N_6211,N_6263);
nor U6437 (N_6437,N_6164,N_6135);
and U6438 (N_6438,N_6004,N_6031);
xnor U6439 (N_6439,N_6254,N_6264);
and U6440 (N_6440,N_6290,N_6103);
nor U6441 (N_6441,N_6053,N_6195);
and U6442 (N_6442,N_6258,N_6208);
and U6443 (N_6443,N_6294,N_6154);
nor U6444 (N_6444,N_6076,N_6156);
or U6445 (N_6445,N_6260,N_6073);
nand U6446 (N_6446,N_6051,N_6094);
nand U6447 (N_6447,N_6012,N_6265);
and U6448 (N_6448,N_6163,N_6289);
nand U6449 (N_6449,N_6252,N_6215);
xnor U6450 (N_6450,N_6206,N_6148);
and U6451 (N_6451,N_6012,N_6189);
or U6452 (N_6452,N_6235,N_6167);
nor U6453 (N_6453,N_6022,N_6279);
xnor U6454 (N_6454,N_6061,N_6056);
and U6455 (N_6455,N_6236,N_6130);
xor U6456 (N_6456,N_6041,N_6018);
and U6457 (N_6457,N_6090,N_6009);
or U6458 (N_6458,N_6233,N_6035);
and U6459 (N_6459,N_6200,N_6089);
nand U6460 (N_6460,N_6061,N_6263);
or U6461 (N_6461,N_6035,N_6152);
nor U6462 (N_6462,N_6145,N_6013);
nand U6463 (N_6463,N_6208,N_6042);
and U6464 (N_6464,N_6129,N_6092);
nor U6465 (N_6465,N_6245,N_6144);
and U6466 (N_6466,N_6215,N_6018);
and U6467 (N_6467,N_6174,N_6017);
or U6468 (N_6468,N_6202,N_6257);
or U6469 (N_6469,N_6000,N_6132);
or U6470 (N_6470,N_6146,N_6070);
xnor U6471 (N_6471,N_6187,N_6236);
xnor U6472 (N_6472,N_6134,N_6143);
nand U6473 (N_6473,N_6032,N_6207);
xor U6474 (N_6474,N_6229,N_6233);
nand U6475 (N_6475,N_6124,N_6012);
nor U6476 (N_6476,N_6111,N_6152);
nor U6477 (N_6477,N_6135,N_6049);
xnor U6478 (N_6478,N_6087,N_6232);
or U6479 (N_6479,N_6264,N_6239);
nand U6480 (N_6480,N_6142,N_6287);
or U6481 (N_6481,N_6011,N_6158);
nor U6482 (N_6482,N_6070,N_6082);
or U6483 (N_6483,N_6154,N_6135);
and U6484 (N_6484,N_6131,N_6277);
or U6485 (N_6485,N_6123,N_6132);
nand U6486 (N_6486,N_6028,N_6099);
xnor U6487 (N_6487,N_6040,N_6111);
and U6488 (N_6488,N_6021,N_6234);
nor U6489 (N_6489,N_6048,N_6102);
nand U6490 (N_6490,N_6126,N_6199);
nand U6491 (N_6491,N_6005,N_6049);
nor U6492 (N_6492,N_6280,N_6038);
nor U6493 (N_6493,N_6152,N_6110);
xor U6494 (N_6494,N_6089,N_6008);
or U6495 (N_6495,N_6063,N_6155);
nor U6496 (N_6496,N_6261,N_6256);
xnor U6497 (N_6497,N_6025,N_6282);
nand U6498 (N_6498,N_6164,N_6069);
and U6499 (N_6499,N_6005,N_6180);
xor U6500 (N_6500,N_6248,N_6036);
nor U6501 (N_6501,N_6152,N_6163);
or U6502 (N_6502,N_6015,N_6041);
nand U6503 (N_6503,N_6173,N_6066);
xnor U6504 (N_6504,N_6157,N_6279);
and U6505 (N_6505,N_6106,N_6080);
xnor U6506 (N_6506,N_6157,N_6237);
or U6507 (N_6507,N_6007,N_6280);
xor U6508 (N_6508,N_6213,N_6141);
xnor U6509 (N_6509,N_6289,N_6122);
xnor U6510 (N_6510,N_6023,N_6071);
xor U6511 (N_6511,N_6090,N_6250);
and U6512 (N_6512,N_6137,N_6158);
xnor U6513 (N_6513,N_6099,N_6050);
nor U6514 (N_6514,N_6052,N_6224);
nor U6515 (N_6515,N_6279,N_6034);
nor U6516 (N_6516,N_6125,N_6134);
nor U6517 (N_6517,N_6147,N_6185);
and U6518 (N_6518,N_6205,N_6068);
or U6519 (N_6519,N_6193,N_6125);
nor U6520 (N_6520,N_6004,N_6141);
xnor U6521 (N_6521,N_6166,N_6130);
nor U6522 (N_6522,N_6286,N_6097);
xor U6523 (N_6523,N_6149,N_6033);
nor U6524 (N_6524,N_6054,N_6241);
xnor U6525 (N_6525,N_6146,N_6267);
and U6526 (N_6526,N_6120,N_6160);
or U6527 (N_6527,N_6286,N_6050);
nand U6528 (N_6528,N_6000,N_6248);
xnor U6529 (N_6529,N_6164,N_6241);
xnor U6530 (N_6530,N_6286,N_6295);
nand U6531 (N_6531,N_6152,N_6003);
nor U6532 (N_6532,N_6012,N_6037);
or U6533 (N_6533,N_6124,N_6277);
xor U6534 (N_6534,N_6177,N_6148);
and U6535 (N_6535,N_6011,N_6090);
nand U6536 (N_6536,N_6148,N_6076);
xnor U6537 (N_6537,N_6188,N_6133);
nor U6538 (N_6538,N_6059,N_6250);
nor U6539 (N_6539,N_6147,N_6191);
nand U6540 (N_6540,N_6290,N_6046);
nand U6541 (N_6541,N_6252,N_6274);
or U6542 (N_6542,N_6117,N_6199);
xor U6543 (N_6543,N_6121,N_6056);
xnor U6544 (N_6544,N_6287,N_6172);
nand U6545 (N_6545,N_6104,N_6198);
nand U6546 (N_6546,N_6105,N_6171);
nor U6547 (N_6547,N_6075,N_6148);
or U6548 (N_6548,N_6107,N_6293);
nand U6549 (N_6549,N_6169,N_6238);
xor U6550 (N_6550,N_6209,N_6181);
nor U6551 (N_6551,N_6153,N_6111);
or U6552 (N_6552,N_6291,N_6231);
nand U6553 (N_6553,N_6079,N_6147);
nand U6554 (N_6554,N_6073,N_6020);
and U6555 (N_6555,N_6030,N_6104);
xnor U6556 (N_6556,N_6122,N_6077);
nand U6557 (N_6557,N_6249,N_6217);
and U6558 (N_6558,N_6127,N_6113);
nor U6559 (N_6559,N_6007,N_6067);
xor U6560 (N_6560,N_6236,N_6115);
or U6561 (N_6561,N_6092,N_6120);
xnor U6562 (N_6562,N_6251,N_6130);
nand U6563 (N_6563,N_6152,N_6285);
nand U6564 (N_6564,N_6083,N_6060);
nor U6565 (N_6565,N_6152,N_6002);
nand U6566 (N_6566,N_6216,N_6173);
or U6567 (N_6567,N_6048,N_6205);
or U6568 (N_6568,N_6231,N_6041);
nand U6569 (N_6569,N_6126,N_6112);
nand U6570 (N_6570,N_6056,N_6018);
and U6571 (N_6571,N_6281,N_6194);
or U6572 (N_6572,N_6042,N_6108);
and U6573 (N_6573,N_6026,N_6045);
or U6574 (N_6574,N_6278,N_6144);
or U6575 (N_6575,N_6241,N_6158);
nand U6576 (N_6576,N_6189,N_6185);
nor U6577 (N_6577,N_6020,N_6185);
xnor U6578 (N_6578,N_6249,N_6012);
xor U6579 (N_6579,N_6291,N_6112);
nor U6580 (N_6580,N_6017,N_6265);
nor U6581 (N_6581,N_6264,N_6141);
nor U6582 (N_6582,N_6117,N_6239);
nand U6583 (N_6583,N_6159,N_6116);
nor U6584 (N_6584,N_6006,N_6169);
nor U6585 (N_6585,N_6250,N_6190);
nand U6586 (N_6586,N_6244,N_6267);
nand U6587 (N_6587,N_6061,N_6114);
or U6588 (N_6588,N_6125,N_6030);
xnor U6589 (N_6589,N_6064,N_6080);
xnor U6590 (N_6590,N_6054,N_6065);
nor U6591 (N_6591,N_6295,N_6040);
nor U6592 (N_6592,N_6114,N_6192);
and U6593 (N_6593,N_6096,N_6266);
nor U6594 (N_6594,N_6123,N_6236);
nor U6595 (N_6595,N_6252,N_6163);
nor U6596 (N_6596,N_6054,N_6279);
xnor U6597 (N_6597,N_6151,N_6223);
xnor U6598 (N_6598,N_6163,N_6067);
and U6599 (N_6599,N_6057,N_6209);
and U6600 (N_6600,N_6447,N_6310);
and U6601 (N_6601,N_6575,N_6594);
and U6602 (N_6602,N_6434,N_6474);
nand U6603 (N_6603,N_6592,N_6438);
or U6604 (N_6604,N_6366,N_6379);
or U6605 (N_6605,N_6329,N_6322);
and U6606 (N_6606,N_6486,N_6497);
nand U6607 (N_6607,N_6303,N_6414);
and U6608 (N_6608,N_6330,N_6503);
nor U6609 (N_6609,N_6335,N_6589);
and U6610 (N_6610,N_6587,N_6467);
or U6611 (N_6611,N_6457,N_6432);
nor U6612 (N_6612,N_6401,N_6358);
nand U6613 (N_6613,N_6495,N_6521);
xor U6614 (N_6614,N_6593,N_6524);
and U6615 (N_6615,N_6378,N_6386);
nand U6616 (N_6616,N_6501,N_6428);
or U6617 (N_6617,N_6542,N_6461);
or U6618 (N_6618,N_6412,N_6558);
nor U6619 (N_6619,N_6563,N_6419);
xor U6620 (N_6620,N_6393,N_6529);
xnor U6621 (N_6621,N_6328,N_6562);
xnor U6622 (N_6622,N_6314,N_6571);
nand U6623 (N_6623,N_6450,N_6327);
nor U6624 (N_6624,N_6312,N_6357);
xnor U6625 (N_6625,N_6370,N_6359);
nand U6626 (N_6626,N_6475,N_6546);
and U6627 (N_6627,N_6406,N_6410);
and U6628 (N_6628,N_6469,N_6554);
nand U6629 (N_6629,N_6363,N_6507);
xor U6630 (N_6630,N_6307,N_6599);
nor U6631 (N_6631,N_6523,N_6400);
xor U6632 (N_6632,N_6548,N_6390);
nor U6633 (N_6633,N_6513,N_6388);
and U6634 (N_6634,N_6527,N_6349);
or U6635 (N_6635,N_6384,N_6308);
and U6636 (N_6636,N_6369,N_6526);
xor U6637 (N_6637,N_6510,N_6361);
xnor U6638 (N_6638,N_6333,N_6586);
and U6639 (N_6639,N_6352,N_6337);
nor U6640 (N_6640,N_6399,N_6397);
and U6641 (N_6641,N_6518,N_6462);
nand U6642 (N_6642,N_6535,N_6415);
or U6643 (N_6643,N_6446,N_6590);
and U6644 (N_6644,N_6568,N_6582);
nand U6645 (N_6645,N_6341,N_6313);
nand U6646 (N_6646,N_6360,N_6392);
nand U6647 (N_6647,N_6413,N_6460);
or U6648 (N_6648,N_6483,N_6347);
or U6649 (N_6649,N_6407,N_6464);
xor U6650 (N_6650,N_6560,N_6383);
xor U6651 (N_6651,N_6455,N_6425);
nor U6652 (N_6652,N_6448,N_6569);
nand U6653 (N_6653,N_6502,N_6519);
nor U6654 (N_6654,N_6319,N_6585);
nand U6655 (N_6655,N_6345,N_6403);
and U6656 (N_6656,N_6520,N_6487);
xor U6657 (N_6657,N_6477,N_6476);
and U6658 (N_6658,N_6334,N_6380);
nor U6659 (N_6659,N_6348,N_6431);
or U6660 (N_6660,N_6488,N_6556);
and U6661 (N_6661,N_6484,N_6325);
nor U6662 (N_6662,N_6496,N_6533);
or U6663 (N_6663,N_6435,N_6444);
and U6664 (N_6664,N_6591,N_6385);
nand U6665 (N_6665,N_6371,N_6433);
or U6666 (N_6666,N_6597,N_6309);
or U6667 (N_6667,N_6317,N_6458);
or U6668 (N_6668,N_6498,N_6387);
or U6669 (N_6669,N_6479,N_6532);
nand U6670 (N_6670,N_6346,N_6511);
nand U6671 (N_6671,N_6342,N_6515);
xnor U6672 (N_6672,N_6367,N_6538);
nor U6673 (N_6673,N_6493,N_6382);
xor U6674 (N_6674,N_6478,N_6408);
or U6675 (N_6675,N_6530,N_6364);
or U6676 (N_6676,N_6417,N_6528);
nor U6677 (N_6677,N_6557,N_6490);
xor U6678 (N_6678,N_6423,N_6445);
and U6679 (N_6679,N_6315,N_6578);
nor U6680 (N_6680,N_6541,N_6581);
nand U6681 (N_6681,N_6429,N_6454);
nand U6682 (N_6682,N_6372,N_6517);
nand U6683 (N_6683,N_6405,N_6453);
or U6684 (N_6684,N_6300,N_6579);
nor U6685 (N_6685,N_6443,N_6340);
nor U6686 (N_6686,N_6394,N_6426);
nand U6687 (N_6687,N_6306,N_6505);
xor U6688 (N_6688,N_6336,N_6540);
and U6689 (N_6689,N_6598,N_6305);
xor U6690 (N_6690,N_6375,N_6343);
and U6691 (N_6691,N_6323,N_6537);
and U6692 (N_6692,N_6427,N_6440);
nand U6693 (N_6693,N_6504,N_6566);
xor U6694 (N_6694,N_6332,N_6583);
and U6695 (N_6695,N_6350,N_6442);
or U6696 (N_6696,N_6588,N_6411);
xnor U6697 (N_6697,N_6574,N_6451);
nand U6698 (N_6698,N_6466,N_6456);
nand U6699 (N_6699,N_6577,N_6356);
xnor U6700 (N_6700,N_6439,N_6355);
xor U6701 (N_6701,N_6320,N_6485);
nand U6702 (N_6702,N_6508,N_6420);
nor U6703 (N_6703,N_6326,N_6559);
xor U6704 (N_6704,N_6351,N_6580);
xnor U6705 (N_6705,N_6304,N_6395);
nor U6706 (N_6706,N_6472,N_6377);
or U6707 (N_6707,N_6573,N_6500);
nor U6708 (N_6708,N_6465,N_6324);
nor U6709 (N_6709,N_6353,N_6381);
and U6710 (N_6710,N_6561,N_6374);
or U6711 (N_6711,N_6522,N_6338);
xnor U6712 (N_6712,N_6489,N_6567);
or U6713 (N_6713,N_6547,N_6549);
nand U6714 (N_6714,N_6316,N_6321);
xnor U6715 (N_6715,N_6301,N_6482);
xor U6716 (N_6716,N_6389,N_6595);
nand U6717 (N_6717,N_6572,N_6553);
nand U6718 (N_6718,N_6514,N_6481);
nor U6719 (N_6719,N_6449,N_6534);
or U6720 (N_6720,N_6565,N_6509);
or U6721 (N_6721,N_6318,N_6402);
xor U6722 (N_6722,N_6362,N_6471);
nor U6723 (N_6723,N_6584,N_6409);
nand U6724 (N_6724,N_6376,N_6550);
and U6725 (N_6725,N_6368,N_6545);
or U6726 (N_6726,N_6516,N_6421);
xnor U6727 (N_6727,N_6552,N_6512);
xnor U6728 (N_6728,N_6441,N_6437);
and U6729 (N_6729,N_6576,N_6422);
nor U6730 (N_6730,N_6452,N_6339);
nand U6731 (N_6731,N_6391,N_6354);
and U6732 (N_6732,N_6544,N_6480);
nand U6733 (N_6733,N_6492,N_6536);
or U6734 (N_6734,N_6365,N_6302);
xnor U6735 (N_6735,N_6398,N_6539);
xor U6736 (N_6736,N_6525,N_6570);
and U6737 (N_6737,N_6416,N_6564);
and U6738 (N_6738,N_6418,N_6468);
and U6739 (N_6739,N_6555,N_6424);
nor U6740 (N_6740,N_6430,N_6499);
xnor U6741 (N_6741,N_6436,N_6470);
and U6742 (N_6742,N_6373,N_6463);
nor U6743 (N_6743,N_6473,N_6331);
nand U6744 (N_6744,N_6344,N_6311);
or U6745 (N_6745,N_6596,N_6494);
or U6746 (N_6746,N_6543,N_6404);
nand U6747 (N_6747,N_6506,N_6396);
nor U6748 (N_6748,N_6491,N_6551);
xor U6749 (N_6749,N_6531,N_6459);
xnor U6750 (N_6750,N_6530,N_6525);
nor U6751 (N_6751,N_6563,N_6331);
and U6752 (N_6752,N_6566,N_6361);
and U6753 (N_6753,N_6492,N_6525);
and U6754 (N_6754,N_6506,N_6457);
xnor U6755 (N_6755,N_6589,N_6308);
nor U6756 (N_6756,N_6318,N_6417);
and U6757 (N_6757,N_6373,N_6548);
or U6758 (N_6758,N_6504,N_6466);
nor U6759 (N_6759,N_6450,N_6547);
nor U6760 (N_6760,N_6455,N_6526);
nand U6761 (N_6761,N_6530,N_6593);
or U6762 (N_6762,N_6352,N_6437);
and U6763 (N_6763,N_6443,N_6472);
or U6764 (N_6764,N_6564,N_6327);
or U6765 (N_6765,N_6375,N_6391);
or U6766 (N_6766,N_6355,N_6595);
and U6767 (N_6767,N_6318,N_6320);
nor U6768 (N_6768,N_6568,N_6481);
or U6769 (N_6769,N_6512,N_6490);
xor U6770 (N_6770,N_6387,N_6493);
nand U6771 (N_6771,N_6401,N_6398);
nand U6772 (N_6772,N_6490,N_6509);
nand U6773 (N_6773,N_6595,N_6520);
and U6774 (N_6774,N_6449,N_6326);
xor U6775 (N_6775,N_6475,N_6395);
nor U6776 (N_6776,N_6587,N_6362);
or U6777 (N_6777,N_6456,N_6546);
or U6778 (N_6778,N_6413,N_6462);
xor U6779 (N_6779,N_6580,N_6471);
and U6780 (N_6780,N_6484,N_6434);
or U6781 (N_6781,N_6515,N_6474);
nand U6782 (N_6782,N_6306,N_6440);
nand U6783 (N_6783,N_6535,N_6356);
or U6784 (N_6784,N_6334,N_6389);
nand U6785 (N_6785,N_6355,N_6370);
nand U6786 (N_6786,N_6583,N_6512);
or U6787 (N_6787,N_6327,N_6521);
xor U6788 (N_6788,N_6513,N_6344);
xor U6789 (N_6789,N_6525,N_6571);
xnor U6790 (N_6790,N_6493,N_6441);
nand U6791 (N_6791,N_6502,N_6353);
or U6792 (N_6792,N_6564,N_6527);
nand U6793 (N_6793,N_6394,N_6403);
or U6794 (N_6794,N_6339,N_6325);
and U6795 (N_6795,N_6580,N_6370);
xnor U6796 (N_6796,N_6570,N_6540);
nor U6797 (N_6797,N_6482,N_6541);
and U6798 (N_6798,N_6582,N_6583);
nor U6799 (N_6799,N_6530,N_6464);
xor U6800 (N_6800,N_6423,N_6553);
nor U6801 (N_6801,N_6580,N_6510);
nand U6802 (N_6802,N_6432,N_6588);
nor U6803 (N_6803,N_6314,N_6561);
xnor U6804 (N_6804,N_6319,N_6494);
nand U6805 (N_6805,N_6438,N_6312);
and U6806 (N_6806,N_6361,N_6413);
nor U6807 (N_6807,N_6424,N_6598);
nand U6808 (N_6808,N_6472,N_6498);
nor U6809 (N_6809,N_6433,N_6458);
xor U6810 (N_6810,N_6585,N_6586);
nand U6811 (N_6811,N_6593,N_6382);
xnor U6812 (N_6812,N_6334,N_6313);
nand U6813 (N_6813,N_6460,N_6555);
nand U6814 (N_6814,N_6532,N_6484);
nand U6815 (N_6815,N_6571,N_6475);
or U6816 (N_6816,N_6418,N_6478);
nand U6817 (N_6817,N_6391,N_6460);
and U6818 (N_6818,N_6596,N_6416);
nand U6819 (N_6819,N_6494,N_6564);
xor U6820 (N_6820,N_6525,N_6593);
nor U6821 (N_6821,N_6397,N_6340);
xnor U6822 (N_6822,N_6535,N_6362);
and U6823 (N_6823,N_6559,N_6563);
or U6824 (N_6824,N_6441,N_6352);
nand U6825 (N_6825,N_6461,N_6387);
nand U6826 (N_6826,N_6494,N_6356);
or U6827 (N_6827,N_6543,N_6507);
nand U6828 (N_6828,N_6585,N_6567);
and U6829 (N_6829,N_6515,N_6452);
and U6830 (N_6830,N_6326,N_6410);
and U6831 (N_6831,N_6433,N_6369);
nor U6832 (N_6832,N_6319,N_6374);
and U6833 (N_6833,N_6599,N_6401);
nor U6834 (N_6834,N_6538,N_6595);
or U6835 (N_6835,N_6440,N_6562);
and U6836 (N_6836,N_6412,N_6518);
nand U6837 (N_6837,N_6380,N_6376);
or U6838 (N_6838,N_6470,N_6350);
xnor U6839 (N_6839,N_6375,N_6422);
or U6840 (N_6840,N_6301,N_6384);
xor U6841 (N_6841,N_6344,N_6534);
nand U6842 (N_6842,N_6343,N_6425);
nor U6843 (N_6843,N_6448,N_6531);
or U6844 (N_6844,N_6365,N_6519);
and U6845 (N_6845,N_6360,N_6425);
and U6846 (N_6846,N_6550,N_6522);
and U6847 (N_6847,N_6429,N_6400);
and U6848 (N_6848,N_6308,N_6425);
or U6849 (N_6849,N_6428,N_6445);
nor U6850 (N_6850,N_6390,N_6582);
nor U6851 (N_6851,N_6513,N_6383);
nor U6852 (N_6852,N_6599,N_6482);
xnor U6853 (N_6853,N_6326,N_6437);
xor U6854 (N_6854,N_6303,N_6460);
or U6855 (N_6855,N_6450,N_6374);
nor U6856 (N_6856,N_6511,N_6529);
or U6857 (N_6857,N_6459,N_6460);
nor U6858 (N_6858,N_6527,N_6496);
xor U6859 (N_6859,N_6528,N_6494);
nand U6860 (N_6860,N_6303,N_6542);
and U6861 (N_6861,N_6593,N_6315);
or U6862 (N_6862,N_6315,N_6590);
nand U6863 (N_6863,N_6399,N_6529);
nor U6864 (N_6864,N_6418,N_6575);
nand U6865 (N_6865,N_6388,N_6551);
and U6866 (N_6866,N_6593,N_6473);
or U6867 (N_6867,N_6394,N_6500);
xor U6868 (N_6868,N_6327,N_6443);
xor U6869 (N_6869,N_6504,N_6370);
and U6870 (N_6870,N_6430,N_6388);
or U6871 (N_6871,N_6344,N_6354);
nand U6872 (N_6872,N_6466,N_6490);
nor U6873 (N_6873,N_6507,N_6334);
or U6874 (N_6874,N_6595,N_6417);
xnor U6875 (N_6875,N_6475,N_6428);
and U6876 (N_6876,N_6511,N_6448);
or U6877 (N_6877,N_6517,N_6391);
xnor U6878 (N_6878,N_6516,N_6538);
or U6879 (N_6879,N_6422,N_6490);
or U6880 (N_6880,N_6474,N_6323);
nand U6881 (N_6881,N_6324,N_6489);
nand U6882 (N_6882,N_6315,N_6520);
nand U6883 (N_6883,N_6562,N_6548);
or U6884 (N_6884,N_6464,N_6482);
nand U6885 (N_6885,N_6394,N_6535);
xnor U6886 (N_6886,N_6351,N_6449);
and U6887 (N_6887,N_6422,N_6318);
nand U6888 (N_6888,N_6375,N_6597);
xnor U6889 (N_6889,N_6521,N_6507);
nor U6890 (N_6890,N_6432,N_6594);
or U6891 (N_6891,N_6321,N_6387);
xor U6892 (N_6892,N_6411,N_6592);
and U6893 (N_6893,N_6386,N_6390);
nor U6894 (N_6894,N_6527,N_6394);
xnor U6895 (N_6895,N_6590,N_6425);
nand U6896 (N_6896,N_6572,N_6493);
xor U6897 (N_6897,N_6441,N_6424);
nand U6898 (N_6898,N_6301,N_6511);
nor U6899 (N_6899,N_6406,N_6402);
nor U6900 (N_6900,N_6886,N_6812);
nor U6901 (N_6901,N_6609,N_6701);
xor U6902 (N_6902,N_6696,N_6602);
nand U6903 (N_6903,N_6712,N_6827);
and U6904 (N_6904,N_6860,N_6797);
nor U6905 (N_6905,N_6615,N_6822);
and U6906 (N_6906,N_6893,N_6695);
or U6907 (N_6907,N_6635,N_6705);
or U6908 (N_6908,N_6662,N_6623);
or U6909 (N_6909,N_6832,N_6698);
and U6910 (N_6910,N_6769,N_6774);
nand U6911 (N_6911,N_6702,N_6835);
xnor U6912 (N_6912,N_6783,N_6888);
nand U6913 (N_6913,N_6803,N_6852);
nand U6914 (N_6914,N_6823,N_6897);
xnor U6915 (N_6915,N_6850,N_6639);
or U6916 (N_6916,N_6829,N_6855);
or U6917 (N_6917,N_6857,N_6826);
xor U6918 (N_6918,N_6776,N_6614);
nor U6919 (N_6919,N_6786,N_6634);
nand U6920 (N_6920,N_6762,N_6805);
or U6921 (N_6921,N_6863,N_6728);
xnor U6922 (N_6922,N_6811,N_6600);
nand U6923 (N_6923,N_6793,N_6646);
xor U6924 (N_6924,N_6645,N_6670);
nor U6925 (N_6925,N_6732,N_6727);
and U6926 (N_6926,N_6664,N_6711);
or U6927 (N_6927,N_6733,N_6633);
xnor U6928 (N_6928,N_6726,N_6881);
and U6929 (N_6929,N_6761,N_6756);
and U6930 (N_6930,N_6757,N_6810);
nand U6931 (N_6931,N_6708,N_6713);
xnor U6932 (N_6932,N_6649,N_6871);
or U6933 (N_6933,N_6661,N_6778);
and U6934 (N_6934,N_6868,N_6741);
nand U6935 (N_6935,N_6692,N_6628);
nor U6936 (N_6936,N_6849,N_6875);
nor U6937 (N_6937,N_6876,N_6874);
or U6938 (N_6938,N_6697,N_6703);
or U6939 (N_6939,N_6854,N_6684);
nand U6940 (N_6940,N_6790,N_6690);
and U6941 (N_6941,N_6714,N_6845);
and U6942 (N_6942,N_6819,N_6869);
nand U6943 (N_6943,N_6770,N_6842);
xnor U6944 (N_6944,N_6848,N_6693);
and U6945 (N_6945,N_6709,N_6794);
or U6946 (N_6946,N_6800,N_6813);
and U6947 (N_6947,N_6867,N_6729);
xor U6948 (N_6948,N_6866,N_6740);
nand U6949 (N_6949,N_6884,N_6608);
nor U6950 (N_6950,N_6706,N_6652);
nor U6951 (N_6951,N_6808,N_6632);
and U6952 (N_6952,N_6744,N_6717);
xor U6953 (N_6953,N_6838,N_6804);
and U6954 (N_6954,N_6704,N_6719);
and U6955 (N_6955,N_6889,N_6840);
and U6956 (N_6956,N_6647,N_6631);
nor U6957 (N_6957,N_6831,N_6636);
or U6958 (N_6958,N_6650,N_6674);
nand U6959 (N_6959,N_6752,N_6643);
nand U6960 (N_6960,N_6616,N_6629);
nand U6961 (N_6961,N_6807,N_6653);
or U6962 (N_6962,N_6681,N_6739);
and U6963 (N_6963,N_6895,N_6809);
xnor U6964 (N_6964,N_6678,N_6675);
and U6965 (N_6965,N_6676,N_6816);
and U6966 (N_6966,N_6766,N_6768);
nand U6967 (N_6967,N_6754,N_6722);
and U6968 (N_6968,N_6802,N_6792);
and U6969 (N_6969,N_6872,N_6689);
xor U6970 (N_6970,N_6742,N_6789);
and U6971 (N_6971,N_6621,N_6753);
nand U6972 (N_6972,N_6891,N_6864);
or U6973 (N_6973,N_6839,N_6718);
and U6974 (N_6974,N_6806,N_6841);
nand U6975 (N_6975,N_6737,N_6767);
or U6976 (N_6976,N_6626,N_6836);
and U6977 (N_6977,N_6777,N_6715);
or U6978 (N_6978,N_6765,N_6755);
xnor U6979 (N_6979,N_6707,N_6673);
nand U6980 (N_6980,N_6782,N_6870);
or U6981 (N_6981,N_6685,N_6736);
xor U6982 (N_6982,N_6773,N_6610);
or U6983 (N_6983,N_6723,N_6892);
xnor U6984 (N_6984,N_6747,N_6825);
or U6985 (N_6985,N_6730,N_6877);
xnor U6986 (N_6986,N_6785,N_6666);
nand U6987 (N_6987,N_6898,N_6873);
and U6988 (N_6988,N_6613,N_6682);
nand U6989 (N_6989,N_6654,N_6680);
or U6990 (N_6990,N_6784,N_6625);
and U6991 (N_6991,N_6688,N_6815);
nand U6992 (N_6992,N_6846,N_6780);
and U6993 (N_6993,N_6856,N_6796);
or U6994 (N_6994,N_6851,N_6878);
and U6995 (N_6995,N_6791,N_6724);
nor U6996 (N_6996,N_6833,N_6894);
and U6997 (N_6997,N_6788,N_6749);
or U6998 (N_6998,N_6882,N_6795);
nand U6999 (N_6999,N_6710,N_6745);
xnor U7000 (N_7000,N_6779,N_6817);
nand U7001 (N_7001,N_6834,N_6772);
nor U7002 (N_7002,N_6801,N_6859);
nor U7003 (N_7003,N_6853,N_6775);
nor U7004 (N_7004,N_6885,N_6735);
nand U7005 (N_7005,N_6843,N_6883);
nand U7006 (N_7006,N_6657,N_6837);
xnor U7007 (N_7007,N_6665,N_6624);
and U7008 (N_7008,N_6659,N_6604);
nand U7009 (N_7009,N_6828,N_6821);
nand U7010 (N_7010,N_6799,N_6830);
or U7011 (N_7011,N_6656,N_6638);
and U7012 (N_7012,N_6763,N_6743);
nor U7013 (N_7013,N_6660,N_6618);
or U7014 (N_7014,N_6686,N_6607);
nor U7015 (N_7015,N_6606,N_6642);
nor U7016 (N_7016,N_6787,N_6865);
xnor U7017 (N_7017,N_6640,N_6691);
nand U7018 (N_7018,N_6637,N_6844);
or U7019 (N_7019,N_6746,N_6824);
xor U7020 (N_7020,N_6687,N_6862);
nand U7021 (N_7021,N_6748,N_6814);
nor U7022 (N_7022,N_6725,N_6820);
nor U7023 (N_7023,N_6896,N_6771);
nor U7024 (N_7024,N_6738,N_6879);
nand U7025 (N_7025,N_6603,N_6671);
and U7026 (N_7026,N_6605,N_6612);
xor U7027 (N_7027,N_6630,N_6699);
nor U7028 (N_7028,N_6663,N_6751);
xnor U7029 (N_7029,N_6734,N_6619);
nor U7030 (N_7030,N_6641,N_6858);
xor U7031 (N_7031,N_6694,N_6861);
xor U7032 (N_7032,N_6764,N_6611);
and U7033 (N_7033,N_6759,N_6716);
or U7034 (N_7034,N_6622,N_6750);
or U7035 (N_7035,N_6601,N_6620);
or U7036 (N_7036,N_6700,N_6720);
and U7037 (N_7037,N_6658,N_6627);
nand U7038 (N_7038,N_6818,N_6760);
xnor U7039 (N_7039,N_6880,N_6644);
nor U7040 (N_7040,N_6617,N_6683);
or U7041 (N_7041,N_6672,N_6887);
and U7042 (N_7042,N_6668,N_6847);
and U7043 (N_7043,N_6890,N_6721);
or U7044 (N_7044,N_6899,N_6798);
xnor U7045 (N_7045,N_6731,N_6667);
nor U7046 (N_7046,N_6655,N_6669);
nand U7047 (N_7047,N_6758,N_6651);
nand U7048 (N_7048,N_6781,N_6677);
or U7049 (N_7049,N_6679,N_6648);
and U7050 (N_7050,N_6862,N_6863);
or U7051 (N_7051,N_6725,N_6861);
and U7052 (N_7052,N_6649,N_6678);
or U7053 (N_7053,N_6748,N_6803);
and U7054 (N_7054,N_6666,N_6743);
nand U7055 (N_7055,N_6825,N_6669);
or U7056 (N_7056,N_6870,N_6793);
or U7057 (N_7057,N_6698,N_6685);
nor U7058 (N_7058,N_6714,N_6805);
nor U7059 (N_7059,N_6774,N_6759);
or U7060 (N_7060,N_6606,N_6637);
nand U7061 (N_7061,N_6631,N_6816);
xor U7062 (N_7062,N_6720,N_6819);
or U7063 (N_7063,N_6676,N_6890);
nor U7064 (N_7064,N_6726,N_6862);
nor U7065 (N_7065,N_6621,N_6840);
nand U7066 (N_7066,N_6630,N_6782);
nor U7067 (N_7067,N_6792,N_6764);
nand U7068 (N_7068,N_6838,N_6734);
and U7069 (N_7069,N_6805,N_6859);
nor U7070 (N_7070,N_6618,N_6711);
or U7071 (N_7071,N_6715,N_6874);
and U7072 (N_7072,N_6720,N_6809);
nand U7073 (N_7073,N_6836,N_6813);
nand U7074 (N_7074,N_6604,N_6769);
or U7075 (N_7075,N_6840,N_6666);
nand U7076 (N_7076,N_6615,N_6883);
or U7077 (N_7077,N_6664,N_6651);
xnor U7078 (N_7078,N_6860,N_6606);
nand U7079 (N_7079,N_6685,N_6815);
or U7080 (N_7080,N_6779,N_6623);
and U7081 (N_7081,N_6777,N_6637);
nor U7082 (N_7082,N_6865,N_6767);
nand U7083 (N_7083,N_6894,N_6826);
xor U7084 (N_7084,N_6792,N_6730);
and U7085 (N_7085,N_6796,N_6697);
nand U7086 (N_7086,N_6696,N_6828);
and U7087 (N_7087,N_6814,N_6680);
nand U7088 (N_7088,N_6885,N_6892);
nor U7089 (N_7089,N_6836,N_6774);
nand U7090 (N_7090,N_6736,N_6634);
or U7091 (N_7091,N_6737,N_6765);
or U7092 (N_7092,N_6711,N_6654);
nand U7093 (N_7093,N_6760,N_6694);
nand U7094 (N_7094,N_6706,N_6658);
nand U7095 (N_7095,N_6745,N_6814);
and U7096 (N_7096,N_6897,N_6867);
nand U7097 (N_7097,N_6608,N_6790);
nand U7098 (N_7098,N_6608,N_6897);
nand U7099 (N_7099,N_6750,N_6760);
xor U7100 (N_7100,N_6809,N_6695);
nand U7101 (N_7101,N_6833,N_6701);
nand U7102 (N_7102,N_6790,N_6655);
nor U7103 (N_7103,N_6881,N_6618);
nor U7104 (N_7104,N_6616,N_6725);
and U7105 (N_7105,N_6775,N_6622);
and U7106 (N_7106,N_6799,N_6728);
xnor U7107 (N_7107,N_6767,N_6841);
and U7108 (N_7108,N_6786,N_6850);
or U7109 (N_7109,N_6673,N_6730);
or U7110 (N_7110,N_6684,N_6609);
nand U7111 (N_7111,N_6832,N_6729);
or U7112 (N_7112,N_6800,N_6674);
or U7113 (N_7113,N_6703,N_6628);
xor U7114 (N_7114,N_6879,N_6615);
and U7115 (N_7115,N_6812,N_6890);
and U7116 (N_7116,N_6830,N_6823);
or U7117 (N_7117,N_6627,N_6886);
or U7118 (N_7118,N_6899,N_6735);
and U7119 (N_7119,N_6741,N_6772);
xor U7120 (N_7120,N_6657,N_6718);
nor U7121 (N_7121,N_6812,N_6751);
and U7122 (N_7122,N_6814,N_6710);
xor U7123 (N_7123,N_6849,N_6657);
nand U7124 (N_7124,N_6717,N_6810);
nand U7125 (N_7125,N_6739,N_6765);
nor U7126 (N_7126,N_6620,N_6667);
nand U7127 (N_7127,N_6680,N_6717);
nor U7128 (N_7128,N_6830,N_6898);
nand U7129 (N_7129,N_6757,N_6744);
nor U7130 (N_7130,N_6831,N_6807);
and U7131 (N_7131,N_6737,N_6646);
nor U7132 (N_7132,N_6623,N_6649);
xor U7133 (N_7133,N_6744,N_6728);
or U7134 (N_7134,N_6722,N_6736);
and U7135 (N_7135,N_6684,N_6886);
nand U7136 (N_7136,N_6774,N_6766);
nand U7137 (N_7137,N_6709,N_6824);
and U7138 (N_7138,N_6726,N_6664);
nand U7139 (N_7139,N_6879,N_6617);
or U7140 (N_7140,N_6768,N_6861);
nand U7141 (N_7141,N_6830,N_6735);
nand U7142 (N_7142,N_6883,N_6622);
or U7143 (N_7143,N_6639,N_6733);
nor U7144 (N_7144,N_6641,N_6834);
nand U7145 (N_7145,N_6662,N_6753);
and U7146 (N_7146,N_6763,N_6610);
xor U7147 (N_7147,N_6713,N_6860);
nand U7148 (N_7148,N_6649,N_6711);
nor U7149 (N_7149,N_6684,N_6855);
or U7150 (N_7150,N_6635,N_6865);
nand U7151 (N_7151,N_6664,N_6771);
or U7152 (N_7152,N_6685,N_6793);
nor U7153 (N_7153,N_6773,N_6657);
xor U7154 (N_7154,N_6714,N_6755);
and U7155 (N_7155,N_6784,N_6871);
and U7156 (N_7156,N_6649,N_6724);
nand U7157 (N_7157,N_6719,N_6666);
nor U7158 (N_7158,N_6703,N_6787);
nand U7159 (N_7159,N_6790,N_6736);
or U7160 (N_7160,N_6782,N_6748);
or U7161 (N_7161,N_6721,N_6735);
nand U7162 (N_7162,N_6612,N_6789);
xor U7163 (N_7163,N_6875,N_6782);
or U7164 (N_7164,N_6802,N_6640);
nand U7165 (N_7165,N_6899,N_6667);
nand U7166 (N_7166,N_6837,N_6895);
nand U7167 (N_7167,N_6749,N_6835);
nor U7168 (N_7168,N_6689,N_6862);
and U7169 (N_7169,N_6717,N_6686);
nand U7170 (N_7170,N_6838,N_6702);
xnor U7171 (N_7171,N_6870,N_6854);
xnor U7172 (N_7172,N_6626,N_6710);
nand U7173 (N_7173,N_6843,N_6677);
or U7174 (N_7174,N_6610,N_6700);
nor U7175 (N_7175,N_6896,N_6818);
nand U7176 (N_7176,N_6794,N_6874);
xor U7177 (N_7177,N_6642,N_6726);
xnor U7178 (N_7178,N_6867,N_6795);
and U7179 (N_7179,N_6791,N_6834);
nand U7180 (N_7180,N_6748,N_6739);
and U7181 (N_7181,N_6650,N_6739);
nor U7182 (N_7182,N_6817,N_6818);
and U7183 (N_7183,N_6780,N_6683);
nand U7184 (N_7184,N_6702,N_6748);
or U7185 (N_7185,N_6840,N_6884);
or U7186 (N_7186,N_6726,N_6768);
nand U7187 (N_7187,N_6803,N_6877);
nor U7188 (N_7188,N_6739,N_6677);
nand U7189 (N_7189,N_6617,N_6730);
nand U7190 (N_7190,N_6602,N_6861);
xnor U7191 (N_7191,N_6620,N_6779);
xnor U7192 (N_7192,N_6877,N_6824);
xor U7193 (N_7193,N_6798,N_6842);
and U7194 (N_7194,N_6755,N_6769);
xor U7195 (N_7195,N_6657,N_6871);
and U7196 (N_7196,N_6824,N_6637);
and U7197 (N_7197,N_6616,N_6670);
or U7198 (N_7198,N_6777,N_6876);
nor U7199 (N_7199,N_6708,N_6675);
or U7200 (N_7200,N_6929,N_6983);
and U7201 (N_7201,N_6915,N_7073);
nand U7202 (N_7202,N_7120,N_7161);
or U7203 (N_7203,N_7066,N_7174);
nor U7204 (N_7204,N_7167,N_7024);
nor U7205 (N_7205,N_6946,N_7124);
and U7206 (N_7206,N_7086,N_6937);
nand U7207 (N_7207,N_7052,N_7096);
and U7208 (N_7208,N_7019,N_7021);
nor U7209 (N_7209,N_6997,N_7043);
and U7210 (N_7210,N_7062,N_7127);
or U7211 (N_7211,N_7103,N_7034);
nor U7212 (N_7212,N_7118,N_7137);
nand U7213 (N_7213,N_6954,N_6994);
xor U7214 (N_7214,N_7033,N_7100);
nor U7215 (N_7215,N_7038,N_7075);
and U7216 (N_7216,N_7087,N_7074);
nand U7217 (N_7217,N_7159,N_6921);
and U7218 (N_7218,N_6973,N_7064);
nor U7219 (N_7219,N_7117,N_6991);
nor U7220 (N_7220,N_7131,N_6999);
or U7221 (N_7221,N_7199,N_6952);
or U7222 (N_7222,N_7029,N_6912);
and U7223 (N_7223,N_7168,N_6988);
and U7224 (N_7224,N_7044,N_7028);
xor U7225 (N_7225,N_7192,N_7015);
nand U7226 (N_7226,N_6942,N_6966);
nand U7227 (N_7227,N_7164,N_6910);
nand U7228 (N_7228,N_6948,N_7008);
and U7229 (N_7229,N_6905,N_6904);
nand U7230 (N_7230,N_7069,N_7187);
or U7231 (N_7231,N_6926,N_6927);
and U7232 (N_7232,N_6964,N_7106);
nand U7233 (N_7233,N_6913,N_7094);
nor U7234 (N_7234,N_6963,N_7101);
or U7235 (N_7235,N_6949,N_7122);
nor U7236 (N_7236,N_6974,N_7182);
nor U7237 (N_7237,N_7047,N_7079);
nand U7238 (N_7238,N_7080,N_7156);
nand U7239 (N_7239,N_7025,N_6982);
or U7240 (N_7240,N_7088,N_6906);
nand U7241 (N_7241,N_7057,N_7102);
and U7242 (N_7242,N_7160,N_7040);
xor U7243 (N_7243,N_6986,N_7000);
xor U7244 (N_7244,N_7185,N_6995);
xnor U7245 (N_7245,N_7145,N_7039);
xor U7246 (N_7246,N_6977,N_7022);
xor U7247 (N_7247,N_7197,N_6924);
nor U7248 (N_7248,N_7179,N_7175);
nor U7249 (N_7249,N_7155,N_7190);
nor U7250 (N_7250,N_7030,N_7129);
nor U7251 (N_7251,N_6944,N_7095);
nor U7252 (N_7252,N_7191,N_7189);
and U7253 (N_7253,N_6993,N_7169);
xor U7254 (N_7254,N_7170,N_7188);
xor U7255 (N_7255,N_7071,N_6928);
and U7256 (N_7256,N_7007,N_7108);
and U7257 (N_7257,N_6950,N_6996);
nand U7258 (N_7258,N_6951,N_7135);
nor U7259 (N_7259,N_7154,N_7054);
and U7260 (N_7260,N_7126,N_6980);
nand U7261 (N_7261,N_7001,N_7140);
nand U7262 (N_7262,N_7026,N_7093);
and U7263 (N_7263,N_7020,N_7051);
or U7264 (N_7264,N_7198,N_7112);
and U7265 (N_7265,N_7076,N_6945);
nor U7266 (N_7266,N_7032,N_7151);
nand U7267 (N_7267,N_6969,N_7107);
nor U7268 (N_7268,N_6958,N_7173);
nand U7269 (N_7269,N_6960,N_7013);
xnor U7270 (N_7270,N_7031,N_7176);
nand U7271 (N_7271,N_6900,N_7009);
xor U7272 (N_7272,N_6919,N_7092);
nand U7273 (N_7273,N_6979,N_7070);
and U7274 (N_7274,N_7050,N_7090);
nand U7275 (N_7275,N_7099,N_7121);
nor U7276 (N_7276,N_7049,N_6943);
and U7277 (N_7277,N_7045,N_7085);
and U7278 (N_7278,N_7068,N_7004);
xor U7279 (N_7279,N_7016,N_7125);
xor U7280 (N_7280,N_7010,N_7149);
or U7281 (N_7281,N_7193,N_7147);
and U7282 (N_7282,N_7035,N_6934);
and U7283 (N_7283,N_7061,N_7110);
nand U7284 (N_7284,N_7132,N_7184);
and U7285 (N_7285,N_7134,N_7158);
xor U7286 (N_7286,N_7183,N_7150);
and U7287 (N_7287,N_6908,N_6976);
and U7288 (N_7288,N_7083,N_6918);
xnor U7289 (N_7289,N_7153,N_7136);
or U7290 (N_7290,N_6978,N_6925);
nor U7291 (N_7291,N_6992,N_6989);
or U7292 (N_7292,N_6968,N_7119);
or U7293 (N_7293,N_7162,N_6940);
nor U7294 (N_7294,N_7114,N_7115);
nand U7295 (N_7295,N_6933,N_6916);
nor U7296 (N_7296,N_7181,N_7005);
nor U7297 (N_7297,N_7078,N_7067);
and U7298 (N_7298,N_7098,N_6959);
xnor U7299 (N_7299,N_6967,N_7065);
nor U7300 (N_7300,N_7037,N_7017);
and U7301 (N_7301,N_6985,N_7081);
xnor U7302 (N_7302,N_7111,N_7186);
xor U7303 (N_7303,N_7053,N_6935);
and U7304 (N_7304,N_7084,N_7058);
nor U7305 (N_7305,N_6909,N_7091);
and U7306 (N_7306,N_7018,N_6975);
nor U7307 (N_7307,N_6917,N_6962);
and U7308 (N_7308,N_6965,N_7060);
and U7309 (N_7309,N_6990,N_7195);
and U7310 (N_7310,N_7163,N_7104);
and U7311 (N_7311,N_6953,N_7027);
nor U7312 (N_7312,N_7089,N_7194);
nor U7313 (N_7313,N_6938,N_7128);
and U7314 (N_7314,N_6947,N_6941);
nand U7315 (N_7315,N_7148,N_7116);
nor U7316 (N_7316,N_7152,N_7138);
and U7317 (N_7317,N_6911,N_6922);
nor U7318 (N_7318,N_6970,N_6998);
nor U7319 (N_7319,N_7109,N_7014);
nor U7320 (N_7320,N_6957,N_6956);
xnor U7321 (N_7321,N_7196,N_6936);
nand U7322 (N_7322,N_6914,N_7059);
nand U7323 (N_7323,N_7063,N_6955);
nand U7324 (N_7324,N_7097,N_7048);
xnor U7325 (N_7325,N_6939,N_6902);
nand U7326 (N_7326,N_7143,N_7142);
and U7327 (N_7327,N_7036,N_7082);
and U7328 (N_7328,N_7157,N_6981);
or U7329 (N_7329,N_6961,N_7177);
or U7330 (N_7330,N_7003,N_7146);
nand U7331 (N_7331,N_7133,N_7113);
and U7332 (N_7332,N_6903,N_7123);
xnor U7333 (N_7333,N_7077,N_6972);
xnor U7334 (N_7334,N_6930,N_7178);
nand U7335 (N_7335,N_7165,N_6920);
and U7336 (N_7336,N_7002,N_7141);
xnor U7337 (N_7337,N_7171,N_6987);
nor U7338 (N_7338,N_6932,N_7105);
nand U7339 (N_7339,N_7023,N_7166);
nor U7340 (N_7340,N_6907,N_7144);
and U7341 (N_7341,N_7072,N_7139);
xnor U7342 (N_7342,N_7006,N_7055);
nand U7343 (N_7343,N_7012,N_7130);
nor U7344 (N_7344,N_6931,N_7042);
and U7345 (N_7345,N_7180,N_6984);
and U7346 (N_7346,N_7056,N_7172);
or U7347 (N_7347,N_6901,N_7011);
xnor U7348 (N_7348,N_7046,N_7041);
nor U7349 (N_7349,N_6923,N_6971);
or U7350 (N_7350,N_6902,N_7110);
nand U7351 (N_7351,N_7007,N_7003);
xor U7352 (N_7352,N_7091,N_7192);
nor U7353 (N_7353,N_7065,N_6966);
and U7354 (N_7354,N_6922,N_6925);
and U7355 (N_7355,N_6912,N_7141);
and U7356 (N_7356,N_7020,N_7027);
xor U7357 (N_7357,N_6979,N_6985);
nor U7358 (N_7358,N_7189,N_6951);
nand U7359 (N_7359,N_6972,N_7054);
nand U7360 (N_7360,N_7186,N_6997);
nand U7361 (N_7361,N_7055,N_7128);
and U7362 (N_7362,N_7061,N_7042);
or U7363 (N_7363,N_7060,N_6941);
and U7364 (N_7364,N_7057,N_6993);
and U7365 (N_7365,N_6993,N_6905);
nand U7366 (N_7366,N_7198,N_7073);
xor U7367 (N_7367,N_7120,N_7150);
xnor U7368 (N_7368,N_7024,N_6999);
and U7369 (N_7369,N_7150,N_6996);
and U7370 (N_7370,N_6921,N_6910);
nor U7371 (N_7371,N_7058,N_6914);
or U7372 (N_7372,N_6975,N_7186);
nor U7373 (N_7373,N_7058,N_7065);
nor U7374 (N_7374,N_7157,N_7166);
and U7375 (N_7375,N_7060,N_7065);
nor U7376 (N_7376,N_7001,N_7087);
and U7377 (N_7377,N_7119,N_6915);
nor U7378 (N_7378,N_7007,N_7144);
nand U7379 (N_7379,N_7067,N_7026);
xor U7380 (N_7380,N_6927,N_7192);
nand U7381 (N_7381,N_7042,N_7027);
nor U7382 (N_7382,N_7197,N_7053);
nand U7383 (N_7383,N_7106,N_7147);
or U7384 (N_7384,N_7068,N_7072);
xor U7385 (N_7385,N_6998,N_7097);
nand U7386 (N_7386,N_7042,N_7068);
xnor U7387 (N_7387,N_7035,N_6946);
xor U7388 (N_7388,N_7179,N_6906);
nand U7389 (N_7389,N_7113,N_7070);
and U7390 (N_7390,N_7093,N_6920);
nor U7391 (N_7391,N_6935,N_7116);
or U7392 (N_7392,N_7043,N_7022);
and U7393 (N_7393,N_6982,N_7000);
and U7394 (N_7394,N_6941,N_7055);
or U7395 (N_7395,N_7012,N_7145);
and U7396 (N_7396,N_6934,N_6959);
nand U7397 (N_7397,N_7046,N_7022);
nand U7398 (N_7398,N_7081,N_7118);
nand U7399 (N_7399,N_7159,N_7129);
xnor U7400 (N_7400,N_7116,N_6955);
nand U7401 (N_7401,N_7061,N_7168);
or U7402 (N_7402,N_6951,N_6929);
xor U7403 (N_7403,N_6936,N_7048);
and U7404 (N_7404,N_6910,N_7028);
or U7405 (N_7405,N_7165,N_7013);
nand U7406 (N_7406,N_7198,N_7032);
and U7407 (N_7407,N_7121,N_7005);
nor U7408 (N_7408,N_6980,N_7102);
nor U7409 (N_7409,N_6908,N_7193);
nor U7410 (N_7410,N_7187,N_6912);
and U7411 (N_7411,N_7138,N_7009);
and U7412 (N_7412,N_7004,N_7101);
xnor U7413 (N_7413,N_7051,N_6951);
nor U7414 (N_7414,N_6981,N_7008);
xnor U7415 (N_7415,N_6928,N_6981);
or U7416 (N_7416,N_6925,N_7019);
nand U7417 (N_7417,N_7020,N_7089);
or U7418 (N_7418,N_7177,N_7192);
or U7419 (N_7419,N_7156,N_7087);
and U7420 (N_7420,N_7166,N_7090);
xnor U7421 (N_7421,N_7146,N_6919);
nand U7422 (N_7422,N_7015,N_6927);
nor U7423 (N_7423,N_7046,N_6930);
xnor U7424 (N_7424,N_6928,N_7111);
nand U7425 (N_7425,N_6974,N_7088);
nor U7426 (N_7426,N_6942,N_7165);
nand U7427 (N_7427,N_7021,N_7076);
or U7428 (N_7428,N_7025,N_7179);
and U7429 (N_7429,N_6950,N_7088);
and U7430 (N_7430,N_7009,N_7034);
or U7431 (N_7431,N_7132,N_6947);
nor U7432 (N_7432,N_6926,N_6975);
or U7433 (N_7433,N_6951,N_6921);
and U7434 (N_7434,N_6900,N_6932);
and U7435 (N_7435,N_7124,N_7050);
or U7436 (N_7436,N_7022,N_7052);
nand U7437 (N_7437,N_6922,N_7128);
or U7438 (N_7438,N_6927,N_7108);
or U7439 (N_7439,N_7168,N_7100);
or U7440 (N_7440,N_6909,N_7055);
nor U7441 (N_7441,N_7170,N_7083);
and U7442 (N_7442,N_7056,N_7020);
nand U7443 (N_7443,N_7108,N_6930);
nand U7444 (N_7444,N_7123,N_6969);
and U7445 (N_7445,N_7091,N_6967);
and U7446 (N_7446,N_7075,N_7192);
nor U7447 (N_7447,N_6901,N_6968);
and U7448 (N_7448,N_7039,N_7130);
and U7449 (N_7449,N_6902,N_7198);
and U7450 (N_7450,N_6953,N_7071);
nand U7451 (N_7451,N_7081,N_7142);
nand U7452 (N_7452,N_7131,N_7060);
nand U7453 (N_7453,N_7163,N_6937);
xnor U7454 (N_7454,N_6942,N_7000);
xor U7455 (N_7455,N_6914,N_7068);
xor U7456 (N_7456,N_7134,N_6932);
or U7457 (N_7457,N_7083,N_7129);
or U7458 (N_7458,N_7028,N_7055);
nand U7459 (N_7459,N_7068,N_6970);
and U7460 (N_7460,N_7178,N_6972);
and U7461 (N_7461,N_7171,N_6950);
or U7462 (N_7462,N_7053,N_7103);
xnor U7463 (N_7463,N_7099,N_6935);
xnor U7464 (N_7464,N_7141,N_6980);
or U7465 (N_7465,N_7141,N_7189);
nor U7466 (N_7466,N_7122,N_7162);
xor U7467 (N_7467,N_7136,N_6926);
nand U7468 (N_7468,N_7110,N_7199);
or U7469 (N_7469,N_6943,N_6902);
and U7470 (N_7470,N_7047,N_7114);
and U7471 (N_7471,N_7055,N_7041);
nor U7472 (N_7472,N_6921,N_7084);
nand U7473 (N_7473,N_6900,N_7128);
and U7474 (N_7474,N_7156,N_7124);
xnor U7475 (N_7475,N_7196,N_7102);
nand U7476 (N_7476,N_6938,N_6971);
nor U7477 (N_7477,N_6968,N_6927);
and U7478 (N_7478,N_7000,N_7030);
and U7479 (N_7479,N_7151,N_7165);
and U7480 (N_7480,N_7087,N_7090);
nor U7481 (N_7481,N_6912,N_7193);
nor U7482 (N_7482,N_6943,N_7057);
or U7483 (N_7483,N_7003,N_6951);
or U7484 (N_7484,N_7013,N_7059);
and U7485 (N_7485,N_6904,N_7035);
and U7486 (N_7486,N_7164,N_7072);
nor U7487 (N_7487,N_7012,N_7112);
xor U7488 (N_7488,N_7117,N_7006);
xnor U7489 (N_7489,N_6974,N_7096);
or U7490 (N_7490,N_7180,N_6983);
or U7491 (N_7491,N_6949,N_6942);
xor U7492 (N_7492,N_6906,N_7085);
xor U7493 (N_7493,N_6961,N_6974);
xor U7494 (N_7494,N_7053,N_7142);
nand U7495 (N_7495,N_7173,N_7002);
nand U7496 (N_7496,N_7149,N_7154);
nor U7497 (N_7497,N_7181,N_7198);
nor U7498 (N_7498,N_6946,N_7126);
xnor U7499 (N_7499,N_6927,N_7171);
nor U7500 (N_7500,N_7285,N_7388);
and U7501 (N_7501,N_7350,N_7490);
nor U7502 (N_7502,N_7299,N_7304);
or U7503 (N_7503,N_7225,N_7264);
nand U7504 (N_7504,N_7426,N_7246);
nand U7505 (N_7505,N_7453,N_7268);
and U7506 (N_7506,N_7408,N_7403);
nand U7507 (N_7507,N_7280,N_7398);
nor U7508 (N_7508,N_7455,N_7283);
and U7509 (N_7509,N_7243,N_7258);
xor U7510 (N_7510,N_7245,N_7241);
nand U7511 (N_7511,N_7282,N_7262);
or U7512 (N_7512,N_7421,N_7306);
nor U7513 (N_7513,N_7332,N_7239);
nor U7514 (N_7514,N_7473,N_7227);
or U7515 (N_7515,N_7308,N_7253);
and U7516 (N_7516,N_7361,N_7499);
xnor U7517 (N_7517,N_7414,N_7444);
nand U7518 (N_7518,N_7357,N_7276);
nand U7519 (N_7519,N_7291,N_7410);
nor U7520 (N_7520,N_7244,N_7437);
or U7521 (N_7521,N_7201,N_7354);
and U7522 (N_7522,N_7396,N_7255);
nand U7523 (N_7523,N_7384,N_7458);
and U7524 (N_7524,N_7335,N_7389);
nor U7525 (N_7525,N_7419,N_7307);
or U7526 (N_7526,N_7395,N_7406);
and U7527 (N_7527,N_7327,N_7247);
nand U7528 (N_7528,N_7294,N_7281);
and U7529 (N_7529,N_7380,N_7325);
nand U7530 (N_7530,N_7234,N_7439);
nand U7531 (N_7531,N_7359,N_7420);
and U7532 (N_7532,N_7373,N_7236);
or U7533 (N_7533,N_7349,N_7256);
and U7534 (N_7534,N_7428,N_7488);
or U7535 (N_7535,N_7411,N_7266);
xor U7536 (N_7536,N_7212,N_7464);
nand U7537 (N_7537,N_7498,N_7219);
and U7538 (N_7538,N_7412,N_7315);
and U7539 (N_7539,N_7339,N_7312);
xnor U7540 (N_7540,N_7237,N_7347);
nand U7541 (N_7541,N_7222,N_7461);
nor U7542 (N_7542,N_7249,N_7269);
nor U7543 (N_7543,N_7487,N_7329);
or U7544 (N_7544,N_7287,N_7353);
and U7545 (N_7545,N_7497,N_7378);
and U7546 (N_7546,N_7360,N_7386);
nand U7547 (N_7547,N_7441,N_7393);
or U7548 (N_7548,N_7479,N_7477);
nor U7549 (N_7549,N_7211,N_7451);
or U7550 (N_7550,N_7338,N_7430);
or U7551 (N_7551,N_7240,N_7209);
nor U7552 (N_7552,N_7427,N_7486);
and U7553 (N_7553,N_7452,N_7480);
or U7554 (N_7554,N_7418,N_7434);
and U7555 (N_7555,N_7213,N_7392);
and U7556 (N_7556,N_7472,N_7333);
xor U7557 (N_7557,N_7460,N_7448);
nand U7558 (N_7558,N_7316,N_7416);
nor U7559 (N_7559,N_7300,N_7336);
xnor U7560 (N_7560,N_7242,N_7491);
or U7561 (N_7561,N_7217,N_7367);
and U7562 (N_7562,N_7492,N_7482);
and U7563 (N_7563,N_7478,N_7371);
nand U7564 (N_7564,N_7407,N_7330);
xor U7565 (N_7565,N_7286,N_7374);
nor U7566 (N_7566,N_7221,N_7485);
nor U7567 (N_7567,N_7443,N_7381);
or U7568 (N_7568,N_7436,N_7214);
nand U7569 (N_7569,N_7385,N_7383);
nor U7570 (N_7570,N_7296,N_7366);
or U7571 (N_7571,N_7224,N_7289);
nor U7572 (N_7572,N_7326,N_7345);
nor U7573 (N_7573,N_7489,N_7334);
nand U7574 (N_7574,N_7376,N_7493);
xnor U7575 (N_7575,N_7409,N_7232);
or U7576 (N_7576,N_7290,N_7405);
xnor U7577 (N_7577,N_7203,N_7404);
and U7578 (N_7578,N_7348,N_7310);
and U7579 (N_7579,N_7252,N_7231);
or U7580 (N_7580,N_7313,N_7302);
xor U7581 (N_7581,N_7394,N_7495);
and U7582 (N_7582,N_7447,N_7228);
xnor U7583 (N_7583,N_7462,N_7362);
nor U7584 (N_7584,N_7220,N_7210);
and U7585 (N_7585,N_7494,N_7440);
xnor U7586 (N_7586,N_7397,N_7295);
and U7587 (N_7587,N_7379,N_7450);
xor U7588 (N_7588,N_7305,N_7230);
or U7589 (N_7589,N_7355,N_7342);
or U7590 (N_7590,N_7496,N_7351);
nor U7591 (N_7591,N_7275,N_7229);
xnor U7592 (N_7592,N_7476,N_7278);
nor U7593 (N_7593,N_7425,N_7352);
xnor U7594 (N_7594,N_7457,N_7320);
and U7595 (N_7595,N_7470,N_7235);
xnor U7596 (N_7596,N_7321,N_7466);
and U7597 (N_7597,N_7288,N_7358);
nand U7598 (N_7598,N_7260,N_7319);
and U7599 (N_7599,N_7233,N_7415);
xnor U7600 (N_7600,N_7206,N_7356);
xor U7601 (N_7601,N_7257,N_7390);
xnor U7602 (N_7602,N_7204,N_7413);
xor U7603 (N_7603,N_7363,N_7469);
nand U7604 (N_7604,N_7277,N_7435);
and U7605 (N_7605,N_7322,N_7271);
nand U7606 (N_7606,N_7422,N_7387);
xnor U7607 (N_7607,N_7433,N_7218);
or U7608 (N_7608,N_7314,N_7454);
xor U7609 (N_7609,N_7442,N_7463);
nand U7610 (N_7610,N_7331,N_7456);
xor U7611 (N_7611,N_7263,N_7250);
nor U7612 (N_7612,N_7446,N_7208);
and U7613 (N_7613,N_7303,N_7216);
nor U7614 (N_7614,N_7270,N_7438);
nor U7615 (N_7615,N_7297,N_7431);
nand U7616 (N_7616,N_7340,N_7267);
nor U7617 (N_7617,N_7292,N_7429);
nand U7618 (N_7618,N_7475,N_7215);
and U7619 (N_7619,N_7324,N_7465);
nor U7620 (N_7620,N_7391,N_7365);
nor U7621 (N_7621,N_7272,N_7223);
nand U7622 (N_7622,N_7474,N_7259);
and U7623 (N_7623,N_7341,N_7207);
or U7624 (N_7624,N_7346,N_7417);
xor U7625 (N_7625,N_7481,N_7254);
or U7626 (N_7626,N_7468,N_7445);
nor U7627 (N_7627,N_7205,N_7200);
nand U7628 (N_7628,N_7328,N_7251);
or U7629 (N_7629,N_7375,N_7471);
xor U7630 (N_7630,N_7226,N_7343);
and U7631 (N_7631,N_7401,N_7424);
or U7632 (N_7632,N_7377,N_7467);
xor U7633 (N_7633,N_7459,N_7202);
and U7634 (N_7634,N_7261,N_7317);
nand U7635 (N_7635,N_7399,N_7344);
xnor U7636 (N_7636,N_7432,N_7293);
or U7637 (N_7637,N_7284,N_7372);
nand U7638 (N_7638,N_7337,N_7309);
and U7639 (N_7639,N_7483,N_7248);
nor U7640 (N_7640,N_7368,N_7265);
nand U7641 (N_7641,N_7369,N_7323);
nand U7642 (N_7642,N_7423,N_7238);
or U7643 (N_7643,N_7449,N_7484);
nand U7644 (N_7644,N_7311,N_7402);
nand U7645 (N_7645,N_7364,N_7318);
nand U7646 (N_7646,N_7273,N_7274);
and U7647 (N_7647,N_7298,N_7382);
xnor U7648 (N_7648,N_7400,N_7301);
or U7649 (N_7649,N_7279,N_7370);
xnor U7650 (N_7650,N_7428,N_7496);
nor U7651 (N_7651,N_7427,N_7275);
nor U7652 (N_7652,N_7432,N_7449);
xor U7653 (N_7653,N_7215,N_7298);
nand U7654 (N_7654,N_7394,N_7372);
xor U7655 (N_7655,N_7230,N_7362);
and U7656 (N_7656,N_7268,N_7327);
or U7657 (N_7657,N_7444,N_7286);
or U7658 (N_7658,N_7454,N_7414);
xnor U7659 (N_7659,N_7451,N_7218);
and U7660 (N_7660,N_7473,N_7343);
nor U7661 (N_7661,N_7405,N_7384);
nor U7662 (N_7662,N_7288,N_7379);
and U7663 (N_7663,N_7485,N_7330);
and U7664 (N_7664,N_7433,N_7223);
and U7665 (N_7665,N_7420,N_7269);
nor U7666 (N_7666,N_7300,N_7258);
nand U7667 (N_7667,N_7275,N_7254);
nor U7668 (N_7668,N_7319,N_7440);
nand U7669 (N_7669,N_7410,N_7292);
or U7670 (N_7670,N_7465,N_7435);
nor U7671 (N_7671,N_7336,N_7237);
and U7672 (N_7672,N_7461,N_7457);
xor U7673 (N_7673,N_7382,N_7241);
nand U7674 (N_7674,N_7455,N_7446);
xnor U7675 (N_7675,N_7436,N_7208);
or U7676 (N_7676,N_7364,N_7296);
nor U7677 (N_7677,N_7356,N_7467);
nor U7678 (N_7678,N_7265,N_7324);
nand U7679 (N_7679,N_7356,N_7355);
nand U7680 (N_7680,N_7260,N_7480);
nand U7681 (N_7681,N_7497,N_7269);
or U7682 (N_7682,N_7471,N_7333);
xnor U7683 (N_7683,N_7291,N_7208);
xor U7684 (N_7684,N_7360,N_7408);
nand U7685 (N_7685,N_7283,N_7424);
nand U7686 (N_7686,N_7313,N_7418);
xor U7687 (N_7687,N_7393,N_7430);
xnor U7688 (N_7688,N_7412,N_7280);
and U7689 (N_7689,N_7304,N_7277);
xor U7690 (N_7690,N_7458,N_7417);
nand U7691 (N_7691,N_7486,N_7431);
and U7692 (N_7692,N_7374,N_7426);
or U7693 (N_7693,N_7365,N_7272);
and U7694 (N_7694,N_7351,N_7396);
xor U7695 (N_7695,N_7401,N_7422);
or U7696 (N_7696,N_7326,N_7263);
or U7697 (N_7697,N_7416,N_7258);
nor U7698 (N_7698,N_7389,N_7442);
and U7699 (N_7699,N_7271,N_7267);
or U7700 (N_7700,N_7367,N_7363);
nor U7701 (N_7701,N_7420,N_7228);
and U7702 (N_7702,N_7205,N_7352);
and U7703 (N_7703,N_7447,N_7493);
and U7704 (N_7704,N_7216,N_7425);
nand U7705 (N_7705,N_7200,N_7468);
nand U7706 (N_7706,N_7334,N_7294);
nor U7707 (N_7707,N_7328,N_7272);
and U7708 (N_7708,N_7476,N_7409);
nor U7709 (N_7709,N_7421,N_7293);
and U7710 (N_7710,N_7420,N_7268);
nor U7711 (N_7711,N_7404,N_7325);
xor U7712 (N_7712,N_7427,N_7210);
nand U7713 (N_7713,N_7392,N_7495);
nor U7714 (N_7714,N_7386,N_7241);
and U7715 (N_7715,N_7373,N_7409);
and U7716 (N_7716,N_7385,N_7489);
nand U7717 (N_7717,N_7432,N_7328);
or U7718 (N_7718,N_7449,N_7257);
nor U7719 (N_7719,N_7372,N_7385);
and U7720 (N_7720,N_7208,N_7237);
nand U7721 (N_7721,N_7453,N_7255);
and U7722 (N_7722,N_7276,N_7351);
and U7723 (N_7723,N_7464,N_7226);
or U7724 (N_7724,N_7490,N_7253);
nor U7725 (N_7725,N_7385,N_7342);
and U7726 (N_7726,N_7256,N_7394);
and U7727 (N_7727,N_7489,N_7453);
nor U7728 (N_7728,N_7361,N_7496);
or U7729 (N_7729,N_7298,N_7293);
or U7730 (N_7730,N_7311,N_7314);
xnor U7731 (N_7731,N_7352,N_7320);
or U7732 (N_7732,N_7328,N_7237);
nand U7733 (N_7733,N_7397,N_7312);
xor U7734 (N_7734,N_7219,N_7470);
and U7735 (N_7735,N_7259,N_7305);
nand U7736 (N_7736,N_7402,N_7416);
nand U7737 (N_7737,N_7410,N_7273);
nand U7738 (N_7738,N_7333,N_7448);
nor U7739 (N_7739,N_7468,N_7309);
nand U7740 (N_7740,N_7450,N_7239);
nand U7741 (N_7741,N_7310,N_7266);
nor U7742 (N_7742,N_7466,N_7250);
and U7743 (N_7743,N_7380,N_7406);
and U7744 (N_7744,N_7214,N_7461);
nor U7745 (N_7745,N_7283,N_7338);
nand U7746 (N_7746,N_7318,N_7376);
nor U7747 (N_7747,N_7449,N_7364);
nand U7748 (N_7748,N_7223,N_7448);
or U7749 (N_7749,N_7295,N_7430);
or U7750 (N_7750,N_7416,N_7205);
and U7751 (N_7751,N_7342,N_7442);
nor U7752 (N_7752,N_7270,N_7304);
or U7753 (N_7753,N_7236,N_7432);
or U7754 (N_7754,N_7237,N_7472);
or U7755 (N_7755,N_7419,N_7473);
or U7756 (N_7756,N_7337,N_7365);
or U7757 (N_7757,N_7287,N_7308);
and U7758 (N_7758,N_7288,N_7344);
and U7759 (N_7759,N_7427,N_7311);
and U7760 (N_7760,N_7435,N_7201);
xnor U7761 (N_7761,N_7424,N_7465);
or U7762 (N_7762,N_7381,N_7245);
and U7763 (N_7763,N_7251,N_7326);
xor U7764 (N_7764,N_7384,N_7455);
or U7765 (N_7765,N_7356,N_7378);
or U7766 (N_7766,N_7349,N_7390);
xor U7767 (N_7767,N_7365,N_7279);
and U7768 (N_7768,N_7272,N_7396);
and U7769 (N_7769,N_7262,N_7344);
xnor U7770 (N_7770,N_7349,N_7303);
nor U7771 (N_7771,N_7231,N_7257);
and U7772 (N_7772,N_7392,N_7228);
xnor U7773 (N_7773,N_7205,N_7373);
or U7774 (N_7774,N_7355,N_7488);
and U7775 (N_7775,N_7330,N_7421);
nand U7776 (N_7776,N_7309,N_7209);
nor U7777 (N_7777,N_7284,N_7380);
nand U7778 (N_7778,N_7287,N_7442);
or U7779 (N_7779,N_7352,N_7393);
and U7780 (N_7780,N_7300,N_7410);
xnor U7781 (N_7781,N_7297,N_7253);
xor U7782 (N_7782,N_7324,N_7475);
nor U7783 (N_7783,N_7246,N_7299);
nand U7784 (N_7784,N_7306,N_7438);
xor U7785 (N_7785,N_7476,N_7491);
nor U7786 (N_7786,N_7377,N_7320);
xnor U7787 (N_7787,N_7305,N_7483);
or U7788 (N_7788,N_7344,N_7333);
xor U7789 (N_7789,N_7237,N_7333);
and U7790 (N_7790,N_7469,N_7346);
xnor U7791 (N_7791,N_7435,N_7473);
xnor U7792 (N_7792,N_7417,N_7214);
nor U7793 (N_7793,N_7400,N_7468);
and U7794 (N_7794,N_7361,N_7213);
and U7795 (N_7795,N_7465,N_7242);
nand U7796 (N_7796,N_7348,N_7488);
and U7797 (N_7797,N_7233,N_7486);
nand U7798 (N_7798,N_7248,N_7237);
xor U7799 (N_7799,N_7481,N_7228);
or U7800 (N_7800,N_7661,N_7564);
or U7801 (N_7801,N_7527,N_7696);
or U7802 (N_7802,N_7655,N_7724);
nand U7803 (N_7803,N_7591,N_7691);
and U7804 (N_7804,N_7702,N_7751);
or U7805 (N_7805,N_7638,N_7662);
nand U7806 (N_7806,N_7504,N_7722);
nand U7807 (N_7807,N_7641,N_7554);
and U7808 (N_7808,N_7573,N_7558);
nand U7809 (N_7809,N_7595,N_7605);
nand U7810 (N_7810,N_7782,N_7594);
xnor U7811 (N_7811,N_7741,N_7673);
or U7812 (N_7812,N_7637,N_7614);
nand U7813 (N_7813,N_7557,N_7509);
xnor U7814 (N_7814,N_7784,N_7787);
or U7815 (N_7815,N_7569,N_7750);
nand U7816 (N_7816,N_7528,N_7779);
nor U7817 (N_7817,N_7508,N_7648);
and U7818 (N_7818,N_7626,N_7664);
or U7819 (N_7819,N_7681,N_7789);
or U7820 (N_7820,N_7596,N_7701);
or U7821 (N_7821,N_7689,N_7560);
nand U7822 (N_7822,N_7600,N_7629);
xnor U7823 (N_7823,N_7721,N_7517);
nor U7824 (N_7824,N_7776,N_7767);
and U7825 (N_7825,N_7777,N_7780);
or U7826 (N_7826,N_7617,N_7778);
xor U7827 (N_7827,N_7618,N_7576);
xnor U7828 (N_7828,N_7511,N_7765);
nand U7829 (N_7829,N_7642,N_7533);
xor U7830 (N_7830,N_7652,N_7633);
and U7831 (N_7831,N_7516,N_7500);
and U7832 (N_7832,N_7530,N_7615);
or U7833 (N_7833,N_7715,N_7717);
and U7834 (N_7834,N_7676,N_7670);
or U7835 (N_7835,N_7773,N_7612);
or U7836 (N_7836,N_7790,N_7797);
and U7837 (N_7837,N_7796,N_7710);
nand U7838 (N_7838,N_7708,N_7669);
nand U7839 (N_7839,N_7674,N_7644);
or U7840 (N_7840,N_7745,N_7513);
or U7841 (N_7841,N_7540,N_7768);
xor U7842 (N_7842,N_7624,N_7622);
nand U7843 (N_7843,N_7623,N_7792);
nand U7844 (N_7844,N_7534,N_7650);
or U7845 (N_7845,N_7526,N_7561);
and U7846 (N_7846,N_7572,N_7593);
nor U7847 (N_7847,N_7603,N_7549);
nand U7848 (N_7848,N_7657,N_7690);
nor U7849 (N_7849,N_7639,N_7791);
xnor U7850 (N_7850,N_7542,N_7544);
nand U7851 (N_7851,N_7758,N_7694);
nor U7852 (N_7852,N_7737,N_7728);
or U7853 (N_7853,N_7720,N_7552);
and U7854 (N_7854,N_7537,N_7551);
or U7855 (N_7855,N_7584,N_7632);
and U7856 (N_7856,N_7733,N_7525);
nand U7857 (N_7857,N_7645,N_7589);
or U7858 (N_7858,N_7760,N_7772);
and U7859 (N_7859,N_7671,N_7601);
and U7860 (N_7860,N_7746,N_7667);
nor U7861 (N_7861,N_7625,N_7620);
and U7862 (N_7862,N_7547,N_7795);
nand U7863 (N_7863,N_7687,N_7518);
xor U7864 (N_7864,N_7683,N_7763);
or U7865 (N_7865,N_7582,N_7535);
xnor U7866 (N_7866,N_7726,N_7666);
and U7867 (N_7867,N_7718,N_7744);
or U7868 (N_7868,N_7581,N_7597);
xnor U7869 (N_7869,N_7672,N_7588);
and U7870 (N_7870,N_7607,N_7586);
or U7871 (N_7871,N_7755,N_7748);
nor U7872 (N_7872,N_7663,N_7677);
nor U7873 (N_7873,N_7538,N_7546);
nor U7874 (N_7874,N_7619,N_7532);
xor U7875 (N_7875,N_7679,N_7501);
and U7876 (N_7876,N_7680,N_7653);
or U7877 (N_7877,N_7568,N_7700);
xor U7878 (N_7878,N_7740,N_7695);
xnor U7879 (N_7879,N_7592,N_7628);
xor U7880 (N_7880,N_7660,N_7602);
or U7881 (N_7881,N_7580,N_7606);
or U7882 (N_7882,N_7685,N_7643);
and U7883 (N_7883,N_7545,N_7523);
nand U7884 (N_7884,N_7735,N_7570);
and U7885 (N_7885,N_7698,N_7522);
nand U7886 (N_7886,N_7736,N_7781);
or U7887 (N_7887,N_7524,N_7775);
nor U7888 (N_7888,N_7719,N_7759);
nand U7889 (N_7889,N_7578,N_7709);
nor U7890 (N_7890,N_7656,N_7684);
or U7891 (N_7891,N_7519,N_7732);
nand U7892 (N_7892,N_7640,N_7598);
or U7893 (N_7893,N_7506,N_7539);
and U7894 (N_7894,N_7565,N_7743);
or U7895 (N_7895,N_7543,N_7766);
and U7896 (N_7896,N_7556,N_7520);
xnor U7897 (N_7897,N_7727,N_7703);
or U7898 (N_7898,N_7675,N_7553);
and U7899 (N_7899,N_7636,N_7630);
nor U7900 (N_7900,N_7716,N_7774);
nand U7901 (N_7901,N_7742,N_7510);
or U7902 (N_7902,N_7608,N_7699);
and U7903 (N_7903,N_7697,N_7668);
or U7904 (N_7904,N_7610,N_7512);
and U7905 (N_7905,N_7713,N_7756);
nor U7906 (N_7906,N_7575,N_7658);
xor U7907 (N_7907,N_7753,N_7514);
xor U7908 (N_7908,N_7665,N_7786);
and U7909 (N_7909,N_7705,N_7646);
xor U7910 (N_7910,N_7686,N_7563);
xnor U7911 (N_7911,N_7788,N_7647);
nor U7912 (N_7912,N_7793,N_7567);
nand U7913 (N_7913,N_7611,N_7529);
nand U7914 (N_7914,N_7574,N_7503);
xor U7915 (N_7915,N_7536,N_7559);
nand U7916 (N_7916,N_7548,N_7585);
nand U7917 (N_7917,N_7616,N_7730);
and U7918 (N_7918,N_7550,N_7723);
or U7919 (N_7919,N_7649,N_7659);
and U7920 (N_7920,N_7785,N_7502);
nand U7921 (N_7921,N_7752,N_7579);
xnor U7922 (N_7922,N_7604,N_7754);
nand U7923 (N_7923,N_7706,N_7729);
and U7924 (N_7924,N_7714,N_7507);
xnor U7925 (N_7925,N_7562,N_7515);
and U7926 (N_7926,N_7731,N_7771);
xnor U7927 (N_7927,N_7505,N_7734);
xor U7928 (N_7928,N_7739,N_7747);
nand U7929 (N_7929,N_7688,N_7599);
or U7930 (N_7930,N_7761,N_7749);
nand U7931 (N_7931,N_7678,N_7634);
nor U7932 (N_7932,N_7692,N_7566);
nand U7933 (N_7933,N_7654,N_7609);
xnor U7934 (N_7934,N_7541,N_7764);
xor U7935 (N_7935,N_7707,N_7712);
nand U7936 (N_7936,N_7635,N_7794);
and U7937 (N_7937,N_7531,N_7693);
nor U7938 (N_7938,N_7590,N_7783);
or U7939 (N_7939,N_7555,N_7631);
or U7940 (N_7940,N_7769,N_7577);
and U7941 (N_7941,N_7799,N_7798);
or U7942 (N_7942,N_7725,N_7704);
or U7943 (N_7943,N_7682,N_7621);
nor U7944 (N_7944,N_7587,N_7770);
xor U7945 (N_7945,N_7627,N_7738);
or U7946 (N_7946,N_7757,N_7651);
or U7947 (N_7947,N_7521,N_7613);
nor U7948 (N_7948,N_7571,N_7711);
nor U7949 (N_7949,N_7762,N_7583);
nor U7950 (N_7950,N_7528,N_7633);
or U7951 (N_7951,N_7790,N_7752);
nand U7952 (N_7952,N_7576,N_7512);
nand U7953 (N_7953,N_7530,N_7603);
or U7954 (N_7954,N_7785,N_7582);
xor U7955 (N_7955,N_7586,N_7568);
xor U7956 (N_7956,N_7589,N_7789);
nor U7957 (N_7957,N_7581,N_7543);
and U7958 (N_7958,N_7738,N_7741);
xnor U7959 (N_7959,N_7542,N_7535);
xnor U7960 (N_7960,N_7621,N_7762);
nor U7961 (N_7961,N_7739,N_7728);
nor U7962 (N_7962,N_7500,N_7644);
nand U7963 (N_7963,N_7514,N_7569);
xnor U7964 (N_7964,N_7678,N_7790);
or U7965 (N_7965,N_7674,N_7565);
or U7966 (N_7966,N_7675,N_7528);
nor U7967 (N_7967,N_7737,N_7669);
or U7968 (N_7968,N_7664,N_7531);
and U7969 (N_7969,N_7680,N_7723);
and U7970 (N_7970,N_7552,N_7701);
nor U7971 (N_7971,N_7790,N_7638);
or U7972 (N_7972,N_7707,N_7670);
and U7973 (N_7973,N_7593,N_7745);
nand U7974 (N_7974,N_7682,N_7664);
nand U7975 (N_7975,N_7643,N_7747);
nor U7976 (N_7976,N_7690,N_7742);
nand U7977 (N_7977,N_7708,N_7620);
and U7978 (N_7978,N_7532,N_7636);
nor U7979 (N_7979,N_7671,N_7517);
nand U7980 (N_7980,N_7776,N_7783);
or U7981 (N_7981,N_7569,N_7742);
nand U7982 (N_7982,N_7710,N_7694);
nand U7983 (N_7983,N_7502,N_7627);
or U7984 (N_7984,N_7678,N_7755);
or U7985 (N_7985,N_7767,N_7744);
nand U7986 (N_7986,N_7672,N_7766);
xnor U7987 (N_7987,N_7544,N_7688);
nand U7988 (N_7988,N_7610,N_7709);
and U7989 (N_7989,N_7736,N_7666);
nand U7990 (N_7990,N_7796,N_7725);
and U7991 (N_7991,N_7703,N_7596);
or U7992 (N_7992,N_7584,N_7567);
nand U7993 (N_7993,N_7688,N_7512);
nor U7994 (N_7994,N_7619,N_7613);
xnor U7995 (N_7995,N_7567,N_7549);
and U7996 (N_7996,N_7703,N_7527);
nor U7997 (N_7997,N_7663,N_7709);
nor U7998 (N_7998,N_7696,N_7775);
and U7999 (N_7999,N_7790,N_7714);
nand U8000 (N_8000,N_7727,N_7595);
xor U8001 (N_8001,N_7637,N_7544);
or U8002 (N_8002,N_7518,N_7675);
nand U8003 (N_8003,N_7661,N_7729);
nand U8004 (N_8004,N_7728,N_7659);
nor U8005 (N_8005,N_7521,N_7704);
nor U8006 (N_8006,N_7754,N_7517);
nand U8007 (N_8007,N_7613,N_7635);
or U8008 (N_8008,N_7602,N_7616);
xnor U8009 (N_8009,N_7577,N_7657);
or U8010 (N_8010,N_7520,N_7654);
xor U8011 (N_8011,N_7753,N_7604);
xor U8012 (N_8012,N_7557,N_7611);
or U8013 (N_8013,N_7679,N_7776);
and U8014 (N_8014,N_7513,N_7721);
nand U8015 (N_8015,N_7731,N_7791);
or U8016 (N_8016,N_7709,N_7699);
or U8017 (N_8017,N_7542,N_7750);
nand U8018 (N_8018,N_7600,N_7709);
nand U8019 (N_8019,N_7626,N_7505);
nand U8020 (N_8020,N_7644,N_7711);
nor U8021 (N_8021,N_7662,N_7560);
or U8022 (N_8022,N_7527,N_7690);
and U8023 (N_8023,N_7766,N_7602);
and U8024 (N_8024,N_7611,N_7790);
nor U8025 (N_8025,N_7755,N_7726);
or U8026 (N_8026,N_7788,N_7666);
xnor U8027 (N_8027,N_7788,N_7736);
and U8028 (N_8028,N_7721,N_7597);
and U8029 (N_8029,N_7759,N_7550);
or U8030 (N_8030,N_7746,N_7712);
and U8031 (N_8031,N_7510,N_7692);
xnor U8032 (N_8032,N_7569,N_7747);
nand U8033 (N_8033,N_7574,N_7530);
nand U8034 (N_8034,N_7786,N_7658);
xor U8035 (N_8035,N_7537,N_7607);
nand U8036 (N_8036,N_7516,N_7679);
and U8037 (N_8037,N_7509,N_7561);
xnor U8038 (N_8038,N_7618,N_7727);
xnor U8039 (N_8039,N_7706,N_7705);
and U8040 (N_8040,N_7557,N_7645);
or U8041 (N_8041,N_7630,N_7698);
nand U8042 (N_8042,N_7527,N_7504);
nand U8043 (N_8043,N_7719,N_7696);
or U8044 (N_8044,N_7589,N_7571);
nor U8045 (N_8045,N_7748,N_7665);
or U8046 (N_8046,N_7632,N_7648);
xnor U8047 (N_8047,N_7585,N_7646);
nor U8048 (N_8048,N_7703,N_7552);
nor U8049 (N_8049,N_7757,N_7527);
and U8050 (N_8050,N_7700,N_7533);
xor U8051 (N_8051,N_7661,N_7574);
xnor U8052 (N_8052,N_7734,N_7710);
xor U8053 (N_8053,N_7716,N_7608);
and U8054 (N_8054,N_7708,N_7606);
nor U8055 (N_8055,N_7510,N_7554);
nor U8056 (N_8056,N_7534,N_7579);
and U8057 (N_8057,N_7606,N_7624);
and U8058 (N_8058,N_7537,N_7502);
nor U8059 (N_8059,N_7710,N_7762);
nor U8060 (N_8060,N_7728,N_7652);
nor U8061 (N_8061,N_7724,N_7529);
and U8062 (N_8062,N_7684,N_7613);
and U8063 (N_8063,N_7692,N_7617);
xor U8064 (N_8064,N_7663,N_7638);
nor U8065 (N_8065,N_7706,N_7754);
or U8066 (N_8066,N_7632,N_7772);
xnor U8067 (N_8067,N_7663,N_7747);
xnor U8068 (N_8068,N_7631,N_7559);
and U8069 (N_8069,N_7579,N_7578);
and U8070 (N_8070,N_7616,N_7525);
and U8071 (N_8071,N_7747,N_7738);
nor U8072 (N_8072,N_7610,N_7533);
or U8073 (N_8073,N_7683,N_7752);
or U8074 (N_8074,N_7641,N_7788);
nor U8075 (N_8075,N_7791,N_7697);
or U8076 (N_8076,N_7753,N_7528);
nor U8077 (N_8077,N_7589,N_7538);
and U8078 (N_8078,N_7594,N_7503);
and U8079 (N_8079,N_7701,N_7686);
nand U8080 (N_8080,N_7760,N_7516);
and U8081 (N_8081,N_7511,N_7633);
xnor U8082 (N_8082,N_7751,N_7712);
or U8083 (N_8083,N_7558,N_7730);
xnor U8084 (N_8084,N_7788,N_7755);
and U8085 (N_8085,N_7610,N_7781);
or U8086 (N_8086,N_7684,N_7665);
and U8087 (N_8087,N_7775,N_7537);
and U8088 (N_8088,N_7622,N_7503);
or U8089 (N_8089,N_7578,N_7673);
nand U8090 (N_8090,N_7534,N_7543);
nand U8091 (N_8091,N_7624,N_7711);
nand U8092 (N_8092,N_7693,N_7564);
nor U8093 (N_8093,N_7592,N_7564);
xor U8094 (N_8094,N_7735,N_7717);
nand U8095 (N_8095,N_7637,N_7543);
nor U8096 (N_8096,N_7620,N_7648);
and U8097 (N_8097,N_7531,N_7660);
and U8098 (N_8098,N_7786,N_7710);
and U8099 (N_8099,N_7783,N_7698);
nor U8100 (N_8100,N_8065,N_7834);
xnor U8101 (N_8101,N_7902,N_7824);
and U8102 (N_8102,N_7841,N_7931);
nand U8103 (N_8103,N_7857,N_7838);
nor U8104 (N_8104,N_8086,N_8073);
xnor U8105 (N_8105,N_7869,N_8071);
nand U8106 (N_8106,N_7949,N_8016);
nand U8107 (N_8107,N_7845,N_7906);
nor U8108 (N_8108,N_7804,N_7870);
nand U8109 (N_8109,N_7843,N_7997);
nor U8110 (N_8110,N_8033,N_7895);
xnor U8111 (N_8111,N_7844,N_8053);
nand U8112 (N_8112,N_7928,N_7907);
xor U8113 (N_8113,N_7863,N_8068);
or U8114 (N_8114,N_8050,N_7876);
xnor U8115 (N_8115,N_7886,N_7871);
or U8116 (N_8116,N_7940,N_7967);
and U8117 (N_8117,N_7964,N_7802);
nand U8118 (N_8118,N_8088,N_7976);
nand U8119 (N_8119,N_8078,N_7889);
xor U8120 (N_8120,N_8080,N_7933);
nand U8121 (N_8121,N_8083,N_8008);
nand U8122 (N_8122,N_8040,N_7956);
nor U8123 (N_8123,N_8061,N_7968);
nor U8124 (N_8124,N_7810,N_7939);
nand U8125 (N_8125,N_7935,N_7842);
and U8126 (N_8126,N_7922,N_7855);
or U8127 (N_8127,N_8044,N_7835);
or U8128 (N_8128,N_7919,N_8001);
nand U8129 (N_8129,N_8049,N_7819);
nand U8130 (N_8130,N_7829,N_8023);
xnor U8131 (N_8131,N_7944,N_8066);
xnor U8132 (N_8132,N_7912,N_8036);
nand U8133 (N_8133,N_8024,N_8019);
or U8134 (N_8134,N_8082,N_7881);
xor U8135 (N_8135,N_7951,N_7884);
or U8136 (N_8136,N_8076,N_8054);
or U8137 (N_8137,N_7822,N_8069);
and U8138 (N_8138,N_7915,N_7960);
nand U8139 (N_8139,N_7962,N_7961);
or U8140 (N_8140,N_7980,N_7850);
or U8141 (N_8141,N_7926,N_7866);
or U8142 (N_8142,N_7836,N_7899);
nand U8143 (N_8143,N_8070,N_7945);
or U8144 (N_8144,N_7830,N_8087);
or U8145 (N_8145,N_8017,N_7882);
and U8146 (N_8146,N_7957,N_7910);
xnor U8147 (N_8147,N_7973,N_7878);
nor U8148 (N_8148,N_8028,N_7809);
or U8149 (N_8149,N_7833,N_7827);
or U8150 (N_8150,N_7904,N_7814);
and U8151 (N_8151,N_8081,N_8022);
and U8152 (N_8152,N_8097,N_7999);
xor U8153 (N_8153,N_7903,N_7990);
and U8154 (N_8154,N_7985,N_7803);
nor U8155 (N_8155,N_7925,N_8005);
nand U8156 (N_8156,N_7891,N_8030);
nand U8157 (N_8157,N_8072,N_7856);
nor U8158 (N_8158,N_7971,N_8095);
nor U8159 (N_8159,N_7894,N_7984);
and U8160 (N_8160,N_8043,N_7879);
nor U8161 (N_8161,N_7888,N_7832);
and U8162 (N_8162,N_8090,N_7821);
xnor U8163 (N_8163,N_8015,N_8037);
nand U8164 (N_8164,N_7986,N_7946);
nor U8165 (N_8165,N_7812,N_7995);
xnor U8166 (N_8166,N_8059,N_8021);
or U8167 (N_8167,N_7828,N_7862);
xnor U8168 (N_8168,N_7996,N_7801);
nand U8169 (N_8169,N_7965,N_7974);
xor U8170 (N_8170,N_7992,N_7911);
xnor U8171 (N_8171,N_8055,N_7848);
or U8172 (N_8172,N_7941,N_7808);
xnor U8173 (N_8173,N_7811,N_8041);
nand U8174 (N_8174,N_7859,N_8047);
xor U8175 (N_8175,N_7916,N_7959);
or U8176 (N_8176,N_7860,N_7813);
xor U8177 (N_8177,N_7937,N_8060);
or U8178 (N_8178,N_8009,N_7938);
xnor U8179 (N_8179,N_7872,N_7849);
nand U8180 (N_8180,N_8056,N_7991);
nor U8181 (N_8181,N_8092,N_7952);
and U8182 (N_8182,N_7924,N_8002);
nor U8183 (N_8183,N_7875,N_8012);
xnor U8184 (N_8184,N_8098,N_7908);
nand U8185 (N_8185,N_7837,N_7988);
nor U8186 (N_8186,N_7818,N_7897);
and U8187 (N_8187,N_7977,N_7918);
and U8188 (N_8188,N_7989,N_7982);
nand U8189 (N_8189,N_7981,N_8099);
nand U8190 (N_8190,N_7913,N_7800);
or U8191 (N_8191,N_8058,N_8062);
nor U8192 (N_8192,N_8013,N_7987);
nand U8193 (N_8193,N_8035,N_7874);
and U8194 (N_8194,N_7994,N_7831);
nor U8195 (N_8195,N_8048,N_7900);
xor U8196 (N_8196,N_7806,N_7825);
nand U8197 (N_8197,N_8074,N_7885);
xor U8198 (N_8198,N_8052,N_7979);
nand U8199 (N_8199,N_7883,N_7815);
and U8200 (N_8200,N_7880,N_7853);
nor U8201 (N_8201,N_7877,N_7953);
or U8202 (N_8202,N_7970,N_7839);
nor U8203 (N_8203,N_7963,N_8026);
or U8204 (N_8204,N_7958,N_7846);
nand U8205 (N_8205,N_7864,N_8034);
nand U8206 (N_8206,N_8011,N_7807);
nand U8207 (N_8207,N_7826,N_7868);
or U8208 (N_8208,N_8018,N_8064);
or U8209 (N_8209,N_8038,N_8067);
or U8210 (N_8210,N_7805,N_8029);
xor U8211 (N_8211,N_8000,N_7873);
or U8212 (N_8212,N_8084,N_8094);
xor U8213 (N_8213,N_7923,N_8057);
or U8214 (N_8214,N_8051,N_8039);
or U8215 (N_8215,N_7993,N_8042);
or U8216 (N_8216,N_7921,N_7887);
or U8217 (N_8217,N_7932,N_7978);
nand U8218 (N_8218,N_7920,N_7947);
nor U8219 (N_8219,N_8032,N_8046);
xor U8220 (N_8220,N_7901,N_7983);
nor U8221 (N_8221,N_8010,N_7927);
nor U8222 (N_8222,N_7954,N_7998);
xor U8223 (N_8223,N_7936,N_7969);
or U8224 (N_8224,N_7861,N_8025);
or U8225 (N_8225,N_7929,N_8031);
nor U8226 (N_8226,N_7865,N_7917);
or U8227 (N_8227,N_7858,N_7905);
nand U8228 (N_8228,N_7930,N_7851);
nor U8229 (N_8229,N_7840,N_8075);
nand U8230 (N_8230,N_8079,N_7942);
or U8231 (N_8231,N_7893,N_7890);
or U8232 (N_8232,N_7975,N_8063);
xnor U8233 (N_8233,N_8006,N_7854);
xnor U8234 (N_8234,N_8014,N_8045);
and U8235 (N_8235,N_8004,N_8077);
and U8236 (N_8236,N_7867,N_7914);
nand U8237 (N_8237,N_8020,N_8085);
nand U8238 (N_8238,N_8091,N_7823);
nand U8239 (N_8239,N_7896,N_7950);
and U8240 (N_8240,N_8007,N_7847);
or U8241 (N_8241,N_7898,N_7817);
nand U8242 (N_8242,N_8093,N_7892);
xor U8243 (N_8243,N_7966,N_7934);
nor U8244 (N_8244,N_7972,N_7943);
nor U8245 (N_8245,N_8096,N_7955);
nand U8246 (N_8246,N_8089,N_7909);
or U8247 (N_8247,N_7816,N_7820);
nor U8248 (N_8248,N_7948,N_7852);
nor U8249 (N_8249,N_8003,N_8027);
or U8250 (N_8250,N_8062,N_8021);
nor U8251 (N_8251,N_8013,N_8099);
nand U8252 (N_8252,N_8011,N_7968);
or U8253 (N_8253,N_7996,N_7979);
or U8254 (N_8254,N_8079,N_7911);
and U8255 (N_8255,N_7925,N_8024);
nor U8256 (N_8256,N_8055,N_7801);
and U8257 (N_8257,N_8065,N_8044);
and U8258 (N_8258,N_8006,N_7909);
xnor U8259 (N_8259,N_7800,N_7848);
nand U8260 (N_8260,N_8043,N_7838);
nand U8261 (N_8261,N_7824,N_8084);
and U8262 (N_8262,N_8061,N_7892);
and U8263 (N_8263,N_7803,N_7816);
nand U8264 (N_8264,N_8095,N_7903);
or U8265 (N_8265,N_8082,N_7888);
xor U8266 (N_8266,N_7948,N_7927);
or U8267 (N_8267,N_7828,N_8029);
or U8268 (N_8268,N_7921,N_7955);
nor U8269 (N_8269,N_8089,N_7915);
nor U8270 (N_8270,N_7958,N_7829);
or U8271 (N_8271,N_7965,N_8037);
xnor U8272 (N_8272,N_8071,N_8085);
nor U8273 (N_8273,N_7803,N_8047);
or U8274 (N_8274,N_7950,N_7907);
nor U8275 (N_8275,N_8062,N_7840);
and U8276 (N_8276,N_7934,N_7978);
nor U8277 (N_8277,N_8098,N_7845);
and U8278 (N_8278,N_8096,N_7980);
nor U8279 (N_8279,N_7832,N_7873);
or U8280 (N_8280,N_7883,N_8097);
or U8281 (N_8281,N_7892,N_7885);
xnor U8282 (N_8282,N_7861,N_8044);
or U8283 (N_8283,N_8084,N_7856);
nand U8284 (N_8284,N_7883,N_8076);
xnor U8285 (N_8285,N_8054,N_8000);
xor U8286 (N_8286,N_8021,N_8011);
or U8287 (N_8287,N_7855,N_8024);
nor U8288 (N_8288,N_7888,N_8043);
and U8289 (N_8289,N_7898,N_7804);
nand U8290 (N_8290,N_7901,N_8004);
nand U8291 (N_8291,N_7868,N_8003);
nand U8292 (N_8292,N_7894,N_7924);
xnor U8293 (N_8293,N_7881,N_8061);
nor U8294 (N_8294,N_7903,N_7997);
nor U8295 (N_8295,N_8061,N_7814);
and U8296 (N_8296,N_7827,N_7840);
or U8297 (N_8297,N_7865,N_8092);
and U8298 (N_8298,N_7904,N_7819);
nor U8299 (N_8299,N_7903,N_7883);
or U8300 (N_8300,N_8031,N_8000);
nor U8301 (N_8301,N_7924,N_7905);
nand U8302 (N_8302,N_7949,N_7958);
or U8303 (N_8303,N_8099,N_7802);
nand U8304 (N_8304,N_7864,N_7883);
and U8305 (N_8305,N_7855,N_7821);
xor U8306 (N_8306,N_7827,N_7854);
nand U8307 (N_8307,N_7997,N_8038);
xnor U8308 (N_8308,N_7872,N_8068);
nand U8309 (N_8309,N_7899,N_7974);
or U8310 (N_8310,N_7985,N_7986);
nand U8311 (N_8311,N_7925,N_7920);
or U8312 (N_8312,N_8079,N_7822);
and U8313 (N_8313,N_8075,N_8038);
and U8314 (N_8314,N_7905,N_7872);
or U8315 (N_8315,N_7909,N_8080);
nor U8316 (N_8316,N_8066,N_8030);
xor U8317 (N_8317,N_8030,N_8048);
nand U8318 (N_8318,N_7971,N_7985);
or U8319 (N_8319,N_7913,N_7835);
nand U8320 (N_8320,N_7821,N_8050);
or U8321 (N_8321,N_7972,N_7820);
and U8322 (N_8322,N_7953,N_8099);
or U8323 (N_8323,N_8098,N_7898);
nand U8324 (N_8324,N_7997,N_8067);
nor U8325 (N_8325,N_8077,N_7955);
xnor U8326 (N_8326,N_8041,N_8086);
nor U8327 (N_8327,N_7889,N_7801);
nand U8328 (N_8328,N_8000,N_7921);
and U8329 (N_8329,N_7895,N_8007);
or U8330 (N_8330,N_7978,N_7966);
nand U8331 (N_8331,N_7860,N_7825);
or U8332 (N_8332,N_7908,N_8099);
nand U8333 (N_8333,N_7846,N_7898);
nand U8334 (N_8334,N_7828,N_7969);
xor U8335 (N_8335,N_7968,N_7939);
nand U8336 (N_8336,N_8004,N_7919);
and U8337 (N_8337,N_7915,N_7854);
nor U8338 (N_8338,N_7893,N_7869);
nand U8339 (N_8339,N_7980,N_8099);
or U8340 (N_8340,N_7864,N_7852);
xnor U8341 (N_8341,N_7847,N_7939);
nand U8342 (N_8342,N_7997,N_7849);
nor U8343 (N_8343,N_8058,N_7917);
xor U8344 (N_8344,N_7998,N_8031);
nand U8345 (N_8345,N_7896,N_8004);
and U8346 (N_8346,N_8097,N_8083);
nand U8347 (N_8347,N_8053,N_7960);
nand U8348 (N_8348,N_8076,N_7952);
and U8349 (N_8349,N_7845,N_7819);
xnor U8350 (N_8350,N_8031,N_7925);
and U8351 (N_8351,N_8066,N_7972);
and U8352 (N_8352,N_7801,N_7976);
and U8353 (N_8353,N_7862,N_7894);
nand U8354 (N_8354,N_7861,N_8005);
or U8355 (N_8355,N_7833,N_7891);
xnor U8356 (N_8356,N_7886,N_7807);
and U8357 (N_8357,N_7907,N_8034);
and U8358 (N_8358,N_7956,N_7885);
xnor U8359 (N_8359,N_7817,N_7837);
or U8360 (N_8360,N_8063,N_7917);
nor U8361 (N_8361,N_7990,N_8055);
nor U8362 (N_8362,N_7807,N_7961);
xor U8363 (N_8363,N_8082,N_8031);
nand U8364 (N_8364,N_7884,N_7905);
nor U8365 (N_8365,N_8045,N_7962);
nor U8366 (N_8366,N_7825,N_7820);
xor U8367 (N_8367,N_7952,N_8037);
nand U8368 (N_8368,N_7841,N_7831);
xor U8369 (N_8369,N_7995,N_8039);
and U8370 (N_8370,N_7917,N_7932);
nand U8371 (N_8371,N_7917,N_7862);
xnor U8372 (N_8372,N_8072,N_8000);
or U8373 (N_8373,N_7886,N_8038);
and U8374 (N_8374,N_7968,N_8007);
nand U8375 (N_8375,N_8033,N_7841);
xnor U8376 (N_8376,N_8088,N_8045);
or U8377 (N_8377,N_8020,N_7805);
xor U8378 (N_8378,N_7953,N_7854);
xor U8379 (N_8379,N_7850,N_7965);
and U8380 (N_8380,N_7820,N_7975);
xor U8381 (N_8381,N_7998,N_7926);
or U8382 (N_8382,N_7962,N_8049);
or U8383 (N_8383,N_7832,N_7974);
and U8384 (N_8384,N_7892,N_7925);
or U8385 (N_8385,N_7959,N_7865);
and U8386 (N_8386,N_7965,N_7812);
xnor U8387 (N_8387,N_8007,N_7912);
xor U8388 (N_8388,N_7864,N_7803);
nor U8389 (N_8389,N_7894,N_8025);
xor U8390 (N_8390,N_8083,N_7978);
nor U8391 (N_8391,N_7813,N_7858);
or U8392 (N_8392,N_7804,N_7830);
and U8393 (N_8393,N_7850,N_7974);
nor U8394 (N_8394,N_7833,N_8059);
and U8395 (N_8395,N_7941,N_8084);
and U8396 (N_8396,N_8026,N_7807);
or U8397 (N_8397,N_7937,N_7816);
and U8398 (N_8398,N_7991,N_7827);
nor U8399 (N_8399,N_7976,N_7879);
xnor U8400 (N_8400,N_8293,N_8265);
nor U8401 (N_8401,N_8239,N_8387);
nand U8402 (N_8402,N_8145,N_8247);
or U8403 (N_8403,N_8328,N_8207);
or U8404 (N_8404,N_8219,N_8297);
nor U8405 (N_8405,N_8267,N_8276);
and U8406 (N_8406,N_8223,N_8237);
and U8407 (N_8407,N_8235,N_8113);
nand U8408 (N_8408,N_8157,N_8316);
nand U8409 (N_8409,N_8136,N_8204);
nand U8410 (N_8410,N_8230,N_8282);
xnor U8411 (N_8411,N_8268,N_8289);
and U8412 (N_8412,N_8137,N_8330);
nor U8413 (N_8413,N_8240,N_8197);
and U8414 (N_8414,N_8349,N_8167);
and U8415 (N_8415,N_8103,N_8324);
xnor U8416 (N_8416,N_8250,N_8149);
or U8417 (N_8417,N_8307,N_8215);
nand U8418 (N_8418,N_8160,N_8394);
nor U8419 (N_8419,N_8181,N_8122);
nor U8420 (N_8420,N_8141,N_8382);
nand U8421 (N_8421,N_8143,N_8308);
and U8422 (N_8422,N_8364,N_8217);
nand U8423 (N_8423,N_8283,N_8298);
and U8424 (N_8424,N_8246,N_8114);
or U8425 (N_8425,N_8363,N_8377);
nor U8426 (N_8426,N_8241,N_8100);
xor U8427 (N_8427,N_8356,N_8198);
nand U8428 (N_8428,N_8390,N_8395);
or U8429 (N_8429,N_8288,N_8168);
nand U8430 (N_8430,N_8211,N_8385);
nor U8431 (N_8431,N_8106,N_8251);
nor U8432 (N_8432,N_8314,N_8109);
xnor U8433 (N_8433,N_8301,N_8108);
and U8434 (N_8434,N_8152,N_8373);
and U8435 (N_8435,N_8111,N_8202);
or U8436 (N_8436,N_8115,N_8337);
nand U8437 (N_8437,N_8357,N_8203);
xor U8438 (N_8438,N_8194,N_8131);
or U8439 (N_8439,N_8279,N_8233);
and U8440 (N_8440,N_8112,N_8275);
xnor U8441 (N_8441,N_8325,N_8124);
nand U8442 (N_8442,N_8133,N_8326);
or U8443 (N_8443,N_8192,N_8266);
and U8444 (N_8444,N_8256,N_8179);
nor U8445 (N_8445,N_8304,N_8205);
and U8446 (N_8446,N_8389,N_8333);
or U8447 (N_8447,N_8173,N_8386);
nor U8448 (N_8448,N_8225,N_8273);
and U8449 (N_8449,N_8105,N_8343);
xnor U8450 (N_8450,N_8370,N_8381);
and U8451 (N_8451,N_8231,N_8185);
xor U8452 (N_8452,N_8163,N_8290);
nor U8453 (N_8453,N_8366,N_8378);
nor U8454 (N_8454,N_8234,N_8208);
xnor U8455 (N_8455,N_8224,N_8148);
nor U8456 (N_8456,N_8201,N_8322);
xor U8457 (N_8457,N_8354,N_8218);
xor U8458 (N_8458,N_8156,N_8399);
xor U8459 (N_8459,N_8362,N_8147);
nor U8460 (N_8460,N_8153,N_8227);
and U8461 (N_8461,N_8398,N_8245);
xnor U8462 (N_8462,N_8269,N_8123);
or U8463 (N_8463,N_8117,N_8161);
xnor U8464 (N_8464,N_8359,N_8249);
nand U8465 (N_8465,N_8294,N_8263);
nand U8466 (N_8466,N_8150,N_8320);
nor U8467 (N_8467,N_8313,N_8391);
or U8468 (N_8468,N_8232,N_8174);
or U8469 (N_8469,N_8261,N_8210);
nor U8470 (N_8470,N_8209,N_8393);
or U8471 (N_8471,N_8158,N_8213);
xor U8472 (N_8472,N_8336,N_8144);
or U8473 (N_8473,N_8258,N_8272);
nor U8474 (N_8474,N_8236,N_8271);
and U8475 (N_8475,N_8396,N_8169);
and U8476 (N_8476,N_8116,N_8120);
xor U8477 (N_8477,N_8214,N_8392);
nor U8478 (N_8478,N_8128,N_8348);
or U8479 (N_8479,N_8342,N_8216);
or U8480 (N_8480,N_8278,N_8340);
xnor U8481 (N_8481,N_8255,N_8350);
xnor U8482 (N_8482,N_8339,N_8353);
nor U8483 (N_8483,N_8270,N_8369);
nor U8484 (N_8484,N_8193,N_8302);
nand U8485 (N_8485,N_8220,N_8196);
or U8486 (N_8486,N_8335,N_8191);
nor U8487 (N_8487,N_8321,N_8257);
and U8488 (N_8488,N_8190,N_8379);
and U8489 (N_8489,N_8332,N_8345);
xnor U8490 (N_8490,N_8125,N_8182);
nand U8491 (N_8491,N_8130,N_8187);
or U8492 (N_8492,N_8121,N_8380);
and U8493 (N_8493,N_8260,N_8281);
and U8494 (N_8494,N_8132,N_8178);
nor U8495 (N_8495,N_8154,N_8284);
or U8496 (N_8496,N_8329,N_8372);
and U8497 (N_8497,N_8368,N_8300);
or U8498 (N_8498,N_8338,N_8295);
and U8499 (N_8499,N_8280,N_8306);
nor U8500 (N_8500,N_8146,N_8129);
nand U8501 (N_8501,N_8311,N_8119);
xnor U8502 (N_8502,N_8199,N_8186);
nor U8503 (N_8503,N_8176,N_8228);
and U8504 (N_8504,N_8151,N_8375);
xor U8505 (N_8505,N_8262,N_8172);
and U8506 (N_8506,N_8101,N_8365);
nand U8507 (N_8507,N_8355,N_8159);
nand U8508 (N_8508,N_8162,N_8351);
xor U8509 (N_8509,N_8376,N_8274);
or U8510 (N_8510,N_8253,N_8110);
and U8511 (N_8511,N_8384,N_8327);
and U8512 (N_8512,N_8171,N_8277);
or U8513 (N_8513,N_8222,N_8102);
and U8514 (N_8514,N_8134,N_8212);
nor U8515 (N_8515,N_8170,N_8341);
or U8516 (N_8516,N_8259,N_8371);
nor U8517 (N_8517,N_8206,N_8286);
nor U8518 (N_8518,N_8383,N_8243);
xor U8519 (N_8519,N_8138,N_8177);
xnor U8520 (N_8520,N_8347,N_8299);
xor U8521 (N_8521,N_8305,N_8315);
xnor U8522 (N_8522,N_8244,N_8309);
and U8523 (N_8523,N_8140,N_8296);
nor U8524 (N_8524,N_8184,N_8226);
nor U8525 (N_8525,N_8254,N_8195);
and U8526 (N_8526,N_8200,N_8367);
nand U8527 (N_8527,N_8165,N_8118);
nand U8528 (N_8528,N_8323,N_8252);
or U8529 (N_8529,N_8318,N_8189);
and U8530 (N_8530,N_8248,N_8242);
nor U8531 (N_8531,N_8238,N_8388);
and U8532 (N_8532,N_8180,N_8107);
or U8533 (N_8533,N_8358,N_8303);
nor U8534 (N_8534,N_8352,N_8317);
nor U8535 (N_8535,N_8164,N_8135);
or U8536 (N_8536,N_8344,N_8175);
nand U8537 (N_8537,N_8319,N_8346);
nor U8538 (N_8538,N_8166,N_8287);
or U8539 (N_8539,N_8397,N_8126);
xor U8540 (N_8540,N_8264,N_8183);
or U8541 (N_8541,N_8331,N_8334);
and U8542 (N_8542,N_8127,N_8155);
and U8543 (N_8543,N_8188,N_8361);
xnor U8544 (N_8544,N_8312,N_8142);
and U8545 (N_8545,N_8139,N_8285);
nor U8546 (N_8546,N_8291,N_8374);
or U8547 (N_8547,N_8310,N_8104);
xnor U8548 (N_8548,N_8221,N_8229);
nor U8549 (N_8549,N_8292,N_8360);
and U8550 (N_8550,N_8230,N_8211);
nor U8551 (N_8551,N_8205,N_8361);
nand U8552 (N_8552,N_8147,N_8359);
and U8553 (N_8553,N_8134,N_8169);
nand U8554 (N_8554,N_8152,N_8200);
nand U8555 (N_8555,N_8286,N_8193);
or U8556 (N_8556,N_8332,N_8394);
nor U8557 (N_8557,N_8234,N_8114);
or U8558 (N_8558,N_8232,N_8357);
or U8559 (N_8559,N_8284,N_8148);
and U8560 (N_8560,N_8222,N_8218);
nand U8561 (N_8561,N_8200,N_8396);
xnor U8562 (N_8562,N_8160,N_8361);
xnor U8563 (N_8563,N_8182,N_8256);
nand U8564 (N_8564,N_8394,N_8241);
nand U8565 (N_8565,N_8257,N_8217);
xor U8566 (N_8566,N_8379,N_8325);
or U8567 (N_8567,N_8303,N_8204);
and U8568 (N_8568,N_8137,N_8196);
and U8569 (N_8569,N_8344,N_8136);
xnor U8570 (N_8570,N_8353,N_8295);
nand U8571 (N_8571,N_8106,N_8131);
nand U8572 (N_8572,N_8332,N_8359);
xor U8573 (N_8573,N_8228,N_8118);
and U8574 (N_8574,N_8169,N_8371);
xnor U8575 (N_8575,N_8309,N_8162);
or U8576 (N_8576,N_8253,N_8158);
nand U8577 (N_8577,N_8206,N_8146);
nand U8578 (N_8578,N_8356,N_8262);
nor U8579 (N_8579,N_8216,N_8360);
xnor U8580 (N_8580,N_8107,N_8235);
nand U8581 (N_8581,N_8298,N_8342);
and U8582 (N_8582,N_8320,N_8275);
and U8583 (N_8583,N_8380,N_8216);
and U8584 (N_8584,N_8189,N_8145);
and U8585 (N_8585,N_8179,N_8399);
nand U8586 (N_8586,N_8319,N_8333);
nor U8587 (N_8587,N_8110,N_8309);
or U8588 (N_8588,N_8263,N_8152);
or U8589 (N_8589,N_8121,N_8213);
nand U8590 (N_8590,N_8152,N_8178);
or U8591 (N_8591,N_8288,N_8304);
nor U8592 (N_8592,N_8397,N_8190);
and U8593 (N_8593,N_8394,N_8374);
nand U8594 (N_8594,N_8166,N_8386);
xor U8595 (N_8595,N_8193,N_8234);
xor U8596 (N_8596,N_8273,N_8390);
nor U8597 (N_8597,N_8180,N_8132);
nor U8598 (N_8598,N_8187,N_8174);
xnor U8599 (N_8599,N_8149,N_8122);
nand U8600 (N_8600,N_8318,N_8198);
or U8601 (N_8601,N_8269,N_8212);
or U8602 (N_8602,N_8300,N_8111);
nand U8603 (N_8603,N_8110,N_8183);
and U8604 (N_8604,N_8205,N_8218);
and U8605 (N_8605,N_8220,N_8360);
xnor U8606 (N_8606,N_8125,N_8374);
and U8607 (N_8607,N_8162,N_8183);
or U8608 (N_8608,N_8152,N_8214);
and U8609 (N_8609,N_8328,N_8166);
xnor U8610 (N_8610,N_8341,N_8295);
xnor U8611 (N_8611,N_8149,N_8354);
nor U8612 (N_8612,N_8388,N_8330);
xnor U8613 (N_8613,N_8376,N_8115);
or U8614 (N_8614,N_8140,N_8384);
nand U8615 (N_8615,N_8150,N_8203);
xnor U8616 (N_8616,N_8214,N_8165);
nor U8617 (N_8617,N_8272,N_8330);
xnor U8618 (N_8618,N_8202,N_8187);
xor U8619 (N_8619,N_8310,N_8247);
and U8620 (N_8620,N_8378,N_8308);
nor U8621 (N_8621,N_8393,N_8292);
and U8622 (N_8622,N_8390,N_8350);
xor U8623 (N_8623,N_8301,N_8182);
nand U8624 (N_8624,N_8324,N_8343);
nor U8625 (N_8625,N_8355,N_8217);
or U8626 (N_8626,N_8207,N_8234);
nand U8627 (N_8627,N_8122,N_8226);
xnor U8628 (N_8628,N_8303,N_8271);
nor U8629 (N_8629,N_8111,N_8266);
xnor U8630 (N_8630,N_8301,N_8308);
nor U8631 (N_8631,N_8223,N_8230);
xnor U8632 (N_8632,N_8161,N_8328);
and U8633 (N_8633,N_8343,N_8148);
nand U8634 (N_8634,N_8350,N_8182);
nor U8635 (N_8635,N_8102,N_8379);
nor U8636 (N_8636,N_8242,N_8387);
nand U8637 (N_8637,N_8251,N_8229);
nand U8638 (N_8638,N_8334,N_8321);
nor U8639 (N_8639,N_8192,N_8173);
or U8640 (N_8640,N_8169,N_8258);
or U8641 (N_8641,N_8102,N_8103);
xnor U8642 (N_8642,N_8291,N_8234);
xor U8643 (N_8643,N_8146,N_8209);
xnor U8644 (N_8644,N_8287,N_8283);
xnor U8645 (N_8645,N_8154,N_8244);
xnor U8646 (N_8646,N_8131,N_8301);
or U8647 (N_8647,N_8198,N_8340);
nor U8648 (N_8648,N_8226,N_8280);
nand U8649 (N_8649,N_8120,N_8113);
nand U8650 (N_8650,N_8302,N_8129);
nor U8651 (N_8651,N_8370,N_8358);
xnor U8652 (N_8652,N_8346,N_8127);
nand U8653 (N_8653,N_8224,N_8388);
nor U8654 (N_8654,N_8319,N_8183);
and U8655 (N_8655,N_8362,N_8112);
or U8656 (N_8656,N_8240,N_8148);
or U8657 (N_8657,N_8285,N_8119);
nor U8658 (N_8658,N_8323,N_8385);
xnor U8659 (N_8659,N_8222,N_8350);
xnor U8660 (N_8660,N_8176,N_8135);
or U8661 (N_8661,N_8378,N_8159);
or U8662 (N_8662,N_8139,N_8289);
nor U8663 (N_8663,N_8165,N_8318);
xor U8664 (N_8664,N_8150,N_8172);
xor U8665 (N_8665,N_8187,N_8157);
or U8666 (N_8666,N_8391,N_8257);
xnor U8667 (N_8667,N_8329,N_8138);
or U8668 (N_8668,N_8395,N_8112);
or U8669 (N_8669,N_8179,N_8190);
and U8670 (N_8670,N_8214,N_8286);
and U8671 (N_8671,N_8379,N_8204);
and U8672 (N_8672,N_8222,N_8229);
nand U8673 (N_8673,N_8333,N_8275);
or U8674 (N_8674,N_8359,N_8309);
and U8675 (N_8675,N_8185,N_8340);
xor U8676 (N_8676,N_8252,N_8104);
nor U8677 (N_8677,N_8146,N_8342);
nor U8678 (N_8678,N_8384,N_8245);
or U8679 (N_8679,N_8242,N_8163);
xor U8680 (N_8680,N_8252,N_8273);
nor U8681 (N_8681,N_8138,N_8224);
xnor U8682 (N_8682,N_8212,N_8337);
and U8683 (N_8683,N_8339,N_8377);
nor U8684 (N_8684,N_8305,N_8300);
nor U8685 (N_8685,N_8144,N_8100);
or U8686 (N_8686,N_8110,N_8232);
and U8687 (N_8687,N_8266,N_8373);
or U8688 (N_8688,N_8346,N_8353);
nor U8689 (N_8689,N_8297,N_8147);
and U8690 (N_8690,N_8157,N_8238);
or U8691 (N_8691,N_8377,N_8168);
or U8692 (N_8692,N_8389,N_8194);
and U8693 (N_8693,N_8169,N_8331);
nor U8694 (N_8694,N_8305,N_8243);
or U8695 (N_8695,N_8174,N_8220);
xor U8696 (N_8696,N_8193,N_8397);
xor U8697 (N_8697,N_8286,N_8290);
and U8698 (N_8698,N_8215,N_8249);
nor U8699 (N_8699,N_8217,N_8226);
or U8700 (N_8700,N_8572,N_8614);
or U8701 (N_8701,N_8639,N_8622);
nor U8702 (N_8702,N_8451,N_8549);
or U8703 (N_8703,N_8441,N_8477);
xor U8704 (N_8704,N_8541,N_8499);
nor U8705 (N_8705,N_8576,N_8450);
xnor U8706 (N_8706,N_8400,N_8519);
xor U8707 (N_8707,N_8508,N_8408);
or U8708 (N_8708,N_8427,N_8438);
xnor U8709 (N_8709,N_8570,N_8442);
and U8710 (N_8710,N_8401,N_8613);
nand U8711 (N_8711,N_8533,N_8555);
or U8712 (N_8712,N_8635,N_8697);
and U8713 (N_8713,N_8542,N_8421);
or U8714 (N_8714,N_8603,N_8654);
nand U8715 (N_8715,N_8470,N_8688);
and U8716 (N_8716,N_8648,N_8534);
nor U8717 (N_8717,N_8678,N_8655);
nand U8718 (N_8718,N_8522,N_8556);
or U8719 (N_8719,N_8406,N_8646);
xor U8720 (N_8720,N_8524,N_8620);
and U8721 (N_8721,N_8457,N_8439);
xnor U8722 (N_8722,N_8590,N_8405);
or U8723 (N_8723,N_8540,N_8568);
or U8724 (N_8724,N_8452,N_8619);
or U8725 (N_8725,N_8559,N_8530);
and U8726 (N_8726,N_8505,N_8504);
nand U8727 (N_8727,N_8604,N_8468);
nor U8728 (N_8728,N_8448,N_8480);
nor U8729 (N_8729,N_8637,N_8666);
or U8730 (N_8730,N_8463,N_8691);
and U8731 (N_8731,N_8511,N_8615);
or U8732 (N_8732,N_8544,N_8523);
and U8733 (N_8733,N_8644,N_8626);
nand U8734 (N_8734,N_8415,N_8445);
and U8735 (N_8735,N_8512,N_8669);
xnor U8736 (N_8736,N_8684,N_8675);
nor U8737 (N_8737,N_8539,N_8548);
and U8738 (N_8738,N_8699,N_8687);
xor U8739 (N_8739,N_8485,N_8643);
nand U8740 (N_8740,N_8492,N_8525);
nor U8741 (N_8741,N_8526,N_8419);
or U8742 (N_8742,N_8591,N_8597);
and U8743 (N_8743,N_8586,N_8612);
xnor U8744 (N_8744,N_8671,N_8552);
nor U8745 (N_8745,N_8589,N_8667);
and U8746 (N_8746,N_8436,N_8564);
xor U8747 (N_8747,N_8455,N_8404);
or U8748 (N_8748,N_8543,N_8513);
nand U8749 (N_8749,N_8469,N_8488);
or U8750 (N_8750,N_8577,N_8449);
nor U8751 (N_8751,N_8690,N_8420);
or U8752 (N_8752,N_8502,N_8453);
nor U8753 (N_8753,N_8557,N_8497);
or U8754 (N_8754,N_8696,N_8633);
or U8755 (N_8755,N_8662,N_8608);
nand U8756 (N_8756,N_8647,N_8661);
xnor U8757 (N_8757,N_8645,N_8573);
and U8758 (N_8758,N_8531,N_8680);
and U8759 (N_8759,N_8514,N_8657);
nor U8760 (N_8760,N_8641,N_8429);
xor U8761 (N_8761,N_8658,N_8506);
nand U8762 (N_8762,N_8430,N_8456);
nor U8763 (N_8763,N_8592,N_8528);
nor U8764 (N_8764,N_8625,N_8536);
xor U8765 (N_8765,N_8414,N_8495);
or U8766 (N_8766,N_8618,N_8546);
or U8767 (N_8767,N_8659,N_8474);
nand U8768 (N_8768,N_8676,N_8407);
or U8769 (N_8769,N_8631,N_8518);
and U8770 (N_8770,N_8493,N_8561);
nor U8771 (N_8771,N_8642,N_8563);
xor U8772 (N_8772,N_8571,N_8607);
xor U8773 (N_8773,N_8532,N_8417);
nand U8774 (N_8774,N_8566,N_8692);
nand U8775 (N_8775,N_8446,N_8464);
xnor U8776 (N_8776,N_8527,N_8550);
or U8777 (N_8777,N_8634,N_8409);
and U8778 (N_8778,N_8670,N_8652);
xor U8779 (N_8779,N_8695,N_8567);
and U8780 (N_8780,N_8594,N_8489);
nor U8781 (N_8781,N_8569,N_8606);
or U8782 (N_8782,N_8616,N_8610);
and U8783 (N_8783,N_8585,N_8593);
nand U8784 (N_8784,N_8412,N_8627);
xor U8785 (N_8785,N_8423,N_8600);
or U8786 (N_8786,N_8459,N_8575);
or U8787 (N_8787,N_8598,N_8458);
xnor U8788 (N_8788,N_8490,N_8460);
and U8789 (N_8789,N_8617,N_8581);
nand U8790 (N_8790,N_8478,N_8413);
xor U8791 (N_8791,N_8596,N_8500);
nor U8792 (N_8792,N_8483,N_8595);
xor U8793 (N_8793,N_8579,N_8694);
xnor U8794 (N_8794,N_8501,N_8698);
nand U8795 (N_8795,N_8447,N_8584);
xor U8796 (N_8796,N_8693,N_8599);
and U8797 (N_8797,N_8624,N_8679);
nor U8798 (N_8798,N_8665,N_8565);
nor U8799 (N_8799,N_8491,N_8481);
xnor U8800 (N_8800,N_8416,N_8580);
or U8801 (N_8801,N_8475,N_8529);
and U8802 (N_8802,N_8686,N_8578);
nand U8803 (N_8803,N_8660,N_8473);
and U8804 (N_8804,N_8547,N_8682);
xnor U8805 (N_8805,N_8560,N_8621);
nor U8806 (N_8806,N_8588,N_8426);
nand U8807 (N_8807,N_8437,N_8486);
or U8808 (N_8808,N_8681,N_8471);
xor U8809 (N_8809,N_8650,N_8515);
nor U8810 (N_8810,N_8444,N_8428);
and U8811 (N_8811,N_8454,N_8602);
xnor U8812 (N_8812,N_8609,N_8461);
nand U8813 (N_8813,N_8443,N_8494);
nand U8814 (N_8814,N_8551,N_8554);
nor U8815 (N_8815,N_8677,N_8465);
nor U8816 (N_8816,N_8663,N_8668);
nand U8817 (N_8817,N_8630,N_8587);
and U8818 (N_8818,N_8418,N_8611);
nor U8819 (N_8819,N_8649,N_8651);
and U8820 (N_8820,N_8664,N_8507);
nor U8821 (N_8821,N_8623,N_8672);
xor U8822 (N_8822,N_8479,N_8435);
and U8823 (N_8823,N_8410,N_8628);
nor U8824 (N_8824,N_8476,N_8520);
and U8825 (N_8825,N_8673,N_8605);
nor U8826 (N_8826,N_8509,N_8640);
or U8827 (N_8827,N_8538,N_8462);
and U8828 (N_8828,N_8403,N_8434);
nor U8829 (N_8829,N_8425,N_8422);
nor U8830 (N_8830,N_8498,N_8601);
nand U8831 (N_8831,N_8482,N_8562);
xnor U8832 (N_8832,N_8685,N_8411);
nor U8833 (N_8833,N_8484,N_8583);
xnor U8834 (N_8834,N_8433,N_8510);
or U8835 (N_8835,N_8632,N_8466);
and U8836 (N_8836,N_8440,N_8402);
and U8837 (N_8837,N_8517,N_8674);
xor U8838 (N_8838,N_8656,N_8521);
xor U8839 (N_8839,N_8545,N_8472);
and U8840 (N_8840,N_8558,N_8537);
nor U8841 (N_8841,N_8467,N_8638);
and U8842 (N_8842,N_8535,N_8582);
or U8843 (N_8843,N_8516,N_8432);
nor U8844 (N_8844,N_8683,N_8689);
xnor U8845 (N_8845,N_8424,N_8653);
xor U8846 (N_8846,N_8503,N_8574);
and U8847 (N_8847,N_8487,N_8431);
nor U8848 (N_8848,N_8496,N_8553);
xor U8849 (N_8849,N_8636,N_8629);
and U8850 (N_8850,N_8664,N_8631);
and U8851 (N_8851,N_8561,N_8617);
and U8852 (N_8852,N_8642,N_8616);
nand U8853 (N_8853,N_8557,N_8595);
nand U8854 (N_8854,N_8574,N_8543);
nand U8855 (N_8855,N_8490,N_8622);
nor U8856 (N_8856,N_8522,N_8428);
or U8857 (N_8857,N_8685,N_8635);
xor U8858 (N_8858,N_8560,N_8427);
and U8859 (N_8859,N_8473,N_8494);
nand U8860 (N_8860,N_8446,N_8682);
and U8861 (N_8861,N_8639,N_8500);
nor U8862 (N_8862,N_8692,N_8509);
and U8863 (N_8863,N_8590,N_8665);
or U8864 (N_8864,N_8415,N_8532);
and U8865 (N_8865,N_8630,N_8453);
or U8866 (N_8866,N_8692,N_8560);
xor U8867 (N_8867,N_8405,N_8685);
nand U8868 (N_8868,N_8654,N_8656);
or U8869 (N_8869,N_8615,N_8648);
nand U8870 (N_8870,N_8492,N_8507);
nand U8871 (N_8871,N_8504,N_8585);
or U8872 (N_8872,N_8574,N_8542);
nor U8873 (N_8873,N_8523,N_8681);
nor U8874 (N_8874,N_8479,N_8641);
or U8875 (N_8875,N_8593,N_8517);
xor U8876 (N_8876,N_8419,N_8546);
xor U8877 (N_8877,N_8542,N_8660);
nand U8878 (N_8878,N_8592,N_8685);
nand U8879 (N_8879,N_8627,N_8626);
nor U8880 (N_8880,N_8570,N_8481);
nand U8881 (N_8881,N_8557,N_8587);
xor U8882 (N_8882,N_8444,N_8511);
or U8883 (N_8883,N_8414,N_8690);
or U8884 (N_8884,N_8695,N_8592);
and U8885 (N_8885,N_8450,N_8669);
xnor U8886 (N_8886,N_8578,N_8442);
nor U8887 (N_8887,N_8636,N_8447);
nor U8888 (N_8888,N_8451,N_8687);
nand U8889 (N_8889,N_8688,N_8427);
xor U8890 (N_8890,N_8688,N_8404);
and U8891 (N_8891,N_8519,N_8595);
and U8892 (N_8892,N_8468,N_8534);
nor U8893 (N_8893,N_8530,N_8516);
nand U8894 (N_8894,N_8424,N_8515);
xnor U8895 (N_8895,N_8401,N_8501);
nor U8896 (N_8896,N_8695,N_8612);
nor U8897 (N_8897,N_8552,N_8622);
nor U8898 (N_8898,N_8449,N_8582);
nor U8899 (N_8899,N_8425,N_8462);
nor U8900 (N_8900,N_8527,N_8696);
nand U8901 (N_8901,N_8540,N_8455);
nand U8902 (N_8902,N_8695,N_8439);
or U8903 (N_8903,N_8544,N_8683);
or U8904 (N_8904,N_8546,N_8520);
or U8905 (N_8905,N_8510,N_8518);
xnor U8906 (N_8906,N_8429,N_8415);
nor U8907 (N_8907,N_8446,N_8496);
nor U8908 (N_8908,N_8414,N_8560);
nor U8909 (N_8909,N_8688,N_8492);
and U8910 (N_8910,N_8577,N_8442);
nor U8911 (N_8911,N_8411,N_8491);
or U8912 (N_8912,N_8584,N_8572);
or U8913 (N_8913,N_8403,N_8602);
and U8914 (N_8914,N_8602,N_8406);
nor U8915 (N_8915,N_8669,N_8457);
nor U8916 (N_8916,N_8677,N_8646);
xor U8917 (N_8917,N_8624,N_8623);
or U8918 (N_8918,N_8648,N_8595);
or U8919 (N_8919,N_8434,N_8541);
xor U8920 (N_8920,N_8403,N_8665);
nand U8921 (N_8921,N_8566,N_8518);
and U8922 (N_8922,N_8422,N_8612);
xor U8923 (N_8923,N_8573,N_8568);
nand U8924 (N_8924,N_8661,N_8434);
nand U8925 (N_8925,N_8455,N_8612);
nor U8926 (N_8926,N_8610,N_8641);
nand U8927 (N_8927,N_8682,N_8641);
nor U8928 (N_8928,N_8444,N_8653);
nand U8929 (N_8929,N_8679,N_8664);
nand U8930 (N_8930,N_8480,N_8587);
xnor U8931 (N_8931,N_8446,N_8640);
nand U8932 (N_8932,N_8620,N_8523);
or U8933 (N_8933,N_8607,N_8532);
nand U8934 (N_8934,N_8404,N_8539);
and U8935 (N_8935,N_8422,N_8539);
and U8936 (N_8936,N_8665,N_8442);
and U8937 (N_8937,N_8479,N_8457);
nand U8938 (N_8938,N_8513,N_8411);
nor U8939 (N_8939,N_8509,N_8413);
nor U8940 (N_8940,N_8452,N_8427);
xnor U8941 (N_8941,N_8510,N_8673);
or U8942 (N_8942,N_8527,N_8611);
nand U8943 (N_8943,N_8674,N_8553);
or U8944 (N_8944,N_8658,N_8641);
nand U8945 (N_8945,N_8591,N_8400);
or U8946 (N_8946,N_8432,N_8665);
nand U8947 (N_8947,N_8685,N_8471);
or U8948 (N_8948,N_8451,N_8672);
nor U8949 (N_8949,N_8510,N_8593);
xnor U8950 (N_8950,N_8500,N_8417);
nor U8951 (N_8951,N_8635,N_8666);
xor U8952 (N_8952,N_8534,N_8636);
or U8953 (N_8953,N_8425,N_8679);
nand U8954 (N_8954,N_8682,N_8455);
nand U8955 (N_8955,N_8593,N_8567);
nor U8956 (N_8956,N_8645,N_8432);
xnor U8957 (N_8957,N_8500,N_8698);
nor U8958 (N_8958,N_8522,N_8503);
nor U8959 (N_8959,N_8402,N_8553);
nor U8960 (N_8960,N_8657,N_8649);
nand U8961 (N_8961,N_8508,N_8421);
xor U8962 (N_8962,N_8555,N_8462);
and U8963 (N_8963,N_8543,N_8559);
nand U8964 (N_8964,N_8545,N_8697);
or U8965 (N_8965,N_8658,N_8527);
and U8966 (N_8966,N_8417,N_8498);
and U8967 (N_8967,N_8439,N_8458);
and U8968 (N_8968,N_8570,N_8468);
nand U8969 (N_8969,N_8604,N_8567);
xor U8970 (N_8970,N_8627,N_8678);
xor U8971 (N_8971,N_8659,N_8499);
and U8972 (N_8972,N_8630,N_8428);
nand U8973 (N_8973,N_8654,N_8437);
nor U8974 (N_8974,N_8441,N_8575);
and U8975 (N_8975,N_8614,N_8427);
xnor U8976 (N_8976,N_8537,N_8471);
nand U8977 (N_8977,N_8454,N_8421);
nor U8978 (N_8978,N_8541,N_8453);
xnor U8979 (N_8979,N_8518,N_8685);
nor U8980 (N_8980,N_8638,N_8432);
xor U8981 (N_8981,N_8404,N_8522);
and U8982 (N_8982,N_8439,N_8553);
or U8983 (N_8983,N_8603,N_8538);
xor U8984 (N_8984,N_8435,N_8533);
or U8985 (N_8985,N_8515,N_8429);
nor U8986 (N_8986,N_8579,N_8578);
xor U8987 (N_8987,N_8664,N_8528);
nand U8988 (N_8988,N_8645,N_8647);
and U8989 (N_8989,N_8583,N_8689);
nor U8990 (N_8990,N_8491,N_8573);
nand U8991 (N_8991,N_8589,N_8556);
or U8992 (N_8992,N_8635,N_8698);
and U8993 (N_8993,N_8445,N_8540);
xnor U8994 (N_8994,N_8443,N_8549);
or U8995 (N_8995,N_8531,N_8643);
nand U8996 (N_8996,N_8690,N_8554);
nand U8997 (N_8997,N_8409,N_8528);
xnor U8998 (N_8998,N_8574,N_8455);
nand U8999 (N_8999,N_8644,N_8683);
nand U9000 (N_9000,N_8833,N_8931);
and U9001 (N_9001,N_8792,N_8707);
nor U9002 (N_9002,N_8969,N_8848);
xnor U9003 (N_9003,N_8800,N_8837);
or U9004 (N_9004,N_8738,N_8722);
nand U9005 (N_9005,N_8902,N_8885);
or U9006 (N_9006,N_8730,N_8739);
nor U9007 (N_9007,N_8899,N_8794);
xnor U9008 (N_9008,N_8727,N_8766);
nand U9009 (N_9009,N_8881,N_8988);
nor U9010 (N_9010,N_8838,N_8767);
and U9011 (N_9011,N_8765,N_8701);
nand U9012 (N_9012,N_8956,N_8940);
nand U9013 (N_9013,N_8753,N_8732);
nand U9014 (N_9014,N_8923,N_8777);
xor U9015 (N_9015,N_8776,N_8803);
and U9016 (N_9016,N_8755,N_8799);
nor U9017 (N_9017,N_8933,N_8890);
xor U9018 (N_9018,N_8895,N_8867);
nor U9019 (N_9019,N_8834,N_8851);
nand U9020 (N_9020,N_8912,N_8966);
and U9021 (N_9021,N_8789,N_8760);
nor U9022 (N_9022,N_8754,N_8712);
or U9023 (N_9023,N_8791,N_8770);
or U9024 (N_9024,N_8886,N_8802);
xor U9025 (N_9025,N_8807,N_8823);
or U9026 (N_9026,N_8728,N_8769);
nor U9027 (N_9027,N_8781,N_8904);
and U9028 (N_9028,N_8909,N_8716);
or U9029 (N_9029,N_8978,N_8845);
xor U9030 (N_9030,N_8897,N_8748);
nor U9031 (N_9031,N_8979,N_8925);
nor U9032 (N_9032,N_8873,N_8758);
xnor U9033 (N_9033,N_8733,N_8872);
xor U9034 (N_9034,N_8962,N_8827);
nand U9035 (N_9035,N_8907,N_8920);
or U9036 (N_9036,N_8945,N_8847);
and U9037 (N_9037,N_8868,N_8718);
nand U9038 (N_9038,N_8968,N_8866);
or U9039 (N_9039,N_8936,N_8939);
nand U9040 (N_9040,N_8858,N_8922);
xnor U9041 (N_9041,N_8926,N_8976);
nor U9042 (N_9042,N_8786,N_8859);
or U9043 (N_9043,N_8999,N_8764);
nand U9044 (N_9044,N_8879,N_8977);
and U9045 (N_9045,N_8793,N_8884);
nand U9046 (N_9046,N_8841,N_8743);
or U9047 (N_9047,N_8970,N_8832);
nor U9048 (N_9048,N_8741,N_8975);
nand U9049 (N_9049,N_8715,N_8842);
and U9050 (N_9050,N_8919,N_8959);
and U9051 (N_9051,N_8856,N_8958);
nand U9052 (N_9052,N_8844,N_8865);
nand U9053 (N_9053,N_8757,N_8759);
and U9054 (N_9054,N_8949,N_8903);
or U9055 (N_9055,N_8729,N_8984);
xor U9056 (N_9056,N_8714,N_8994);
nor U9057 (N_9057,N_8952,N_8773);
or U9058 (N_9058,N_8982,N_8960);
nand U9059 (N_9059,N_8908,N_8826);
xnor U9060 (N_9060,N_8702,N_8893);
nor U9061 (N_9061,N_8849,N_8916);
or U9062 (N_9062,N_8756,N_8947);
nand U9063 (N_9063,N_8888,N_8783);
nor U9064 (N_9064,N_8967,N_8915);
nor U9065 (N_9065,N_8941,N_8705);
xor U9066 (N_9066,N_8991,N_8804);
and U9067 (N_9067,N_8942,N_8986);
nor U9068 (N_9068,N_8906,N_8708);
nand U9069 (N_9069,N_8911,N_8980);
nand U9070 (N_9070,N_8700,N_8752);
nand U9071 (N_9071,N_8720,N_8948);
and U9072 (N_9072,N_8735,N_8882);
nor U9073 (N_9073,N_8816,N_8726);
nand U9074 (N_9074,N_8955,N_8734);
xnor U9075 (N_9075,N_8921,N_8954);
nor U9076 (N_9076,N_8957,N_8820);
nand U9077 (N_9077,N_8853,N_8987);
nand U9078 (N_9078,N_8742,N_8993);
or U9079 (N_9079,N_8740,N_8787);
nand U9080 (N_9080,N_8717,N_8796);
or U9081 (N_9081,N_8905,N_8703);
and U9082 (N_9082,N_8883,N_8965);
nor U9083 (N_9083,N_8797,N_8749);
and U9084 (N_9084,N_8795,N_8953);
and U9085 (N_9085,N_8724,N_8710);
nor U9086 (N_9086,N_8798,N_8812);
nand U9087 (N_9087,N_8736,N_8721);
or U9088 (N_9088,N_8778,N_8870);
nand U9089 (N_9089,N_8857,N_8854);
nand U9090 (N_9090,N_8861,N_8963);
nand U9091 (N_9091,N_8880,N_8863);
xor U9092 (N_9092,N_8896,N_8917);
or U9093 (N_9093,N_8995,N_8788);
nor U9094 (N_9094,N_8779,N_8864);
or U9095 (N_9095,N_8876,N_8985);
and U9096 (N_9096,N_8805,N_8889);
or U9097 (N_9097,N_8981,N_8846);
nor U9098 (N_9098,N_8815,N_8709);
and U9099 (N_9099,N_8898,N_8747);
nor U9100 (N_9100,N_8725,N_8819);
nor U9101 (N_9101,N_8751,N_8871);
and U9102 (N_9102,N_8840,N_8943);
nand U9103 (N_9103,N_8768,N_8887);
or U9104 (N_9104,N_8964,N_8878);
and U9105 (N_9105,N_8811,N_8744);
and U9106 (N_9106,N_8813,N_8763);
nor U9107 (N_9107,N_8824,N_8998);
and U9108 (N_9108,N_8713,N_8852);
or U9109 (N_9109,N_8706,N_8737);
nor U9110 (N_9110,N_8996,N_8782);
nand U9111 (N_9111,N_8875,N_8771);
xor U9112 (N_9112,N_8900,N_8990);
or U9113 (N_9113,N_8946,N_8892);
nand U9114 (N_9114,N_8828,N_8901);
nand U9115 (N_9115,N_8938,N_8806);
nand U9116 (N_9116,N_8830,N_8731);
xor U9117 (N_9117,N_8814,N_8809);
nor U9118 (N_9118,N_8997,N_8790);
or U9119 (N_9119,N_8745,N_8989);
xor U9120 (N_9120,N_8932,N_8808);
and U9121 (N_9121,N_8704,N_8860);
or U9122 (N_9122,N_8924,N_8877);
nand U9123 (N_9123,N_8821,N_8831);
nand U9124 (N_9124,N_8874,N_8850);
and U9125 (N_9125,N_8910,N_8918);
xor U9126 (N_9126,N_8891,N_8855);
nand U9127 (N_9127,N_8974,N_8930);
or U9128 (N_9128,N_8972,N_8784);
and U9129 (N_9129,N_8762,N_8914);
and U9130 (N_9130,N_8934,N_8927);
xor U9131 (N_9131,N_8810,N_8818);
or U9132 (N_9132,N_8775,N_8913);
and U9133 (N_9133,N_8774,N_8822);
nand U9134 (N_9134,N_8973,N_8983);
and U9135 (N_9135,N_8817,N_8825);
nand U9136 (N_9136,N_8835,N_8894);
nor U9137 (N_9137,N_8935,N_8992);
and U9138 (N_9138,N_8711,N_8929);
or U9139 (N_9139,N_8843,N_8761);
or U9140 (N_9140,N_8723,N_8869);
or U9141 (N_9141,N_8937,N_8961);
or U9142 (N_9142,N_8839,N_8836);
xnor U9143 (N_9143,N_8829,N_8772);
and U9144 (N_9144,N_8971,N_8785);
or U9145 (N_9145,N_8951,N_8862);
or U9146 (N_9146,N_8780,N_8944);
and U9147 (N_9147,N_8928,N_8801);
nand U9148 (N_9148,N_8950,N_8750);
and U9149 (N_9149,N_8719,N_8746);
nand U9150 (N_9150,N_8914,N_8893);
or U9151 (N_9151,N_8761,N_8759);
xnor U9152 (N_9152,N_8927,N_8903);
nor U9153 (N_9153,N_8854,N_8745);
or U9154 (N_9154,N_8874,N_8898);
nand U9155 (N_9155,N_8895,N_8728);
xor U9156 (N_9156,N_8808,N_8969);
nand U9157 (N_9157,N_8935,N_8752);
nor U9158 (N_9158,N_8976,N_8717);
nor U9159 (N_9159,N_8847,N_8711);
and U9160 (N_9160,N_8733,N_8738);
xor U9161 (N_9161,N_8783,N_8983);
nand U9162 (N_9162,N_8913,N_8971);
xor U9163 (N_9163,N_8711,N_8899);
nor U9164 (N_9164,N_8957,N_8789);
nand U9165 (N_9165,N_8951,N_8999);
nor U9166 (N_9166,N_8946,N_8790);
nand U9167 (N_9167,N_8925,N_8976);
and U9168 (N_9168,N_8761,N_8818);
xnor U9169 (N_9169,N_8772,N_8927);
and U9170 (N_9170,N_8905,N_8881);
nor U9171 (N_9171,N_8914,N_8701);
or U9172 (N_9172,N_8908,N_8882);
nor U9173 (N_9173,N_8732,N_8830);
nand U9174 (N_9174,N_8898,N_8818);
or U9175 (N_9175,N_8845,N_8702);
nor U9176 (N_9176,N_8879,N_8947);
nor U9177 (N_9177,N_8969,N_8998);
and U9178 (N_9178,N_8848,N_8981);
xnor U9179 (N_9179,N_8876,N_8964);
and U9180 (N_9180,N_8789,N_8903);
or U9181 (N_9181,N_8747,N_8845);
or U9182 (N_9182,N_8709,N_8706);
nor U9183 (N_9183,N_8897,N_8709);
nand U9184 (N_9184,N_8890,N_8796);
or U9185 (N_9185,N_8987,N_8966);
nand U9186 (N_9186,N_8889,N_8874);
nor U9187 (N_9187,N_8720,N_8826);
xnor U9188 (N_9188,N_8835,N_8918);
or U9189 (N_9189,N_8760,N_8917);
nand U9190 (N_9190,N_8904,N_8744);
and U9191 (N_9191,N_8857,N_8751);
nand U9192 (N_9192,N_8881,N_8737);
nor U9193 (N_9193,N_8776,N_8857);
xor U9194 (N_9194,N_8916,N_8754);
xor U9195 (N_9195,N_8887,N_8931);
xor U9196 (N_9196,N_8755,N_8813);
nand U9197 (N_9197,N_8809,N_8813);
nor U9198 (N_9198,N_8722,N_8880);
xnor U9199 (N_9199,N_8786,N_8838);
nand U9200 (N_9200,N_8859,N_8966);
and U9201 (N_9201,N_8723,N_8978);
or U9202 (N_9202,N_8997,N_8951);
nor U9203 (N_9203,N_8833,N_8786);
nor U9204 (N_9204,N_8777,N_8738);
and U9205 (N_9205,N_8732,N_8799);
or U9206 (N_9206,N_8858,N_8925);
nor U9207 (N_9207,N_8759,N_8843);
nand U9208 (N_9208,N_8997,N_8877);
or U9209 (N_9209,N_8837,N_8925);
and U9210 (N_9210,N_8832,N_8737);
nor U9211 (N_9211,N_8873,N_8973);
nand U9212 (N_9212,N_8798,N_8711);
and U9213 (N_9213,N_8933,N_8797);
and U9214 (N_9214,N_8819,N_8708);
nand U9215 (N_9215,N_8943,N_8947);
or U9216 (N_9216,N_8873,N_8809);
and U9217 (N_9217,N_8948,N_8916);
and U9218 (N_9218,N_8905,N_8946);
xor U9219 (N_9219,N_8998,N_8999);
xnor U9220 (N_9220,N_8984,N_8919);
xor U9221 (N_9221,N_8750,N_8900);
and U9222 (N_9222,N_8895,N_8845);
and U9223 (N_9223,N_8701,N_8703);
or U9224 (N_9224,N_8980,N_8837);
nand U9225 (N_9225,N_8812,N_8771);
xor U9226 (N_9226,N_8875,N_8911);
nand U9227 (N_9227,N_8742,N_8924);
or U9228 (N_9228,N_8770,N_8906);
nor U9229 (N_9229,N_8997,N_8724);
and U9230 (N_9230,N_8727,N_8946);
or U9231 (N_9231,N_8787,N_8798);
nor U9232 (N_9232,N_8702,N_8915);
and U9233 (N_9233,N_8949,N_8856);
or U9234 (N_9234,N_8932,N_8987);
nor U9235 (N_9235,N_8981,N_8821);
xor U9236 (N_9236,N_8940,N_8777);
nor U9237 (N_9237,N_8950,N_8713);
and U9238 (N_9238,N_8760,N_8812);
xor U9239 (N_9239,N_8908,N_8890);
nor U9240 (N_9240,N_8738,N_8729);
nor U9241 (N_9241,N_8825,N_8822);
nand U9242 (N_9242,N_8713,N_8884);
nand U9243 (N_9243,N_8955,N_8874);
nand U9244 (N_9244,N_8795,N_8979);
nand U9245 (N_9245,N_8777,N_8842);
nor U9246 (N_9246,N_8973,N_8803);
xor U9247 (N_9247,N_8733,N_8744);
nor U9248 (N_9248,N_8756,N_8856);
or U9249 (N_9249,N_8991,N_8952);
or U9250 (N_9250,N_8973,N_8855);
nor U9251 (N_9251,N_8732,N_8875);
and U9252 (N_9252,N_8849,N_8747);
nand U9253 (N_9253,N_8961,N_8846);
nand U9254 (N_9254,N_8968,N_8732);
nor U9255 (N_9255,N_8998,N_8843);
or U9256 (N_9256,N_8755,N_8893);
nand U9257 (N_9257,N_8810,N_8853);
nor U9258 (N_9258,N_8903,N_8958);
and U9259 (N_9259,N_8750,N_8909);
and U9260 (N_9260,N_8920,N_8863);
or U9261 (N_9261,N_8715,N_8894);
xor U9262 (N_9262,N_8803,N_8805);
and U9263 (N_9263,N_8803,N_8863);
and U9264 (N_9264,N_8741,N_8707);
nor U9265 (N_9265,N_8750,N_8720);
and U9266 (N_9266,N_8732,N_8982);
nor U9267 (N_9267,N_8877,N_8880);
xnor U9268 (N_9268,N_8833,N_8797);
xor U9269 (N_9269,N_8712,N_8898);
or U9270 (N_9270,N_8872,N_8969);
nor U9271 (N_9271,N_8819,N_8945);
nor U9272 (N_9272,N_8704,N_8920);
xnor U9273 (N_9273,N_8738,N_8833);
nor U9274 (N_9274,N_8960,N_8807);
nor U9275 (N_9275,N_8740,N_8841);
nor U9276 (N_9276,N_8826,N_8725);
and U9277 (N_9277,N_8750,N_8942);
nor U9278 (N_9278,N_8723,N_8936);
xnor U9279 (N_9279,N_8803,N_8787);
nand U9280 (N_9280,N_8818,N_8835);
xnor U9281 (N_9281,N_8859,N_8985);
and U9282 (N_9282,N_8742,N_8766);
xor U9283 (N_9283,N_8922,N_8979);
xnor U9284 (N_9284,N_8949,N_8800);
and U9285 (N_9285,N_8828,N_8753);
and U9286 (N_9286,N_8735,N_8839);
xor U9287 (N_9287,N_8707,N_8829);
xnor U9288 (N_9288,N_8790,N_8815);
or U9289 (N_9289,N_8987,N_8927);
nor U9290 (N_9290,N_8703,N_8935);
nand U9291 (N_9291,N_8864,N_8968);
and U9292 (N_9292,N_8732,N_8787);
nand U9293 (N_9293,N_8938,N_8990);
or U9294 (N_9294,N_8785,N_8711);
xor U9295 (N_9295,N_8868,N_8864);
and U9296 (N_9296,N_8870,N_8789);
nand U9297 (N_9297,N_8987,N_8986);
xor U9298 (N_9298,N_8860,N_8917);
or U9299 (N_9299,N_8721,N_8767);
nor U9300 (N_9300,N_9013,N_9214);
nor U9301 (N_9301,N_9097,N_9117);
nand U9302 (N_9302,N_9271,N_9202);
xor U9303 (N_9303,N_9121,N_9055);
and U9304 (N_9304,N_9032,N_9099);
xnor U9305 (N_9305,N_9212,N_9056);
xor U9306 (N_9306,N_9018,N_9232);
nand U9307 (N_9307,N_9141,N_9112);
nand U9308 (N_9308,N_9186,N_9125);
and U9309 (N_9309,N_9225,N_9113);
nor U9310 (N_9310,N_9154,N_9098);
nand U9311 (N_9311,N_9175,N_9131);
xor U9312 (N_9312,N_9031,N_9253);
nor U9313 (N_9313,N_9206,N_9181);
and U9314 (N_9314,N_9240,N_9058);
nor U9315 (N_9315,N_9241,N_9020);
xnor U9316 (N_9316,N_9027,N_9156);
nand U9317 (N_9317,N_9219,N_9015);
nor U9318 (N_9318,N_9163,N_9143);
and U9319 (N_9319,N_9092,N_9268);
xnor U9320 (N_9320,N_9235,N_9289);
nor U9321 (N_9321,N_9093,N_9286);
xnor U9322 (N_9322,N_9223,N_9216);
nand U9323 (N_9323,N_9201,N_9274);
xor U9324 (N_9324,N_9010,N_9057);
or U9325 (N_9325,N_9108,N_9078);
or U9326 (N_9326,N_9278,N_9101);
nor U9327 (N_9327,N_9244,N_9280);
or U9328 (N_9328,N_9066,N_9245);
nand U9329 (N_9329,N_9034,N_9155);
nor U9330 (N_9330,N_9046,N_9148);
or U9331 (N_9331,N_9257,N_9177);
or U9332 (N_9332,N_9072,N_9256);
xor U9333 (N_9333,N_9009,N_9000);
nor U9334 (N_9334,N_9264,N_9248);
nand U9335 (N_9335,N_9224,N_9254);
and U9336 (N_9336,N_9048,N_9153);
or U9337 (N_9337,N_9085,N_9115);
nor U9338 (N_9338,N_9127,N_9218);
xor U9339 (N_9339,N_9063,N_9067);
or U9340 (N_9340,N_9238,N_9060);
or U9341 (N_9341,N_9139,N_9227);
xnor U9342 (N_9342,N_9123,N_9190);
and U9343 (N_9343,N_9135,N_9045);
and U9344 (N_9344,N_9069,N_9091);
nand U9345 (N_9345,N_9221,N_9088);
nor U9346 (N_9346,N_9061,N_9267);
nor U9347 (N_9347,N_9052,N_9180);
xnor U9348 (N_9348,N_9166,N_9124);
nor U9349 (N_9349,N_9172,N_9295);
xnor U9350 (N_9350,N_9059,N_9262);
xor U9351 (N_9351,N_9208,N_9263);
and U9352 (N_9352,N_9205,N_9176);
and U9353 (N_9353,N_9026,N_9287);
nand U9354 (N_9354,N_9265,N_9251);
nor U9355 (N_9355,N_9179,N_9193);
and U9356 (N_9356,N_9173,N_9076);
nor U9357 (N_9357,N_9041,N_9182);
xnor U9358 (N_9358,N_9142,N_9003);
nand U9359 (N_9359,N_9270,N_9298);
nor U9360 (N_9360,N_9087,N_9035);
nor U9361 (N_9361,N_9294,N_9169);
nor U9362 (N_9362,N_9284,N_9033);
nor U9363 (N_9363,N_9100,N_9090);
xor U9364 (N_9364,N_9114,N_9037);
nand U9365 (N_9365,N_9165,N_9188);
or U9366 (N_9366,N_9203,N_9189);
xnor U9367 (N_9367,N_9200,N_9158);
nand U9368 (N_9368,N_9239,N_9122);
or U9369 (N_9369,N_9102,N_9126);
or U9370 (N_9370,N_9044,N_9084);
nand U9371 (N_9371,N_9081,N_9011);
nor U9372 (N_9372,N_9006,N_9001);
xor U9373 (N_9373,N_9028,N_9259);
or U9374 (N_9374,N_9290,N_9247);
nor U9375 (N_9375,N_9082,N_9174);
nand U9376 (N_9376,N_9283,N_9120);
xnor U9377 (N_9377,N_9103,N_9104);
nand U9378 (N_9378,N_9002,N_9183);
xor U9379 (N_9379,N_9252,N_9133);
xnor U9380 (N_9380,N_9222,N_9211);
nand U9381 (N_9381,N_9288,N_9297);
and U9382 (N_9382,N_9054,N_9255);
nand U9383 (N_9383,N_9207,N_9276);
nor U9384 (N_9384,N_9261,N_9043);
nor U9385 (N_9385,N_9049,N_9147);
xor U9386 (N_9386,N_9249,N_9149);
and U9387 (N_9387,N_9016,N_9168);
xnor U9388 (N_9388,N_9215,N_9146);
nor U9389 (N_9389,N_9277,N_9137);
xor U9390 (N_9390,N_9150,N_9164);
nor U9391 (N_9391,N_9075,N_9167);
nand U9392 (N_9392,N_9089,N_9136);
and U9393 (N_9393,N_9110,N_9030);
nor U9394 (N_9394,N_9138,N_9079);
nand U9395 (N_9395,N_9275,N_9230);
nor U9396 (N_9396,N_9272,N_9210);
nor U9397 (N_9397,N_9038,N_9039);
or U9398 (N_9398,N_9152,N_9184);
nor U9399 (N_9399,N_9291,N_9233);
nor U9400 (N_9400,N_9296,N_9226);
and U9401 (N_9401,N_9070,N_9129);
nand U9402 (N_9402,N_9246,N_9106);
xnor U9403 (N_9403,N_9229,N_9051);
and U9404 (N_9404,N_9021,N_9132);
or U9405 (N_9405,N_9014,N_9134);
and U9406 (N_9406,N_9064,N_9118);
xor U9407 (N_9407,N_9105,N_9077);
or U9408 (N_9408,N_9116,N_9192);
and U9409 (N_9409,N_9074,N_9022);
or U9410 (N_9410,N_9217,N_9005);
nand U9411 (N_9411,N_9086,N_9040);
xnor U9412 (N_9412,N_9273,N_9231);
xor U9413 (N_9413,N_9008,N_9053);
nor U9414 (N_9414,N_9292,N_9236);
nor U9415 (N_9415,N_9228,N_9029);
nor U9416 (N_9416,N_9242,N_9160);
and U9417 (N_9417,N_9145,N_9017);
xnor U9418 (N_9418,N_9197,N_9237);
or U9419 (N_9419,N_9243,N_9194);
and U9420 (N_9420,N_9128,N_9250);
and U9421 (N_9421,N_9073,N_9065);
or U9422 (N_9422,N_9130,N_9285);
nand U9423 (N_9423,N_9107,N_9161);
nand U9424 (N_9424,N_9119,N_9050);
and U9425 (N_9425,N_9209,N_9220);
or U9426 (N_9426,N_9004,N_9109);
nor U9427 (N_9427,N_9213,N_9080);
or U9428 (N_9428,N_9171,N_9071);
xor U9429 (N_9429,N_9094,N_9269);
and U9430 (N_9430,N_9162,N_9042);
or U9431 (N_9431,N_9234,N_9204);
nand U9432 (N_9432,N_9293,N_9258);
or U9433 (N_9433,N_9151,N_9199);
nand U9434 (N_9434,N_9279,N_9170);
or U9435 (N_9435,N_9260,N_9195);
or U9436 (N_9436,N_9178,N_9024);
and U9437 (N_9437,N_9023,N_9159);
nand U9438 (N_9438,N_9266,N_9012);
or U9439 (N_9439,N_9007,N_9281);
nor U9440 (N_9440,N_9036,N_9019);
and U9441 (N_9441,N_9140,N_9282);
or U9442 (N_9442,N_9187,N_9191);
xor U9443 (N_9443,N_9144,N_9196);
xnor U9444 (N_9444,N_9095,N_9198);
nor U9445 (N_9445,N_9111,N_9047);
nor U9446 (N_9446,N_9299,N_9096);
or U9447 (N_9447,N_9062,N_9157);
xnor U9448 (N_9448,N_9083,N_9185);
and U9449 (N_9449,N_9025,N_9068);
nor U9450 (N_9450,N_9131,N_9098);
xnor U9451 (N_9451,N_9161,N_9167);
xor U9452 (N_9452,N_9084,N_9275);
xnor U9453 (N_9453,N_9108,N_9012);
or U9454 (N_9454,N_9045,N_9035);
and U9455 (N_9455,N_9157,N_9261);
xor U9456 (N_9456,N_9231,N_9216);
xnor U9457 (N_9457,N_9293,N_9055);
and U9458 (N_9458,N_9051,N_9211);
nor U9459 (N_9459,N_9128,N_9151);
and U9460 (N_9460,N_9011,N_9129);
xor U9461 (N_9461,N_9021,N_9017);
and U9462 (N_9462,N_9121,N_9144);
nand U9463 (N_9463,N_9288,N_9224);
nand U9464 (N_9464,N_9094,N_9081);
or U9465 (N_9465,N_9219,N_9051);
and U9466 (N_9466,N_9077,N_9089);
xnor U9467 (N_9467,N_9112,N_9144);
nand U9468 (N_9468,N_9078,N_9115);
or U9469 (N_9469,N_9252,N_9059);
or U9470 (N_9470,N_9253,N_9057);
or U9471 (N_9471,N_9269,N_9174);
and U9472 (N_9472,N_9232,N_9148);
xnor U9473 (N_9473,N_9109,N_9050);
xor U9474 (N_9474,N_9160,N_9054);
and U9475 (N_9475,N_9132,N_9086);
nand U9476 (N_9476,N_9277,N_9211);
and U9477 (N_9477,N_9028,N_9142);
or U9478 (N_9478,N_9216,N_9054);
nand U9479 (N_9479,N_9116,N_9130);
and U9480 (N_9480,N_9016,N_9029);
nor U9481 (N_9481,N_9219,N_9198);
and U9482 (N_9482,N_9248,N_9077);
and U9483 (N_9483,N_9241,N_9080);
nor U9484 (N_9484,N_9220,N_9286);
or U9485 (N_9485,N_9278,N_9138);
and U9486 (N_9486,N_9296,N_9215);
nor U9487 (N_9487,N_9239,N_9132);
nand U9488 (N_9488,N_9047,N_9125);
xor U9489 (N_9489,N_9103,N_9258);
xor U9490 (N_9490,N_9031,N_9287);
or U9491 (N_9491,N_9238,N_9117);
nor U9492 (N_9492,N_9056,N_9220);
or U9493 (N_9493,N_9211,N_9098);
nor U9494 (N_9494,N_9235,N_9010);
nor U9495 (N_9495,N_9296,N_9000);
or U9496 (N_9496,N_9284,N_9270);
and U9497 (N_9497,N_9246,N_9092);
or U9498 (N_9498,N_9080,N_9255);
nand U9499 (N_9499,N_9141,N_9168);
xnor U9500 (N_9500,N_9188,N_9229);
xnor U9501 (N_9501,N_9261,N_9053);
xor U9502 (N_9502,N_9113,N_9010);
nand U9503 (N_9503,N_9144,N_9087);
nor U9504 (N_9504,N_9276,N_9280);
and U9505 (N_9505,N_9151,N_9109);
or U9506 (N_9506,N_9188,N_9169);
xnor U9507 (N_9507,N_9245,N_9140);
nand U9508 (N_9508,N_9135,N_9261);
nand U9509 (N_9509,N_9212,N_9197);
nand U9510 (N_9510,N_9085,N_9202);
or U9511 (N_9511,N_9003,N_9290);
nand U9512 (N_9512,N_9079,N_9001);
or U9513 (N_9513,N_9262,N_9129);
nor U9514 (N_9514,N_9033,N_9296);
nor U9515 (N_9515,N_9127,N_9080);
and U9516 (N_9516,N_9225,N_9294);
nor U9517 (N_9517,N_9213,N_9116);
or U9518 (N_9518,N_9164,N_9178);
nor U9519 (N_9519,N_9181,N_9083);
nand U9520 (N_9520,N_9199,N_9259);
xnor U9521 (N_9521,N_9155,N_9289);
xor U9522 (N_9522,N_9089,N_9076);
or U9523 (N_9523,N_9113,N_9297);
xor U9524 (N_9524,N_9138,N_9099);
or U9525 (N_9525,N_9082,N_9183);
or U9526 (N_9526,N_9049,N_9001);
or U9527 (N_9527,N_9027,N_9218);
xor U9528 (N_9528,N_9103,N_9013);
nand U9529 (N_9529,N_9246,N_9008);
xor U9530 (N_9530,N_9001,N_9120);
nand U9531 (N_9531,N_9159,N_9059);
nand U9532 (N_9532,N_9043,N_9297);
xor U9533 (N_9533,N_9152,N_9067);
xor U9534 (N_9534,N_9087,N_9231);
or U9535 (N_9535,N_9284,N_9101);
nor U9536 (N_9536,N_9048,N_9113);
xor U9537 (N_9537,N_9183,N_9167);
or U9538 (N_9538,N_9253,N_9206);
xnor U9539 (N_9539,N_9257,N_9157);
nor U9540 (N_9540,N_9231,N_9100);
nand U9541 (N_9541,N_9010,N_9206);
or U9542 (N_9542,N_9052,N_9024);
xor U9543 (N_9543,N_9201,N_9212);
nor U9544 (N_9544,N_9215,N_9195);
or U9545 (N_9545,N_9000,N_9049);
nand U9546 (N_9546,N_9051,N_9279);
and U9547 (N_9547,N_9217,N_9240);
xnor U9548 (N_9548,N_9060,N_9192);
nor U9549 (N_9549,N_9275,N_9047);
or U9550 (N_9550,N_9056,N_9007);
and U9551 (N_9551,N_9162,N_9168);
and U9552 (N_9552,N_9100,N_9217);
or U9553 (N_9553,N_9179,N_9108);
nor U9554 (N_9554,N_9229,N_9293);
xnor U9555 (N_9555,N_9270,N_9132);
nor U9556 (N_9556,N_9099,N_9013);
xor U9557 (N_9557,N_9128,N_9256);
xnor U9558 (N_9558,N_9042,N_9256);
and U9559 (N_9559,N_9140,N_9049);
nor U9560 (N_9560,N_9104,N_9016);
or U9561 (N_9561,N_9242,N_9273);
and U9562 (N_9562,N_9266,N_9272);
or U9563 (N_9563,N_9164,N_9279);
and U9564 (N_9564,N_9127,N_9230);
nand U9565 (N_9565,N_9202,N_9049);
xnor U9566 (N_9566,N_9244,N_9126);
nor U9567 (N_9567,N_9298,N_9049);
nor U9568 (N_9568,N_9168,N_9194);
nor U9569 (N_9569,N_9079,N_9060);
and U9570 (N_9570,N_9291,N_9234);
nor U9571 (N_9571,N_9200,N_9260);
xnor U9572 (N_9572,N_9159,N_9189);
or U9573 (N_9573,N_9007,N_9009);
xnor U9574 (N_9574,N_9210,N_9023);
nor U9575 (N_9575,N_9237,N_9144);
and U9576 (N_9576,N_9124,N_9223);
nand U9577 (N_9577,N_9173,N_9145);
nand U9578 (N_9578,N_9186,N_9188);
xor U9579 (N_9579,N_9098,N_9195);
nand U9580 (N_9580,N_9267,N_9256);
and U9581 (N_9581,N_9030,N_9215);
or U9582 (N_9582,N_9152,N_9107);
nand U9583 (N_9583,N_9250,N_9294);
nor U9584 (N_9584,N_9133,N_9224);
nor U9585 (N_9585,N_9202,N_9025);
and U9586 (N_9586,N_9133,N_9169);
xor U9587 (N_9587,N_9127,N_9158);
or U9588 (N_9588,N_9253,N_9230);
or U9589 (N_9589,N_9269,N_9228);
nor U9590 (N_9590,N_9196,N_9238);
nand U9591 (N_9591,N_9179,N_9258);
nor U9592 (N_9592,N_9093,N_9282);
xor U9593 (N_9593,N_9048,N_9241);
and U9594 (N_9594,N_9213,N_9249);
or U9595 (N_9595,N_9200,N_9192);
xnor U9596 (N_9596,N_9019,N_9051);
nand U9597 (N_9597,N_9284,N_9107);
or U9598 (N_9598,N_9067,N_9074);
or U9599 (N_9599,N_9230,N_9248);
nand U9600 (N_9600,N_9491,N_9534);
or U9601 (N_9601,N_9500,N_9504);
nand U9602 (N_9602,N_9484,N_9468);
xor U9603 (N_9603,N_9446,N_9532);
xor U9604 (N_9604,N_9336,N_9367);
nor U9605 (N_9605,N_9330,N_9577);
nand U9606 (N_9606,N_9392,N_9308);
xnor U9607 (N_9607,N_9584,N_9545);
nor U9608 (N_9608,N_9320,N_9544);
nor U9609 (N_9609,N_9561,N_9307);
or U9610 (N_9610,N_9485,N_9474);
xnor U9611 (N_9611,N_9448,N_9475);
nand U9612 (N_9612,N_9497,N_9573);
and U9613 (N_9613,N_9439,N_9355);
xor U9614 (N_9614,N_9562,N_9456);
nand U9615 (N_9615,N_9376,N_9323);
or U9616 (N_9616,N_9520,N_9536);
or U9617 (N_9617,N_9481,N_9319);
nor U9618 (N_9618,N_9597,N_9315);
or U9619 (N_9619,N_9337,N_9524);
xor U9620 (N_9620,N_9507,N_9440);
xnor U9621 (N_9621,N_9342,N_9457);
xor U9622 (N_9622,N_9382,N_9362);
xor U9623 (N_9623,N_9385,N_9451);
xor U9624 (N_9624,N_9384,N_9419);
or U9625 (N_9625,N_9450,N_9310);
xor U9626 (N_9626,N_9370,N_9329);
and U9627 (N_9627,N_9334,N_9430);
and U9628 (N_9628,N_9361,N_9306);
or U9629 (N_9629,N_9333,N_9574);
or U9630 (N_9630,N_9452,N_9543);
or U9631 (N_9631,N_9348,N_9447);
and U9632 (N_9632,N_9332,N_9346);
nor U9633 (N_9633,N_9441,N_9453);
and U9634 (N_9634,N_9403,N_9565);
nor U9635 (N_9635,N_9381,N_9483);
and U9636 (N_9636,N_9445,N_9391);
nor U9637 (N_9637,N_9321,N_9486);
and U9638 (N_9638,N_9414,N_9581);
nor U9639 (N_9639,N_9404,N_9428);
nand U9640 (N_9640,N_9371,N_9575);
and U9641 (N_9641,N_9579,N_9592);
or U9642 (N_9642,N_9469,N_9402);
and U9643 (N_9643,N_9425,N_9488);
and U9644 (N_9644,N_9585,N_9501);
and U9645 (N_9645,N_9454,N_9596);
or U9646 (N_9646,N_9422,N_9525);
nand U9647 (N_9647,N_9519,N_9487);
xor U9648 (N_9648,N_9398,N_9318);
nor U9649 (N_9649,N_9350,N_9528);
and U9650 (N_9650,N_9435,N_9311);
nand U9651 (N_9651,N_9570,N_9477);
and U9652 (N_9652,N_9563,N_9427);
and U9653 (N_9653,N_9364,N_9541);
nand U9654 (N_9654,N_9369,N_9399);
xnor U9655 (N_9655,N_9314,N_9359);
nor U9656 (N_9656,N_9464,N_9499);
nor U9657 (N_9657,N_9530,N_9328);
nor U9658 (N_9658,N_9401,N_9415);
or U9659 (N_9659,N_9313,N_9358);
xnor U9660 (N_9660,N_9508,N_9305);
xor U9661 (N_9661,N_9316,N_9303);
nand U9662 (N_9662,N_9365,N_9537);
nand U9663 (N_9663,N_9503,N_9394);
xnor U9664 (N_9664,N_9416,N_9523);
or U9665 (N_9665,N_9400,N_9552);
or U9666 (N_9666,N_9521,N_9312);
xnor U9667 (N_9667,N_9331,N_9409);
or U9668 (N_9668,N_9423,N_9309);
nand U9669 (N_9669,N_9588,N_9568);
nor U9670 (N_9670,N_9433,N_9405);
nand U9671 (N_9671,N_9513,N_9458);
and U9672 (N_9672,N_9438,N_9397);
xor U9673 (N_9673,N_9571,N_9304);
or U9674 (N_9674,N_9515,N_9495);
xor U9675 (N_9675,N_9449,N_9300);
and U9676 (N_9676,N_9412,N_9480);
nor U9677 (N_9677,N_9366,N_9436);
and U9678 (N_9678,N_9388,N_9529);
nand U9679 (N_9679,N_9443,N_9374);
nor U9680 (N_9680,N_9408,N_9482);
and U9681 (N_9681,N_9465,N_9599);
nand U9682 (N_9682,N_9302,N_9420);
nor U9683 (N_9683,N_9442,N_9535);
and U9684 (N_9684,N_9533,N_9527);
or U9685 (N_9685,N_9353,N_9595);
or U9686 (N_9686,N_9411,N_9470);
and U9687 (N_9687,N_9569,N_9572);
and U9688 (N_9688,N_9496,N_9531);
xor U9689 (N_9689,N_9548,N_9386);
xnor U9690 (N_9690,N_9357,N_9340);
nor U9691 (N_9691,N_9378,N_9550);
nand U9692 (N_9692,N_9512,N_9406);
xnor U9693 (N_9693,N_9338,N_9559);
and U9694 (N_9694,N_9476,N_9356);
or U9695 (N_9695,N_9522,N_9461);
nand U9696 (N_9696,N_9557,N_9418);
xnor U9697 (N_9697,N_9322,N_9553);
xor U9698 (N_9698,N_9466,N_9349);
nand U9699 (N_9699,N_9551,N_9554);
xnor U9700 (N_9700,N_9372,N_9327);
xnor U9701 (N_9701,N_9510,N_9383);
nand U9702 (N_9702,N_9493,N_9434);
and U9703 (N_9703,N_9343,N_9344);
and U9704 (N_9704,N_9437,N_9432);
nor U9705 (N_9705,N_9410,N_9345);
nand U9706 (N_9706,N_9377,N_9455);
nand U9707 (N_9707,N_9444,N_9594);
and U9708 (N_9708,N_9335,N_9556);
or U9709 (N_9709,N_9549,N_9472);
xor U9710 (N_9710,N_9429,N_9478);
nor U9711 (N_9711,N_9462,N_9375);
and U9712 (N_9712,N_9360,N_9301);
or U9713 (N_9713,N_9593,N_9317);
and U9714 (N_9714,N_9326,N_9560);
and U9715 (N_9715,N_9517,N_9490);
and U9716 (N_9716,N_9598,N_9539);
or U9717 (N_9717,N_9538,N_9516);
xor U9718 (N_9718,N_9542,N_9583);
nor U9719 (N_9719,N_9586,N_9591);
and U9720 (N_9720,N_9354,N_9511);
or U9721 (N_9721,N_9479,N_9502);
and U9722 (N_9722,N_9540,N_9471);
nor U9723 (N_9723,N_9380,N_9580);
xor U9724 (N_9724,N_9341,N_9339);
and U9725 (N_9725,N_9363,N_9387);
xor U9726 (N_9726,N_9546,N_9492);
xnor U9727 (N_9727,N_9558,N_9379);
xnor U9728 (N_9728,N_9396,N_9351);
or U9729 (N_9729,N_9373,N_9390);
nor U9730 (N_9730,N_9324,N_9567);
xor U9731 (N_9731,N_9413,N_9566);
or U9732 (N_9732,N_9494,N_9325);
nand U9733 (N_9733,N_9489,N_9463);
xnor U9734 (N_9734,N_9578,N_9587);
xor U9735 (N_9735,N_9590,N_9589);
nand U9736 (N_9736,N_9426,N_9582);
or U9737 (N_9737,N_9459,N_9389);
xor U9738 (N_9738,N_9514,N_9460);
nor U9739 (N_9739,N_9473,N_9506);
or U9740 (N_9740,N_9505,N_9395);
xnor U9741 (N_9741,N_9368,N_9347);
nand U9742 (N_9742,N_9526,N_9509);
nand U9743 (N_9743,N_9352,N_9393);
xnor U9744 (N_9744,N_9421,N_9547);
or U9745 (N_9745,N_9498,N_9467);
or U9746 (N_9746,N_9518,N_9431);
and U9747 (N_9747,N_9407,N_9576);
and U9748 (N_9748,N_9417,N_9555);
and U9749 (N_9749,N_9424,N_9564);
nand U9750 (N_9750,N_9513,N_9492);
nor U9751 (N_9751,N_9355,N_9528);
nor U9752 (N_9752,N_9493,N_9545);
or U9753 (N_9753,N_9426,N_9495);
xor U9754 (N_9754,N_9362,N_9548);
or U9755 (N_9755,N_9392,N_9418);
nand U9756 (N_9756,N_9309,N_9389);
or U9757 (N_9757,N_9401,N_9339);
nand U9758 (N_9758,N_9395,N_9312);
nor U9759 (N_9759,N_9518,N_9426);
nor U9760 (N_9760,N_9562,N_9498);
xor U9761 (N_9761,N_9304,N_9488);
nor U9762 (N_9762,N_9520,N_9387);
nand U9763 (N_9763,N_9525,N_9479);
nand U9764 (N_9764,N_9551,N_9452);
nand U9765 (N_9765,N_9448,N_9325);
nor U9766 (N_9766,N_9470,N_9351);
xnor U9767 (N_9767,N_9595,N_9313);
and U9768 (N_9768,N_9475,N_9512);
xor U9769 (N_9769,N_9589,N_9492);
xor U9770 (N_9770,N_9415,N_9378);
or U9771 (N_9771,N_9551,N_9581);
and U9772 (N_9772,N_9448,N_9408);
nand U9773 (N_9773,N_9445,N_9519);
or U9774 (N_9774,N_9300,N_9346);
nand U9775 (N_9775,N_9344,N_9441);
nand U9776 (N_9776,N_9583,N_9444);
or U9777 (N_9777,N_9580,N_9348);
xnor U9778 (N_9778,N_9519,N_9518);
xor U9779 (N_9779,N_9328,N_9407);
xnor U9780 (N_9780,N_9329,N_9558);
and U9781 (N_9781,N_9593,N_9407);
or U9782 (N_9782,N_9561,N_9376);
nand U9783 (N_9783,N_9542,N_9310);
nor U9784 (N_9784,N_9417,N_9418);
and U9785 (N_9785,N_9575,N_9541);
and U9786 (N_9786,N_9347,N_9556);
and U9787 (N_9787,N_9558,N_9556);
or U9788 (N_9788,N_9464,N_9559);
or U9789 (N_9789,N_9412,N_9492);
or U9790 (N_9790,N_9520,N_9395);
xnor U9791 (N_9791,N_9535,N_9550);
and U9792 (N_9792,N_9422,N_9453);
xnor U9793 (N_9793,N_9358,N_9329);
xor U9794 (N_9794,N_9529,N_9568);
nor U9795 (N_9795,N_9528,N_9365);
or U9796 (N_9796,N_9315,N_9320);
nor U9797 (N_9797,N_9519,N_9324);
and U9798 (N_9798,N_9418,N_9519);
nor U9799 (N_9799,N_9519,N_9452);
and U9800 (N_9800,N_9550,N_9329);
and U9801 (N_9801,N_9582,N_9438);
and U9802 (N_9802,N_9367,N_9322);
and U9803 (N_9803,N_9478,N_9469);
nor U9804 (N_9804,N_9330,N_9509);
nand U9805 (N_9805,N_9394,N_9575);
nand U9806 (N_9806,N_9374,N_9307);
nand U9807 (N_9807,N_9535,N_9415);
xnor U9808 (N_9808,N_9363,N_9320);
nor U9809 (N_9809,N_9382,N_9566);
or U9810 (N_9810,N_9347,N_9400);
and U9811 (N_9811,N_9547,N_9484);
xnor U9812 (N_9812,N_9434,N_9398);
nand U9813 (N_9813,N_9344,N_9307);
xnor U9814 (N_9814,N_9395,N_9435);
and U9815 (N_9815,N_9367,N_9469);
and U9816 (N_9816,N_9557,N_9539);
nor U9817 (N_9817,N_9449,N_9527);
or U9818 (N_9818,N_9587,N_9540);
nand U9819 (N_9819,N_9576,N_9593);
xor U9820 (N_9820,N_9575,N_9500);
or U9821 (N_9821,N_9446,N_9566);
xnor U9822 (N_9822,N_9460,N_9315);
nor U9823 (N_9823,N_9440,N_9333);
xor U9824 (N_9824,N_9385,N_9346);
and U9825 (N_9825,N_9512,N_9449);
xor U9826 (N_9826,N_9375,N_9511);
xnor U9827 (N_9827,N_9500,N_9356);
nand U9828 (N_9828,N_9375,N_9556);
or U9829 (N_9829,N_9407,N_9398);
nor U9830 (N_9830,N_9582,N_9316);
or U9831 (N_9831,N_9449,N_9434);
and U9832 (N_9832,N_9334,N_9568);
nor U9833 (N_9833,N_9485,N_9411);
nand U9834 (N_9834,N_9352,N_9305);
and U9835 (N_9835,N_9529,N_9439);
nor U9836 (N_9836,N_9490,N_9458);
xor U9837 (N_9837,N_9532,N_9380);
nor U9838 (N_9838,N_9410,N_9443);
or U9839 (N_9839,N_9584,N_9445);
and U9840 (N_9840,N_9440,N_9364);
nand U9841 (N_9841,N_9373,N_9509);
nor U9842 (N_9842,N_9491,N_9514);
and U9843 (N_9843,N_9510,N_9450);
and U9844 (N_9844,N_9438,N_9300);
or U9845 (N_9845,N_9418,N_9342);
nand U9846 (N_9846,N_9451,N_9338);
and U9847 (N_9847,N_9337,N_9466);
nor U9848 (N_9848,N_9311,N_9559);
nand U9849 (N_9849,N_9326,N_9423);
and U9850 (N_9850,N_9414,N_9395);
nor U9851 (N_9851,N_9531,N_9560);
xnor U9852 (N_9852,N_9520,N_9360);
and U9853 (N_9853,N_9382,N_9329);
and U9854 (N_9854,N_9527,N_9325);
nand U9855 (N_9855,N_9420,N_9447);
nor U9856 (N_9856,N_9490,N_9320);
or U9857 (N_9857,N_9482,N_9322);
nand U9858 (N_9858,N_9420,N_9464);
xor U9859 (N_9859,N_9506,N_9407);
nor U9860 (N_9860,N_9487,N_9329);
xor U9861 (N_9861,N_9381,N_9523);
nand U9862 (N_9862,N_9337,N_9527);
xor U9863 (N_9863,N_9540,N_9365);
xor U9864 (N_9864,N_9356,N_9386);
and U9865 (N_9865,N_9533,N_9430);
nor U9866 (N_9866,N_9518,N_9333);
nor U9867 (N_9867,N_9378,N_9438);
or U9868 (N_9868,N_9379,N_9499);
and U9869 (N_9869,N_9395,N_9574);
xor U9870 (N_9870,N_9526,N_9534);
nor U9871 (N_9871,N_9496,N_9473);
nand U9872 (N_9872,N_9586,N_9462);
nor U9873 (N_9873,N_9420,N_9303);
or U9874 (N_9874,N_9560,N_9517);
nor U9875 (N_9875,N_9513,N_9436);
or U9876 (N_9876,N_9405,N_9459);
xor U9877 (N_9877,N_9442,N_9443);
or U9878 (N_9878,N_9357,N_9477);
and U9879 (N_9879,N_9597,N_9499);
nor U9880 (N_9880,N_9384,N_9564);
nand U9881 (N_9881,N_9503,N_9465);
nand U9882 (N_9882,N_9543,N_9369);
and U9883 (N_9883,N_9353,N_9374);
or U9884 (N_9884,N_9433,N_9482);
or U9885 (N_9885,N_9362,N_9546);
nor U9886 (N_9886,N_9516,N_9498);
nand U9887 (N_9887,N_9314,N_9516);
and U9888 (N_9888,N_9475,N_9311);
or U9889 (N_9889,N_9525,N_9402);
or U9890 (N_9890,N_9468,N_9378);
and U9891 (N_9891,N_9525,N_9384);
xor U9892 (N_9892,N_9590,N_9454);
and U9893 (N_9893,N_9590,N_9535);
or U9894 (N_9894,N_9483,N_9421);
and U9895 (N_9895,N_9302,N_9536);
or U9896 (N_9896,N_9301,N_9466);
or U9897 (N_9897,N_9367,N_9464);
xor U9898 (N_9898,N_9367,N_9470);
or U9899 (N_9899,N_9468,N_9469);
xor U9900 (N_9900,N_9858,N_9642);
nand U9901 (N_9901,N_9802,N_9765);
xor U9902 (N_9902,N_9748,N_9777);
or U9903 (N_9903,N_9878,N_9884);
nand U9904 (N_9904,N_9856,N_9654);
nor U9905 (N_9905,N_9874,N_9789);
nor U9906 (N_9906,N_9625,N_9804);
or U9907 (N_9907,N_9863,N_9619);
and U9908 (N_9908,N_9681,N_9702);
nor U9909 (N_9909,N_9883,N_9656);
nor U9910 (N_9910,N_9790,N_9690);
nor U9911 (N_9911,N_9658,N_9800);
xor U9912 (N_9912,N_9742,N_9627);
or U9913 (N_9913,N_9771,N_9859);
and U9914 (N_9914,N_9749,N_9734);
nand U9915 (N_9915,N_9674,N_9780);
nor U9916 (N_9916,N_9728,N_9626);
nor U9917 (N_9917,N_9847,N_9823);
or U9918 (N_9918,N_9840,N_9822);
and U9919 (N_9919,N_9620,N_9692);
xor U9920 (N_9920,N_9752,N_9875);
or U9921 (N_9921,N_9796,N_9854);
nand U9922 (N_9922,N_9757,N_9631);
and U9923 (N_9923,N_9716,N_9662);
xnor U9924 (N_9924,N_9704,N_9645);
and U9925 (N_9925,N_9705,N_9851);
nand U9926 (N_9926,N_9613,N_9809);
or U9927 (N_9927,N_9652,N_9871);
nor U9928 (N_9928,N_9678,N_9798);
nand U9929 (N_9929,N_9653,N_9684);
or U9930 (N_9930,N_9829,N_9755);
nor U9931 (N_9931,N_9865,N_9675);
nor U9932 (N_9932,N_9892,N_9853);
and U9933 (N_9933,N_9710,N_9621);
nand U9934 (N_9934,N_9737,N_9778);
or U9935 (N_9935,N_9766,N_9870);
and U9936 (N_9936,N_9651,N_9609);
xnor U9937 (N_9937,N_9806,N_9751);
or U9938 (N_9938,N_9608,N_9744);
nand U9939 (N_9939,N_9836,N_9786);
nor U9940 (N_9940,N_9896,N_9719);
xnor U9941 (N_9941,N_9826,N_9723);
or U9942 (N_9942,N_9827,N_9876);
nand U9943 (N_9943,N_9696,N_9667);
or U9944 (N_9944,N_9830,N_9747);
nand U9945 (N_9945,N_9890,N_9741);
or U9946 (N_9946,N_9717,N_9797);
or U9947 (N_9947,N_9888,N_9808);
or U9948 (N_9948,N_9849,N_9756);
and U9949 (N_9949,N_9616,N_9779);
nand U9950 (N_9950,N_9724,N_9894);
xnor U9951 (N_9951,N_9699,N_9818);
nand U9952 (N_9952,N_9610,N_9671);
nand U9953 (N_9953,N_9623,N_9782);
xor U9954 (N_9954,N_9686,N_9636);
nand U9955 (N_9955,N_9688,N_9770);
xnor U9956 (N_9956,N_9739,N_9868);
and U9957 (N_9957,N_9731,N_9810);
or U9958 (N_9958,N_9655,N_9828);
nor U9959 (N_9959,N_9709,N_9793);
nand U9960 (N_9960,N_9657,N_9601);
xnor U9961 (N_9961,N_9821,N_9711);
xnor U9962 (N_9962,N_9861,N_9899);
and U9963 (N_9963,N_9791,N_9722);
and U9964 (N_9964,N_9857,N_9689);
or U9965 (N_9965,N_9834,N_9708);
xnor U9966 (N_9966,N_9841,N_9832);
xor U9967 (N_9967,N_9727,N_9641);
or U9968 (N_9968,N_9817,N_9781);
and U9969 (N_9969,N_9885,N_9666);
and U9970 (N_9970,N_9738,N_9605);
and U9971 (N_9971,N_9694,N_9735);
nor U9972 (N_9972,N_9783,N_9611);
xnor U9973 (N_9973,N_9635,N_9837);
or U9974 (N_9974,N_9669,N_9624);
and U9975 (N_9975,N_9839,N_9887);
xor U9976 (N_9976,N_9816,N_9762);
or U9977 (N_9977,N_9638,N_9649);
or U9978 (N_9978,N_9672,N_9615);
nand U9979 (N_9979,N_9824,N_9603);
nand U9980 (N_9980,N_9882,N_9763);
or U9981 (N_9981,N_9864,N_9693);
nor U9982 (N_9982,N_9866,N_9873);
nand U9983 (N_9983,N_9776,N_9803);
and U9984 (N_9984,N_9707,N_9761);
and U9985 (N_9985,N_9842,N_9644);
or U9986 (N_9986,N_9607,N_9880);
or U9987 (N_9987,N_9785,N_9895);
nor U9988 (N_9988,N_9814,N_9881);
nand U9989 (N_9989,N_9805,N_9740);
xnor U9990 (N_9990,N_9617,N_9665);
xnor U9991 (N_9991,N_9787,N_9637);
nand U9992 (N_9992,N_9732,N_9813);
nand U9993 (N_9993,N_9773,N_9713);
nor U9994 (N_9994,N_9768,N_9618);
nor U9995 (N_9995,N_9898,N_9893);
xnor U9996 (N_9996,N_9646,N_9753);
and U9997 (N_9997,N_9758,N_9784);
nor U9998 (N_9998,N_9820,N_9661);
nor U9999 (N_9999,N_9715,N_9845);
nor U10000 (N_10000,N_9676,N_9663);
nand U10001 (N_10001,N_9628,N_9691);
nand U10002 (N_10002,N_9819,N_9680);
nor U10003 (N_10003,N_9639,N_9759);
or U10004 (N_10004,N_9687,N_9677);
nor U10005 (N_10005,N_9685,N_9721);
xor U10006 (N_10006,N_9604,N_9659);
xor U10007 (N_10007,N_9774,N_9750);
nand U10008 (N_10008,N_9633,N_9729);
and U10009 (N_10009,N_9668,N_9640);
xnor U10010 (N_10010,N_9825,N_9643);
and U10011 (N_10011,N_9760,N_9862);
xnor U10012 (N_10012,N_9852,N_9647);
nor U10013 (N_10013,N_9835,N_9600);
and U10014 (N_10014,N_9889,N_9650);
nor U10015 (N_10015,N_9788,N_9673);
nand U10016 (N_10016,N_9701,N_9879);
or U10017 (N_10017,N_9794,N_9877);
nand U10018 (N_10018,N_9754,N_9695);
or U10019 (N_10019,N_9886,N_9670);
nor U10020 (N_10020,N_9869,N_9746);
and U10021 (N_10021,N_9714,N_9745);
xnor U10022 (N_10022,N_9855,N_9831);
nor U10023 (N_10023,N_9860,N_9614);
nor U10024 (N_10024,N_9718,N_9767);
nor U10025 (N_10025,N_9630,N_9772);
or U10026 (N_10026,N_9811,N_9850);
nand U10027 (N_10027,N_9602,N_9799);
or U10028 (N_10028,N_9632,N_9736);
or U10029 (N_10029,N_9634,N_9698);
and U10030 (N_10030,N_9730,N_9897);
nand U10031 (N_10031,N_9843,N_9612);
nor U10032 (N_10032,N_9706,N_9697);
or U10033 (N_10033,N_9648,N_9801);
nand U10034 (N_10034,N_9743,N_9712);
xor U10035 (N_10035,N_9838,N_9725);
or U10036 (N_10036,N_9812,N_9867);
nor U10037 (N_10037,N_9775,N_9815);
or U10038 (N_10038,N_9720,N_9733);
nor U10039 (N_10039,N_9764,N_9872);
and U10040 (N_10040,N_9629,N_9700);
nor U10041 (N_10041,N_9726,N_9703);
and U10042 (N_10042,N_9664,N_9679);
xor U10043 (N_10043,N_9846,N_9683);
nand U10044 (N_10044,N_9833,N_9769);
and U10045 (N_10045,N_9682,N_9606);
xor U10046 (N_10046,N_9807,N_9660);
nand U10047 (N_10047,N_9795,N_9792);
and U10048 (N_10048,N_9622,N_9844);
and U10049 (N_10049,N_9848,N_9891);
xor U10050 (N_10050,N_9754,N_9843);
nor U10051 (N_10051,N_9818,N_9793);
nand U10052 (N_10052,N_9854,N_9662);
and U10053 (N_10053,N_9625,N_9851);
xor U10054 (N_10054,N_9642,N_9663);
or U10055 (N_10055,N_9806,N_9870);
xor U10056 (N_10056,N_9809,N_9679);
nand U10057 (N_10057,N_9615,N_9714);
nand U10058 (N_10058,N_9860,N_9795);
or U10059 (N_10059,N_9653,N_9696);
nand U10060 (N_10060,N_9717,N_9894);
xor U10061 (N_10061,N_9708,N_9836);
or U10062 (N_10062,N_9859,N_9635);
and U10063 (N_10063,N_9720,N_9673);
and U10064 (N_10064,N_9801,N_9815);
and U10065 (N_10065,N_9823,N_9711);
and U10066 (N_10066,N_9666,N_9614);
and U10067 (N_10067,N_9858,N_9750);
nand U10068 (N_10068,N_9795,N_9644);
nand U10069 (N_10069,N_9712,N_9803);
and U10070 (N_10070,N_9719,N_9632);
or U10071 (N_10071,N_9773,N_9655);
and U10072 (N_10072,N_9751,N_9817);
or U10073 (N_10073,N_9616,N_9696);
xor U10074 (N_10074,N_9827,N_9801);
xor U10075 (N_10075,N_9714,N_9628);
xnor U10076 (N_10076,N_9873,N_9794);
or U10077 (N_10077,N_9640,N_9769);
and U10078 (N_10078,N_9709,N_9833);
xnor U10079 (N_10079,N_9685,N_9758);
xor U10080 (N_10080,N_9803,N_9625);
nand U10081 (N_10081,N_9705,N_9743);
or U10082 (N_10082,N_9762,N_9688);
nor U10083 (N_10083,N_9655,N_9726);
or U10084 (N_10084,N_9841,N_9764);
xnor U10085 (N_10085,N_9664,N_9844);
nor U10086 (N_10086,N_9847,N_9874);
and U10087 (N_10087,N_9728,N_9862);
or U10088 (N_10088,N_9822,N_9706);
nand U10089 (N_10089,N_9791,N_9829);
and U10090 (N_10090,N_9658,N_9836);
xor U10091 (N_10091,N_9846,N_9770);
nor U10092 (N_10092,N_9828,N_9759);
nand U10093 (N_10093,N_9605,N_9601);
nand U10094 (N_10094,N_9805,N_9703);
nor U10095 (N_10095,N_9741,N_9817);
xor U10096 (N_10096,N_9770,N_9786);
nand U10097 (N_10097,N_9898,N_9614);
or U10098 (N_10098,N_9805,N_9643);
or U10099 (N_10099,N_9614,N_9742);
xnor U10100 (N_10100,N_9666,N_9836);
xnor U10101 (N_10101,N_9671,N_9857);
or U10102 (N_10102,N_9704,N_9780);
and U10103 (N_10103,N_9875,N_9774);
nand U10104 (N_10104,N_9672,N_9726);
nand U10105 (N_10105,N_9898,N_9820);
xor U10106 (N_10106,N_9780,N_9658);
nand U10107 (N_10107,N_9798,N_9603);
nor U10108 (N_10108,N_9726,N_9646);
or U10109 (N_10109,N_9648,N_9690);
and U10110 (N_10110,N_9639,N_9805);
nor U10111 (N_10111,N_9749,N_9822);
xnor U10112 (N_10112,N_9731,N_9869);
xnor U10113 (N_10113,N_9728,N_9687);
nor U10114 (N_10114,N_9822,N_9630);
xnor U10115 (N_10115,N_9769,N_9728);
or U10116 (N_10116,N_9628,N_9649);
nand U10117 (N_10117,N_9854,N_9788);
nand U10118 (N_10118,N_9801,N_9694);
nand U10119 (N_10119,N_9684,N_9882);
and U10120 (N_10120,N_9602,N_9601);
nand U10121 (N_10121,N_9833,N_9676);
xor U10122 (N_10122,N_9617,N_9697);
and U10123 (N_10123,N_9738,N_9720);
nand U10124 (N_10124,N_9706,N_9708);
nor U10125 (N_10125,N_9837,N_9639);
or U10126 (N_10126,N_9710,N_9809);
nand U10127 (N_10127,N_9837,N_9802);
or U10128 (N_10128,N_9829,N_9647);
and U10129 (N_10129,N_9862,N_9730);
and U10130 (N_10130,N_9620,N_9771);
or U10131 (N_10131,N_9674,N_9722);
and U10132 (N_10132,N_9735,N_9843);
nor U10133 (N_10133,N_9758,N_9855);
nand U10134 (N_10134,N_9715,N_9777);
or U10135 (N_10135,N_9747,N_9825);
or U10136 (N_10136,N_9738,N_9817);
nor U10137 (N_10137,N_9786,N_9803);
nor U10138 (N_10138,N_9848,N_9874);
xor U10139 (N_10139,N_9762,N_9606);
nor U10140 (N_10140,N_9851,N_9760);
and U10141 (N_10141,N_9896,N_9830);
nand U10142 (N_10142,N_9760,N_9615);
xnor U10143 (N_10143,N_9815,N_9627);
nor U10144 (N_10144,N_9864,N_9734);
nand U10145 (N_10145,N_9621,N_9607);
xnor U10146 (N_10146,N_9650,N_9601);
and U10147 (N_10147,N_9829,N_9628);
and U10148 (N_10148,N_9669,N_9827);
nor U10149 (N_10149,N_9716,N_9837);
nor U10150 (N_10150,N_9685,N_9791);
or U10151 (N_10151,N_9798,N_9844);
nor U10152 (N_10152,N_9626,N_9789);
and U10153 (N_10153,N_9629,N_9812);
nand U10154 (N_10154,N_9618,N_9635);
or U10155 (N_10155,N_9735,N_9793);
nand U10156 (N_10156,N_9765,N_9803);
or U10157 (N_10157,N_9665,N_9721);
xor U10158 (N_10158,N_9885,N_9756);
and U10159 (N_10159,N_9868,N_9671);
nand U10160 (N_10160,N_9632,N_9600);
and U10161 (N_10161,N_9885,N_9622);
nor U10162 (N_10162,N_9726,N_9890);
or U10163 (N_10163,N_9802,N_9701);
or U10164 (N_10164,N_9737,N_9860);
nand U10165 (N_10165,N_9612,N_9687);
and U10166 (N_10166,N_9783,N_9786);
nand U10167 (N_10167,N_9676,N_9891);
nand U10168 (N_10168,N_9697,N_9878);
nor U10169 (N_10169,N_9690,N_9824);
nor U10170 (N_10170,N_9793,N_9613);
or U10171 (N_10171,N_9764,N_9826);
nand U10172 (N_10172,N_9809,N_9754);
xor U10173 (N_10173,N_9849,N_9843);
nor U10174 (N_10174,N_9628,N_9819);
nand U10175 (N_10175,N_9699,N_9833);
nor U10176 (N_10176,N_9635,N_9721);
nand U10177 (N_10177,N_9898,N_9803);
nand U10178 (N_10178,N_9612,N_9882);
nor U10179 (N_10179,N_9735,N_9710);
and U10180 (N_10180,N_9629,N_9670);
xnor U10181 (N_10181,N_9888,N_9719);
and U10182 (N_10182,N_9629,N_9736);
xnor U10183 (N_10183,N_9801,N_9716);
or U10184 (N_10184,N_9719,N_9853);
and U10185 (N_10185,N_9786,N_9883);
nand U10186 (N_10186,N_9847,N_9761);
and U10187 (N_10187,N_9685,N_9669);
nor U10188 (N_10188,N_9685,N_9810);
or U10189 (N_10189,N_9824,N_9607);
and U10190 (N_10190,N_9673,N_9751);
nor U10191 (N_10191,N_9795,N_9726);
and U10192 (N_10192,N_9688,N_9649);
nand U10193 (N_10193,N_9873,N_9782);
nand U10194 (N_10194,N_9803,N_9797);
and U10195 (N_10195,N_9624,N_9740);
nand U10196 (N_10196,N_9693,N_9654);
and U10197 (N_10197,N_9773,N_9649);
xnor U10198 (N_10198,N_9621,N_9675);
and U10199 (N_10199,N_9716,N_9735);
and U10200 (N_10200,N_10170,N_9905);
xor U10201 (N_10201,N_9967,N_10079);
nor U10202 (N_10202,N_10029,N_9919);
or U10203 (N_10203,N_10113,N_10050);
nand U10204 (N_10204,N_10056,N_10104);
nor U10205 (N_10205,N_10039,N_9960);
and U10206 (N_10206,N_9952,N_10008);
and U10207 (N_10207,N_10100,N_10054);
nor U10208 (N_10208,N_9998,N_10180);
or U10209 (N_10209,N_10147,N_10002);
xnor U10210 (N_10210,N_10169,N_9913);
and U10211 (N_10211,N_10138,N_9947);
xor U10212 (N_10212,N_10165,N_10181);
xnor U10213 (N_10213,N_9937,N_10073);
nor U10214 (N_10214,N_10193,N_10115);
xor U10215 (N_10215,N_9944,N_10091);
or U10216 (N_10216,N_10040,N_9971);
and U10217 (N_10217,N_10037,N_10199);
and U10218 (N_10218,N_10101,N_10148);
nand U10219 (N_10219,N_10108,N_9916);
xnor U10220 (N_10220,N_9974,N_10190);
or U10221 (N_10221,N_10175,N_10015);
and U10222 (N_10222,N_10048,N_10127);
or U10223 (N_10223,N_10025,N_10195);
nor U10224 (N_10224,N_10109,N_10159);
xnor U10225 (N_10225,N_9982,N_9959);
nand U10226 (N_10226,N_9909,N_9924);
nand U10227 (N_10227,N_10131,N_9938);
nand U10228 (N_10228,N_9997,N_10125);
and U10229 (N_10229,N_10005,N_9953);
or U10230 (N_10230,N_9958,N_10064);
or U10231 (N_10231,N_9999,N_10173);
nor U10232 (N_10232,N_10088,N_10179);
nand U10233 (N_10233,N_10007,N_10076);
xnor U10234 (N_10234,N_10185,N_9976);
nand U10235 (N_10235,N_9934,N_10126);
nor U10236 (N_10236,N_9908,N_9981);
nor U10237 (N_10237,N_10060,N_10086);
or U10238 (N_10238,N_9964,N_10102);
xor U10239 (N_10239,N_10003,N_10132);
or U10240 (N_10240,N_9918,N_9943);
and U10241 (N_10241,N_10160,N_10186);
xnor U10242 (N_10242,N_9992,N_10106);
nor U10243 (N_10243,N_10046,N_10083);
nand U10244 (N_10244,N_9901,N_10153);
nand U10245 (N_10245,N_10090,N_10082);
or U10246 (N_10246,N_9903,N_10158);
or U10247 (N_10247,N_9923,N_10033);
and U10248 (N_10248,N_10028,N_9926);
xor U10249 (N_10249,N_10198,N_9989);
or U10250 (N_10250,N_10062,N_9948);
and U10251 (N_10251,N_9950,N_10096);
xor U10252 (N_10252,N_9925,N_10000);
nand U10253 (N_10253,N_10045,N_10098);
nand U10254 (N_10254,N_10194,N_10011);
and U10255 (N_10255,N_10116,N_9973);
nand U10256 (N_10256,N_10023,N_10168);
nand U10257 (N_10257,N_10192,N_10051);
nor U10258 (N_10258,N_9990,N_10140);
and U10259 (N_10259,N_10187,N_9911);
or U10260 (N_10260,N_10154,N_10097);
nand U10261 (N_10261,N_10103,N_10157);
or U10262 (N_10262,N_10026,N_9979);
nor U10263 (N_10263,N_10178,N_10013);
and U10264 (N_10264,N_10123,N_10119);
or U10265 (N_10265,N_10156,N_10139);
nor U10266 (N_10266,N_10164,N_10152);
nand U10267 (N_10267,N_9929,N_9980);
nor U10268 (N_10268,N_10174,N_10141);
nand U10269 (N_10269,N_10093,N_10110);
nor U10270 (N_10270,N_9942,N_9921);
or U10271 (N_10271,N_10124,N_9983);
xnor U10272 (N_10272,N_9957,N_10134);
or U10273 (N_10273,N_9932,N_10171);
and U10274 (N_10274,N_10032,N_10117);
xor U10275 (N_10275,N_10092,N_9966);
or U10276 (N_10276,N_10105,N_9935);
xnor U10277 (N_10277,N_9955,N_10120);
or U10278 (N_10278,N_9945,N_10068);
and U10279 (N_10279,N_10111,N_10089);
and U10280 (N_10280,N_10167,N_10020);
xor U10281 (N_10281,N_10112,N_9946);
and U10282 (N_10282,N_9969,N_9920);
nand U10283 (N_10283,N_9991,N_9972);
or U10284 (N_10284,N_10144,N_9987);
and U10285 (N_10285,N_9963,N_10004);
and U10286 (N_10286,N_9930,N_10183);
and U10287 (N_10287,N_9975,N_9954);
and U10288 (N_10288,N_9927,N_10075);
xnor U10289 (N_10289,N_9941,N_10043);
or U10290 (N_10290,N_10069,N_10063);
or U10291 (N_10291,N_10024,N_10049);
xnor U10292 (N_10292,N_10122,N_10053);
nor U10293 (N_10293,N_9965,N_10145);
nor U10294 (N_10294,N_10143,N_10071);
nand U10295 (N_10295,N_9994,N_10099);
and U10296 (N_10296,N_10166,N_9986);
nor U10297 (N_10297,N_10107,N_10066);
and U10298 (N_10298,N_10016,N_10085);
nor U10299 (N_10299,N_10095,N_10018);
nand U10300 (N_10300,N_10010,N_10135);
xnor U10301 (N_10301,N_9956,N_9984);
nor U10302 (N_10302,N_9931,N_10163);
nand U10303 (N_10303,N_10009,N_10042);
nand U10304 (N_10304,N_10162,N_10021);
xor U10305 (N_10305,N_9902,N_10155);
nor U10306 (N_10306,N_10177,N_10114);
or U10307 (N_10307,N_10038,N_9914);
or U10308 (N_10308,N_9936,N_10118);
and U10309 (N_10309,N_10057,N_9922);
nand U10310 (N_10310,N_9996,N_10133);
or U10311 (N_10311,N_10172,N_10196);
or U10312 (N_10312,N_10151,N_10142);
or U10313 (N_10313,N_10078,N_10137);
and U10314 (N_10314,N_10197,N_10121);
nand U10315 (N_10315,N_9910,N_9988);
nand U10316 (N_10316,N_9928,N_10059);
or U10317 (N_10317,N_10094,N_9907);
nor U10318 (N_10318,N_10047,N_10030);
xor U10319 (N_10319,N_10041,N_10072);
or U10320 (N_10320,N_9906,N_10189);
nor U10321 (N_10321,N_10014,N_10188);
nand U10322 (N_10322,N_10161,N_10061);
xnor U10323 (N_10323,N_10087,N_9933);
or U10324 (N_10324,N_9970,N_10084);
nand U10325 (N_10325,N_9985,N_9917);
nand U10326 (N_10326,N_10022,N_10017);
xor U10327 (N_10327,N_10129,N_10182);
nand U10328 (N_10328,N_9904,N_10031);
xnor U10329 (N_10329,N_9940,N_10176);
or U10330 (N_10330,N_9978,N_10019);
nand U10331 (N_10331,N_10044,N_9977);
and U10332 (N_10332,N_9915,N_9968);
and U10333 (N_10333,N_9962,N_10070);
xnor U10334 (N_10334,N_10001,N_10136);
nor U10335 (N_10335,N_10149,N_10065);
and U10336 (N_10336,N_10081,N_10012);
or U10337 (N_10337,N_9993,N_10077);
xor U10338 (N_10338,N_9939,N_10006);
xnor U10339 (N_10339,N_10052,N_10067);
or U10340 (N_10340,N_9995,N_10034);
xor U10341 (N_10341,N_10184,N_10191);
nand U10342 (N_10342,N_10128,N_9951);
nor U10343 (N_10343,N_10036,N_10146);
xor U10344 (N_10344,N_10035,N_9900);
nand U10345 (N_10345,N_10074,N_10150);
and U10346 (N_10346,N_9949,N_10080);
xnor U10347 (N_10347,N_10058,N_9912);
nor U10348 (N_10348,N_10055,N_10027);
nor U10349 (N_10349,N_9961,N_10130);
or U10350 (N_10350,N_10077,N_9979);
nor U10351 (N_10351,N_10097,N_10041);
nand U10352 (N_10352,N_9936,N_10192);
nand U10353 (N_10353,N_10112,N_9995);
nor U10354 (N_10354,N_9997,N_10175);
nor U10355 (N_10355,N_9924,N_9935);
nand U10356 (N_10356,N_9955,N_10041);
or U10357 (N_10357,N_9995,N_10123);
xnor U10358 (N_10358,N_9925,N_9919);
xnor U10359 (N_10359,N_9965,N_9998);
nand U10360 (N_10360,N_10110,N_10066);
or U10361 (N_10361,N_10057,N_9975);
nor U10362 (N_10362,N_10078,N_10063);
and U10363 (N_10363,N_10162,N_9999);
and U10364 (N_10364,N_10023,N_10021);
nand U10365 (N_10365,N_9991,N_10110);
nand U10366 (N_10366,N_10100,N_10078);
nand U10367 (N_10367,N_9934,N_9921);
and U10368 (N_10368,N_9948,N_9966);
and U10369 (N_10369,N_10094,N_9987);
and U10370 (N_10370,N_9952,N_9976);
or U10371 (N_10371,N_10034,N_10163);
nand U10372 (N_10372,N_10145,N_10093);
or U10373 (N_10373,N_10040,N_10102);
and U10374 (N_10374,N_9919,N_10104);
or U10375 (N_10375,N_10061,N_10048);
and U10376 (N_10376,N_9901,N_10029);
nor U10377 (N_10377,N_9973,N_10043);
nand U10378 (N_10378,N_10095,N_10179);
nand U10379 (N_10379,N_9953,N_10154);
nor U10380 (N_10380,N_9947,N_10176);
and U10381 (N_10381,N_10148,N_10174);
and U10382 (N_10382,N_9947,N_10175);
or U10383 (N_10383,N_9969,N_10121);
and U10384 (N_10384,N_9971,N_10189);
xor U10385 (N_10385,N_9939,N_9920);
nand U10386 (N_10386,N_10138,N_10165);
nor U10387 (N_10387,N_10180,N_9976);
nand U10388 (N_10388,N_10182,N_10027);
or U10389 (N_10389,N_10106,N_10014);
or U10390 (N_10390,N_9923,N_10039);
nand U10391 (N_10391,N_9979,N_10099);
nor U10392 (N_10392,N_10120,N_9908);
xor U10393 (N_10393,N_9992,N_10155);
xor U10394 (N_10394,N_10142,N_10194);
xor U10395 (N_10395,N_10148,N_9974);
xor U10396 (N_10396,N_9992,N_9961);
and U10397 (N_10397,N_10069,N_10133);
and U10398 (N_10398,N_10061,N_10066);
and U10399 (N_10399,N_9985,N_9970);
and U10400 (N_10400,N_10164,N_10197);
or U10401 (N_10401,N_9987,N_9908);
and U10402 (N_10402,N_10021,N_10003);
nor U10403 (N_10403,N_10055,N_9927);
nand U10404 (N_10404,N_10019,N_9943);
and U10405 (N_10405,N_10193,N_10118);
nor U10406 (N_10406,N_10061,N_10077);
nor U10407 (N_10407,N_10124,N_10158);
or U10408 (N_10408,N_9985,N_10114);
nor U10409 (N_10409,N_10163,N_9901);
or U10410 (N_10410,N_10077,N_9968);
nor U10411 (N_10411,N_10109,N_10091);
nand U10412 (N_10412,N_9911,N_10142);
and U10413 (N_10413,N_9998,N_10115);
or U10414 (N_10414,N_10013,N_9968);
or U10415 (N_10415,N_10152,N_10180);
or U10416 (N_10416,N_10122,N_10095);
nand U10417 (N_10417,N_9904,N_10145);
nand U10418 (N_10418,N_10052,N_10145);
and U10419 (N_10419,N_9958,N_10018);
nor U10420 (N_10420,N_10187,N_10076);
or U10421 (N_10421,N_9946,N_10069);
or U10422 (N_10422,N_10117,N_10161);
xor U10423 (N_10423,N_10097,N_9978);
or U10424 (N_10424,N_10035,N_10107);
xor U10425 (N_10425,N_10086,N_9949);
nand U10426 (N_10426,N_9902,N_10195);
and U10427 (N_10427,N_10171,N_9995);
nor U10428 (N_10428,N_9978,N_10139);
nand U10429 (N_10429,N_10057,N_9987);
nand U10430 (N_10430,N_10188,N_10030);
nand U10431 (N_10431,N_10041,N_9967);
nand U10432 (N_10432,N_10037,N_9942);
nor U10433 (N_10433,N_10074,N_10049);
xor U10434 (N_10434,N_10084,N_10053);
nor U10435 (N_10435,N_9920,N_10147);
xor U10436 (N_10436,N_10173,N_10097);
nand U10437 (N_10437,N_10103,N_10099);
or U10438 (N_10438,N_9952,N_10012);
and U10439 (N_10439,N_10120,N_9953);
and U10440 (N_10440,N_10084,N_9932);
nand U10441 (N_10441,N_10193,N_10015);
and U10442 (N_10442,N_10182,N_9975);
and U10443 (N_10443,N_9953,N_10043);
nand U10444 (N_10444,N_10094,N_10165);
or U10445 (N_10445,N_10104,N_9930);
or U10446 (N_10446,N_9955,N_10170);
xor U10447 (N_10447,N_10148,N_9969);
xnor U10448 (N_10448,N_10174,N_10158);
nor U10449 (N_10449,N_9954,N_9995);
or U10450 (N_10450,N_10068,N_10177);
nor U10451 (N_10451,N_10086,N_9904);
xnor U10452 (N_10452,N_9919,N_9930);
nor U10453 (N_10453,N_9932,N_10063);
or U10454 (N_10454,N_10136,N_10079);
nand U10455 (N_10455,N_10127,N_10123);
nor U10456 (N_10456,N_9904,N_10115);
nand U10457 (N_10457,N_10024,N_10166);
nand U10458 (N_10458,N_10023,N_10198);
xor U10459 (N_10459,N_10163,N_10056);
nand U10460 (N_10460,N_10142,N_9932);
xor U10461 (N_10461,N_9946,N_10115);
and U10462 (N_10462,N_9921,N_9923);
and U10463 (N_10463,N_10074,N_10100);
and U10464 (N_10464,N_9910,N_10109);
xnor U10465 (N_10465,N_10090,N_10137);
or U10466 (N_10466,N_9942,N_10065);
nor U10467 (N_10467,N_10040,N_10094);
or U10468 (N_10468,N_9921,N_10028);
nand U10469 (N_10469,N_10151,N_9952);
and U10470 (N_10470,N_10176,N_10150);
and U10471 (N_10471,N_10121,N_10072);
nand U10472 (N_10472,N_9914,N_10161);
or U10473 (N_10473,N_9960,N_9994);
or U10474 (N_10474,N_9903,N_10046);
and U10475 (N_10475,N_10119,N_10127);
nor U10476 (N_10476,N_9916,N_10034);
nor U10477 (N_10477,N_9947,N_10099);
xor U10478 (N_10478,N_10067,N_10090);
nand U10479 (N_10479,N_10185,N_9915);
or U10480 (N_10480,N_10184,N_9983);
nor U10481 (N_10481,N_10084,N_10162);
nand U10482 (N_10482,N_9918,N_9958);
and U10483 (N_10483,N_9987,N_10127);
or U10484 (N_10484,N_10102,N_9926);
nand U10485 (N_10485,N_10082,N_10191);
or U10486 (N_10486,N_10177,N_9970);
nor U10487 (N_10487,N_9916,N_10020);
nand U10488 (N_10488,N_9929,N_10102);
and U10489 (N_10489,N_9923,N_9928);
nand U10490 (N_10490,N_10194,N_9928);
or U10491 (N_10491,N_10167,N_9971);
nor U10492 (N_10492,N_9990,N_10183);
xnor U10493 (N_10493,N_9991,N_10122);
and U10494 (N_10494,N_10135,N_10061);
and U10495 (N_10495,N_10114,N_10134);
nor U10496 (N_10496,N_10169,N_10029);
nand U10497 (N_10497,N_9961,N_9910);
or U10498 (N_10498,N_10162,N_10170);
nand U10499 (N_10499,N_9985,N_9926);
xnor U10500 (N_10500,N_10405,N_10343);
or U10501 (N_10501,N_10445,N_10346);
or U10502 (N_10502,N_10418,N_10288);
xor U10503 (N_10503,N_10248,N_10218);
nor U10504 (N_10504,N_10320,N_10252);
or U10505 (N_10505,N_10460,N_10254);
nor U10506 (N_10506,N_10373,N_10419);
and U10507 (N_10507,N_10358,N_10206);
and U10508 (N_10508,N_10241,N_10387);
nand U10509 (N_10509,N_10340,N_10426);
or U10510 (N_10510,N_10287,N_10223);
or U10511 (N_10511,N_10214,N_10407);
and U10512 (N_10512,N_10285,N_10383);
xnor U10513 (N_10513,N_10303,N_10388);
nand U10514 (N_10514,N_10255,N_10441);
nor U10515 (N_10515,N_10447,N_10274);
nand U10516 (N_10516,N_10294,N_10203);
and U10517 (N_10517,N_10385,N_10275);
nand U10518 (N_10518,N_10257,N_10456);
nand U10519 (N_10519,N_10327,N_10313);
nor U10520 (N_10520,N_10415,N_10413);
and U10521 (N_10521,N_10236,N_10348);
or U10522 (N_10522,N_10310,N_10264);
nor U10523 (N_10523,N_10361,N_10446);
or U10524 (N_10524,N_10334,N_10448);
or U10525 (N_10525,N_10300,N_10296);
xor U10526 (N_10526,N_10490,N_10424);
nand U10527 (N_10527,N_10462,N_10484);
and U10528 (N_10528,N_10459,N_10495);
xnor U10529 (N_10529,N_10216,N_10307);
nor U10530 (N_10530,N_10399,N_10375);
nand U10531 (N_10531,N_10233,N_10226);
or U10532 (N_10532,N_10457,N_10379);
and U10533 (N_10533,N_10369,N_10243);
xnor U10534 (N_10534,N_10440,N_10409);
and U10535 (N_10535,N_10488,N_10208);
and U10536 (N_10536,N_10434,N_10472);
and U10537 (N_10537,N_10229,N_10230);
xor U10538 (N_10538,N_10325,N_10240);
nand U10539 (N_10539,N_10332,N_10353);
or U10540 (N_10540,N_10271,N_10485);
or U10541 (N_10541,N_10480,N_10266);
nand U10542 (N_10542,N_10333,N_10256);
xor U10543 (N_10543,N_10272,N_10225);
nor U10544 (N_10544,N_10464,N_10468);
nand U10545 (N_10545,N_10279,N_10481);
or U10546 (N_10546,N_10444,N_10317);
nor U10547 (N_10547,N_10276,N_10473);
and U10548 (N_10548,N_10471,N_10262);
nor U10549 (N_10549,N_10319,N_10431);
xnor U10550 (N_10550,N_10304,N_10258);
xor U10551 (N_10551,N_10430,N_10368);
or U10552 (N_10552,N_10392,N_10224);
and U10553 (N_10553,N_10377,N_10253);
and U10554 (N_10554,N_10284,N_10416);
xnor U10555 (N_10555,N_10278,N_10398);
nand U10556 (N_10556,N_10268,N_10201);
and U10557 (N_10557,N_10466,N_10302);
nor U10558 (N_10558,N_10357,N_10293);
nand U10559 (N_10559,N_10492,N_10234);
and U10560 (N_10560,N_10386,N_10267);
and U10561 (N_10561,N_10299,N_10238);
nor U10562 (N_10562,N_10423,N_10259);
nand U10563 (N_10563,N_10232,N_10382);
and U10564 (N_10564,N_10401,N_10378);
xnor U10565 (N_10565,N_10482,N_10355);
nand U10566 (N_10566,N_10298,N_10396);
or U10567 (N_10567,N_10371,N_10433);
or U10568 (N_10568,N_10207,N_10328);
and U10569 (N_10569,N_10393,N_10477);
nand U10570 (N_10570,N_10350,N_10443);
nand U10571 (N_10571,N_10273,N_10402);
nand U10572 (N_10572,N_10452,N_10250);
xnor U10573 (N_10573,N_10360,N_10221);
or U10574 (N_10574,N_10322,N_10364);
and U10575 (N_10575,N_10499,N_10367);
xor U10576 (N_10576,N_10394,N_10412);
and U10577 (N_10577,N_10289,N_10458);
or U10578 (N_10578,N_10249,N_10493);
nand U10579 (N_10579,N_10395,N_10404);
and U10580 (N_10580,N_10354,N_10215);
xnor U10581 (N_10581,N_10269,N_10261);
nor U10582 (N_10582,N_10479,N_10245);
and U10583 (N_10583,N_10321,N_10489);
nor U10584 (N_10584,N_10366,N_10453);
xor U10585 (N_10585,N_10345,N_10370);
nand U10586 (N_10586,N_10376,N_10421);
nand U10587 (N_10587,N_10432,N_10389);
and U10588 (N_10588,N_10309,N_10286);
xnor U10589 (N_10589,N_10292,N_10380);
nand U10590 (N_10590,N_10403,N_10295);
nand U10591 (N_10591,N_10429,N_10476);
xnor U10592 (N_10592,N_10384,N_10372);
nand U10593 (N_10593,N_10204,N_10239);
xor U10594 (N_10594,N_10474,N_10342);
nand U10595 (N_10595,N_10242,N_10437);
xnor U10596 (N_10596,N_10337,N_10381);
and U10597 (N_10597,N_10470,N_10314);
nor U10598 (N_10598,N_10335,N_10222);
nor U10599 (N_10599,N_10455,N_10359);
nor U10600 (N_10600,N_10246,N_10281);
or U10601 (N_10601,N_10260,N_10497);
nor U10602 (N_10602,N_10341,N_10263);
nand U10603 (N_10603,N_10220,N_10291);
and U10604 (N_10604,N_10491,N_10330);
or U10605 (N_10605,N_10283,N_10211);
nand U10606 (N_10606,N_10237,N_10280);
nand U10607 (N_10607,N_10217,N_10465);
nand U10608 (N_10608,N_10339,N_10336);
xnor U10609 (N_10609,N_10362,N_10420);
nor U10610 (N_10610,N_10200,N_10391);
and U10611 (N_10611,N_10410,N_10406);
nor U10612 (N_10612,N_10311,N_10270);
and U10613 (N_10613,N_10439,N_10247);
and U10614 (N_10614,N_10400,N_10265);
nand U10615 (N_10615,N_10352,N_10312);
xor U10616 (N_10616,N_10228,N_10483);
nor U10617 (N_10617,N_10210,N_10351);
and U10618 (N_10618,N_10486,N_10449);
nand U10619 (N_10619,N_10251,N_10344);
xnor U10620 (N_10620,N_10338,N_10463);
nand U10621 (N_10621,N_10306,N_10475);
nor U10622 (N_10622,N_10451,N_10305);
nor U10623 (N_10623,N_10478,N_10390);
nand U10624 (N_10624,N_10467,N_10202);
and U10625 (N_10625,N_10212,N_10301);
nor U10626 (N_10626,N_10326,N_10435);
or U10627 (N_10627,N_10454,N_10417);
xor U10628 (N_10628,N_10461,N_10408);
and U10629 (N_10629,N_10244,N_10496);
nand U10630 (N_10630,N_10277,N_10469);
nor U10631 (N_10631,N_10323,N_10315);
or U10632 (N_10632,N_10290,N_10428);
xnor U10633 (N_10633,N_10494,N_10318);
or U10634 (N_10634,N_10487,N_10329);
nand U10635 (N_10635,N_10347,N_10414);
nand U10636 (N_10636,N_10436,N_10308);
and U10637 (N_10637,N_10213,N_10282);
nand U10638 (N_10638,N_10450,N_10411);
nand U10639 (N_10639,N_10297,N_10442);
xnor U10640 (N_10640,N_10363,N_10331);
xor U10641 (N_10641,N_10365,N_10498);
or U10642 (N_10642,N_10316,N_10219);
or U10643 (N_10643,N_10205,N_10227);
and U10644 (N_10644,N_10324,N_10374);
and U10645 (N_10645,N_10397,N_10438);
nand U10646 (N_10646,N_10235,N_10422);
xor U10647 (N_10647,N_10231,N_10356);
and U10648 (N_10648,N_10427,N_10209);
and U10649 (N_10649,N_10349,N_10425);
nor U10650 (N_10650,N_10242,N_10381);
and U10651 (N_10651,N_10464,N_10329);
nand U10652 (N_10652,N_10361,N_10226);
or U10653 (N_10653,N_10315,N_10424);
nor U10654 (N_10654,N_10209,N_10498);
nor U10655 (N_10655,N_10222,N_10327);
xor U10656 (N_10656,N_10296,N_10445);
and U10657 (N_10657,N_10297,N_10411);
or U10658 (N_10658,N_10220,N_10319);
or U10659 (N_10659,N_10290,N_10423);
nor U10660 (N_10660,N_10324,N_10208);
xor U10661 (N_10661,N_10437,N_10356);
nor U10662 (N_10662,N_10476,N_10425);
and U10663 (N_10663,N_10440,N_10365);
or U10664 (N_10664,N_10468,N_10299);
nand U10665 (N_10665,N_10259,N_10323);
xor U10666 (N_10666,N_10265,N_10353);
or U10667 (N_10667,N_10399,N_10223);
and U10668 (N_10668,N_10247,N_10433);
nor U10669 (N_10669,N_10418,N_10454);
nand U10670 (N_10670,N_10378,N_10200);
nor U10671 (N_10671,N_10421,N_10292);
and U10672 (N_10672,N_10271,N_10362);
or U10673 (N_10673,N_10401,N_10279);
xnor U10674 (N_10674,N_10229,N_10346);
nand U10675 (N_10675,N_10442,N_10441);
and U10676 (N_10676,N_10485,N_10281);
xnor U10677 (N_10677,N_10368,N_10379);
and U10678 (N_10678,N_10308,N_10218);
and U10679 (N_10679,N_10459,N_10286);
nand U10680 (N_10680,N_10271,N_10371);
nor U10681 (N_10681,N_10370,N_10415);
xnor U10682 (N_10682,N_10448,N_10499);
nand U10683 (N_10683,N_10251,N_10346);
nor U10684 (N_10684,N_10455,N_10289);
or U10685 (N_10685,N_10225,N_10236);
or U10686 (N_10686,N_10238,N_10213);
nand U10687 (N_10687,N_10263,N_10488);
nand U10688 (N_10688,N_10395,N_10385);
and U10689 (N_10689,N_10493,N_10385);
nand U10690 (N_10690,N_10366,N_10441);
xor U10691 (N_10691,N_10443,N_10338);
or U10692 (N_10692,N_10371,N_10340);
and U10693 (N_10693,N_10418,N_10408);
and U10694 (N_10694,N_10356,N_10367);
or U10695 (N_10695,N_10360,N_10317);
and U10696 (N_10696,N_10449,N_10325);
and U10697 (N_10697,N_10246,N_10478);
or U10698 (N_10698,N_10335,N_10468);
nor U10699 (N_10699,N_10388,N_10493);
or U10700 (N_10700,N_10424,N_10207);
nor U10701 (N_10701,N_10312,N_10244);
xor U10702 (N_10702,N_10493,N_10239);
nor U10703 (N_10703,N_10322,N_10296);
or U10704 (N_10704,N_10393,N_10469);
and U10705 (N_10705,N_10322,N_10430);
xnor U10706 (N_10706,N_10466,N_10496);
xor U10707 (N_10707,N_10207,N_10420);
and U10708 (N_10708,N_10315,N_10475);
xnor U10709 (N_10709,N_10250,N_10352);
xor U10710 (N_10710,N_10316,N_10206);
or U10711 (N_10711,N_10225,N_10279);
nand U10712 (N_10712,N_10308,N_10397);
xor U10713 (N_10713,N_10391,N_10216);
and U10714 (N_10714,N_10296,N_10275);
nor U10715 (N_10715,N_10451,N_10212);
or U10716 (N_10716,N_10269,N_10481);
nor U10717 (N_10717,N_10396,N_10368);
or U10718 (N_10718,N_10319,N_10238);
or U10719 (N_10719,N_10416,N_10403);
nor U10720 (N_10720,N_10420,N_10337);
and U10721 (N_10721,N_10348,N_10363);
nor U10722 (N_10722,N_10279,N_10324);
or U10723 (N_10723,N_10309,N_10473);
xor U10724 (N_10724,N_10444,N_10403);
nor U10725 (N_10725,N_10210,N_10308);
nor U10726 (N_10726,N_10410,N_10341);
nand U10727 (N_10727,N_10303,N_10286);
or U10728 (N_10728,N_10327,N_10362);
nand U10729 (N_10729,N_10297,N_10359);
or U10730 (N_10730,N_10236,N_10361);
nor U10731 (N_10731,N_10222,N_10415);
nand U10732 (N_10732,N_10301,N_10282);
and U10733 (N_10733,N_10264,N_10447);
or U10734 (N_10734,N_10405,N_10344);
xor U10735 (N_10735,N_10356,N_10428);
nand U10736 (N_10736,N_10455,N_10452);
nor U10737 (N_10737,N_10353,N_10263);
xnor U10738 (N_10738,N_10491,N_10250);
and U10739 (N_10739,N_10377,N_10224);
or U10740 (N_10740,N_10430,N_10431);
and U10741 (N_10741,N_10379,N_10314);
or U10742 (N_10742,N_10240,N_10472);
and U10743 (N_10743,N_10331,N_10237);
or U10744 (N_10744,N_10374,N_10288);
nor U10745 (N_10745,N_10333,N_10465);
or U10746 (N_10746,N_10450,N_10293);
or U10747 (N_10747,N_10384,N_10469);
xnor U10748 (N_10748,N_10354,N_10444);
nand U10749 (N_10749,N_10272,N_10206);
nor U10750 (N_10750,N_10385,N_10323);
or U10751 (N_10751,N_10484,N_10496);
nor U10752 (N_10752,N_10409,N_10427);
nand U10753 (N_10753,N_10362,N_10436);
and U10754 (N_10754,N_10220,N_10257);
xnor U10755 (N_10755,N_10366,N_10497);
nand U10756 (N_10756,N_10482,N_10453);
nand U10757 (N_10757,N_10288,N_10404);
and U10758 (N_10758,N_10270,N_10490);
nor U10759 (N_10759,N_10260,N_10437);
xor U10760 (N_10760,N_10395,N_10367);
or U10761 (N_10761,N_10345,N_10266);
or U10762 (N_10762,N_10434,N_10284);
and U10763 (N_10763,N_10292,N_10383);
and U10764 (N_10764,N_10347,N_10221);
nor U10765 (N_10765,N_10338,N_10425);
nor U10766 (N_10766,N_10348,N_10220);
nand U10767 (N_10767,N_10478,N_10499);
xnor U10768 (N_10768,N_10281,N_10268);
nand U10769 (N_10769,N_10462,N_10315);
xnor U10770 (N_10770,N_10252,N_10490);
and U10771 (N_10771,N_10318,N_10372);
xnor U10772 (N_10772,N_10469,N_10322);
nand U10773 (N_10773,N_10346,N_10434);
or U10774 (N_10774,N_10499,N_10275);
nor U10775 (N_10775,N_10461,N_10427);
xnor U10776 (N_10776,N_10358,N_10340);
nand U10777 (N_10777,N_10257,N_10216);
and U10778 (N_10778,N_10382,N_10485);
nand U10779 (N_10779,N_10496,N_10234);
nor U10780 (N_10780,N_10352,N_10440);
xor U10781 (N_10781,N_10362,N_10335);
nor U10782 (N_10782,N_10210,N_10341);
nand U10783 (N_10783,N_10464,N_10305);
nor U10784 (N_10784,N_10319,N_10369);
or U10785 (N_10785,N_10337,N_10318);
xnor U10786 (N_10786,N_10490,N_10275);
or U10787 (N_10787,N_10438,N_10247);
or U10788 (N_10788,N_10493,N_10294);
and U10789 (N_10789,N_10314,N_10394);
and U10790 (N_10790,N_10448,N_10266);
or U10791 (N_10791,N_10318,N_10303);
and U10792 (N_10792,N_10332,N_10272);
xor U10793 (N_10793,N_10312,N_10332);
and U10794 (N_10794,N_10380,N_10439);
and U10795 (N_10795,N_10221,N_10447);
and U10796 (N_10796,N_10318,N_10348);
xnor U10797 (N_10797,N_10292,N_10217);
xnor U10798 (N_10798,N_10322,N_10332);
nor U10799 (N_10799,N_10479,N_10465);
nor U10800 (N_10800,N_10541,N_10623);
xor U10801 (N_10801,N_10653,N_10567);
and U10802 (N_10802,N_10558,N_10589);
nand U10803 (N_10803,N_10610,N_10678);
and U10804 (N_10804,N_10578,N_10507);
nand U10805 (N_10805,N_10561,N_10745);
nand U10806 (N_10806,N_10786,N_10620);
nand U10807 (N_10807,N_10570,N_10532);
and U10808 (N_10808,N_10650,N_10547);
nor U10809 (N_10809,N_10714,N_10711);
or U10810 (N_10810,N_10764,N_10528);
or U10811 (N_10811,N_10747,N_10503);
nand U10812 (N_10812,N_10624,N_10735);
nor U10813 (N_10813,N_10577,N_10562);
nor U10814 (N_10814,N_10795,N_10686);
xnor U10815 (N_10815,N_10593,N_10749);
or U10816 (N_10816,N_10613,N_10753);
nand U10817 (N_10817,N_10664,N_10649);
nor U10818 (N_10818,N_10693,N_10515);
and U10819 (N_10819,N_10676,N_10603);
nor U10820 (N_10820,N_10772,N_10658);
xnor U10821 (N_10821,N_10571,N_10703);
nand U10822 (N_10822,N_10636,N_10672);
nor U10823 (N_10823,N_10796,N_10778);
nand U10824 (N_10824,N_10768,N_10504);
and U10825 (N_10825,N_10712,N_10557);
or U10826 (N_10826,N_10677,N_10596);
nand U10827 (N_10827,N_10704,N_10709);
and U10828 (N_10828,N_10741,N_10725);
and U10829 (N_10829,N_10523,N_10780);
nor U10830 (N_10830,N_10595,N_10785);
xnor U10831 (N_10831,N_10627,N_10536);
or U10832 (N_10832,N_10534,N_10537);
xor U10833 (N_10833,N_10614,N_10789);
or U10834 (N_10834,N_10581,N_10750);
xor U10835 (N_10835,N_10621,N_10584);
and U10836 (N_10836,N_10628,N_10645);
nand U10837 (N_10837,N_10544,N_10533);
nand U10838 (N_10838,N_10759,N_10762);
and U10839 (N_10839,N_10654,N_10739);
and U10840 (N_10840,N_10530,N_10667);
xnor U10841 (N_10841,N_10559,N_10738);
xor U10842 (N_10842,N_10708,N_10661);
xnor U10843 (N_10843,N_10788,N_10763);
nand U10844 (N_10844,N_10542,N_10767);
xor U10845 (N_10845,N_10692,N_10553);
nand U10846 (N_10846,N_10682,N_10619);
and U10847 (N_10847,N_10668,N_10510);
xnor U10848 (N_10848,N_10638,N_10605);
nand U10849 (N_10849,N_10520,N_10582);
or U10850 (N_10850,N_10509,N_10508);
nand U10851 (N_10851,N_10666,N_10773);
or U10852 (N_10852,N_10798,N_10500);
nor U10853 (N_10853,N_10643,N_10782);
nor U10854 (N_10854,N_10684,N_10646);
xnor U10855 (N_10855,N_10514,N_10512);
nor U10856 (N_10856,N_10794,N_10549);
and U10857 (N_10857,N_10572,N_10550);
and U10858 (N_10858,N_10531,N_10642);
nor U10859 (N_10859,N_10633,N_10560);
nor U10860 (N_10860,N_10612,N_10580);
nor U10861 (N_10861,N_10784,N_10518);
and U10862 (N_10862,N_10710,N_10724);
nor U10863 (N_10863,N_10591,N_10565);
nand U10864 (N_10864,N_10715,N_10700);
nand U10865 (N_10865,N_10742,N_10607);
xor U10866 (N_10866,N_10630,N_10655);
xor U10867 (N_10867,N_10594,N_10637);
and U10868 (N_10868,N_10616,N_10790);
nand U10869 (N_10869,N_10516,N_10679);
xor U10870 (N_10870,N_10727,N_10617);
nand U10871 (N_10871,N_10644,N_10588);
nand U10872 (N_10872,N_10718,N_10635);
nand U10873 (N_10873,N_10583,N_10760);
nand U10874 (N_10874,N_10662,N_10733);
nor U10875 (N_10875,N_10699,N_10587);
and U10876 (N_10876,N_10713,N_10652);
nand U10877 (N_10877,N_10506,N_10706);
and U10878 (N_10878,N_10698,N_10761);
and U10879 (N_10879,N_10629,N_10511);
or U10880 (N_10880,N_10774,N_10600);
and U10881 (N_10881,N_10769,N_10543);
nand U10882 (N_10882,N_10740,N_10590);
nand U10883 (N_10883,N_10669,N_10721);
or U10884 (N_10884,N_10770,N_10746);
or U10885 (N_10885,N_10731,N_10564);
nand U10886 (N_10886,N_10674,N_10734);
nor U10887 (N_10887,N_10601,N_10576);
xor U10888 (N_10888,N_10728,N_10551);
or U10889 (N_10889,N_10639,N_10556);
nor U10890 (N_10890,N_10793,N_10688);
xnor U10891 (N_10891,N_10680,N_10776);
nand U10892 (N_10892,N_10615,N_10502);
and U10893 (N_10893,N_10690,N_10701);
xnor U10894 (N_10894,N_10597,N_10573);
xor U10895 (N_10895,N_10548,N_10771);
and U10896 (N_10896,N_10799,N_10640);
nor U10897 (N_10897,N_10505,N_10729);
or U10898 (N_10898,N_10566,N_10694);
xnor U10899 (N_10899,N_10608,N_10719);
or U10900 (N_10900,N_10775,N_10632);
or U10901 (N_10901,N_10579,N_10585);
and U10902 (N_10902,N_10797,N_10671);
nor U10903 (N_10903,N_10501,N_10622);
nand U10904 (N_10904,N_10602,N_10681);
nand U10905 (N_10905,N_10777,N_10521);
nor U10906 (N_10906,N_10540,N_10670);
xnor U10907 (N_10907,N_10525,N_10609);
nor U10908 (N_10908,N_10513,N_10598);
nor U10909 (N_10909,N_10683,N_10611);
nand U10910 (N_10910,N_10522,N_10535);
xor U10911 (N_10911,N_10563,N_10604);
or U10912 (N_10912,N_10569,N_10779);
and U10913 (N_10913,N_10791,N_10575);
nand U10914 (N_10914,N_10527,N_10765);
nor U10915 (N_10915,N_10618,N_10730);
or U10916 (N_10916,N_10631,N_10599);
xor U10917 (N_10917,N_10526,N_10647);
or U10918 (N_10918,N_10552,N_10758);
and U10919 (N_10919,N_10783,N_10545);
xnor U10920 (N_10920,N_10720,N_10687);
or U10921 (N_10921,N_10722,N_10625);
or U10922 (N_10922,N_10660,N_10754);
or U10923 (N_10923,N_10695,N_10539);
nand U10924 (N_10924,N_10751,N_10648);
nand U10925 (N_10925,N_10781,N_10787);
or U10926 (N_10926,N_10606,N_10726);
nor U10927 (N_10927,N_10685,N_10675);
and U10928 (N_10928,N_10524,N_10691);
nand U10929 (N_10929,N_10519,N_10574);
xnor U10930 (N_10930,N_10736,N_10656);
or U10931 (N_10931,N_10529,N_10752);
or U10932 (N_10932,N_10568,N_10517);
or U10933 (N_10933,N_10546,N_10657);
xnor U10934 (N_10934,N_10744,N_10716);
and U10935 (N_10935,N_10689,N_10766);
xnor U10936 (N_10936,N_10641,N_10792);
xnor U10937 (N_10937,N_10756,N_10697);
and U10938 (N_10938,N_10665,N_10696);
or U10939 (N_10939,N_10673,N_10743);
and U10940 (N_10940,N_10634,N_10651);
or U10941 (N_10941,N_10717,N_10757);
xor U10942 (N_10942,N_10538,N_10554);
and U10943 (N_10943,N_10755,N_10555);
and U10944 (N_10944,N_10705,N_10732);
xor U10945 (N_10945,N_10663,N_10626);
nor U10946 (N_10946,N_10748,N_10723);
xor U10947 (N_10947,N_10702,N_10592);
xor U10948 (N_10948,N_10586,N_10737);
nand U10949 (N_10949,N_10659,N_10707);
or U10950 (N_10950,N_10751,N_10511);
xnor U10951 (N_10951,N_10643,N_10699);
xor U10952 (N_10952,N_10759,N_10649);
nand U10953 (N_10953,N_10649,N_10556);
nand U10954 (N_10954,N_10750,N_10672);
xor U10955 (N_10955,N_10650,N_10638);
nor U10956 (N_10956,N_10540,N_10577);
or U10957 (N_10957,N_10558,N_10746);
xor U10958 (N_10958,N_10779,N_10775);
and U10959 (N_10959,N_10774,N_10563);
or U10960 (N_10960,N_10615,N_10738);
or U10961 (N_10961,N_10602,N_10551);
and U10962 (N_10962,N_10721,N_10716);
or U10963 (N_10963,N_10697,N_10572);
nor U10964 (N_10964,N_10713,N_10710);
or U10965 (N_10965,N_10523,N_10542);
xor U10966 (N_10966,N_10689,N_10656);
xnor U10967 (N_10967,N_10655,N_10782);
nor U10968 (N_10968,N_10686,N_10584);
or U10969 (N_10969,N_10609,N_10593);
and U10970 (N_10970,N_10667,N_10678);
and U10971 (N_10971,N_10792,N_10566);
and U10972 (N_10972,N_10675,N_10703);
or U10973 (N_10973,N_10555,N_10551);
or U10974 (N_10974,N_10560,N_10669);
nand U10975 (N_10975,N_10564,N_10576);
nor U10976 (N_10976,N_10651,N_10520);
nor U10977 (N_10977,N_10526,N_10776);
nand U10978 (N_10978,N_10515,N_10686);
or U10979 (N_10979,N_10575,N_10706);
or U10980 (N_10980,N_10516,N_10755);
nand U10981 (N_10981,N_10565,N_10787);
or U10982 (N_10982,N_10640,N_10743);
and U10983 (N_10983,N_10590,N_10684);
nand U10984 (N_10984,N_10502,N_10671);
and U10985 (N_10985,N_10716,N_10532);
and U10986 (N_10986,N_10564,N_10683);
or U10987 (N_10987,N_10585,N_10783);
xnor U10988 (N_10988,N_10611,N_10735);
or U10989 (N_10989,N_10753,N_10686);
nor U10990 (N_10990,N_10675,N_10761);
nand U10991 (N_10991,N_10790,N_10718);
or U10992 (N_10992,N_10507,N_10670);
nor U10993 (N_10993,N_10634,N_10699);
and U10994 (N_10994,N_10537,N_10724);
nor U10995 (N_10995,N_10672,N_10678);
xnor U10996 (N_10996,N_10621,N_10503);
nor U10997 (N_10997,N_10773,N_10525);
and U10998 (N_10998,N_10588,N_10548);
and U10999 (N_10999,N_10758,N_10598);
nor U11000 (N_11000,N_10639,N_10762);
or U11001 (N_11001,N_10668,N_10521);
xor U11002 (N_11002,N_10644,N_10668);
nor U11003 (N_11003,N_10595,N_10782);
xnor U11004 (N_11004,N_10750,N_10566);
or U11005 (N_11005,N_10501,N_10730);
and U11006 (N_11006,N_10678,N_10541);
nand U11007 (N_11007,N_10506,N_10756);
nor U11008 (N_11008,N_10625,N_10642);
and U11009 (N_11009,N_10673,N_10573);
or U11010 (N_11010,N_10652,N_10529);
nor U11011 (N_11011,N_10698,N_10620);
nand U11012 (N_11012,N_10561,N_10661);
nor U11013 (N_11013,N_10531,N_10730);
xor U11014 (N_11014,N_10621,N_10502);
and U11015 (N_11015,N_10717,N_10731);
or U11016 (N_11016,N_10619,N_10615);
and U11017 (N_11017,N_10506,N_10555);
nand U11018 (N_11018,N_10500,N_10674);
and U11019 (N_11019,N_10573,N_10636);
nor U11020 (N_11020,N_10557,N_10711);
nor U11021 (N_11021,N_10503,N_10651);
and U11022 (N_11022,N_10693,N_10691);
nor U11023 (N_11023,N_10683,N_10706);
nor U11024 (N_11024,N_10782,N_10615);
nor U11025 (N_11025,N_10758,N_10575);
xor U11026 (N_11026,N_10752,N_10559);
or U11027 (N_11027,N_10655,N_10671);
or U11028 (N_11028,N_10623,N_10754);
nand U11029 (N_11029,N_10562,N_10762);
and U11030 (N_11030,N_10531,N_10529);
or U11031 (N_11031,N_10656,N_10731);
and U11032 (N_11032,N_10684,N_10522);
xor U11033 (N_11033,N_10650,N_10642);
and U11034 (N_11034,N_10730,N_10650);
or U11035 (N_11035,N_10524,N_10783);
and U11036 (N_11036,N_10698,N_10592);
or U11037 (N_11037,N_10727,N_10698);
xor U11038 (N_11038,N_10653,N_10680);
or U11039 (N_11039,N_10687,N_10690);
and U11040 (N_11040,N_10757,N_10644);
or U11041 (N_11041,N_10552,N_10676);
nor U11042 (N_11042,N_10558,N_10586);
nor U11043 (N_11043,N_10537,N_10524);
and U11044 (N_11044,N_10513,N_10684);
or U11045 (N_11045,N_10611,N_10659);
nor U11046 (N_11046,N_10619,N_10700);
and U11047 (N_11047,N_10666,N_10767);
nand U11048 (N_11048,N_10734,N_10579);
nand U11049 (N_11049,N_10701,N_10587);
and U11050 (N_11050,N_10623,N_10716);
or U11051 (N_11051,N_10721,N_10588);
xor U11052 (N_11052,N_10730,N_10620);
or U11053 (N_11053,N_10629,N_10532);
xnor U11054 (N_11054,N_10513,N_10602);
xor U11055 (N_11055,N_10734,N_10638);
and U11056 (N_11056,N_10798,N_10527);
nor U11057 (N_11057,N_10608,N_10721);
nor U11058 (N_11058,N_10532,N_10696);
nor U11059 (N_11059,N_10791,N_10538);
or U11060 (N_11060,N_10688,N_10775);
nand U11061 (N_11061,N_10691,N_10743);
and U11062 (N_11062,N_10768,N_10542);
nor U11063 (N_11063,N_10595,N_10552);
or U11064 (N_11064,N_10736,N_10550);
or U11065 (N_11065,N_10568,N_10503);
xor U11066 (N_11066,N_10753,N_10566);
xnor U11067 (N_11067,N_10550,N_10515);
and U11068 (N_11068,N_10700,N_10580);
nor U11069 (N_11069,N_10745,N_10559);
nor U11070 (N_11070,N_10551,N_10789);
nand U11071 (N_11071,N_10776,N_10563);
or U11072 (N_11072,N_10758,N_10522);
nand U11073 (N_11073,N_10569,N_10682);
xnor U11074 (N_11074,N_10677,N_10659);
nand U11075 (N_11075,N_10623,N_10711);
nor U11076 (N_11076,N_10723,N_10746);
or U11077 (N_11077,N_10647,N_10788);
nor U11078 (N_11078,N_10585,N_10653);
and U11079 (N_11079,N_10720,N_10773);
xor U11080 (N_11080,N_10590,N_10517);
nor U11081 (N_11081,N_10653,N_10736);
or U11082 (N_11082,N_10776,N_10523);
nand U11083 (N_11083,N_10754,N_10520);
nand U11084 (N_11084,N_10509,N_10572);
xnor U11085 (N_11085,N_10739,N_10563);
and U11086 (N_11086,N_10570,N_10704);
and U11087 (N_11087,N_10738,N_10747);
nand U11088 (N_11088,N_10774,N_10776);
or U11089 (N_11089,N_10563,N_10644);
nand U11090 (N_11090,N_10500,N_10789);
or U11091 (N_11091,N_10627,N_10587);
nand U11092 (N_11092,N_10634,N_10612);
nand U11093 (N_11093,N_10798,N_10614);
nand U11094 (N_11094,N_10744,N_10712);
nand U11095 (N_11095,N_10566,N_10515);
and U11096 (N_11096,N_10774,N_10645);
nand U11097 (N_11097,N_10741,N_10765);
nand U11098 (N_11098,N_10785,N_10612);
or U11099 (N_11099,N_10721,N_10607);
and U11100 (N_11100,N_10819,N_10863);
and U11101 (N_11101,N_10996,N_10939);
and U11102 (N_11102,N_10812,N_10831);
or U11103 (N_11103,N_11027,N_10985);
nor U11104 (N_11104,N_10884,N_10937);
nand U11105 (N_11105,N_10967,N_10981);
xor U11106 (N_11106,N_10908,N_11005);
xnor U11107 (N_11107,N_10961,N_11032);
xor U11108 (N_11108,N_10933,N_10929);
and U11109 (N_11109,N_11003,N_10823);
nor U11110 (N_11110,N_10916,N_10962);
and U11111 (N_11111,N_11076,N_11039);
nand U11112 (N_11112,N_11019,N_11068);
or U11113 (N_11113,N_11020,N_11085);
or U11114 (N_11114,N_11061,N_10803);
xnor U11115 (N_11115,N_10953,N_10815);
nor U11116 (N_11116,N_10903,N_10988);
or U11117 (N_11117,N_11035,N_10851);
and U11118 (N_11118,N_10820,N_10972);
nor U11119 (N_11119,N_11052,N_10817);
nand U11120 (N_11120,N_10917,N_11042);
nor U11121 (N_11121,N_10942,N_11016);
or U11122 (N_11122,N_10915,N_11098);
nand U11123 (N_11123,N_10970,N_11021);
or U11124 (N_11124,N_10881,N_10880);
nand U11125 (N_11125,N_10842,N_10906);
nand U11126 (N_11126,N_10926,N_10836);
nand U11127 (N_11127,N_10801,N_10810);
nor U11128 (N_11128,N_10847,N_10922);
and U11129 (N_11129,N_10832,N_11075);
nor U11130 (N_11130,N_11022,N_10844);
and U11131 (N_11131,N_10954,N_10934);
nor U11132 (N_11132,N_10945,N_10809);
and U11133 (N_11133,N_10867,N_10982);
nor U11134 (N_11134,N_10857,N_10833);
nor U11135 (N_11135,N_10897,N_11009);
nor U11136 (N_11136,N_10856,N_11093);
nor U11137 (N_11137,N_11092,N_11072);
or U11138 (N_11138,N_11034,N_11063);
nor U11139 (N_11139,N_11018,N_10913);
and U11140 (N_11140,N_11007,N_11053);
and U11141 (N_11141,N_11049,N_10840);
or U11142 (N_11142,N_11082,N_10925);
xnor U11143 (N_11143,N_10993,N_10886);
nand U11144 (N_11144,N_11046,N_10907);
xnor U11145 (N_11145,N_11028,N_10923);
nand U11146 (N_11146,N_10814,N_10931);
and U11147 (N_11147,N_11004,N_10861);
nor U11148 (N_11148,N_11074,N_11000);
or U11149 (N_11149,N_11064,N_10980);
and U11150 (N_11150,N_10888,N_10860);
or U11151 (N_11151,N_10892,N_11081);
nor U11152 (N_11152,N_11090,N_10914);
nor U11153 (N_11153,N_10966,N_10850);
xor U11154 (N_11154,N_10887,N_11045);
and U11155 (N_11155,N_11030,N_10994);
and U11156 (N_11156,N_10987,N_11070);
and U11157 (N_11157,N_10895,N_11083);
nor U11158 (N_11158,N_11040,N_11038);
nand U11159 (N_11159,N_11036,N_11023);
or U11160 (N_11160,N_10870,N_10885);
nand U11161 (N_11161,N_10998,N_11033);
nor U11162 (N_11162,N_10991,N_10979);
and U11163 (N_11163,N_10873,N_10841);
or U11164 (N_11164,N_10955,N_10855);
nor U11165 (N_11165,N_11008,N_10944);
and U11166 (N_11166,N_10992,N_10859);
xnor U11167 (N_11167,N_10977,N_11065);
nand U11168 (N_11168,N_10893,N_10806);
nor U11169 (N_11169,N_10986,N_10997);
nor U11170 (N_11170,N_10865,N_10968);
nor U11171 (N_11171,N_11060,N_10858);
and U11172 (N_11172,N_10808,N_10894);
nand U11173 (N_11173,N_11043,N_10930);
and U11174 (N_11174,N_10989,N_11071);
nand U11175 (N_11175,N_10825,N_10956);
xnor U11176 (N_11176,N_10990,N_10800);
nor U11177 (N_11177,N_11086,N_10898);
xor U11178 (N_11178,N_10843,N_10862);
nand U11179 (N_11179,N_10951,N_10837);
nand U11180 (N_11180,N_11062,N_11015);
nor U11181 (N_11181,N_11026,N_11044);
nand U11182 (N_11182,N_11094,N_10868);
xor U11183 (N_11183,N_10901,N_10973);
nor U11184 (N_11184,N_10950,N_10821);
or U11185 (N_11185,N_10811,N_10941);
nor U11186 (N_11186,N_10827,N_10984);
or U11187 (N_11187,N_10995,N_11088);
xnor U11188 (N_11188,N_10872,N_10902);
xor U11189 (N_11189,N_10804,N_10975);
and U11190 (N_11190,N_10957,N_11097);
xnor U11191 (N_11191,N_11056,N_10802);
or U11192 (N_11192,N_10932,N_10935);
xnor U11193 (N_11193,N_11017,N_10871);
nand U11194 (N_11194,N_10849,N_11002);
xor U11195 (N_11195,N_11067,N_11078);
xor U11196 (N_11196,N_10852,N_10826);
xnor U11197 (N_11197,N_10876,N_10835);
or U11198 (N_11198,N_10924,N_11050);
nand U11199 (N_11199,N_11091,N_10905);
nor U11200 (N_11200,N_10940,N_10952);
nor U11201 (N_11201,N_10877,N_11014);
nor U11202 (N_11202,N_11073,N_10936);
nor U11203 (N_11203,N_10999,N_11041);
and U11204 (N_11204,N_10829,N_10976);
nor U11205 (N_11205,N_10864,N_11006);
xor U11206 (N_11206,N_11077,N_11037);
and U11207 (N_11207,N_10912,N_10813);
nor U11208 (N_11208,N_10900,N_11087);
nor U11209 (N_11209,N_10818,N_10963);
nand U11210 (N_11210,N_10899,N_11058);
and U11211 (N_11211,N_11079,N_10816);
xor U11212 (N_11212,N_11011,N_10910);
and U11213 (N_11213,N_11013,N_11069);
nor U11214 (N_11214,N_10866,N_10882);
xnor U11215 (N_11215,N_11029,N_10890);
and U11216 (N_11216,N_10964,N_10838);
or U11217 (N_11217,N_10848,N_11057);
or U11218 (N_11218,N_10920,N_11001);
or U11219 (N_11219,N_10971,N_10946);
nor U11220 (N_11220,N_10822,N_10828);
nand U11221 (N_11221,N_10978,N_11084);
and U11222 (N_11222,N_11055,N_10943);
xnor U11223 (N_11223,N_10921,N_11025);
nand U11224 (N_11224,N_10947,N_10918);
or U11225 (N_11225,N_10878,N_11031);
or U11226 (N_11226,N_11010,N_10969);
nor U11227 (N_11227,N_11096,N_10927);
or U11228 (N_11228,N_10889,N_10928);
nor U11229 (N_11229,N_11012,N_11054);
xnor U11230 (N_11230,N_10883,N_10805);
or U11231 (N_11231,N_10879,N_10983);
and U11232 (N_11232,N_10909,N_10807);
nor U11233 (N_11233,N_10830,N_10845);
or U11234 (N_11234,N_10853,N_10948);
nor U11235 (N_11235,N_11095,N_11099);
nand U11236 (N_11236,N_10919,N_10959);
and U11237 (N_11237,N_10974,N_10834);
and U11238 (N_11238,N_11089,N_10958);
and U11239 (N_11239,N_10839,N_11048);
nand U11240 (N_11240,N_10854,N_10869);
or U11241 (N_11241,N_11047,N_10896);
or U11242 (N_11242,N_10846,N_10911);
and U11243 (N_11243,N_11051,N_10965);
nand U11244 (N_11244,N_11066,N_10875);
nor U11245 (N_11245,N_10904,N_10960);
or U11246 (N_11246,N_10938,N_11059);
xnor U11247 (N_11247,N_10824,N_11080);
nor U11248 (N_11248,N_10891,N_10949);
nor U11249 (N_11249,N_11024,N_10874);
xor U11250 (N_11250,N_10894,N_10973);
and U11251 (N_11251,N_10866,N_10898);
nand U11252 (N_11252,N_10884,N_10810);
xnor U11253 (N_11253,N_10879,N_11074);
nand U11254 (N_11254,N_10887,N_11040);
or U11255 (N_11255,N_10980,N_10944);
or U11256 (N_11256,N_10847,N_10842);
nand U11257 (N_11257,N_11074,N_10945);
nand U11258 (N_11258,N_11068,N_10841);
or U11259 (N_11259,N_10835,N_11041);
nor U11260 (N_11260,N_10947,N_10816);
and U11261 (N_11261,N_10870,N_10922);
nand U11262 (N_11262,N_10825,N_10850);
or U11263 (N_11263,N_11041,N_10932);
nand U11264 (N_11264,N_10942,N_10993);
xor U11265 (N_11265,N_10820,N_10827);
and U11266 (N_11266,N_10880,N_10969);
and U11267 (N_11267,N_11072,N_10893);
nor U11268 (N_11268,N_10801,N_10817);
and U11269 (N_11269,N_10964,N_10870);
nor U11270 (N_11270,N_11007,N_11058);
nand U11271 (N_11271,N_10912,N_10951);
or U11272 (N_11272,N_11093,N_10927);
or U11273 (N_11273,N_10863,N_11081);
or U11274 (N_11274,N_10922,N_10936);
and U11275 (N_11275,N_11097,N_10839);
nand U11276 (N_11276,N_10800,N_10817);
nor U11277 (N_11277,N_11091,N_10944);
or U11278 (N_11278,N_10868,N_10905);
or U11279 (N_11279,N_10889,N_11063);
nand U11280 (N_11280,N_11010,N_11030);
or U11281 (N_11281,N_10963,N_10834);
and U11282 (N_11282,N_10801,N_11056);
xor U11283 (N_11283,N_10805,N_11031);
and U11284 (N_11284,N_10804,N_11035);
and U11285 (N_11285,N_11017,N_10815);
nand U11286 (N_11286,N_10881,N_11096);
nand U11287 (N_11287,N_11009,N_10921);
and U11288 (N_11288,N_11085,N_11054);
nand U11289 (N_11289,N_10862,N_11062);
or U11290 (N_11290,N_10832,N_10950);
nand U11291 (N_11291,N_10982,N_10955);
xor U11292 (N_11292,N_10951,N_10918);
and U11293 (N_11293,N_10979,N_10929);
or U11294 (N_11294,N_10866,N_10981);
nand U11295 (N_11295,N_10818,N_10990);
nor U11296 (N_11296,N_10875,N_10824);
xnor U11297 (N_11297,N_11036,N_11038);
and U11298 (N_11298,N_10846,N_11071);
xnor U11299 (N_11299,N_10980,N_10908);
nor U11300 (N_11300,N_10903,N_10928);
and U11301 (N_11301,N_11078,N_10881);
xor U11302 (N_11302,N_10893,N_11033);
and U11303 (N_11303,N_10888,N_10850);
nand U11304 (N_11304,N_10996,N_11008);
nor U11305 (N_11305,N_10891,N_10873);
nand U11306 (N_11306,N_11009,N_11044);
or U11307 (N_11307,N_11033,N_10980);
nor U11308 (N_11308,N_11075,N_10972);
nor U11309 (N_11309,N_10970,N_11095);
and U11310 (N_11310,N_10816,N_10913);
xor U11311 (N_11311,N_10848,N_10879);
nor U11312 (N_11312,N_10936,N_11047);
nor U11313 (N_11313,N_10854,N_11097);
and U11314 (N_11314,N_10879,N_10820);
nor U11315 (N_11315,N_10989,N_11061);
xnor U11316 (N_11316,N_11087,N_10980);
and U11317 (N_11317,N_11063,N_10949);
or U11318 (N_11318,N_11009,N_10870);
or U11319 (N_11319,N_10955,N_11001);
or U11320 (N_11320,N_10836,N_10979);
nand U11321 (N_11321,N_10945,N_10922);
nand U11322 (N_11322,N_11030,N_11018);
nor U11323 (N_11323,N_11072,N_10860);
nand U11324 (N_11324,N_10883,N_10807);
and U11325 (N_11325,N_11014,N_10809);
and U11326 (N_11326,N_10863,N_11018);
or U11327 (N_11327,N_10845,N_11064);
and U11328 (N_11328,N_10867,N_10945);
xnor U11329 (N_11329,N_10883,N_10916);
nor U11330 (N_11330,N_10950,N_11078);
nor U11331 (N_11331,N_11034,N_10909);
xnor U11332 (N_11332,N_11067,N_10834);
and U11333 (N_11333,N_11047,N_11080);
or U11334 (N_11334,N_10809,N_11003);
nor U11335 (N_11335,N_10858,N_10851);
or U11336 (N_11336,N_10944,N_11034);
xnor U11337 (N_11337,N_10810,N_10825);
xor U11338 (N_11338,N_11007,N_10870);
nor U11339 (N_11339,N_10857,N_11085);
nor U11340 (N_11340,N_10933,N_11008);
xnor U11341 (N_11341,N_10913,N_11077);
xnor U11342 (N_11342,N_10850,N_10886);
nor U11343 (N_11343,N_11074,N_10894);
or U11344 (N_11344,N_11042,N_11079);
nand U11345 (N_11345,N_10913,N_10845);
xnor U11346 (N_11346,N_11071,N_10867);
or U11347 (N_11347,N_10969,N_10862);
and U11348 (N_11348,N_10877,N_10829);
and U11349 (N_11349,N_10873,N_10952);
and U11350 (N_11350,N_10815,N_10826);
or U11351 (N_11351,N_10911,N_10899);
or U11352 (N_11352,N_10916,N_10837);
nor U11353 (N_11353,N_10972,N_10848);
and U11354 (N_11354,N_11072,N_10867);
nor U11355 (N_11355,N_10952,N_11030);
and U11356 (N_11356,N_11013,N_10929);
and U11357 (N_11357,N_10802,N_10836);
nor U11358 (N_11358,N_11019,N_11046);
nor U11359 (N_11359,N_10964,N_10981);
nor U11360 (N_11360,N_10864,N_11021);
or U11361 (N_11361,N_10823,N_10847);
xor U11362 (N_11362,N_11045,N_10999);
xor U11363 (N_11363,N_10859,N_10833);
nand U11364 (N_11364,N_10943,N_10926);
and U11365 (N_11365,N_11011,N_10871);
and U11366 (N_11366,N_11085,N_10848);
or U11367 (N_11367,N_11066,N_11015);
or U11368 (N_11368,N_10850,N_10904);
or U11369 (N_11369,N_10858,N_10917);
nor U11370 (N_11370,N_10831,N_11001);
and U11371 (N_11371,N_10805,N_10956);
or U11372 (N_11372,N_11029,N_10895);
nand U11373 (N_11373,N_11040,N_10807);
and U11374 (N_11374,N_11025,N_10981);
or U11375 (N_11375,N_11079,N_10955);
xnor U11376 (N_11376,N_10972,N_10891);
or U11377 (N_11377,N_10990,N_11061);
nor U11378 (N_11378,N_11057,N_11088);
or U11379 (N_11379,N_10951,N_10910);
or U11380 (N_11380,N_10970,N_10817);
and U11381 (N_11381,N_11033,N_11040);
or U11382 (N_11382,N_11028,N_10979);
nand U11383 (N_11383,N_10979,N_10985);
and U11384 (N_11384,N_10898,N_10877);
nor U11385 (N_11385,N_11010,N_10985);
nand U11386 (N_11386,N_10867,N_11067);
or U11387 (N_11387,N_10989,N_10847);
nand U11388 (N_11388,N_10849,N_10947);
nor U11389 (N_11389,N_10878,N_11022);
or U11390 (N_11390,N_10852,N_10937);
nor U11391 (N_11391,N_10910,N_10950);
and U11392 (N_11392,N_10823,N_10920);
nand U11393 (N_11393,N_10971,N_10959);
xnor U11394 (N_11394,N_10867,N_11034);
or U11395 (N_11395,N_11046,N_10959);
and U11396 (N_11396,N_10963,N_11023);
xnor U11397 (N_11397,N_10912,N_10937);
and U11398 (N_11398,N_11077,N_11038);
and U11399 (N_11399,N_10943,N_11076);
xnor U11400 (N_11400,N_11185,N_11171);
and U11401 (N_11401,N_11356,N_11186);
nor U11402 (N_11402,N_11313,N_11328);
xnor U11403 (N_11403,N_11170,N_11224);
nor U11404 (N_11404,N_11152,N_11271);
nand U11405 (N_11405,N_11108,N_11383);
or U11406 (N_11406,N_11306,N_11105);
and U11407 (N_11407,N_11123,N_11348);
nor U11408 (N_11408,N_11134,N_11245);
and U11409 (N_11409,N_11110,N_11154);
nand U11410 (N_11410,N_11203,N_11228);
nor U11411 (N_11411,N_11133,N_11270);
nor U11412 (N_11412,N_11158,N_11294);
nand U11413 (N_11413,N_11194,N_11213);
or U11414 (N_11414,N_11309,N_11126);
nand U11415 (N_11415,N_11188,N_11243);
nand U11416 (N_11416,N_11218,N_11274);
or U11417 (N_11417,N_11260,N_11304);
and U11418 (N_11418,N_11236,N_11193);
nor U11419 (N_11419,N_11192,N_11241);
nand U11420 (N_11420,N_11148,N_11317);
nor U11421 (N_11421,N_11181,N_11381);
nor U11422 (N_11422,N_11139,N_11182);
xor U11423 (N_11423,N_11297,N_11262);
nor U11424 (N_11424,N_11337,N_11330);
or U11425 (N_11425,N_11321,N_11265);
xor U11426 (N_11426,N_11173,N_11372);
and U11427 (N_11427,N_11232,N_11142);
or U11428 (N_11428,N_11353,N_11167);
xnor U11429 (N_11429,N_11131,N_11362);
nor U11430 (N_11430,N_11174,N_11157);
xor U11431 (N_11431,N_11264,N_11135);
nor U11432 (N_11432,N_11367,N_11275);
and U11433 (N_11433,N_11258,N_11128);
nor U11434 (N_11434,N_11252,N_11384);
xnor U11435 (N_11435,N_11333,N_11375);
nor U11436 (N_11436,N_11263,N_11206);
nand U11437 (N_11437,N_11240,N_11360);
nand U11438 (N_11438,N_11251,N_11341);
xor U11439 (N_11439,N_11197,N_11310);
or U11440 (N_11440,N_11136,N_11298);
nand U11441 (N_11441,N_11184,N_11222);
or U11442 (N_11442,N_11201,N_11121);
nor U11443 (N_11443,N_11389,N_11172);
xnor U11444 (N_11444,N_11103,N_11278);
nor U11445 (N_11445,N_11180,N_11279);
xnor U11446 (N_11446,N_11215,N_11102);
nand U11447 (N_11447,N_11351,N_11354);
nor U11448 (N_11448,N_11364,N_11178);
or U11449 (N_11449,N_11151,N_11376);
nor U11450 (N_11450,N_11221,N_11334);
and U11451 (N_11451,N_11371,N_11144);
and U11452 (N_11452,N_11100,N_11385);
nor U11453 (N_11453,N_11155,N_11244);
and U11454 (N_11454,N_11207,N_11387);
nand U11455 (N_11455,N_11250,N_11390);
or U11456 (N_11456,N_11303,N_11374);
nor U11457 (N_11457,N_11106,N_11233);
xnor U11458 (N_11458,N_11277,N_11209);
and U11459 (N_11459,N_11322,N_11166);
or U11460 (N_11460,N_11269,N_11220);
xor U11461 (N_11461,N_11146,N_11379);
and U11462 (N_11462,N_11225,N_11299);
nand U11463 (N_11463,N_11268,N_11204);
nor U11464 (N_11464,N_11287,N_11141);
or U11465 (N_11465,N_11281,N_11346);
nand U11466 (N_11466,N_11234,N_11125);
xor U11467 (N_11467,N_11153,N_11257);
and U11468 (N_11468,N_11329,N_11202);
xor U11469 (N_11469,N_11179,N_11111);
and U11470 (N_11470,N_11326,N_11124);
xnor U11471 (N_11471,N_11164,N_11340);
nand U11472 (N_11472,N_11261,N_11301);
or U11473 (N_11473,N_11284,N_11331);
xor U11474 (N_11474,N_11104,N_11377);
xnor U11475 (N_11475,N_11120,N_11343);
and U11476 (N_11476,N_11370,N_11266);
nor U11477 (N_11477,N_11117,N_11116);
or U11478 (N_11478,N_11373,N_11237);
and U11479 (N_11479,N_11357,N_11249);
nand U11480 (N_11480,N_11253,N_11363);
nand U11481 (N_11481,N_11160,N_11352);
xor U11482 (N_11482,N_11259,N_11292);
nor U11483 (N_11483,N_11288,N_11312);
xor U11484 (N_11484,N_11189,N_11359);
or U11485 (N_11485,N_11183,N_11311);
nor U11486 (N_11486,N_11314,N_11210);
or U11487 (N_11487,N_11280,N_11332);
nor U11488 (N_11488,N_11190,N_11238);
and U11489 (N_11489,N_11256,N_11229);
nand U11490 (N_11490,N_11365,N_11386);
and U11491 (N_11491,N_11289,N_11199);
and U11492 (N_11492,N_11368,N_11395);
nor U11493 (N_11493,N_11388,N_11338);
nor U11494 (N_11494,N_11114,N_11198);
xnor U11495 (N_11495,N_11196,N_11187);
xnor U11496 (N_11496,N_11195,N_11235);
or U11497 (N_11497,N_11169,N_11137);
nor U11498 (N_11498,N_11254,N_11216);
xor U11499 (N_11499,N_11378,N_11226);
nor U11500 (N_11500,N_11349,N_11350);
and U11501 (N_11501,N_11319,N_11159);
and U11502 (N_11502,N_11130,N_11286);
and U11503 (N_11503,N_11361,N_11272);
xnor U11504 (N_11504,N_11344,N_11122);
and U11505 (N_11505,N_11211,N_11369);
xnor U11506 (N_11506,N_11382,N_11161);
or U11507 (N_11507,N_11366,N_11293);
nor U11508 (N_11508,N_11140,N_11101);
or U11509 (N_11509,N_11247,N_11230);
or U11510 (N_11510,N_11318,N_11308);
xor U11511 (N_11511,N_11165,N_11118);
and U11512 (N_11512,N_11119,N_11168);
xnor U11513 (N_11513,N_11358,N_11282);
nand U11514 (N_11514,N_11143,N_11342);
nand U11515 (N_11515,N_11325,N_11212);
or U11516 (N_11516,N_11394,N_11315);
nor U11517 (N_11517,N_11392,N_11112);
or U11518 (N_11518,N_11231,N_11276);
nor U11519 (N_11519,N_11296,N_11335);
xnor U11520 (N_11520,N_11156,N_11107);
xnor U11521 (N_11521,N_11327,N_11205);
nor U11522 (N_11522,N_11132,N_11217);
or U11523 (N_11523,N_11295,N_11399);
nand U11524 (N_11524,N_11176,N_11145);
nor U11525 (N_11525,N_11175,N_11291);
and U11526 (N_11526,N_11191,N_11113);
or U11527 (N_11527,N_11115,N_11177);
nand U11528 (N_11528,N_11208,N_11147);
nand U11529 (N_11529,N_11290,N_11391);
or U11530 (N_11530,N_11302,N_11355);
xor U11531 (N_11531,N_11339,N_11149);
or U11532 (N_11532,N_11345,N_11163);
nand U11533 (N_11533,N_11324,N_11129);
nor U11534 (N_11534,N_11347,N_11200);
xnor U11535 (N_11535,N_11380,N_11393);
or U11536 (N_11536,N_11283,N_11138);
and U11537 (N_11537,N_11307,N_11336);
and U11538 (N_11538,N_11246,N_11320);
xnor U11539 (N_11539,N_11109,N_11162);
or U11540 (N_11540,N_11273,N_11397);
nand U11541 (N_11541,N_11255,N_11127);
nor U11542 (N_11542,N_11300,N_11239);
or U11543 (N_11543,N_11398,N_11323);
and U11544 (N_11544,N_11150,N_11227);
xor U11545 (N_11545,N_11285,N_11396);
nor U11546 (N_11546,N_11305,N_11267);
or U11547 (N_11547,N_11248,N_11242);
xor U11548 (N_11548,N_11214,N_11223);
xor U11549 (N_11549,N_11219,N_11316);
nand U11550 (N_11550,N_11261,N_11270);
nor U11551 (N_11551,N_11192,N_11230);
or U11552 (N_11552,N_11189,N_11233);
nand U11553 (N_11553,N_11156,N_11201);
nand U11554 (N_11554,N_11214,N_11102);
and U11555 (N_11555,N_11159,N_11324);
nand U11556 (N_11556,N_11224,N_11146);
nor U11557 (N_11557,N_11261,N_11155);
xnor U11558 (N_11558,N_11279,N_11340);
nor U11559 (N_11559,N_11200,N_11343);
xnor U11560 (N_11560,N_11164,N_11324);
nor U11561 (N_11561,N_11171,N_11395);
or U11562 (N_11562,N_11148,N_11228);
or U11563 (N_11563,N_11322,N_11190);
nor U11564 (N_11564,N_11219,N_11145);
and U11565 (N_11565,N_11174,N_11219);
nand U11566 (N_11566,N_11227,N_11195);
xor U11567 (N_11567,N_11342,N_11230);
or U11568 (N_11568,N_11146,N_11341);
nor U11569 (N_11569,N_11110,N_11325);
nor U11570 (N_11570,N_11354,N_11275);
or U11571 (N_11571,N_11196,N_11327);
or U11572 (N_11572,N_11215,N_11362);
xor U11573 (N_11573,N_11270,N_11343);
nor U11574 (N_11574,N_11307,N_11136);
nor U11575 (N_11575,N_11108,N_11260);
nor U11576 (N_11576,N_11363,N_11272);
nand U11577 (N_11577,N_11203,N_11281);
xnor U11578 (N_11578,N_11189,N_11263);
nor U11579 (N_11579,N_11142,N_11341);
nor U11580 (N_11580,N_11147,N_11327);
nand U11581 (N_11581,N_11334,N_11202);
and U11582 (N_11582,N_11150,N_11317);
xor U11583 (N_11583,N_11138,N_11125);
and U11584 (N_11584,N_11301,N_11292);
nor U11585 (N_11585,N_11162,N_11343);
nand U11586 (N_11586,N_11387,N_11216);
or U11587 (N_11587,N_11187,N_11382);
xor U11588 (N_11588,N_11329,N_11353);
and U11589 (N_11589,N_11201,N_11329);
nand U11590 (N_11590,N_11347,N_11362);
nand U11591 (N_11591,N_11230,N_11293);
nor U11592 (N_11592,N_11179,N_11370);
or U11593 (N_11593,N_11301,N_11363);
and U11594 (N_11594,N_11333,N_11239);
or U11595 (N_11595,N_11372,N_11184);
xor U11596 (N_11596,N_11216,N_11381);
nand U11597 (N_11597,N_11192,N_11116);
nand U11598 (N_11598,N_11216,N_11282);
nor U11599 (N_11599,N_11123,N_11323);
xor U11600 (N_11600,N_11209,N_11297);
xnor U11601 (N_11601,N_11392,N_11395);
xnor U11602 (N_11602,N_11130,N_11325);
xnor U11603 (N_11603,N_11378,N_11161);
xor U11604 (N_11604,N_11313,N_11144);
or U11605 (N_11605,N_11153,N_11314);
nor U11606 (N_11606,N_11361,N_11356);
nor U11607 (N_11607,N_11155,N_11229);
nor U11608 (N_11608,N_11240,N_11128);
and U11609 (N_11609,N_11122,N_11325);
and U11610 (N_11610,N_11287,N_11397);
nor U11611 (N_11611,N_11201,N_11107);
or U11612 (N_11612,N_11264,N_11180);
xnor U11613 (N_11613,N_11183,N_11376);
nor U11614 (N_11614,N_11167,N_11121);
and U11615 (N_11615,N_11113,N_11213);
xnor U11616 (N_11616,N_11290,N_11139);
xnor U11617 (N_11617,N_11246,N_11219);
or U11618 (N_11618,N_11141,N_11303);
and U11619 (N_11619,N_11149,N_11146);
xnor U11620 (N_11620,N_11310,N_11386);
nand U11621 (N_11621,N_11217,N_11343);
and U11622 (N_11622,N_11338,N_11387);
or U11623 (N_11623,N_11162,N_11165);
or U11624 (N_11624,N_11262,N_11180);
nor U11625 (N_11625,N_11330,N_11169);
nand U11626 (N_11626,N_11228,N_11128);
xor U11627 (N_11627,N_11102,N_11210);
nand U11628 (N_11628,N_11285,N_11349);
or U11629 (N_11629,N_11243,N_11121);
or U11630 (N_11630,N_11161,N_11389);
xor U11631 (N_11631,N_11251,N_11220);
and U11632 (N_11632,N_11343,N_11293);
xnor U11633 (N_11633,N_11185,N_11190);
nor U11634 (N_11634,N_11166,N_11280);
and U11635 (N_11635,N_11326,N_11267);
or U11636 (N_11636,N_11136,N_11266);
and U11637 (N_11637,N_11206,N_11230);
xnor U11638 (N_11638,N_11229,N_11304);
nor U11639 (N_11639,N_11109,N_11140);
nand U11640 (N_11640,N_11220,N_11113);
nand U11641 (N_11641,N_11347,N_11306);
or U11642 (N_11642,N_11356,N_11355);
nand U11643 (N_11643,N_11231,N_11364);
and U11644 (N_11644,N_11310,N_11385);
xor U11645 (N_11645,N_11342,N_11275);
or U11646 (N_11646,N_11390,N_11245);
nand U11647 (N_11647,N_11341,N_11277);
nand U11648 (N_11648,N_11171,N_11327);
xor U11649 (N_11649,N_11351,N_11217);
nand U11650 (N_11650,N_11310,N_11323);
nor U11651 (N_11651,N_11351,N_11221);
nand U11652 (N_11652,N_11392,N_11319);
nor U11653 (N_11653,N_11347,N_11330);
and U11654 (N_11654,N_11169,N_11295);
nor U11655 (N_11655,N_11186,N_11326);
or U11656 (N_11656,N_11254,N_11152);
nand U11657 (N_11657,N_11388,N_11309);
xor U11658 (N_11658,N_11105,N_11358);
or U11659 (N_11659,N_11397,N_11166);
and U11660 (N_11660,N_11285,N_11206);
nor U11661 (N_11661,N_11110,N_11346);
xnor U11662 (N_11662,N_11240,N_11148);
xor U11663 (N_11663,N_11101,N_11344);
nand U11664 (N_11664,N_11344,N_11136);
or U11665 (N_11665,N_11303,N_11248);
nor U11666 (N_11666,N_11389,N_11210);
nor U11667 (N_11667,N_11340,N_11182);
or U11668 (N_11668,N_11226,N_11199);
nor U11669 (N_11669,N_11303,N_11277);
or U11670 (N_11670,N_11103,N_11359);
and U11671 (N_11671,N_11105,N_11326);
nor U11672 (N_11672,N_11275,N_11183);
nand U11673 (N_11673,N_11342,N_11155);
xor U11674 (N_11674,N_11391,N_11366);
nor U11675 (N_11675,N_11138,N_11186);
xnor U11676 (N_11676,N_11227,N_11155);
nor U11677 (N_11677,N_11203,N_11100);
and U11678 (N_11678,N_11230,N_11259);
xor U11679 (N_11679,N_11191,N_11220);
nand U11680 (N_11680,N_11197,N_11204);
and U11681 (N_11681,N_11188,N_11295);
nor U11682 (N_11682,N_11156,N_11135);
nor U11683 (N_11683,N_11298,N_11300);
or U11684 (N_11684,N_11187,N_11316);
nor U11685 (N_11685,N_11162,N_11268);
xnor U11686 (N_11686,N_11177,N_11359);
and U11687 (N_11687,N_11121,N_11213);
and U11688 (N_11688,N_11228,N_11323);
and U11689 (N_11689,N_11365,N_11308);
nand U11690 (N_11690,N_11390,N_11157);
nand U11691 (N_11691,N_11116,N_11316);
nor U11692 (N_11692,N_11398,N_11273);
or U11693 (N_11693,N_11171,N_11250);
xor U11694 (N_11694,N_11329,N_11151);
nand U11695 (N_11695,N_11390,N_11243);
nand U11696 (N_11696,N_11265,N_11315);
xor U11697 (N_11697,N_11300,N_11345);
nand U11698 (N_11698,N_11310,N_11387);
nand U11699 (N_11699,N_11102,N_11197);
xnor U11700 (N_11700,N_11642,N_11648);
and U11701 (N_11701,N_11469,N_11413);
and U11702 (N_11702,N_11529,N_11617);
nor U11703 (N_11703,N_11549,N_11645);
nand U11704 (N_11704,N_11504,N_11538);
or U11705 (N_11705,N_11521,N_11672);
nand U11706 (N_11706,N_11455,N_11693);
nor U11707 (N_11707,N_11593,N_11687);
or U11708 (N_11708,N_11561,N_11406);
nand U11709 (N_11709,N_11546,N_11475);
nand U11710 (N_11710,N_11472,N_11582);
or U11711 (N_11711,N_11612,N_11614);
xnor U11712 (N_11712,N_11500,N_11516);
xnor U11713 (N_11713,N_11497,N_11664);
nand U11714 (N_11714,N_11487,N_11608);
nor U11715 (N_11715,N_11429,N_11552);
and U11716 (N_11716,N_11410,N_11501);
nor U11717 (N_11717,N_11692,N_11613);
xnor U11718 (N_11718,N_11668,N_11584);
xor U11719 (N_11719,N_11626,N_11451);
xor U11720 (N_11720,N_11467,N_11559);
and U11721 (N_11721,N_11573,N_11481);
nand U11722 (N_11722,N_11685,N_11462);
nand U11723 (N_11723,N_11667,N_11418);
nor U11724 (N_11724,N_11651,N_11426);
and U11725 (N_11725,N_11615,N_11661);
xnor U11726 (N_11726,N_11646,N_11464);
nand U11727 (N_11727,N_11486,N_11545);
xor U11728 (N_11728,N_11641,N_11402);
nand U11729 (N_11729,N_11473,N_11405);
xnor U11730 (N_11730,N_11601,N_11659);
nor U11731 (N_11731,N_11490,N_11586);
or U11732 (N_11732,N_11630,N_11621);
or U11733 (N_11733,N_11689,N_11499);
nand U11734 (N_11734,N_11677,N_11430);
xor U11735 (N_11735,N_11474,N_11530);
xor U11736 (N_11736,N_11511,N_11673);
nand U11737 (N_11737,N_11539,N_11638);
xnor U11738 (N_11738,N_11698,N_11512);
nand U11739 (N_11739,N_11611,N_11407);
nand U11740 (N_11740,N_11409,N_11571);
or U11741 (N_11741,N_11569,N_11565);
and U11742 (N_11742,N_11604,N_11543);
and U11743 (N_11743,N_11619,N_11631);
nand U11744 (N_11744,N_11653,N_11633);
or U11745 (N_11745,N_11566,N_11400);
or U11746 (N_11746,N_11595,N_11610);
or U11747 (N_11747,N_11544,N_11656);
nand U11748 (N_11748,N_11507,N_11477);
and U11749 (N_11749,N_11463,N_11423);
nand U11750 (N_11750,N_11449,N_11435);
nand U11751 (N_11751,N_11562,N_11597);
xnor U11752 (N_11752,N_11457,N_11520);
nor U11753 (N_11753,N_11515,N_11574);
xor U11754 (N_11754,N_11422,N_11417);
xnor U11755 (N_11755,N_11583,N_11527);
nand U11756 (N_11756,N_11678,N_11632);
and U11757 (N_11757,N_11528,N_11686);
nor U11758 (N_11758,N_11421,N_11438);
nand U11759 (N_11759,N_11534,N_11436);
nor U11760 (N_11760,N_11437,N_11403);
xor U11761 (N_11761,N_11498,N_11551);
and U11762 (N_11762,N_11697,N_11695);
and U11763 (N_11763,N_11665,N_11494);
nor U11764 (N_11764,N_11588,N_11542);
or U11765 (N_11765,N_11624,N_11427);
and U11766 (N_11766,N_11627,N_11669);
and U11767 (N_11767,N_11446,N_11629);
or U11768 (N_11768,N_11658,N_11680);
xnor U11769 (N_11769,N_11514,N_11452);
or U11770 (N_11770,N_11460,N_11666);
or U11771 (N_11771,N_11591,N_11688);
nand U11772 (N_11772,N_11594,N_11547);
nand U11773 (N_11773,N_11576,N_11606);
and U11774 (N_11774,N_11570,N_11442);
or U11775 (N_11775,N_11690,N_11699);
nor U11776 (N_11776,N_11478,N_11683);
nor U11777 (N_11777,N_11408,N_11577);
xor U11778 (N_11778,N_11556,N_11523);
and U11779 (N_11779,N_11639,N_11696);
nand U11780 (N_11780,N_11517,N_11640);
nor U11781 (N_11781,N_11411,N_11505);
or U11782 (N_11782,N_11404,N_11550);
nor U11783 (N_11783,N_11649,N_11628);
or U11784 (N_11784,N_11682,N_11532);
xor U11785 (N_11785,N_11420,N_11623);
nand U11786 (N_11786,N_11605,N_11581);
or U11787 (N_11787,N_11691,N_11483);
and U11788 (N_11788,N_11489,N_11684);
nand U11789 (N_11789,N_11454,N_11479);
nor U11790 (N_11790,N_11518,N_11548);
and U11791 (N_11791,N_11654,N_11599);
nor U11792 (N_11792,N_11480,N_11424);
nand U11793 (N_11793,N_11652,N_11671);
and U11794 (N_11794,N_11589,N_11635);
nor U11795 (N_11795,N_11575,N_11655);
xor U11796 (N_11796,N_11524,N_11443);
nand U11797 (N_11797,N_11564,N_11603);
nor U11798 (N_11798,N_11681,N_11647);
xor U11799 (N_11799,N_11488,N_11441);
and U11800 (N_11800,N_11419,N_11513);
nand U11801 (N_11801,N_11596,N_11468);
or U11802 (N_11802,N_11412,N_11445);
xnor U11803 (N_11803,N_11465,N_11414);
nor U11804 (N_11804,N_11509,N_11416);
xnor U11805 (N_11805,N_11496,N_11526);
and U11806 (N_11806,N_11415,N_11458);
or U11807 (N_11807,N_11470,N_11440);
xnor U11808 (N_11808,N_11522,N_11568);
nand U11809 (N_11809,N_11491,N_11448);
nand U11810 (N_11810,N_11634,N_11502);
and U11811 (N_11811,N_11618,N_11670);
xor U11812 (N_11812,N_11622,N_11482);
xnor U11813 (N_11813,N_11637,N_11592);
xnor U11814 (N_11814,N_11555,N_11531);
nand U11815 (N_11815,N_11456,N_11663);
or U11816 (N_11816,N_11428,N_11434);
or U11817 (N_11817,N_11662,N_11537);
nand U11818 (N_11818,N_11439,N_11536);
nand U11819 (N_11819,N_11540,N_11471);
nor U11820 (N_11820,N_11650,N_11554);
xnor U11821 (N_11821,N_11625,N_11484);
and U11822 (N_11822,N_11510,N_11572);
nor U11823 (N_11823,N_11508,N_11620);
and U11824 (N_11824,N_11425,N_11607);
xnor U11825 (N_11825,N_11675,N_11679);
or U11826 (N_11826,N_11590,N_11525);
nor U11827 (N_11827,N_11558,N_11461);
xnor U11828 (N_11828,N_11466,N_11495);
nor U11829 (N_11829,N_11578,N_11657);
nand U11830 (N_11830,N_11444,N_11447);
or U11831 (N_11831,N_11432,N_11616);
or U11832 (N_11832,N_11602,N_11560);
xnor U11833 (N_11833,N_11694,N_11476);
nand U11834 (N_11834,N_11587,N_11563);
and U11835 (N_11835,N_11485,N_11506);
nand U11836 (N_11836,N_11636,N_11676);
nor U11837 (N_11837,N_11533,N_11453);
nor U11838 (N_11838,N_11557,N_11433);
nand U11839 (N_11839,N_11643,N_11459);
nor U11840 (N_11840,N_11660,N_11644);
and U11841 (N_11841,N_11598,N_11553);
nor U11842 (N_11842,N_11535,N_11600);
nor U11843 (N_11843,N_11492,N_11567);
and U11844 (N_11844,N_11450,N_11579);
nand U11845 (N_11845,N_11674,N_11503);
and U11846 (N_11846,N_11580,N_11541);
nand U11847 (N_11847,N_11493,N_11401);
nor U11848 (N_11848,N_11431,N_11519);
and U11849 (N_11849,N_11609,N_11585);
or U11850 (N_11850,N_11423,N_11694);
nand U11851 (N_11851,N_11485,N_11404);
nor U11852 (N_11852,N_11479,N_11616);
and U11853 (N_11853,N_11604,N_11461);
nor U11854 (N_11854,N_11479,N_11453);
nand U11855 (N_11855,N_11467,N_11402);
xnor U11856 (N_11856,N_11678,N_11542);
xor U11857 (N_11857,N_11430,N_11621);
xnor U11858 (N_11858,N_11514,N_11564);
and U11859 (N_11859,N_11611,N_11536);
and U11860 (N_11860,N_11682,N_11555);
nor U11861 (N_11861,N_11617,N_11592);
and U11862 (N_11862,N_11676,N_11581);
or U11863 (N_11863,N_11616,N_11699);
xnor U11864 (N_11864,N_11680,N_11471);
nor U11865 (N_11865,N_11411,N_11690);
or U11866 (N_11866,N_11483,N_11430);
nand U11867 (N_11867,N_11433,N_11529);
nand U11868 (N_11868,N_11559,N_11437);
nor U11869 (N_11869,N_11479,N_11669);
xnor U11870 (N_11870,N_11535,N_11408);
nor U11871 (N_11871,N_11519,N_11420);
nor U11872 (N_11872,N_11405,N_11493);
or U11873 (N_11873,N_11560,N_11633);
nand U11874 (N_11874,N_11600,N_11422);
nand U11875 (N_11875,N_11624,N_11640);
or U11876 (N_11876,N_11666,N_11570);
nand U11877 (N_11877,N_11438,N_11454);
nor U11878 (N_11878,N_11458,N_11424);
or U11879 (N_11879,N_11646,N_11638);
nor U11880 (N_11880,N_11535,N_11654);
or U11881 (N_11881,N_11546,N_11656);
nand U11882 (N_11882,N_11585,N_11639);
and U11883 (N_11883,N_11601,N_11536);
or U11884 (N_11884,N_11497,N_11598);
nor U11885 (N_11885,N_11505,N_11410);
and U11886 (N_11886,N_11474,N_11426);
or U11887 (N_11887,N_11458,N_11679);
nor U11888 (N_11888,N_11656,N_11682);
nor U11889 (N_11889,N_11632,N_11681);
xor U11890 (N_11890,N_11530,N_11585);
and U11891 (N_11891,N_11607,N_11688);
nor U11892 (N_11892,N_11510,N_11616);
or U11893 (N_11893,N_11540,N_11572);
xor U11894 (N_11894,N_11532,N_11436);
nand U11895 (N_11895,N_11475,N_11649);
xor U11896 (N_11896,N_11693,N_11526);
or U11897 (N_11897,N_11656,N_11687);
nor U11898 (N_11898,N_11555,N_11489);
or U11899 (N_11899,N_11522,N_11689);
and U11900 (N_11900,N_11488,N_11668);
nand U11901 (N_11901,N_11618,N_11557);
xor U11902 (N_11902,N_11447,N_11524);
xor U11903 (N_11903,N_11462,N_11528);
and U11904 (N_11904,N_11408,N_11449);
xor U11905 (N_11905,N_11451,N_11438);
nand U11906 (N_11906,N_11620,N_11522);
nand U11907 (N_11907,N_11425,N_11612);
and U11908 (N_11908,N_11593,N_11640);
nand U11909 (N_11909,N_11664,N_11641);
or U11910 (N_11910,N_11660,N_11649);
and U11911 (N_11911,N_11416,N_11510);
nand U11912 (N_11912,N_11524,N_11572);
nand U11913 (N_11913,N_11667,N_11498);
and U11914 (N_11914,N_11516,N_11532);
xor U11915 (N_11915,N_11551,N_11605);
xnor U11916 (N_11916,N_11583,N_11425);
or U11917 (N_11917,N_11650,N_11528);
and U11918 (N_11918,N_11422,N_11406);
and U11919 (N_11919,N_11560,N_11559);
xnor U11920 (N_11920,N_11654,N_11526);
or U11921 (N_11921,N_11528,N_11632);
xnor U11922 (N_11922,N_11694,N_11624);
nand U11923 (N_11923,N_11462,N_11574);
xnor U11924 (N_11924,N_11577,N_11421);
and U11925 (N_11925,N_11516,N_11544);
xor U11926 (N_11926,N_11449,N_11533);
nor U11927 (N_11927,N_11672,N_11474);
xnor U11928 (N_11928,N_11494,N_11406);
or U11929 (N_11929,N_11606,N_11452);
nor U11930 (N_11930,N_11501,N_11597);
and U11931 (N_11931,N_11537,N_11437);
and U11932 (N_11932,N_11497,N_11486);
xor U11933 (N_11933,N_11406,N_11633);
xor U11934 (N_11934,N_11484,N_11572);
or U11935 (N_11935,N_11418,N_11658);
nand U11936 (N_11936,N_11453,N_11641);
and U11937 (N_11937,N_11642,N_11624);
or U11938 (N_11938,N_11693,N_11411);
or U11939 (N_11939,N_11401,N_11402);
and U11940 (N_11940,N_11472,N_11665);
nor U11941 (N_11941,N_11506,N_11681);
and U11942 (N_11942,N_11660,N_11516);
xnor U11943 (N_11943,N_11526,N_11481);
xor U11944 (N_11944,N_11465,N_11451);
and U11945 (N_11945,N_11574,N_11586);
or U11946 (N_11946,N_11568,N_11533);
nand U11947 (N_11947,N_11459,N_11692);
nand U11948 (N_11948,N_11608,N_11685);
or U11949 (N_11949,N_11449,N_11578);
and U11950 (N_11950,N_11520,N_11577);
and U11951 (N_11951,N_11415,N_11593);
xnor U11952 (N_11952,N_11450,N_11649);
xor U11953 (N_11953,N_11629,N_11671);
or U11954 (N_11954,N_11557,N_11431);
xnor U11955 (N_11955,N_11633,N_11417);
or U11956 (N_11956,N_11645,N_11498);
xnor U11957 (N_11957,N_11549,N_11621);
or U11958 (N_11958,N_11503,N_11619);
xor U11959 (N_11959,N_11424,N_11407);
and U11960 (N_11960,N_11631,N_11406);
nand U11961 (N_11961,N_11487,N_11647);
xor U11962 (N_11962,N_11616,N_11576);
or U11963 (N_11963,N_11591,N_11538);
nand U11964 (N_11964,N_11509,N_11472);
xor U11965 (N_11965,N_11425,N_11454);
and U11966 (N_11966,N_11576,N_11670);
or U11967 (N_11967,N_11608,N_11643);
xnor U11968 (N_11968,N_11643,N_11465);
nand U11969 (N_11969,N_11514,N_11419);
and U11970 (N_11970,N_11445,N_11535);
and U11971 (N_11971,N_11414,N_11674);
nor U11972 (N_11972,N_11682,N_11408);
xor U11973 (N_11973,N_11665,N_11633);
nor U11974 (N_11974,N_11469,N_11432);
nor U11975 (N_11975,N_11537,N_11687);
nor U11976 (N_11976,N_11646,N_11444);
xnor U11977 (N_11977,N_11423,N_11574);
nor U11978 (N_11978,N_11638,N_11634);
and U11979 (N_11979,N_11518,N_11509);
xor U11980 (N_11980,N_11596,N_11661);
xnor U11981 (N_11981,N_11485,N_11573);
nor U11982 (N_11982,N_11465,N_11680);
xnor U11983 (N_11983,N_11613,N_11595);
nand U11984 (N_11984,N_11523,N_11670);
and U11985 (N_11985,N_11507,N_11626);
xnor U11986 (N_11986,N_11461,N_11638);
xnor U11987 (N_11987,N_11531,N_11438);
nand U11988 (N_11988,N_11510,N_11428);
and U11989 (N_11989,N_11609,N_11548);
and U11990 (N_11990,N_11456,N_11499);
or U11991 (N_11991,N_11670,N_11450);
or U11992 (N_11992,N_11486,N_11595);
nand U11993 (N_11993,N_11427,N_11537);
nor U11994 (N_11994,N_11662,N_11519);
nor U11995 (N_11995,N_11643,N_11633);
nand U11996 (N_11996,N_11602,N_11679);
nand U11997 (N_11997,N_11622,N_11433);
nand U11998 (N_11998,N_11473,N_11542);
nor U11999 (N_11999,N_11421,N_11589);
nand U12000 (N_12000,N_11840,N_11748);
or U12001 (N_12001,N_11972,N_11985);
nor U12002 (N_12002,N_11796,N_11821);
or U12003 (N_12003,N_11783,N_11953);
or U12004 (N_12004,N_11815,N_11722);
nand U12005 (N_12005,N_11829,N_11827);
and U12006 (N_12006,N_11775,N_11993);
xnor U12007 (N_12007,N_11798,N_11915);
nor U12008 (N_12008,N_11854,N_11744);
xnor U12009 (N_12009,N_11835,N_11992);
xor U12010 (N_12010,N_11776,N_11864);
and U12011 (N_12011,N_11949,N_11974);
nor U12012 (N_12012,N_11879,N_11961);
xnor U12013 (N_12013,N_11936,N_11842);
or U12014 (N_12014,N_11717,N_11981);
and U12015 (N_12015,N_11782,N_11742);
xor U12016 (N_12016,N_11866,N_11923);
nand U12017 (N_12017,N_11794,N_11767);
and U12018 (N_12018,N_11705,N_11955);
xnor U12019 (N_12019,N_11839,N_11817);
and U12020 (N_12020,N_11807,N_11982);
or U12021 (N_12021,N_11917,N_11819);
or U12022 (N_12022,N_11938,N_11797);
or U12023 (N_12023,N_11712,N_11701);
nand U12024 (N_12024,N_11778,N_11940);
nand U12025 (N_12025,N_11905,N_11820);
xnor U12026 (N_12026,N_11838,N_11723);
or U12027 (N_12027,N_11979,N_11777);
xnor U12028 (N_12028,N_11709,N_11929);
xor U12029 (N_12029,N_11735,N_11912);
or U12030 (N_12030,N_11920,N_11870);
or U12031 (N_12031,N_11728,N_11769);
nor U12032 (N_12032,N_11909,N_11884);
or U12033 (N_12033,N_11889,N_11947);
nor U12034 (N_12034,N_11881,N_11813);
nor U12035 (N_12035,N_11721,N_11738);
and U12036 (N_12036,N_11977,N_11983);
nor U12037 (N_12037,N_11745,N_11795);
xor U12038 (N_12038,N_11800,N_11894);
nand U12039 (N_12039,N_11998,N_11726);
and U12040 (N_12040,N_11809,N_11890);
and U12041 (N_12041,N_11946,N_11826);
and U12042 (N_12042,N_11868,N_11948);
or U12043 (N_12043,N_11828,N_11924);
nand U12044 (N_12044,N_11850,N_11845);
xor U12045 (N_12045,N_11885,N_11927);
nor U12046 (N_12046,N_11968,N_11987);
or U12047 (N_12047,N_11847,N_11824);
nand U12048 (N_12048,N_11724,N_11932);
xor U12049 (N_12049,N_11770,N_11861);
nor U12050 (N_12050,N_11888,N_11956);
and U12051 (N_12051,N_11846,N_11843);
or U12052 (N_12052,N_11755,N_11700);
xor U12053 (N_12053,N_11916,N_11822);
nor U12054 (N_12054,N_11832,N_11950);
and U12055 (N_12055,N_11789,N_11867);
and U12056 (N_12056,N_11954,N_11971);
nand U12057 (N_12057,N_11706,N_11814);
and U12058 (N_12058,N_11862,N_11959);
nor U12059 (N_12059,N_11988,N_11967);
nand U12060 (N_12060,N_11743,N_11823);
nor U12061 (N_12061,N_11973,N_11939);
nand U12062 (N_12062,N_11825,N_11740);
xnor U12063 (N_12063,N_11871,N_11785);
nor U12064 (N_12064,N_11880,N_11739);
xor U12065 (N_12065,N_11873,N_11986);
xor U12066 (N_12066,N_11964,N_11966);
or U12067 (N_12067,N_11758,N_11902);
and U12068 (N_12068,N_11749,N_11754);
or U12069 (N_12069,N_11812,N_11720);
and U12070 (N_12070,N_11863,N_11747);
or U12071 (N_12071,N_11810,N_11714);
and U12072 (N_12072,N_11801,N_11976);
and U12073 (N_12073,N_11852,N_11907);
or U12074 (N_12074,N_11962,N_11930);
xor U12075 (N_12075,N_11757,N_11764);
and U12076 (N_12076,N_11765,N_11997);
or U12077 (N_12077,N_11841,N_11787);
nor U12078 (N_12078,N_11803,N_11773);
or U12079 (N_12079,N_11844,N_11969);
nor U12080 (N_12080,N_11816,N_11848);
nor U12081 (N_12081,N_11802,N_11791);
xor U12082 (N_12082,N_11899,N_11704);
nor U12083 (N_12083,N_11965,N_11996);
xor U12084 (N_12084,N_11859,N_11913);
nor U12085 (N_12085,N_11718,N_11872);
xnor U12086 (N_12086,N_11837,N_11865);
nor U12087 (N_12087,N_11804,N_11780);
nand U12088 (N_12088,N_11937,N_11926);
nor U12089 (N_12089,N_11897,N_11708);
xnor U12090 (N_12090,N_11741,N_11732);
or U12091 (N_12091,N_11849,N_11901);
or U12092 (N_12092,N_11934,N_11855);
nand U12093 (N_12093,N_11792,N_11702);
nor U12094 (N_12094,N_11896,N_11990);
and U12095 (N_12095,N_11922,N_11910);
xor U12096 (N_12096,N_11761,N_11918);
or U12097 (N_12097,N_11942,N_11994);
or U12098 (N_12098,N_11811,N_11928);
xor U12099 (N_12099,N_11727,N_11991);
or U12100 (N_12100,N_11921,N_11892);
xnor U12101 (N_12101,N_11808,N_11887);
nor U12102 (N_12102,N_11790,N_11799);
nand U12103 (N_12103,N_11752,N_11713);
nor U12104 (N_12104,N_11883,N_11995);
or U12105 (N_12105,N_11898,N_11836);
or U12106 (N_12106,N_11857,N_11958);
xnor U12107 (N_12107,N_11874,N_11750);
and U12108 (N_12108,N_11725,N_11763);
nor U12109 (N_12109,N_11970,N_11779);
xnor U12110 (N_12110,N_11906,N_11925);
and U12111 (N_12111,N_11753,N_11933);
xnor U12112 (N_12112,N_11895,N_11781);
or U12113 (N_12113,N_11914,N_11833);
and U12114 (N_12114,N_11853,N_11893);
or U12115 (N_12115,N_11734,N_11960);
nor U12116 (N_12116,N_11737,N_11900);
and U12117 (N_12117,N_11882,N_11784);
or U12118 (N_12118,N_11805,N_11788);
and U12119 (N_12119,N_11771,N_11707);
nand U12120 (N_12120,N_11856,N_11768);
xor U12121 (N_12121,N_11952,N_11731);
xnor U12122 (N_12122,N_11774,N_11766);
and U12123 (N_12123,N_11984,N_11951);
xnor U12124 (N_12124,N_11886,N_11831);
nor U12125 (N_12125,N_11945,N_11786);
or U12126 (N_12126,N_11751,N_11730);
or U12127 (N_12127,N_11978,N_11830);
nand U12128 (N_12128,N_11878,N_11729);
nand U12129 (N_12129,N_11746,N_11943);
xnor U12130 (N_12130,N_11806,N_11904);
xor U12131 (N_12131,N_11963,N_11851);
or U12132 (N_12132,N_11719,N_11756);
or U12133 (N_12133,N_11935,N_11716);
xor U12134 (N_12134,N_11877,N_11919);
or U12135 (N_12135,N_11875,N_11760);
nor U12136 (N_12136,N_11710,N_11762);
nand U12137 (N_12137,N_11931,N_11858);
xnor U12138 (N_12138,N_11711,N_11759);
or U12139 (N_12139,N_11944,N_11975);
xnor U12140 (N_12140,N_11891,N_11736);
or U12141 (N_12141,N_11860,N_11876);
xnor U12142 (N_12142,N_11772,N_11980);
xor U12143 (N_12143,N_11703,N_11715);
nand U12144 (N_12144,N_11834,N_11869);
xor U12145 (N_12145,N_11911,N_11793);
xnor U12146 (N_12146,N_11818,N_11999);
nor U12147 (N_12147,N_11908,N_11989);
nand U12148 (N_12148,N_11941,N_11957);
nor U12149 (N_12149,N_11733,N_11903);
or U12150 (N_12150,N_11895,N_11941);
and U12151 (N_12151,N_11850,N_11790);
nor U12152 (N_12152,N_11795,N_11741);
nor U12153 (N_12153,N_11838,N_11926);
or U12154 (N_12154,N_11836,N_11755);
xnor U12155 (N_12155,N_11956,N_11982);
and U12156 (N_12156,N_11735,N_11885);
or U12157 (N_12157,N_11897,N_11866);
nand U12158 (N_12158,N_11762,N_11814);
and U12159 (N_12159,N_11793,N_11764);
nor U12160 (N_12160,N_11854,N_11960);
xnor U12161 (N_12161,N_11823,N_11718);
and U12162 (N_12162,N_11833,N_11835);
xnor U12163 (N_12163,N_11828,N_11903);
xor U12164 (N_12164,N_11984,N_11969);
xor U12165 (N_12165,N_11954,N_11902);
and U12166 (N_12166,N_11952,N_11890);
or U12167 (N_12167,N_11896,N_11975);
and U12168 (N_12168,N_11945,N_11739);
and U12169 (N_12169,N_11797,N_11735);
nor U12170 (N_12170,N_11924,N_11703);
or U12171 (N_12171,N_11789,N_11837);
nor U12172 (N_12172,N_11708,N_11728);
xor U12173 (N_12173,N_11901,N_11986);
xnor U12174 (N_12174,N_11925,N_11788);
nor U12175 (N_12175,N_11795,N_11800);
or U12176 (N_12176,N_11991,N_11748);
and U12177 (N_12177,N_11975,N_11899);
xnor U12178 (N_12178,N_11918,N_11798);
nor U12179 (N_12179,N_11960,N_11919);
nor U12180 (N_12180,N_11835,N_11870);
xnor U12181 (N_12181,N_11813,N_11889);
nor U12182 (N_12182,N_11981,N_11863);
nand U12183 (N_12183,N_11753,N_11878);
nor U12184 (N_12184,N_11939,N_11807);
or U12185 (N_12185,N_11911,N_11715);
or U12186 (N_12186,N_11728,N_11998);
nand U12187 (N_12187,N_11834,N_11961);
and U12188 (N_12188,N_11787,N_11816);
nand U12189 (N_12189,N_11934,N_11837);
or U12190 (N_12190,N_11948,N_11862);
nand U12191 (N_12191,N_11973,N_11704);
nor U12192 (N_12192,N_11958,N_11873);
or U12193 (N_12193,N_11919,N_11726);
or U12194 (N_12194,N_11732,N_11802);
or U12195 (N_12195,N_11977,N_11879);
nor U12196 (N_12196,N_11888,N_11765);
and U12197 (N_12197,N_11752,N_11791);
and U12198 (N_12198,N_11727,N_11930);
nor U12199 (N_12199,N_11762,N_11819);
nor U12200 (N_12200,N_11870,N_11972);
and U12201 (N_12201,N_11701,N_11928);
nor U12202 (N_12202,N_11783,N_11743);
nor U12203 (N_12203,N_11853,N_11799);
or U12204 (N_12204,N_11700,N_11918);
nor U12205 (N_12205,N_11913,N_11955);
and U12206 (N_12206,N_11704,N_11785);
or U12207 (N_12207,N_11802,N_11898);
nor U12208 (N_12208,N_11794,N_11821);
xor U12209 (N_12209,N_11717,N_11789);
nand U12210 (N_12210,N_11774,N_11720);
and U12211 (N_12211,N_11961,N_11744);
xor U12212 (N_12212,N_11761,N_11862);
and U12213 (N_12213,N_11938,N_11828);
xnor U12214 (N_12214,N_11754,N_11984);
xor U12215 (N_12215,N_11782,N_11981);
nand U12216 (N_12216,N_11796,N_11930);
or U12217 (N_12217,N_11968,N_11963);
nor U12218 (N_12218,N_11880,N_11888);
and U12219 (N_12219,N_11840,N_11821);
nand U12220 (N_12220,N_11898,N_11930);
nand U12221 (N_12221,N_11884,N_11977);
nand U12222 (N_12222,N_11844,N_11714);
nand U12223 (N_12223,N_11828,N_11988);
nand U12224 (N_12224,N_11801,N_11947);
or U12225 (N_12225,N_11854,N_11907);
and U12226 (N_12226,N_11716,N_11934);
or U12227 (N_12227,N_11909,N_11836);
or U12228 (N_12228,N_11848,N_11962);
and U12229 (N_12229,N_11742,N_11776);
or U12230 (N_12230,N_11767,N_11747);
and U12231 (N_12231,N_11758,N_11846);
nor U12232 (N_12232,N_11868,N_11884);
nand U12233 (N_12233,N_11815,N_11987);
or U12234 (N_12234,N_11797,N_11978);
or U12235 (N_12235,N_11779,N_11764);
xnor U12236 (N_12236,N_11862,N_11776);
xor U12237 (N_12237,N_11949,N_11996);
nand U12238 (N_12238,N_11990,N_11801);
and U12239 (N_12239,N_11906,N_11949);
nor U12240 (N_12240,N_11787,N_11754);
nand U12241 (N_12241,N_11870,N_11788);
nand U12242 (N_12242,N_11988,N_11721);
nor U12243 (N_12243,N_11881,N_11740);
and U12244 (N_12244,N_11981,N_11757);
or U12245 (N_12245,N_11729,N_11731);
xor U12246 (N_12246,N_11879,N_11971);
or U12247 (N_12247,N_11915,N_11950);
or U12248 (N_12248,N_11776,N_11888);
nor U12249 (N_12249,N_11910,N_11756);
and U12250 (N_12250,N_11820,N_11784);
or U12251 (N_12251,N_11954,N_11929);
xnor U12252 (N_12252,N_11803,N_11944);
xor U12253 (N_12253,N_11840,N_11999);
or U12254 (N_12254,N_11814,N_11951);
nor U12255 (N_12255,N_11881,N_11824);
xnor U12256 (N_12256,N_11789,N_11859);
nand U12257 (N_12257,N_11832,N_11965);
nor U12258 (N_12258,N_11905,N_11889);
or U12259 (N_12259,N_11799,N_11994);
xnor U12260 (N_12260,N_11771,N_11703);
and U12261 (N_12261,N_11716,N_11986);
nor U12262 (N_12262,N_11907,N_11707);
nand U12263 (N_12263,N_11768,N_11782);
and U12264 (N_12264,N_11797,N_11996);
xnor U12265 (N_12265,N_11939,N_11911);
and U12266 (N_12266,N_11795,N_11702);
nor U12267 (N_12267,N_11701,N_11790);
nand U12268 (N_12268,N_11720,N_11741);
nor U12269 (N_12269,N_11825,N_11737);
and U12270 (N_12270,N_11899,N_11737);
xnor U12271 (N_12271,N_11741,N_11958);
nand U12272 (N_12272,N_11944,N_11712);
nor U12273 (N_12273,N_11861,N_11778);
xor U12274 (N_12274,N_11804,N_11845);
or U12275 (N_12275,N_11967,N_11761);
and U12276 (N_12276,N_11717,N_11972);
nor U12277 (N_12277,N_11801,N_11956);
and U12278 (N_12278,N_11740,N_11949);
and U12279 (N_12279,N_11882,N_11765);
or U12280 (N_12280,N_11888,N_11910);
and U12281 (N_12281,N_11754,N_11853);
or U12282 (N_12282,N_11743,N_11749);
or U12283 (N_12283,N_11846,N_11971);
and U12284 (N_12284,N_11931,N_11915);
nor U12285 (N_12285,N_11826,N_11955);
xnor U12286 (N_12286,N_11867,N_11929);
nor U12287 (N_12287,N_11927,N_11705);
nor U12288 (N_12288,N_11773,N_11833);
or U12289 (N_12289,N_11978,N_11994);
and U12290 (N_12290,N_11770,N_11829);
or U12291 (N_12291,N_11747,N_11721);
xor U12292 (N_12292,N_11802,N_11799);
nor U12293 (N_12293,N_11942,N_11850);
or U12294 (N_12294,N_11919,N_11799);
nor U12295 (N_12295,N_11704,N_11984);
or U12296 (N_12296,N_11912,N_11773);
and U12297 (N_12297,N_11770,N_11851);
nand U12298 (N_12298,N_11856,N_11779);
nor U12299 (N_12299,N_11858,N_11821);
nor U12300 (N_12300,N_12208,N_12048);
nand U12301 (N_12301,N_12109,N_12039);
nor U12302 (N_12302,N_12050,N_12059);
nor U12303 (N_12303,N_12106,N_12092);
and U12304 (N_12304,N_12250,N_12297);
or U12305 (N_12305,N_12196,N_12282);
nor U12306 (N_12306,N_12190,N_12067);
or U12307 (N_12307,N_12139,N_12075);
nor U12308 (N_12308,N_12099,N_12084);
nor U12309 (N_12309,N_12178,N_12021);
nand U12310 (N_12310,N_12188,N_12136);
and U12311 (N_12311,N_12058,N_12223);
nand U12312 (N_12312,N_12160,N_12291);
or U12313 (N_12313,N_12226,N_12210);
and U12314 (N_12314,N_12085,N_12133);
xnor U12315 (N_12315,N_12045,N_12126);
nor U12316 (N_12316,N_12063,N_12049);
or U12317 (N_12317,N_12254,N_12060);
nand U12318 (N_12318,N_12009,N_12014);
and U12319 (N_12319,N_12164,N_12241);
xnor U12320 (N_12320,N_12203,N_12184);
and U12321 (N_12321,N_12137,N_12266);
and U12322 (N_12322,N_12015,N_12248);
nor U12323 (N_12323,N_12125,N_12120);
and U12324 (N_12324,N_12197,N_12234);
nand U12325 (N_12325,N_12166,N_12138);
or U12326 (N_12326,N_12230,N_12276);
or U12327 (N_12327,N_12065,N_12228);
and U12328 (N_12328,N_12013,N_12259);
xor U12329 (N_12329,N_12274,N_12119);
nand U12330 (N_12330,N_12217,N_12219);
nand U12331 (N_12331,N_12244,N_12082);
xnor U12332 (N_12332,N_12174,N_12182);
and U12333 (N_12333,N_12054,N_12239);
and U12334 (N_12334,N_12224,N_12261);
xor U12335 (N_12335,N_12071,N_12135);
nor U12336 (N_12336,N_12128,N_12105);
nor U12337 (N_12337,N_12279,N_12212);
xnor U12338 (N_12338,N_12189,N_12131);
or U12339 (N_12339,N_12095,N_12235);
nand U12340 (N_12340,N_12094,N_12107);
nor U12341 (N_12341,N_12143,N_12245);
or U12342 (N_12342,N_12149,N_12218);
nor U12343 (N_12343,N_12167,N_12155);
or U12344 (N_12344,N_12031,N_12114);
nand U12345 (N_12345,N_12242,N_12030);
xnor U12346 (N_12346,N_12025,N_12018);
nand U12347 (N_12347,N_12117,N_12225);
nand U12348 (N_12348,N_12086,N_12298);
or U12349 (N_12349,N_12124,N_12080);
nor U12350 (N_12350,N_12122,N_12170);
or U12351 (N_12351,N_12098,N_12186);
and U12352 (N_12352,N_12079,N_12087);
nand U12353 (N_12353,N_12134,N_12206);
xor U12354 (N_12354,N_12003,N_12193);
and U12355 (N_12355,N_12293,N_12100);
or U12356 (N_12356,N_12007,N_12281);
and U12357 (N_12357,N_12264,N_12011);
and U12358 (N_12358,N_12043,N_12019);
nor U12359 (N_12359,N_12200,N_12033);
or U12360 (N_12360,N_12077,N_12012);
nor U12361 (N_12361,N_12140,N_12026);
nand U12362 (N_12362,N_12294,N_12199);
nor U12363 (N_12363,N_12081,N_12284);
xor U12364 (N_12364,N_12295,N_12076);
or U12365 (N_12365,N_12110,N_12004);
and U12366 (N_12366,N_12161,N_12187);
xor U12367 (N_12367,N_12042,N_12256);
nor U12368 (N_12368,N_12127,N_12195);
nand U12369 (N_12369,N_12185,N_12061);
nor U12370 (N_12370,N_12068,N_12260);
nor U12371 (N_12371,N_12157,N_12090);
xor U12372 (N_12372,N_12118,N_12129);
nand U12373 (N_12373,N_12093,N_12289);
and U12374 (N_12374,N_12057,N_12156);
nand U12375 (N_12375,N_12024,N_12147);
and U12376 (N_12376,N_12258,N_12168);
and U12377 (N_12377,N_12027,N_12097);
xor U12378 (N_12378,N_12038,N_12113);
nor U12379 (N_12379,N_12191,N_12102);
xnor U12380 (N_12380,N_12263,N_12202);
nor U12381 (N_12381,N_12028,N_12069);
nand U12382 (N_12382,N_12269,N_12051);
nor U12383 (N_12383,N_12088,N_12180);
nor U12384 (N_12384,N_12035,N_12290);
or U12385 (N_12385,N_12243,N_12267);
or U12386 (N_12386,N_12292,N_12146);
and U12387 (N_12387,N_12141,N_12052);
xor U12388 (N_12388,N_12176,N_12022);
xnor U12389 (N_12389,N_12229,N_12232);
or U12390 (N_12390,N_12236,N_12271);
nor U12391 (N_12391,N_12121,N_12016);
xnor U12392 (N_12392,N_12159,N_12123);
or U12393 (N_12393,N_12103,N_12183);
nand U12394 (N_12394,N_12002,N_12017);
nand U12395 (N_12395,N_12008,N_12020);
nor U12396 (N_12396,N_12181,N_12233);
nor U12397 (N_12397,N_12207,N_12029);
or U12398 (N_12398,N_12154,N_12287);
or U12399 (N_12399,N_12270,N_12177);
nand U12400 (N_12400,N_12053,N_12213);
or U12401 (N_12401,N_12257,N_12044);
nor U12402 (N_12402,N_12116,N_12251);
nand U12403 (N_12403,N_12192,N_12055);
nand U12404 (N_12404,N_12280,N_12249);
xnor U12405 (N_12405,N_12246,N_12142);
nand U12406 (N_12406,N_12096,N_12046);
xnor U12407 (N_12407,N_12062,N_12091);
xnor U12408 (N_12408,N_12252,N_12222);
nor U12409 (N_12409,N_12201,N_12037);
xnor U12410 (N_12410,N_12227,N_12240);
and U12411 (N_12411,N_12072,N_12272);
xor U12412 (N_12412,N_12238,N_12288);
or U12413 (N_12413,N_12247,N_12036);
xor U12414 (N_12414,N_12144,N_12047);
or U12415 (N_12415,N_12194,N_12173);
nor U12416 (N_12416,N_12171,N_12296);
and U12417 (N_12417,N_12286,N_12153);
nand U12418 (N_12418,N_12073,N_12006);
and U12419 (N_12419,N_12214,N_12163);
and U12420 (N_12420,N_12273,N_12148);
or U12421 (N_12421,N_12132,N_12089);
and U12422 (N_12422,N_12083,N_12150);
nand U12423 (N_12423,N_12040,N_12172);
or U12424 (N_12424,N_12130,N_12204);
or U12425 (N_12425,N_12064,N_12010);
nand U12426 (N_12426,N_12151,N_12275);
xor U12427 (N_12427,N_12231,N_12005);
xor U12428 (N_12428,N_12104,N_12255);
or U12429 (N_12429,N_12112,N_12237);
xor U12430 (N_12430,N_12078,N_12299);
and U12431 (N_12431,N_12179,N_12034);
or U12432 (N_12432,N_12175,N_12209);
or U12433 (N_12433,N_12145,N_12056);
nand U12434 (N_12434,N_12198,N_12221);
or U12435 (N_12435,N_12115,N_12211);
nand U12436 (N_12436,N_12101,N_12285);
or U12437 (N_12437,N_12023,N_12152);
xnor U12438 (N_12438,N_12066,N_12070);
nor U12439 (N_12439,N_12268,N_12032);
nor U12440 (N_12440,N_12277,N_12262);
or U12441 (N_12441,N_12169,N_12265);
or U12442 (N_12442,N_12220,N_12165);
xor U12443 (N_12443,N_12158,N_12283);
and U12444 (N_12444,N_12253,N_12000);
nand U12445 (N_12445,N_12041,N_12108);
nor U12446 (N_12446,N_12215,N_12111);
nor U12447 (N_12447,N_12205,N_12278);
nor U12448 (N_12448,N_12162,N_12001);
xnor U12449 (N_12449,N_12074,N_12216);
and U12450 (N_12450,N_12027,N_12202);
xnor U12451 (N_12451,N_12240,N_12076);
nor U12452 (N_12452,N_12056,N_12069);
or U12453 (N_12453,N_12264,N_12133);
and U12454 (N_12454,N_12105,N_12251);
and U12455 (N_12455,N_12236,N_12077);
nand U12456 (N_12456,N_12251,N_12119);
or U12457 (N_12457,N_12201,N_12297);
or U12458 (N_12458,N_12217,N_12191);
or U12459 (N_12459,N_12013,N_12216);
and U12460 (N_12460,N_12077,N_12000);
nand U12461 (N_12461,N_12143,N_12036);
xnor U12462 (N_12462,N_12080,N_12001);
or U12463 (N_12463,N_12192,N_12147);
nor U12464 (N_12464,N_12193,N_12196);
xor U12465 (N_12465,N_12223,N_12114);
nand U12466 (N_12466,N_12211,N_12175);
xnor U12467 (N_12467,N_12162,N_12048);
and U12468 (N_12468,N_12130,N_12291);
or U12469 (N_12469,N_12052,N_12114);
or U12470 (N_12470,N_12123,N_12295);
nand U12471 (N_12471,N_12131,N_12182);
nor U12472 (N_12472,N_12127,N_12153);
nand U12473 (N_12473,N_12107,N_12124);
and U12474 (N_12474,N_12140,N_12150);
or U12475 (N_12475,N_12241,N_12230);
and U12476 (N_12476,N_12011,N_12293);
or U12477 (N_12477,N_12115,N_12164);
nand U12478 (N_12478,N_12242,N_12294);
xor U12479 (N_12479,N_12044,N_12188);
xnor U12480 (N_12480,N_12026,N_12097);
or U12481 (N_12481,N_12069,N_12100);
or U12482 (N_12482,N_12110,N_12156);
xor U12483 (N_12483,N_12164,N_12065);
or U12484 (N_12484,N_12087,N_12242);
or U12485 (N_12485,N_12263,N_12029);
nand U12486 (N_12486,N_12174,N_12023);
or U12487 (N_12487,N_12249,N_12159);
xnor U12488 (N_12488,N_12083,N_12028);
nor U12489 (N_12489,N_12193,N_12032);
xor U12490 (N_12490,N_12059,N_12094);
nand U12491 (N_12491,N_12141,N_12234);
and U12492 (N_12492,N_12222,N_12017);
nor U12493 (N_12493,N_12126,N_12070);
nand U12494 (N_12494,N_12103,N_12131);
nand U12495 (N_12495,N_12126,N_12277);
and U12496 (N_12496,N_12069,N_12053);
xnor U12497 (N_12497,N_12172,N_12280);
or U12498 (N_12498,N_12178,N_12013);
xor U12499 (N_12499,N_12170,N_12162);
or U12500 (N_12500,N_12187,N_12088);
nor U12501 (N_12501,N_12234,N_12094);
xnor U12502 (N_12502,N_12072,N_12034);
nor U12503 (N_12503,N_12073,N_12282);
nor U12504 (N_12504,N_12069,N_12093);
xnor U12505 (N_12505,N_12298,N_12274);
or U12506 (N_12506,N_12226,N_12229);
and U12507 (N_12507,N_12012,N_12088);
nor U12508 (N_12508,N_12129,N_12164);
xnor U12509 (N_12509,N_12195,N_12014);
xor U12510 (N_12510,N_12218,N_12188);
nor U12511 (N_12511,N_12258,N_12139);
xor U12512 (N_12512,N_12157,N_12018);
or U12513 (N_12513,N_12143,N_12094);
nand U12514 (N_12514,N_12072,N_12053);
nand U12515 (N_12515,N_12286,N_12056);
nand U12516 (N_12516,N_12182,N_12222);
nor U12517 (N_12517,N_12064,N_12113);
nor U12518 (N_12518,N_12000,N_12220);
xor U12519 (N_12519,N_12205,N_12193);
nand U12520 (N_12520,N_12255,N_12237);
nor U12521 (N_12521,N_12097,N_12020);
xnor U12522 (N_12522,N_12213,N_12108);
and U12523 (N_12523,N_12248,N_12080);
or U12524 (N_12524,N_12162,N_12245);
nor U12525 (N_12525,N_12253,N_12199);
nand U12526 (N_12526,N_12145,N_12009);
and U12527 (N_12527,N_12218,N_12154);
or U12528 (N_12528,N_12237,N_12297);
nand U12529 (N_12529,N_12097,N_12294);
nor U12530 (N_12530,N_12291,N_12120);
or U12531 (N_12531,N_12060,N_12257);
nor U12532 (N_12532,N_12111,N_12226);
and U12533 (N_12533,N_12054,N_12031);
nor U12534 (N_12534,N_12034,N_12198);
nor U12535 (N_12535,N_12184,N_12130);
nand U12536 (N_12536,N_12002,N_12236);
and U12537 (N_12537,N_12016,N_12012);
nand U12538 (N_12538,N_12029,N_12223);
or U12539 (N_12539,N_12284,N_12200);
nand U12540 (N_12540,N_12087,N_12246);
xor U12541 (N_12541,N_12256,N_12238);
or U12542 (N_12542,N_12193,N_12020);
nand U12543 (N_12543,N_12227,N_12091);
and U12544 (N_12544,N_12269,N_12201);
and U12545 (N_12545,N_12124,N_12094);
nor U12546 (N_12546,N_12218,N_12137);
or U12547 (N_12547,N_12097,N_12165);
nand U12548 (N_12548,N_12067,N_12177);
xnor U12549 (N_12549,N_12065,N_12238);
and U12550 (N_12550,N_12269,N_12232);
nor U12551 (N_12551,N_12130,N_12038);
and U12552 (N_12552,N_12189,N_12091);
nand U12553 (N_12553,N_12072,N_12168);
xnor U12554 (N_12554,N_12152,N_12134);
or U12555 (N_12555,N_12012,N_12142);
xor U12556 (N_12556,N_12074,N_12137);
xnor U12557 (N_12557,N_12136,N_12075);
or U12558 (N_12558,N_12143,N_12248);
xnor U12559 (N_12559,N_12016,N_12276);
nand U12560 (N_12560,N_12205,N_12123);
or U12561 (N_12561,N_12139,N_12058);
nor U12562 (N_12562,N_12177,N_12153);
xnor U12563 (N_12563,N_12291,N_12182);
xor U12564 (N_12564,N_12259,N_12080);
or U12565 (N_12565,N_12282,N_12002);
nor U12566 (N_12566,N_12219,N_12078);
or U12567 (N_12567,N_12030,N_12240);
nand U12568 (N_12568,N_12226,N_12110);
and U12569 (N_12569,N_12107,N_12169);
and U12570 (N_12570,N_12281,N_12299);
and U12571 (N_12571,N_12018,N_12058);
xor U12572 (N_12572,N_12216,N_12298);
xor U12573 (N_12573,N_12019,N_12187);
or U12574 (N_12574,N_12255,N_12169);
and U12575 (N_12575,N_12203,N_12146);
and U12576 (N_12576,N_12118,N_12208);
and U12577 (N_12577,N_12178,N_12071);
or U12578 (N_12578,N_12053,N_12115);
nand U12579 (N_12579,N_12177,N_12114);
xor U12580 (N_12580,N_12204,N_12039);
nor U12581 (N_12581,N_12129,N_12198);
nand U12582 (N_12582,N_12157,N_12107);
or U12583 (N_12583,N_12092,N_12232);
nor U12584 (N_12584,N_12157,N_12053);
and U12585 (N_12585,N_12141,N_12184);
and U12586 (N_12586,N_12008,N_12022);
nor U12587 (N_12587,N_12210,N_12061);
nor U12588 (N_12588,N_12214,N_12102);
nand U12589 (N_12589,N_12237,N_12282);
nor U12590 (N_12590,N_12097,N_12247);
nand U12591 (N_12591,N_12213,N_12075);
nand U12592 (N_12592,N_12102,N_12062);
and U12593 (N_12593,N_12112,N_12260);
nor U12594 (N_12594,N_12151,N_12255);
and U12595 (N_12595,N_12070,N_12087);
nand U12596 (N_12596,N_12157,N_12049);
xnor U12597 (N_12597,N_12009,N_12037);
xnor U12598 (N_12598,N_12249,N_12000);
and U12599 (N_12599,N_12032,N_12222);
and U12600 (N_12600,N_12375,N_12543);
xnor U12601 (N_12601,N_12515,N_12542);
nand U12602 (N_12602,N_12537,N_12523);
nand U12603 (N_12603,N_12541,N_12569);
or U12604 (N_12604,N_12554,N_12453);
and U12605 (N_12605,N_12528,N_12565);
or U12606 (N_12606,N_12438,N_12317);
nor U12607 (N_12607,N_12427,N_12586);
xor U12608 (N_12608,N_12574,N_12402);
or U12609 (N_12609,N_12324,N_12477);
nand U12610 (N_12610,N_12325,N_12355);
or U12611 (N_12611,N_12481,N_12545);
nor U12612 (N_12612,N_12422,N_12464);
nand U12613 (N_12613,N_12327,N_12424);
or U12614 (N_12614,N_12492,N_12465);
nand U12615 (N_12615,N_12524,N_12535);
nor U12616 (N_12616,N_12352,N_12412);
nor U12617 (N_12617,N_12437,N_12447);
or U12618 (N_12618,N_12517,N_12564);
and U12619 (N_12619,N_12457,N_12360);
nor U12620 (N_12620,N_12416,N_12561);
xnor U12621 (N_12621,N_12445,N_12527);
nand U12622 (N_12622,N_12467,N_12534);
nor U12623 (N_12623,N_12566,N_12559);
nand U12624 (N_12624,N_12451,N_12429);
xnor U12625 (N_12625,N_12332,N_12425);
or U12626 (N_12626,N_12343,N_12480);
nand U12627 (N_12627,N_12333,N_12518);
and U12628 (N_12628,N_12419,N_12318);
or U12629 (N_12629,N_12468,N_12345);
and U12630 (N_12630,N_12370,N_12501);
and U12631 (N_12631,N_12516,N_12322);
or U12632 (N_12632,N_12571,N_12396);
and U12633 (N_12633,N_12366,N_12529);
or U12634 (N_12634,N_12488,N_12364);
nand U12635 (N_12635,N_12514,N_12588);
or U12636 (N_12636,N_12404,N_12544);
or U12637 (N_12637,N_12507,N_12315);
nor U12638 (N_12638,N_12374,N_12496);
or U12639 (N_12639,N_12576,N_12335);
nor U12640 (N_12640,N_12472,N_12446);
or U12641 (N_12641,N_12432,N_12369);
xnor U12642 (N_12642,N_12475,N_12338);
nand U12643 (N_12643,N_12577,N_12557);
and U12644 (N_12644,N_12593,N_12428);
and U12645 (N_12645,N_12594,N_12525);
xnor U12646 (N_12646,N_12484,N_12340);
and U12647 (N_12647,N_12431,N_12334);
nor U12648 (N_12648,N_12474,N_12313);
and U12649 (N_12649,N_12392,N_12582);
nor U12650 (N_12650,N_12376,N_12356);
xnor U12651 (N_12651,N_12595,N_12538);
nor U12652 (N_12652,N_12420,N_12367);
and U12653 (N_12653,N_12526,N_12418);
or U12654 (N_12654,N_12407,N_12430);
nor U12655 (N_12655,N_12359,N_12540);
or U12656 (N_12656,N_12456,N_12382);
nand U12657 (N_12657,N_12316,N_12441);
xnor U12658 (N_12658,N_12466,N_12532);
and U12659 (N_12659,N_12377,N_12521);
or U12660 (N_12660,N_12579,N_12556);
and U12661 (N_12661,N_12572,N_12354);
xnor U12662 (N_12662,N_12575,N_12597);
and U12663 (N_12663,N_12387,N_12581);
nand U12664 (N_12664,N_12450,N_12505);
nor U12665 (N_12665,N_12589,N_12336);
nand U12666 (N_12666,N_12536,N_12362);
and U12667 (N_12667,N_12510,N_12469);
and U12668 (N_12668,N_12371,N_12388);
and U12669 (N_12669,N_12341,N_12300);
nor U12670 (N_12670,N_12331,N_12500);
and U12671 (N_12671,N_12573,N_12405);
and U12672 (N_12672,N_12372,N_12596);
xor U12673 (N_12673,N_12379,N_12323);
xor U12674 (N_12674,N_12321,N_12530);
nor U12675 (N_12675,N_12443,N_12381);
nand U12676 (N_12676,N_12478,N_12494);
xor U12677 (N_12677,N_12460,N_12353);
or U12678 (N_12678,N_12319,N_12444);
nand U12679 (N_12679,N_12455,N_12384);
nand U12680 (N_12680,N_12567,N_12358);
nor U12681 (N_12681,N_12351,N_12308);
nor U12682 (N_12682,N_12395,N_12583);
xor U12683 (N_12683,N_12499,N_12433);
nand U12684 (N_12684,N_12533,N_12504);
nand U12685 (N_12685,N_12378,N_12487);
xor U12686 (N_12686,N_12311,N_12421);
nor U12687 (N_12687,N_12549,N_12304);
and U12688 (N_12688,N_12309,N_12479);
and U12689 (N_12689,N_12578,N_12442);
nand U12690 (N_12690,N_12350,N_12326);
xor U12691 (N_12691,N_12509,N_12415);
and U12692 (N_12692,N_12386,N_12417);
or U12693 (N_12693,N_12310,N_12403);
and U12694 (N_12694,N_12346,N_12344);
or U12695 (N_12695,N_12423,N_12495);
nand U12696 (N_12696,N_12539,N_12552);
nor U12697 (N_12697,N_12568,N_12513);
nor U12698 (N_12698,N_12302,N_12411);
or U12699 (N_12699,N_12461,N_12305);
or U12700 (N_12700,N_12587,N_12591);
nand U12701 (N_12701,N_12361,N_12391);
or U12702 (N_12702,N_12368,N_12401);
and U12703 (N_12703,N_12490,N_12476);
nand U12704 (N_12704,N_12506,N_12497);
xor U12705 (N_12705,N_12337,N_12400);
and U12706 (N_12706,N_12555,N_12440);
nand U12707 (N_12707,N_12482,N_12454);
xor U12708 (N_12708,N_12558,N_12531);
and U12709 (N_12709,N_12328,N_12519);
nand U12710 (N_12710,N_12512,N_12398);
or U12711 (N_12711,N_12584,N_12448);
xor U12712 (N_12712,N_12390,N_12397);
nor U12713 (N_12713,N_12491,N_12522);
xnor U12714 (N_12714,N_12473,N_12329);
nand U12715 (N_12715,N_12485,N_12409);
and U12716 (N_12716,N_12449,N_12434);
or U12717 (N_12717,N_12347,N_12590);
nand U12718 (N_12718,N_12503,N_12560);
nor U12719 (N_12719,N_12330,N_12349);
xor U12720 (N_12720,N_12547,N_12303);
xnor U12721 (N_12721,N_12307,N_12342);
and U12722 (N_12722,N_12383,N_12312);
xor U12723 (N_12723,N_12511,N_12562);
or U12724 (N_12724,N_12548,N_12585);
and U12725 (N_12725,N_12580,N_12486);
nor U12726 (N_12726,N_12520,N_12363);
xnor U12727 (N_12727,N_12550,N_12598);
or U12728 (N_12728,N_12551,N_12306);
nand U12729 (N_12729,N_12399,N_12599);
xor U12730 (N_12730,N_12385,N_12348);
xor U12731 (N_12731,N_12498,N_12471);
or U12732 (N_12732,N_12463,N_12426);
or U12733 (N_12733,N_12436,N_12380);
nor U12734 (N_12734,N_12452,N_12439);
xnor U12735 (N_12735,N_12413,N_12458);
or U12736 (N_12736,N_12435,N_12546);
xnor U12737 (N_12737,N_12414,N_12553);
and U12738 (N_12738,N_12462,N_12365);
or U12739 (N_12739,N_12357,N_12393);
nand U12740 (N_12740,N_12389,N_12493);
and U12741 (N_12741,N_12314,N_12320);
and U12742 (N_12742,N_12408,N_12301);
nor U12743 (N_12743,N_12459,N_12508);
xnor U12744 (N_12744,N_12339,N_12470);
nor U12745 (N_12745,N_12394,N_12502);
or U12746 (N_12746,N_12373,N_12483);
nand U12747 (N_12747,N_12570,N_12410);
nand U12748 (N_12748,N_12563,N_12489);
and U12749 (N_12749,N_12592,N_12406);
or U12750 (N_12750,N_12331,N_12558);
or U12751 (N_12751,N_12539,N_12533);
and U12752 (N_12752,N_12460,N_12358);
and U12753 (N_12753,N_12312,N_12448);
nor U12754 (N_12754,N_12315,N_12392);
nand U12755 (N_12755,N_12414,N_12328);
nand U12756 (N_12756,N_12309,N_12526);
nor U12757 (N_12757,N_12455,N_12503);
nor U12758 (N_12758,N_12308,N_12475);
xor U12759 (N_12759,N_12438,N_12470);
or U12760 (N_12760,N_12331,N_12576);
xor U12761 (N_12761,N_12479,N_12513);
or U12762 (N_12762,N_12405,N_12348);
xnor U12763 (N_12763,N_12344,N_12367);
or U12764 (N_12764,N_12432,N_12345);
nand U12765 (N_12765,N_12558,N_12423);
nor U12766 (N_12766,N_12363,N_12590);
nor U12767 (N_12767,N_12430,N_12405);
and U12768 (N_12768,N_12394,N_12441);
nor U12769 (N_12769,N_12432,N_12503);
xnor U12770 (N_12770,N_12459,N_12419);
nand U12771 (N_12771,N_12549,N_12412);
nor U12772 (N_12772,N_12561,N_12425);
or U12773 (N_12773,N_12588,N_12570);
xor U12774 (N_12774,N_12566,N_12352);
or U12775 (N_12775,N_12495,N_12482);
or U12776 (N_12776,N_12446,N_12402);
nand U12777 (N_12777,N_12498,N_12387);
and U12778 (N_12778,N_12437,N_12425);
or U12779 (N_12779,N_12517,N_12573);
nand U12780 (N_12780,N_12443,N_12360);
nand U12781 (N_12781,N_12510,N_12357);
and U12782 (N_12782,N_12568,N_12345);
nor U12783 (N_12783,N_12432,N_12322);
xnor U12784 (N_12784,N_12332,N_12487);
and U12785 (N_12785,N_12559,N_12456);
nor U12786 (N_12786,N_12576,N_12593);
nand U12787 (N_12787,N_12435,N_12379);
nand U12788 (N_12788,N_12546,N_12557);
xor U12789 (N_12789,N_12546,N_12328);
or U12790 (N_12790,N_12370,N_12532);
or U12791 (N_12791,N_12353,N_12432);
and U12792 (N_12792,N_12324,N_12525);
or U12793 (N_12793,N_12408,N_12522);
nor U12794 (N_12794,N_12420,N_12355);
nand U12795 (N_12795,N_12521,N_12372);
xor U12796 (N_12796,N_12562,N_12438);
xnor U12797 (N_12797,N_12389,N_12322);
nor U12798 (N_12798,N_12425,N_12362);
nand U12799 (N_12799,N_12348,N_12523);
and U12800 (N_12800,N_12354,N_12520);
nor U12801 (N_12801,N_12479,N_12380);
nor U12802 (N_12802,N_12432,N_12338);
or U12803 (N_12803,N_12547,N_12580);
nor U12804 (N_12804,N_12317,N_12554);
or U12805 (N_12805,N_12569,N_12599);
nor U12806 (N_12806,N_12307,N_12321);
nand U12807 (N_12807,N_12553,N_12583);
or U12808 (N_12808,N_12349,N_12545);
and U12809 (N_12809,N_12466,N_12581);
nor U12810 (N_12810,N_12341,N_12472);
nor U12811 (N_12811,N_12477,N_12366);
xor U12812 (N_12812,N_12563,N_12305);
nor U12813 (N_12813,N_12427,N_12358);
nor U12814 (N_12814,N_12598,N_12340);
xnor U12815 (N_12815,N_12506,N_12442);
or U12816 (N_12816,N_12592,N_12328);
nand U12817 (N_12817,N_12585,N_12453);
nand U12818 (N_12818,N_12473,N_12450);
nand U12819 (N_12819,N_12340,N_12476);
or U12820 (N_12820,N_12472,N_12358);
and U12821 (N_12821,N_12369,N_12400);
nor U12822 (N_12822,N_12522,N_12476);
nand U12823 (N_12823,N_12306,N_12429);
xnor U12824 (N_12824,N_12509,N_12524);
nand U12825 (N_12825,N_12476,N_12328);
and U12826 (N_12826,N_12454,N_12453);
nor U12827 (N_12827,N_12370,N_12547);
nor U12828 (N_12828,N_12330,N_12476);
and U12829 (N_12829,N_12597,N_12594);
and U12830 (N_12830,N_12455,N_12327);
xor U12831 (N_12831,N_12308,N_12405);
nand U12832 (N_12832,N_12552,N_12598);
nor U12833 (N_12833,N_12490,N_12449);
or U12834 (N_12834,N_12477,N_12378);
or U12835 (N_12835,N_12369,N_12592);
nand U12836 (N_12836,N_12307,N_12446);
nor U12837 (N_12837,N_12347,N_12577);
and U12838 (N_12838,N_12464,N_12573);
and U12839 (N_12839,N_12401,N_12482);
xnor U12840 (N_12840,N_12444,N_12569);
xor U12841 (N_12841,N_12345,N_12455);
and U12842 (N_12842,N_12441,N_12306);
and U12843 (N_12843,N_12344,N_12414);
nor U12844 (N_12844,N_12574,N_12362);
xor U12845 (N_12845,N_12588,N_12376);
or U12846 (N_12846,N_12387,N_12315);
nor U12847 (N_12847,N_12311,N_12388);
or U12848 (N_12848,N_12529,N_12379);
and U12849 (N_12849,N_12393,N_12482);
or U12850 (N_12850,N_12473,N_12326);
nor U12851 (N_12851,N_12320,N_12308);
xnor U12852 (N_12852,N_12384,N_12477);
nor U12853 (N_12853,N_12390,N_12408);
and U12854 (N_12854,N_12441,N_12538);
nand U12855 (N_12855,N_12535,N_12526);
and U12856 (N_12856,N_12484,N_12542);
nand U12857 (N_12857,N_12327,N_12427);
xnor U12858 (N_12858,N_12556,N_12328);
or U12859 (N_12859,N_12463,N_12491);
or U12860 (N_12860,N_12377,N_12362);
nand U12861 (N_12861,N_12374,N_12418);
and U12862 (N_12862,N_12523,N_12568);
and U12863 (N_12863,N_12397,N_12304);
nor U12864 (N_12864,N_12499,N_12459);
and U12865 (N_12865,N_12425,N_12322);
nor U12866 (N_12866,N_12593,N_12398);
or U12867 (N_12867,N_12412,N_12567);
and U12868 (N_12868,N_12530,N_12310);
nor U12869 (N_12869,N_12573,N_12428);
nand U12870 (N_12870,N_12303,N_12441);
or U12871 (N_12871,N_12372,N_12509);
nand U12872 (N_12872,N_12334,N_12507);
nand U12873 (N_12873,N_12511,N_12311);
nand U12874 (N_12874,N_12436,N_12445);
xnor U12875 (N_12875,N_12305,N_12344);
and U12876 (N_12876,N_12565,N_12339);
or U12877 (N_12877,N_12573,N_12542);
nand U12878 (N_12878,N_12585,N_12423);
or U12879 (N_12879,N_12386,N_12457);
nand U12880 (N_12880,N_12398,N_12530);
nand U12881 (N_12881,N_12386,N_12421);
and U12882 (N_12882,N_12562,N_12359);
or U12883 (N_12883,N_12579,N_12467);
nor U12884 (N_12884,N_12332,N_12521);
or U12885 (N_12885,N_12376,N_12335);
xor U12886 (N_12886,N_12398,N_12376);
and U12887 (N_12887,N_12412,N_12553);
nand U12888 (N_12888,N_12563,N_12374);
nand U12889 (N_12889,N_12418,N_12417);
or U12890 (N_12890,N_12443,N_12563);
and U12891 (N_12891,N_12398,N_12563);
nor U12892 (N_12892,N_12336,N_12393);
nand U12893 (N_12893,N_12300,N_12324);
nor U12894 (N_12894,N_12567,N_12476);
and U12895 (N_12895,N_12456,N_12398);
nor U12896 (N_12896,N_12567,N_12454);
nand U12897 (N_12897,N_12497,N_12579);
xor U12898 (N_12898,N_12442,N_12307);
nand U12899 (N_12899,N_12499,N_12432);
and U12900 (N_12900,N_12621,N_12737);
nand U12901 (N_12901,N_12648,N_12710);
xnor U12902 (N_12902,N_12851,N_12610);
nor U12903 (N_12903,N_12662,N_12617);
and U12904 (N_12904,N_12808,N_12891);
xnor U12905 (N_12905,N_12858,N_12714);
and U12906 (N_12906,N_12600,N_12601);
xnor U12907 (N_12907,N_12668,N_12639);
and U12908 (N_12908,N_12734,N_12672);
and U12909 (N_12909,N_12745,N_12711);
or U12910 (N_12910,N_12791,N_12763);
nand U12911 (N_12911,N_12661,N_12762);
xor U12912 (N_12912,N_12814,N_12832);
nand U12913 (N_12913,N_12837,N_12818);
xnor U12914 (N_12914,N_12782,N_12831);
nor U12915 (N_12915,N_12874,N_12728);
nor U12916 (N_12916,N_12602,N_12766);
nand U12917 (N_12917,N_12660,N_12690);
nand U12918 (N_12918,N_12704,N_12868);
nor U12919 (N_12919,N_12893,N_12720);
nor U12920 (N_12920,N_12828,N_12765);
nor U12921 (N_12921,N_12702,N_12681);
or U12922 (N_12922,N_12616,N_12844);
nor U12923 (N_12923,N_12667,N_12856);
nor U12924 (N_12924,N_12877,N_12742);
and U12925 (N_12925,N_12817,N_12693);
nor U12926 (N_12926,N_12747,N_12718);
nor U12927 (N_12927,N_12725,N_12786);
and U12928 (N_12928,N_12756,N_12700);
nand U12929 (N_12929,N_12835,N_12848);
nor U12930 (N_12930,N_12754,N_12875);
xor U12931 (N_12931,N_12675,N_12803);
or U12932 (N_12932,N_12845,N_12883);
xnor U12933 (N_12933,N_12819,N_12859);
and U12934 (N_12934,N_12774,N_12611);
nand U12935 (N_12935,N_12655,N_12836);
nand U12936 (N_12936,N_12801,N_12638);
nor U12937 (N_12937,N_12794,N_12643);
nand U12938 (N_12938,N_12854,N_12838);
nor U12939 (N_12939,N_12771,N_12876);
nand U12940 (N_12940,N_12820,N_12862);
and U12941 (N_12941,N_12824,N_12841);
and U12942 (N_12942,N_12815,N_12634);
nor U12943 (N_12943,N_12863,N_12671);
nor U12944 (N_12944,N_12707,N_12767);
and U12945 (N_12945,N_12618,N_12659);
xnor U12946 (N_12946,N_12726,N_12688);
nand U12947 (N_12947,N_12785,N_12624);
nand U12948 (N_12948,N_12805,N_12649);
xnor U12949 (N_12949,N_12676,N_12789);
or U12950 (N_12950,N_12733,N_12698);
or U12951 (N_12951,N_12846,N_12669);
nand U12952 (N_12952,N_12653,N_12800);
nor U12953 (N_12953,N_12871,N_12886);
xnor U12954 (N_12954,N_12783,N_12810);
nor U12955 (N_12955,N_12899,N_12760);
nor U12956 (N_12956,N_12657,N_12722);
nor U12957 (N_12957,N_12750,N_12646);
xnor U12958 (N_12958,N_12713,N_12879);
nand U12959 (N_12959,N_12853,N_12833);
xor U12960 (N_12960,N_12677,N_12642);
xnor U12961 (N_12961,N_12806,N_12687);
and U12962 (N_12962,N_12855,N_12723);
or U12963 (N_12963,N_12705,N_12701);
nand U12964 (N_12964,N_12622,N_12788);
or U12965 (N_12965,N_12894,N_12694);
and U12966 (N_12966,N_12603,N_12864);
and U12967 (N_12967,N_12829,N_12843);
xnor U12968 (N_12968,N_12682,N_12764);
and U12969 (N_12969,N_12647,N_12708);
xor U12970 (N_12970,N_12790,N_12867);
xor U12971 (N_12971,N_12703,N_12839);
nand U12972 (N_12972,N_12813,N_12697);
nand U12973 (N_12973,N_12768,N_12746);
nor U12974 (N_12974,N_12679,N_12613);
xor U12975 (N_12975,N_12840,N_12873);
and U12976 (N_12976,N_12673,N_12898);
nand U12977 (N_12977,N_12896,N_12888);
nor U12978 (N_12978,N_12881,N_12717);
nor U12979 (N_12979,N_12731,N_12827);
or U12980 (N_12980,N_12842,N_12799);
nor U12981 (N_12981,N_12758,N_12811);
xnor U12982 (N_12982,N_12680,N_12684);
nor U12983 (N_12983,N_12628,N_12644);
xnor U12984 (N_12984,N_12666,N_12890);
or U12985 (N_12985,N_12753,N_12870);
xor U12986 (N_12986,N_12645,N_12732);
xor U12987 (N_12987,N_12619,N_12884);
nor U12988 (N_12988,N_12683,N_12607);
or U12989 (N_12989,N_12626,N_12632);
nor U12990 (N_12990,N_12614,N_12866);
xor U12991 (N_12991,N_12885,N_12685);
nand U12992 (N_12992,N_12847,N_12654);
nand U12993 (N_12993,N_12691,N_12887);
nand U12994 (N_12994,N_12604,N_12777);
and U12995 (N_12995,N_12809,N_12755);
and U12996 (N_12996,N_12736,N_12743);
or U12997 (N_12997,N_12796,N_12757);
and U12998 (N_12998,N_12807,N_12678);
or U12999 (N_12999,N_12686,N_12781);
or U13000 (N_13000,N_12787,N_12608);
and U13001 (N_13001,N_12889,N_12861);
nor U13002 (N_13002,N_12670,N_12625);
or U13003 (N_13003,N_12778,N_12741);
or U13004 (N_13004,N_12878,N_12696);
or U13005 (N_13005,N_12719,N_12752);
xor U13006 (N_13006,N_12739,N_12772);
nand U13007 (N_13007,N_12729,N_12759);
or U13008 (N_13008,N_12651,N_12636);
nor U13009 (N_13009,N_12656,N_12605);
or U13010 (N_13010,N_12735,N_12849);
xor U13011 (N_13011,N_12822,N_12872);
nor U13012 (N_13012,N_12664,N_12712);
nor U13013 (N_13013,N_12804,N_12615);
and U13014 (N_13014,N_12857,N_12612);
nor U13015 (N_13015,N_12620,N_12740);
and U13016 (N_13016,N_12895,N_12709);
nor U13017 (N_13017,N_12738,N_12880);
and U13018 (N_13018,N_12674,N_12770);
and U13019 (N_13019,N_12658,N_12629);
or U13020 (N_13020,N_12716,N_12724);
or U13021 (N_13021,N_12869,N_12623);
or U13022 (N_13022,N_12761,N_12692);
xor U13023 (N_13023,N_12812,N_12830);
or U13024 (N_13024,N_12606,N_12730);
or U13025 (N_13025,N_12850,N_12779);
or U13026 (N_13026,N_12826,N_12792);
or U13027 (N_13027,N_12706,N_12637);
nand U13028 (N_13028,N_12780,N_12821);
xnor U13029 (N_13029,N_12773,N_12609);
nor U13030 (N_13030,N_12665,N_12793);
nor U13031 (N_13031,N_12795,N_12650);
nor U13032 (N_13032,N_12631,N_12751);
and U13033 (N_13033,N_12652,N_12769);
nand U13034 (N_13034,N_12749,N_12699);
nand U13035 (N_13035,N_12695,N_12852);
nand U13036 (N_13036,N_12797,N_12825);
nand U13037 (N_13037,N_12630,N_12627);
xnor U13038 (N_13038,N_12892,N_12640);
or U13039 (N_13039,N_12633,N_12715);
nand U13040 (N_13040,N_12727,N_12689);
and U13041 (N_13041,N_12744,N_12860);
or U13042 (N_13042,N_12784,N_12748);
and U13043 (N_13043,N_12802,N_12897);
or U13044 (N_13044,N_12775,N_12823);
xnor U13045 (N_13045,N_12776,N_12663);
nor U13046 (N_13046,N_12635,N_12834);
xnor U13047 (N_13047,N_12798,N_12882);
or U13048 (N_13048,N_12865,N_12641);
nand U13049 (N_13049,N_12721,N_12816);
nand U13050 (N_13050,N_12836,N_12848);
or U13051 (N_13051,N_12738,N_12850);
nand U13052 (N_13052,N_12705,N_12820);
xor U13053 (N_13053,N_12888,N_12761);
nand U13054 (N_13054,N_12882,N_12817);
or U13055 (N_13055,N_12898,N_12818);
or U13056 (N_13056,N_12874,N_12872);
xnor U13057 (N_13057,N_12749,N_12893);
or U13058 (N_13058,N_12806,N_12788);
or U13059 (N_13059,N_12836,N_12792);
xnor U13060 (N_13060,N_12649,N_12704);
xor U13061 (N_13061,N_12656,N_12719);
and U13062 (N_13062,N_12683,N_12674);
and U13063 (N_13063,N_12809,N_12601);
nand U13064 (N_13064,N_12814,N_12681);
nor U13065 (N_13065,N_12808,N_12623);
nand U13066 (N_13066,N_12625,N_12877);
and U13067 (N_13067,N_12641,N_12701);
and U13068 (N_13068,N_12674,N_12667);
and U13069 (N_13069,N_12651,N_12745);
xor U13070 (N_13070,N_12608,N_12700);
xor U13071 (N_13071,N_12806,N_12864);
xnor U13072 (N_13072,N_12646,N_12603);
and U13073 (N_13073,N_12718,N_12839);
xnor U13074 (N_13074,N_12704,N_12806);
xnor U13075 (N_13075,N_12753,N_12871);
nand U13076 (N_13076,N_12681,N_12758);
nor U13077 (N_13077,N_12638,N_12852);
and U13078 (N_13078,N_12621,N_12791);
xnor U13079 (N_13079,N_12852,N_12765);
nor U13080 (N_13080,N_12606,N_12800);
and U13081 (N_13081,N_12743,N_12710);
xor U13082 (N_13082,N_12755,N_12866);
or U13083 (N_13083,N_12716,N_12758);
xor U13084 (N_13084,N_12721,N_12739);
nand U13085 (N_13085,N_12685,N_12756);
xor U13086 (N_13086,N_12876,N_12779);
nor U13087 (N_13087,N_12699,N_12793);
and U13088 (N_13088,N_12760,N_12670);
nand U13089 (N_13089,N_12610,N_12613);
nor U13090 (N_13090,N_12746,N_12682);
and U13091 (N_13091,N_12798,N_12885);
nand U13092 (N_13092,N_12899,N_12846);
nor U13093 (N_13093,N_12776,N_12814);
or U13094 (N_13094,N_12664,N_12655);
xor U13095 (N_13095,N_12868,N_12636);
nand U13096 (N_13096,N_12616,N_12625);
nor U13097 (N_13097,N_12776,N_12847);
or U13098 (N_13098,N_12685,N_12838);
and U13099 (N_13099,N_12647,N_12774);
or U13100 (N_13100,N_12690,N_12773);
or U13101 (N_13101,N_12783,N_12658);
nand U13102 (N_13102,N_12855,N_12798);
nand U13103 (N_13103,N_12652,N_12656);
nand U13104 (N_13104,N_12715,N_12710);
or U13105 (N_13105,N_12759,N_12683);
xor U13106 (N_13106,N_12870,N_12696);
xnor U13107 (N_13107,N_12826,N_12814);
xor U13108 (N_13108,N_12679,N_12711);
nor U13109 (N_13109,N_12600,N_12685);
nand U13110 (N_13110,N_12810,N_12858);
or U13111 (N_13111,N_12747,N_12687);
and U13112 (N_13112,N_12601,N_12720);
nor U13113 (N_13113,N_12613,N_12622);
nand U13114 (N_13114,N_12606,N_12778);
xor U13115 (N_13115,N_12804,N_12898);
and U13116 (N_13116,N_12604,N_12618);
nor U13117 (N_13117,N_12650,N_12660);
nor U13118 (N_13118,N_12675,N_12611);
and U13119 (N_13119,N_12671,N_12627);
and U13120 (N_13120,N_12632,N_12800);
nor U13121 (N_13121,N_12746,N_12767);
nor U13122 (N_13122,N_12718,N_12860);
xnor U13123 (N_13123,N_12701,N_12673);
nor U13124 (N_13124,N_12889,N_12629);
or U13125 (N_13125,N_12843,N_12658);
xnor U13126 (N_13126,N_12835,N_12843);
nand U13127 (N_13127,N_12698,N_12797);
xnor U13128 (N_13128,N_12864,N_12646);
or U13129 (N_13129,N_12720,N_12651);
nor U13130 (N_13130,N_12684,N_12647);
nand U13131 (N_13131,N_12698,N_12643);
or U13132 (N_13132,N_12676,N_12863);
nor U13133 (N_13133,N_12773,N_12727);
nor U13134 (N_13134,N_12644,N_12685);
and U13135 (N_13135,N_12776,N_12757);
nand U13136 (N_13136,N_12643,N_12751);
or U13137 (N_13137,N_12691,N_12722);
nand U13138 (N_13138,N_12657,N_12679);
and U13139 (N_13139,N_12602,N_12675);
and U13140 (N_13140,N_12614,N_12755);
or U13141 (N_13141,N_12705,N_12696);
or U13142 (N_13142,N_12751,N_12752);
nor U13143 (N_13143,N_12809,N_12708);
and U13144 (N_13144,N_12600,N_12657);
nand U13145 (N_13145,N_12781,N_12613);
xnor U13146 (N_13146,N_12874,N_12835);
xnor U13147 (N_13147,N_12890,N_12717);
xor U13148 (N_13148,N_12688,N_12700);
nand U13149 (N_13149,N_12800,N_12689);
nand U13150 (N_13150,N_12671,N_12801);
and U13151 (N_13151,N_12835,N_12808);
xor U13152 (N_13152,N_12614,N_12819);
or U13153 (N_13153,N_12876,N_12610);
nor U13154 (N_13154,N_12755,N_12847);
nand U13155 (N_13155,N_12891,N_12732);
and U13156 (N_13156,N_12860,N_12707);
nor U13157 (N_13157,N_12644,N_12642);
xor U13158 (N_13158,N_12834,N_12655);
and U13159 (N_13159,N_12722,N_12776);
or U13160 (N_13160,N_12613,N_12649);
nor U13161 (N_13161,N_12632,N_12893);
nor U13162 (N_13162,N_12685,N_12741);
nand U13163 (N_13163,N_12745,N_12640);
xnor U13164 (N_13164,N_12730,N_12893);
nor U13165 (N_13165,N_12862,N_12882);
nor U13166 (N_13166,N_12849,N_12788);
and U13167 (N_13167,N_12668,N_12623);
nand U13168 (N_13168,N_12824,N_12657);
and U13169 (N_13169,N_12797,N_12692);
nand U13170 (N_13170,N_12855,N_12664);
and U13171 (N_13171,N_12778,N_12686);
nand U13172 (N_13172,N_12875,N_12871);
nand U13173 (N_13173,N_12611,N_12615);
xnor U13174 (N_13174,N_12606,N_12715);
nor U13175 (N_13175,N_12851,N_12714);
xnor U13176 (N_13176,N_12767,N_12681);
nor U13177 (N_13177,N_12704,N_12675);
or U13178 (N_13178,N_12780,N_12839);
nand U13179 (N_13179,N_12680,N_12806);
or U13180 (N_13180,N_12615,N_12687);
nand U13181 (N_13181,N_12683,N_12768);
and U13182 (N_13182,N_12619,N_12714);
nor U13183 (N_13183,N_12675,N_12865);
and U13184 (N_13184,N_12665,N_12829);
or U13185 (N_13185,N_12895,N_12795);
and U13186 (N_13186,N_12749,N_12662);
and U13187 (N_13187,N_12729,N_12818);
nand U13188 (N_13188,N_12897,N_12697);
nor U13189 (N_13189,N_12831,N_12657);
xnor U13190 (N_13190,N_12805,N_12875);
nand U13191 (N_13191,N_12767,N_12755);
xor U13192 (N_13192,N_12717,N_12839);
and U13193 (N_13193,N_12871,N_12788);
or U13194 (N_13194,N_12731,N_12600);
nor U13195 (N_13195,N_12627,N_12631);
xor U13196 (N_13196,N_12653,N_12716);
and U13197 (N_13197,N_12744,N_12896);
or U13198 (N_13198,N_12605,N_12634);
nand U13199 (N_13199,N_12623,N_12896);
and U13200 (N_13200,N_12928,N_13008);
nand U13201 (N_13201,N_12940,N_13038);
nand U13202 (N_13202,N_12965,N_13062);
or U13203 (N_13203,N_13033,N_13148);
or U13204 (N_13204,N_12932,N_12971);
xnor U13205 (N_13205,N_12964,N_12995);
nor U13206 (N_13206,N_13144,N_13133);
nor U13207 (N_13207,N_12930,N_12920);
nor U13208 (N_13208,N_12917,N_13034);
xnor U13209 (N_13209,N_13183,N_12931);
nor U13210 (N_13210,N_12956,N_13054);
nand U13211 (N_13211,N_12985,N_13177);
and U13212 (N_13212,N_13128,N_13103);
xnor U13213 (N_13213,N_12982,N_13086);
nor U13214 (N_13214,N_13190,N_12915);
xor U13215 (N_13215,N_13136,N_13021);
and U13216 (N_13216,N_12904,N_13124);
or U13217 (N_13217,N_12970,N_13149);
xor U13218 (N_13218,N_12979,N_13053);
nand U13219 (N_13219,N_13041,N_13057);
or U13220 (N_13220,N_13173,N_13096);
nand U13221 (N_13221,N_13058,N_13176);
xnor U13222 (N_13222,N_12968,N_13055);
xor U13223 (N_13223,N_13040,N_13090);
and U13224 (N_13224,N_13078,N_12903);
xor U13225 (N_13225,N_13016,N_12951);
and U13226 (N_13226,N_12955,N_12948);
or U13227 (N_13227,N_13023,N_13061);
nor U13228 (N_13228,N_13032,N_13025);
nand U13229 (N_13229,N_13168,N_13093);
xor U13230 (N_13230,N_13115,N_13001);
and U13231 (N_13231,N_12952,N_12937);
and U13232 (N_13232,N_13044,N_13082);
and U13233 (N_13233,N_13091,N_13153);
xor U13234 (N_13234,N_13046,N_13026);
xor U13235 (N_13235,N_13193,N_13106);
or U13236 (N_13236,N_12991,N_13129);
xor U13237 (N_13237,N_12916,N_12913);
nand U13238 (N_13238,N_13101,N_13151);
and U13239 (N_13239,N_13035,N_13198);
xnor U13240 (N_13240,N_13045,N_13050);
xnor U13241 (N_13241,N_13126,N_12962);
and U13242 (N_13242,N_12901,N_13132);
nor U13243 (N_13243,N_13105,N_12933);
nand U13244 (N_13244,N_12973,N_13108);
nand U13245 (N_13245,N_12925,N_12987);
or U13246 (N_13246,N_13157,N_12997);
nand U13247 (N_13247,N_12988,N_13127);
and U13248 (N_13248,N_13150,N_12963);
nor U13249 (N_13249,N_13083,N_13122);
and U13250 (N_13250,N_12954,N_12939);
or U13251 (N_13251,N_13161,N_13039);
or U13252 (N_13252,N_13068,N_13081);
or U13253 (N_13253,N_13043,N_13158);
or U13254 (N_13254,N_12953,N_13194);
and U13255 (N_13255,N_13002,N_12942);
and U13256 (N_13256,N_12958,N_12992);
nand U13257 (N_13257,N_12934,N_12935);
or U13258 (N_13258,N_13175,N_12900);
nand U13259 (N_13259,N_13130,N_13089);
or U13260 (N_13260,N_13165,N_13195);
nor U13261 (N_13261,N_12922,N_13007);
or U13262 (N_13262,N_13010,N_13042);
xor U13263 (N_13263,N_12906,N_13076);
nand U13264 (N_13264,N_12936,N_13072);
and U13265 (N_13265,N_12957,N_12912);
and U13266 (N_13266,N_13020,N_13135);
nor U13267 (N_13267,N_13013,N_13147);
nand U13268 (N_13268,N_13169,N_13174);
nand U13269 (N_13269,N_12924,N_13167);
and U13270 (N_13270,N_13071,N_13030);
nand U13271 (N_13271,N_13067,N_12946);
and U13272 (N_13272,N_13180,N_13199);
or U13273 (N_13273,N_13065,N_12918);
nand U13274 (N_13274,N_13184,N_13029);
nand U13275 (N_13275,N_13171,N_12908);
or U13276 (N_13276,N_12984,N_13100);
xnor U13277 (N_13277,N_12910,N_13121);
and U13278 (N_13278,N_13185,N_13036);
nand U13279 (N_13279,N_12977,N_13017);
or U13280 (N_13280,N_13181,N_13162);
and U13281 (N_13281,N_13024,N_13156);
or U13282 (N_13282,N_13085,N_13154);
and U13283 (N_13283,N_13170,N_12950);
nor U13284 (N_13284,N_13131,N_13070);
xor U13285 (N_13285,N_13004,N_13123);
xnor U13286 (N_13286,N_13074,N_13116);
or U13287 (N_13287,N_13117,N_13143);
xor U13288 (N_13288,N_13139,N_13092);
or U13289 (N_13289,N_13012,N_13107);
nor U13290 (N_13290,N_12996,N_13052);
nor U13291 (N_13291,N_13178,N_13060);
or U13292 (N_13292,N_13075,N_12949);
nand U13293 (N_13293,N_13087,N_13189);
or U13294 (N_13294,N_13112,N_12981);
nor U13295 (N_13295,N_13159,N_12907);
nand U13296 (N_13296,N_13006,N_13099);
nor U13297 (N_13297,N_12967,N_12975);
and U13298 (N_13298,N_13137,N_13119);
nand U13299 (N_13299,N_13152,N_13186);
nor U13300 (N_13300,N_12919,N_13097);
xor U13301 (N_13301,N_13003,N_13164);
or U13302 (N_13302,N_13118,N_13109);
nor U13303 (N_13303,N_13037,N_12993);
nor U13304 (N_13304,N_13179,N_12990);
nand U13305 (N_13305,N_13094,N_13048);
nand U13306 (N_13306,N_12944,N_13011);
nor U13307 (N_13307,N_13192,N_12914);
and U13308 (N_13308,N_12983,N_13142);
and U13309 (N_13309,N_12960,N_13166);
or U13310 (N_13310,N_13015,N_12974);
or U13311 (N_13311,N_13120,N_13146);
and U13312 (N_13312,N_13069,N_13073);
xnor U13313 (N_13313,N_13172,N_13114);
xnor U13314 (N_13314,N_13028,N_12989);
and U13315 (N_13315,N_13080,N_13051);
xnor U13316 (N_13316,N_13188,N_12943);
or U13317 (N_13317,N_13187,N_13000);
and U13318 (N_13318,N_13019,N_13104);
nand U13319 (N_13319,N_13056,N_12921);
nand U13320 (N_13320,N_13088,N_13022);
nor U13321 (N_13321,N_12978,N_12911);
xor U13322 (N_13322,N_12961,N_13098);
nand U13323 (N_13323,N_12947,N_13077);
and U13324 (N_13324,N_12969,N_13138);
nor U13325 (N_13325,N_12994,N_12923);
nor U13326 (N_13326,N_12938,N_13182);
nand U13327 (N_13327,N_12929,N_12926);
nor U13328 (N_13328,N_13155,N_13064);
xor U13329 (N_13329,N_13111,N_13160);
and U13330 (N_13330,N_13196,N_13014);
and U13331 (N_13331,N_12945,N_12999);
and U13332 (N_13332,N_13005,N_13145);
xor U13333 (N_13333,N_13140,N_12927);
and U13334 (N_13334,N_13191,N_12905);
and U13335 (N_13335,N_13102,N_13009);
nand U13336 (N_13336,N_12959,N_13066);
nor U13337 (N_13337,N_13018,N_13059);
nand U13338 (N_13338,N_13141,N_12976);
and U13339 (N_13339,N_13084,N_13031);
or U13340 (N_13340,N_12902,N_13095);
nand U13341 (N_13341,N_12909,N_12966);
and U13342 (N_13342,N_13110,N_12998);
nand U13343 (N_13343,N_13047,N_12980);
or U13344 (N_13344,N_13027,N_13079);
nand U13345 (N_13345,N_13049,N_12986);
or U13346 (N_13346,N_13163,N_13125);
nor U13347 (N_13347,N_13134,N_13113);
nand U13348 (N_13348,N_13197,N_12972);
and U13349 (N_13349,N_12941,N_13063);
nor U13350 (N_13350,N_13119,N_13169);
nand U13351 (N_13351,N_13167,N_13138);
nand U13352 (N_13352,N_13195,N_13158);
or U13353 (N_13353,N_13057,N_13087);
and U13354 (N_13354,N_12939,N_12965);
nand U13355 (N_13355,N_13016,N_13163);
or U13356 (N_13356,N_12950,N_13143);
nand U13357 (N_13357,N_13103,N_12987);
xor U13358 (N_13358,N_13161,N_13186);
nor U13359 (N_13359,N_12913,N_12979);
nor U13360 (N_13360,N_13022,N_13124);
xnor U13361 (N_13361,N_13093,N_12977);
and U13362 (N_13362,N_12947,N_13085);
nand U13363 (N_13363,N_12960,N_12916);
and U13364 (N_13364,N_13142,N_13083);
nor U13365 (N_13365,N_13134,N_13044);
nor U13366 (N_13366,N_13101,N_13199);
or U13367 (N_13367,N_13143,N_12930);
and U13368 (N_13368,N_12956,N_13196);
nand U13369 (N_13369,N_12928,N_13115);
and U13370 (N_13370,N_12924,N_13078);
xnor U13371 (N_13371,N_12964,N_13018);
and U13372 (N_13372,N_12908,N_13066);
or U13373 (N_13373,N_12996,N_12904);
nand U13374 (N_13374,N_13050,N_13187);
or U13375 (N_13375,N_13111,N_12952);
and U13376 (N_13376,N_12919,N_13123);
xnor U13377 (N_13377,N_13055,N_13030);
and U13378 (N_13378,N_13047,N_13111);
xor U13379 (N_13379,N_13088,N_12920);
nor U13380 (N_13380,N_13002,N_13087);
nand U13381 (N_13381,N_13038,N_12985);
or U13382 (N_13382,N_13169,N_13160);
and U13383 (N_13383,N_13090,N_12968);
or U13384 (N_13384,N_13162,N_12951);
nand U13385 (N_13385,N_12988,N_12993);
or U13386 (N_13386,N_13002,N_13003);
or U13387 (N_13387,N_13125,N_13112);
nor U13388 (N_13388,N_12980,N_12905);
and U13389 (N_13389,N_12947,N_12992);
nand U13390 (N_13390,N_13073,N_12954);
xnor U13391 (N_13391,N_13185,N_13139);
nor U13392 (N_13392,N_12988,N_13077);
and U13393 (N_13393,N_13171,N_12935);
nand U13394 (N_13394,N_13041,N_12928);
or U13395 (N_13395,N_13125,N_12949);
and U13396 (N_13396,N_13084,N_12918);
and U13397 (N_13397,N_13074,N_13014);
or U13398 (N_13398,N_13183,N_13079);
and U13399 (N_13399,N_13065,N_12901);
xnor U13400 (N_13400,N_13052,N_13117);
or U13401 (N_13401,N_12947,N_13185);
nor U13402 (N_13402,N_12981,N_13072);
and U13403 (N_13403,N_13089,N_13075);
nor U13404 (N_13404,N_13068,N_12998);
and U13405 (N_13405,N_12939,N_13028);
and U13406 (N_13406,N_13135,N_13057);
xor U13407 (N_13407,N_13024,N_13007);
nand U13408 (N_13408,N_13016,N_13073);
and U13409 (N_13409,N_13041,N_13081);
xnor U13410 (N_13410,N_12960,N_12918);
nor U13411 (N_13411,N_13067,N_12959);
and U13412 (N_13412,N_12909,N_12940);
xor U13413 (N_13413,N_12986,N_13067);
nand U13414 (N_13414,N_13145,N_12919);
nand U13415 (N_13415,N_13148,N_13184);
and U13416 (N_13416,N_12937,N_13173);
and U13417 (N_13417,N_13155,N_13096);
and U13418 (N_13418,N_13099,N_13199);
nor U13419 (N_13419,N_13186,N_13009);
nor U13420 (N_13420,N_13009,N_13139);
nor U13421 (N_13421,N_12940,N_12900);
xnor U13422 (N_13422,N_13171,N_12929);
nand U13423 (N_13423,N_12955,N_13190);
and U13424 (N_13424,N_13001,N_13154);
or U13425 (N_13425,N_13047,N_13149);
nor U13426 (N_13426,N_13126,N_12981);
xor U13427 (N_13427,N_13004,N_13021);
or U13428 (N_13428,N_12976,N_13036);
nor U13429 (N_13429,N_12923,N_13053);
xor U13430 (N_13430,N_12960,N_13130);
nand U13431 (N_13431,N_13111,N_12953);
nor U13432 (N_13432,N_13109,N_13065);
xnor U13433 (N_13433,N_13196,N_13030);
or U13434 (N_13434,N_12948,N_12903);
xor U13435 (N_13435,N_13075,N_13194);
nor U13436 (N_13436,N_13156,N_13199);
and U13437 (N_13437,N_13072,N_12999);
or U13438 (N_13438,N_13069,N_13190);
xor U13439 (N_13439,N_13126,N_13178);
and U13440 (N_13440,N_12925,N_13159);
nand U13441 (N_13441,N_13159,N_13051);
and U13442 (N_13442,N_12971,N_13054);
or U13443 (N_13443,N_12934,N_12975);
or U13444 (N_13444,N_13189,N_12949);
and U13445 (N_13445,N_13048,N_12949);
xor U13446 (N_13446,N_13165,N_12957);
xnor U13447 (N_13447,N_13060,N_13101);
or U13448 (N_13448,N_13182,N_13033);
nand U13449 (N_13449,N_13134,N_12929);
nor U13450 (N_13450,N_13132,N_12958);
or U13451 (N_13451,N_12964,N_13069);
or U13452 (N_13452,N_12964,N_13146);
nor U13453 (N_13453,N_13106,N_13052);
or U13454 (N_13454,N_13051,N_13107);
or U13455 (N_13455,N_12962,N_13071);
nand U13456 (N_13456,N_13028,N_13096);
or U13457 (N_13457,N_13138,N_13019);
and U13458 (N_13458,N_13072,N_13082);
nor U13459 (N_13459,N_13038,N_12943);
or U13460 (N_13460,N_13154,N_13087);
and U13461 (N_13461,N_13076,N_12935);
and U13462 (N_13462,N_13128,N_13190);
xnor U13463 (N_13463,N_12944,N_13143);
and U13464 (N_13464,N_13166,N_13118);
or U13465 (N_13465,N_13166,N_13109);
nand U13466 (N_13466,N_13107,N_12945);
and U13467 (N_13467,N_12993,N_13121);
xnor U13468 (N_13468,N_12931,N_13155);
xor U13469 (N_13469,N_12934,N_13046);
nand U13470 (N_13470,N_13111,N_13061);
and U13471 (N_13471,N_13102,N_13112);
and U13472 (N_13472,N_12984,N_13101);
and U13473 (N_13473,N_13053,N_12907);
xor U13474 (N_13474,N_13170,N_13040);
and U13475 (N_13475,N_12932,N_12931);
or U13476 (N_13476,N_13003,N_13193);
nand U13477 (N_13477,N_13112,N_12992);
and U13478 (N_13478,N_13005,N_12954);
xor U13479 (N_13479,N_12998,N_12936);
nand U13480 (N_13480,N_13085,N_12927);
and U13481 (N_13481,N_12916,N_13021);
nand U13482 (N_13482,N_13065,N_12922);
nor U13483 (N_13483,N_13122,N_13151);
xnor U13484 (N_13484,N_12954,N_13086);
or U13485 (N_13485,N_13069,N_13047);
nor U13486 (N_13486,N_13006,N_13008);
or U13487 (N_13487,N_13088,N_12935);
xor U13488 (N_13488,N_13192,N_13141);
or U13489 (N_13489,N_13092,N_12980);
nand U13490 (N_13490,N_13031,N_12994);
xor U13491 (N_13491,N_13033,N_13045);
xnor U13492 (N_13492,N_13085,N_13050);
or U13493 (N_13493,N_12930,N_13074);
nand U13494 (N_13494,N_13193,N_13131);
or U13495 (N_13495,N_13007,N_13034);
nand U13496 (N_13496,N_13015,N_12981);
xor U13497 (N_13497,N_12950,N_13176);
or U13498 (N_13498,N_12931,N_13056);
or U13499 (N_13499,N_13080,N_13158);
and U13500 (N_13500,N_13223,N_13435);
xnor U13501 (N_13501,N_13438,N_13332);
or U13502 (N_13502,N_13497,N_13443);
nand U13503 (N_13503,N_13246,N_13401);
nand U13504 (N_13504,N_13292,N_13330);
xnor U13505 (N_13505,N_13200,N_13300);
nand U13506 (N_13506,N_13262,N_13203);
xnor U13507 (N_13507,N_13419,N_13375);
nor U13508 (N_13508,N_13467,N_13368);
or U13509 (N_13509,N_13316,N_13477);
or U13510 (N_13510,N_13301,N_13232);
nand U13511 (N_13511,N_13282,N_13221);
xnor U13512 (N_13512,N_13474,N_13204);
nand U13513 (N_13513,N_13354,N_13385);
nand U13514 (N_13514,N_13257,N_13266);
xnor U13515 (N_13515,N_13289,N_13376);
nand U13516 (N_13516,N_13444,N_13413);
nor U13517 (N_13517,N_13455,N_13346);
or U13518 (N_13518,N_13270,N_13422);
or U13519 (N_13519,N_13338,N_13358);
nand U13520 (N_13520,N_13252,N_13233);
nand U13521 (N_13521,N_13320,N_13388);
nand U13522 (N_13522,N_13315,N_13234);
nor U13523 (N_13523,N_13275,N_13253);
or U13524 (N_13524,N_13243,N_13420);
or U13525 (N_13525,N_13448,N_13302);
xnor U13526 (N_13526,N_13441,N_13475);
nand U13527 (N_13527,N_13206,N_13484);
nand U13528 (N_13528,N_13481,N_13260);
or U13529 (N_13529,N_13407,N_13214);
xor U13530 (N_13530,N_13499,N_13294);
or U13531 (N_13531,N_13344,N_13361);
nand U13532 (N_13532,N_13379,N_13331);
or U13533 (N_13533,N_13416,N_13212);
nand U13534 (N_13534,N_13390,N_13482);
xor U13535 (N_13535,N_13210,N_13264);
nand U13536 (N_13536,N_13363,N_13383);
nor U13537 (N_13537,N_13318,N_13319);
xnor U13538 (N_13538,N_13227,N_13498);
and U13539 (N_13539,N_13213,N_13286);
and U13540 (N_13540,N_13433,N_13360);
xnor U13541 (N_13541,N_13340,N_13327);
or U13542 (N_13542,N_13237,N_13485);
or U13543 (N_13543,N_13201,N_13426);
and U13544 (N_13544,N_13312,N_13272);
or U13545 (N_13545,N_13391,N_13347);
or U13546 (N_13546,N_13240,N_13290);
nor U13547 (N_13547,N_13356,N_13269);
or U13548 (N_13548,N_13392,N_13247);
or U13549 (N_13549,N_13487,N_13215);
and U13550 (N_13550,N_13350,N_13271);
or U13551 (N_13551,N_13362,N_13397);
nand U13552 (N_13552,N_13229,N_13295);
nor U13553 (N_13553,N_13235,N_13418);
nand U13554 (N_13554,N_13406,N_13461);
and U13555 (N_13555,N_13445,N_13472);
xor U13556 (N_13556,N_13447,N_13432);
or U13557 (N_13557,N_13216,N_13408);
nor U13558 (N_13558,N_13403,N_13278);
or U13559 (N_13559,N_13274,N_13249);
or U13560 (N_13560,N_13202,N_13491);
and U13561 (N_13561,N_13304,N_13226);
or U13562 (N_13562,N_13306,N_13337);
nor U13563 (N_13563,N_13369,N_13393);
nor U13564 (N_13564,N_13440,N_13421);
nor U13565 (N_13565,N_13409,N_13373);
nor U13566 (N_13566,N_13458,N_13366);
nand U13567 (N_13567,N_13353,N_13483);
nor U13568 (N_13568,N_13277,N_13329);
nor U13569 (N_13569,N_13322,N_13317);
and U13570 (N_13570,N_13244,N_13311);
nand U13571 (N_13571,N_13470,N_13450);
nor U13572 (N_13572,N_13442,N_13449);
or U13573 (N_13573,N_13381,N_13384);
nand U13574 (N_13574,N_13281,N_13374);
xor U13575 (N_13575,N_13211,N_13417);
nor U13576 (N_13576,N_13446,N_13437);
or U13577 (N_13577,N_13427,N_13410);
nand U13578 (N_13578,N_13325,N_13411);
xnor U13579 (N_13579,N_13267,N_13473);
and U13580 (N_13580,N_13434,N_13404);
or U13581 (N_13581,N_13241,N_13280);
and U13582 (N_13582,N_13464,N_13298);
nand U13583 (N_13583,N_13256,N_13231);
nor U13584 (N_13584,N_13238,N_13293);
and U13585 (N_13585,N_13396,N_13465);
nand U13586 (N_13586,N_13326,N_13299);
or U13587 (N_13587,N_13323,N_13400);
and U13588 (N_13588,N_13310,N_13431);
nand U13589 (N_13589,N_13436,N_13335);
or U13590 (N_13590,N_13398,N_13394);
or U13591 (N_13591,N_13334,N_13314);
nor U13592 (N_13592,N_13424,N_13205);
and U13593 (N_13593,N_13471,N_13288);
xor U13594 (N_13594,N_13251,N_13462);
or U13595 (N_13595,N_13222,N_13415);
xor U13596 (N_13596,N_13218,N_13254);
xor U13597 (N_13597,N_13261,N_13248);
and U13598 (N_13598,N_13342,N_13303);
xor U13599 (N_13599,N_13242,N_13452);
and U13600 (N_13600,N_13328,N_13297);
or U13601 (N_13601,N_13495,N_13307);
nand U13602 (N_13602,N_13245,N_13490);
xor U13603 (N_13603,N_13460,N_13469);
nand U13604 (N_13604,N_13339,N_13321);
or U13605 (N_13605,N_13333,N_13228);
and U13606 (N_13606,N_13486,N_13456);
or U13607 (N_13607,N_13355,N_13402);
and U13608 (N_13608,N_13341,N_13287);
nor U13609 (N_13609,N_13428,N_13479);
nor U13610 (N_13610,N_13225,N_13208);
nor U13611 (N_13611,N_13496,N_13305);
nand U13612 (N_13612,N_13259,N_13258);
or U13613 (N_13613,N_13357,N_13367);
or U13614 (N_13614,N_13364,N_13453);
or U13615 (N_13615,N_13352,N_13399);
nor U13616 (N_13616,N_13239,N_13372);
xor U13617 (N_13617,N_13273,N_13359);
nand U13618 (N_13618,N_13389,N_13351);
nor U13619 (N_13619,N_13425,N_13378);
or U13620 (N_13620,N_13412,N_13429);
and U13621 (N_13621,N_13336,N_13370);
nor U13622 (N_13622,N_13387,N_13349);
and U13623 (N_13623,N_13459,N_13457);
or U13624 (N_13624,N_13296,N_13377);
xor U13625 (N_13625,N_13492,N_13324);
or U13626 (N_13626,N_13309,N_13430);
xor U13627 (N_13627,N_13494,N_13466);
or U13628 (N_13628,N_13283,N_13439);
nand U13629 (N_13629,N_13284,N_13454);
xnor U13630 (N_13630,N_13268,N_13343);
xor U13631 (N_13631,N_13285,N_13476);
nand U13632 (N_13632,N_13365,N_13217);
xor U13633 (N_13633,N_13308,N_13348);
nor U13634 (N_13634,N_13395,N_13423);
nor U13635 (N_13635,N_13279,N_13451);
nor U13636 (N_13636,N_13313,N_13463);
xnor U13637 (N_13637,N_13386,N_13224);
nor U13638 (N_13638,N_13414,N_13493);
nor U13639 (N_13639,N_13265,N_13255);
nand U13640 (N_13640,N_13219,N_13405);
xnor U13641 (N_13641,N_13380,N_13220);
xor U13642 (N_13642,N_13276,N_13207);
and U13643 (N_13643,N_13345,N_13480);
nand U13644 (N_13644,N_13291,N_13209);
or U13645 (N_13645,N_13468,N_13263);
and U13646 (N_13646,N_13488,N_13382);
and U13647 (N_13647,N_13478,N_13489);
xor U13648 (N_13648,N_13230,N_13236);
xor U13649 (N_13649,N_13250,N_13371);
nand U13650 (N_13650,N_13312,N_13473);
xnor U13651 (N_13651,N_13368,N_13287);
or U13652 (N_13652,N_13274,N_13327);
and U13653 (N_13653,N_13445,N_13433);
nor U13654 (N_13654,N_13326,N_13362);
nand U13655 (N_13655,N_13441,N_13411);
nand U13656 (N_13656,N_13468,N_13274);
or U13657 (N_13657,N_13395,N_13250);
and U13658 (N_13658,N_13436,N_13255);
nor U13659 (N_13659,N_13262,N_13456);
and U13660 (N_13660,N_13413,N_13327);
or U13661 (N_13661,N_13472,N_13455);
or U13662 (N_13662,N_13270,N_13313);
nand U13663 (N_13663,N_13321,N_13212);
or U13664 (N_13664,N_13273,N_13239);
or U13665 (N_13665,N_13265,N_13398);
and U13666 (N_13666,N_13237,N_13423);
xnor U13667 (N_13667,N_13233,N_13208);
xnor U13668 (N_13668,N_13359,N_13223);
xor U13669 (N_13669,N_13276,N_13397);
and U13670 (N_13670,N_13235,N_13283);
and U13671 (N_13671,N_13405,N_13358);
or U13672 (N_13672,N_13255,N_13486);
or U13673 (N_13673,N_13202,N_13242);
xnor U13674 (N_13674,N_13456,N_13404);
nor U13675 (N_13675,N_13306,N_13454);
nor U13676 (N_13676,N_13448,N_13436);
and U13677 (N_13677,N_13366,N_13360);
or U13678 (N_13678,N_13288,N_13269);
or U13679 (N_13679,N_13360,N_13420);
or U13680 (N_13680,N_13205,N_13364);
nand U13681 (N_13681,N_13315,N_13259);
nor U13682 (N_13682,N_13414,N_13449);
or U13683 (N_13683,N_13291,N_13269);
or U13684 (N_13684,N_13208,N_13487);
and U13685 (N_13685,N_13474,N_13212);
or U13686 (N_13686,N_13477,N_13344);
and U13687 (N_13687,N_13289,N_13464);
or U13688 (N_13688,N_13209,N_13476);
nor U13689 (N_13689,N_13342,N_13333);
and U13690 (N_13690,N_13229,N_13271);
and U13691 (N_13691,N_13253,N_13395);
or U13692 (N_13692,N_13369,N_13365);
nor U13693 (N_13693,N_13273,N_13263);
nand U13694 (N_13694,N_13382,N_13448);
or U13695 (N_13695,N_13415,N_13409);
xor U13696 (N_13696,N_13443,N_13269);
or U13697 (N_13697,N_13301,N_13488);
xnor U13698 (N_13698,N_13251,N_13456);
xnor U13699 (N_13699,N_13313,N_13271);
nor U13700 (N_13700,N_13306,N_13422);
nor U13701 (N_13701,N_13351,N_13241);
nor U13702 (N_13702,N_13221,N_13245);
nand U13703 (N_13703,N_13393,N_13240);
nor U13704 (N_13704,N_13224,N_13221);
or U13705 (N_13705,N_13322,N_13483);
xnor U13706 (N_13706,N_13351,N_13361);
and U13707 (N_13707,N_13435,N_13424);
nand U13708 (N_13708,N_13481,N_13203);
nand U13709 (N_13709,N_13236,N_13429);
nor U13710 (N_13710,N_13322,N_13315);
xnor U13711 (N_13711,N_13238,N_13377);
nand U13712 (N_13712,N_13263,N_13318);
or U13713 (N_13713,N_13342,N_13270);
or U13714 (N_13714,N_13292,N_13464);
xor U13715 (N_13715,N_13244,N_13433);
or U13716 (N_13716,N_13440,N_13362);
or U13717 (N_13717,N_13499,N_13363);
nor U13718 (N_13718,N_13346,N_13495);
or U13719 (N_13719,N_13247,N_13461);
xor U13720 (N_13720,N_13209,N_13292);
nand U13721 (N_13721,N_13385,N_13474);
nor U13722 (N_13722,N_13457,N_13380);
nor U13723 (N_13723,N_13412,N_13484);
or U13724 (N_13724,N_13369,N_13450);
or U13725 (N_13725,N_13369,N_13305);
and U13726 (N_13726,N_13296,N_13354);
nand U13727 (N_13727,N_13389,N_13279);
and U13728 (N_13728,N_13476,N_13404);
nor U13729 (N_13729,N_13236,N_13297);
xor U13730 (N_13730,N_13345,N_13288);
or U13731 (N_13731,N_13262,N_13463);
xnor U13732 (N_13732,N_13349,N_13362);
nand U13733 (N_13733,N_13480,N_13253);
or U13734 (N_13734,N_13286,N_13400);
xor U13735 (N_13735,N_13243,N_13405);
nand U13736 (N_13736,N_13368,N_13355);
or U13737 (N_13737,N_13488,N_13403);
and U13738 (N_13738,N_13294,N_13366);
xor U13739 (N_13739,N_13237,N_13373);
nand U13740 (N_13740,N_13423,N_13405);
nor U13741 (N_13741,N_13218,N_13333);
or U13742 (N_13742,N_13290,N_13337);
nand U13743 (N_13743,N_13386,N_13481);
xnor U13744 (N_13744,N_13482,N_13284);
xor U13745 (N_13745,N_13473,N_13451);
nand U13746 (N_13746,N_13252,N_13487);
nor U13747 (N_13747,N_13240,N_13281);
nor U13748 (N_13748,N_13252,N_13492);
xor U13749 (N_13749,N_13366,N_13461);
xnor U13750 (N_13750,N_13410,N_13391);
nor U13751 (N_13751,N_13488,N_13383);
nand U13752 (N_13752,N_13387,N_13248);
or U13753 (N_13753,N_13414,N_13386);
or U13754 (N_13754,N_13226,N_13288);
or U13755 (N_13755,N_13347,N_13302);
and U13756 (N_13756,N_13283,N_13272);
xor U13757 (N_13757,N_13348,N_13265);
and U13758 (N_13758,N_13238,N_13218);
nand U13759 (N_13759,N_13450,N_13466);
nand U13760 (N_13760,N_13205,N_13432);
or U13761 (N_13761,N_13226,N_13261);
or U13762 (N_13762,N_13252,N_13288);
nand U13763 (N_13763,N_13402,N_13366);
xnor U13764 (N_13764,N_13285,N_13395);
nand U13765 (N_13765,N_13454,N_13404);
nand U13766 (N_13766,N_13499,N_13470);
nor U13767 (N_13767,N_13221,N_13271);
or U13768 (N_13768,N_13230,N_13234);
nand U13769 (N_13769,N_13271,N_13317);
or U13770 (N_13770,N_13404,N_13314);
nor U13771 (N_13771,N_13246,N_13299);
nand U13772 (N_13772,N_13331,N_13245);
and U13773 (N_13773,N_13267,N_13416);
xor U13774 (N_13774,N_13241,N_13292);
and U13775 (N_13775,N_13494,N_13284);
nand U13776 (N_13776,N_13476,N_13272);
nor U13777 (N_13777,N_13226,N_13361);
or U13778 (N_13778,N_13382,N_13227);
xnor U13779 (N_13779,N_13415,N_13446);
and U13780 (N_13780,N_13453,N_13354);
and U13781 (N_13781,N_13416,N_13324);
or U13782 (N_13782,N_13202,N_13458);
nor U13783 (N_13783,N_13342,N_13365);
nor U13784 (N_13784,N_13490,N_13357);
xor U13785 (N_13785,N_13218,N_13235);
nor U13786 (N_13786,N_13477,N_13359);
and U13787 (N_13787,N_13362,N_13377);
nand U13788 (N_13788,N_13244,N_13330);
nor U13789 (N_13789,N_13285,N_13220);
or U13790 (N_13790,N_13341,N_13210);
xor U13791 (N_13791,N_13464,N_13433);
nand U13792 (N_13792,N_13425,N_13265);
and U13793 (N_13793,N_13272,N_13306);
nor U13794 (N_13794,N_13428,N_13315);
xor U13795 (N_13795,N_13382,N_13251);
xnor U13796 (N_13796,N_13286,N_13282);
nor U13797 (N_13797,N_13245,N_13378);
nand U13798 (N_13798,N_13316,N_13270);
nand U13799 (N_13799,N_13393,N_13454);
and U13800 (N_13800,N_13522,N_13658);
nand U13801 (N_13801,N_13757,N_13562);
nand U13802 (N_13802,N_13755,N_13544);
xor U13803 (N_13803,N_13785,N_13670);
or U13804 (N_13804,N_13756,N_13650);
nand U13805 (N_13805,N_13586,N_13768);
and U13806 (N_13806,N_13682,N_13604);
nand U13807 (N_13807,N_13551,N_13745);
nor U13808 (N_13808,N_13517,N_13719);
nor U13809 (N_13809,N_13587,N_13527);
and U13810 (N_13810,N_13655,N_13644);
or U13811 (N_13811,N_13634,N_13704);
or U13812 (N_13812,N_13537,N_13688);
or U13813 (N_13813,N_13631,N_13573);
nor U13814 (N_13814,N_13730,N_13507);
and U13815 (N_13815,N_13572,N_13525);
nor U13816 (N_13816,N_13596,N_13740);
nor U13817 (N_13817,N_13514,N_13707);
xor U13818 (N_13818,N_13718,N_13541);
nor U13819 (N_13819,N_13524,N_13649);
nor U13820 (N_13820,N_13590,N_13646);
or U13821 (N_13821,N_13593,N_13619);
nor U13822 (N_13822,N_13661,N_13558);
xnor U13823 (N_13823,N_13595,N_13510);
nand U13824 (N_13824,N_13647,N_13766);
nor U13825 (N_13825,N_13518,N_13735);
xor U13826 (N_13826,N_13712,N_13615);
nor U13827 (N_13827,N_13648,N_13702);
nand U13828 (N_13828,N_13599,N_13790);
nor U13829 (N_13829,N_13552,N_13761);
nor U13830 (N_13830,N_13511,N_13577);
nand U13831 (N_13831,N_13654,N_13501);
nand U13832 (N_13832,N_13538,N_13695);
nand U13833 (N_13833,N_13564,N_13606);
or U13834 (N_13834,N_13771,N_13559);
or U13835 (N_13835,N_13721,N_13554);
nor U13836 (N_13836,N_13546,N_13685);
and U13837 (N_13837,N_13747,N_13767);
or U13838 (N_13838,N_13779,N_13513);
or U13839 (N_13839,N_13660,N_13545);
xor U13840 (N_13840,N_13502,N_13509);
nor U13841 (N_13841,N_13762,N_13746);
xnor U13842 (N_13842,N_13629,N_13722);
xnor U13843 (N_13843,N_13777,N_13597);
and U13844 (N_13844,N_13774,N_13549);
xor U13845 (N_13845,N_13673,N_13607);
and U13846 (N_13846,N_13582,N_13504);
nor U13847 (N_13847,N_13732,N_13625);
nor U13848 (N_13848,N_13679,N_13567);
xnor U13849 (N_13849,N_13566,N_13734);
nand U13850 (N_13850,N_13711,N_13754);
nor U13851 (N_13851,N_13653,N_13742);
nand U13852 (N_13852,N_13609,N_13640);
nand U13853 (N_13853,N_13556,N_13641);
nor U13854 (N_13854,N_13782,N_13540);
or U13855 (N_13855,N_13557,N_13716);
and U13856 (N_13856,N_13693,N_13781);
nand U13857 (N_13857,N_13612,N_13584);
and U13858 (N_13858,N_13605,N_13600);
nor U13859 (N_13859,N_13610,N_13713);
or U13860 (N_13860,N_13737,N_13548);
and U13861 (N_13861,N_13776,N_13698);
nor U13862 (N_13862,N_13534,N_13798);
xor U13863 (N_13863,N_13645,N_13733);
or U13864 (N_13864,N_13638,N_13555);
xnor U13865 (N_13865,N_13576,N_13611);
xnor U13866 (N_13866,N_13613,N_13731);
or U13867 (N_13867,N_13519,N_13563);
nand U13868 (N_13868,N_13694,N_13516);
nor U13869 (N_13869,N_13635,N_13775);
nor U13870 (N_13870,N_13784,N_13715);
or U13871 (N_13871,N_13574,N_13791);
nand U13872 (N_13872,N_13749,N_13750);
nand U13873 (N_13873,N_13580,N_13568);
nor U13874 (N_13874,N_13789,N_13575);
nand U13875 (N_13875,N_13520,N_13668);
or U13876 (N_13876,N_13748,N_13736);
nand U13877 (N_13877,N_13521,N_13585);
and U13878 (N_13878,N_13758,N_13508);
nand U13879 (N_13879,N_13724,N_13530);
xnor U13880 (N_13880,N_13594,N_13643);
xnor U13881 (N_13881,N_13793,N_13616);
nand U13882 (N_13882,N_13662,N_13583);
nand U13883 (N_13883,N_13536,N_13717);
or U13884 (N_13884,N_13759,N_13783);
nor U13885 (N_13885,N_13659,N_13651);
and U13886 (N_13886,N_13743,N_13739);
xnor U13887 (N_13887,N_13671,N_13760);
nor U13888 (N_13888,N_13681,N_13726);
nand U13889 (N_13889,N_13543,N_13669);
nor U13890 (N_13890,N_13565,N_13503);
or U13891 (N_13891,N_13656,N_13686);
nor U13892 (N_13892,N_13764,N_13778);
nand U13893 (N_13893,N_13687,N_13795);
nor U13894 (N_13894,N_13617,N_13531);
nand U13895 (N_13895,N_13710,N_13728);
nor U13896 (N_13896,N_13672,N_13684);
nor U13897 (N_13897,N_13677,N_13547);
or U13898 (N_13898,N_13592,N_13792);
or U13899 (N_13899,N_13633,N_13601);
nor U13900 (N_13900,N_13515,N_13751);
xnor U13901 (N_13901,N_13709,N_13788);
or U13902 (N_13902,N_13614,N_13680);
xnor U13903 (N_13903,N_13697,N_13720);
or U13904 (N_13904,N_13689,N_13787);
and U13905 (N_13905,N_13765,N_13512);
xnor U13906 (N_13906,N_13579,N_13744);
xor U13907 (N_13907,N_13570,N_13701);
nand U13908 (N_13908,N_13589,N_13523);
xor U13909 (N_13909,N_13786,N_13622);
nor U13910 (N_13910,N_13569,N_13591);
nand U13911 (N_13911,N_13618,N_13621);
xor U13912 (N_13912,N_13627,N_13636);
xnor U13913 (N_13913,N_13675,N_13578);
and U13914 (N_13914,N_13729,N_13657);
or U13915 (N_13915,N_13581,N_13620);
and U13916 (N_13916,N_13797,N_13553);
xnor U13917 (N_13917,N_13526,N_13630);
or U13918 (N_13918,N_13741,N_13706);
xnor U13919 (N_13919,N_13794,N_13505);
nand U13920 (N_13920,N_13666,N_13678);
and U13921 (N_13921,N_13738,N_13770);
nand U13922 (N_13922,N_13663,N_13674);
xnor U13923 (N_13923,N_13691,N_13752);
or U13924 (N_13924,N_13769,N_13632);
nand U13925 (N_13925,N_13626,N_13705);
nand U13926 (N_13926,N_13714,N_13598);
and U13927 (N_13927,N_13725,N_13528);
nor U13928 (N_13928,N_13773,N_13571);
nor U13929 (N_13929,N_13628,N_13763);
or U13930 (N_13930,N_13665,N_13550);
nor U13931 (N_13931,N_13699,N_13703);
and U13932 (N_13932,N_13723,N_13700);
and U13933 (N_13933,N_13753,N_13560);
and U13934 (N_13934,N_13772,N_13588);
or U13935 (N_13935,N_13532,N_13637);
nand U13936 (N_13936,N_13506,N_13539);
or U13937 (N_13937,N_13692,N_13533);
nor U13938 (N_13938,N_13602,N_13603);
nor U13939 (N_13939,N_13780,N_13690);
nand U13940 (N_13940,N_13708,N_13529);
xnor U13941 (N_13941,N_13727,N_13799);
or U13942 (N_13942,N_13683,N_13624);
xnor U13943 (N_13943,N_13667,N_13542);
or U13944 (N_13944,N_13642,N_13796);
or U13945 (N_13945,N_13664,N_13535);
nor U13946 (N_13946,N_13561,N_13696);
nor U13947 (N_13947,N_13676,N_13500);
nor U13948 (N_13948,N_13639,N_13623);
nand U13949 (N_13949,N_13652,N_13608);
xnor U13950 (N_13950,N_13517,N_13568);
nand U13951 (N_13951,N_13550,N_13716);
xnor U13952 (N_13952,N_13547,N_13734);
nand U13953 (N_13953,N_13684,N_13565);
and U13954 (N_13954,N_13670,N_13540);
nor U13955 (N_13955,N_13525,N_13677);
xnor U13956 (N_13956,N_13779,N_13687);
or U13957 (N_13957,N_13601,N_13759);
or U13958 (N_13958,N_13749,N_13561);
nand U13959 (N_13959,N_13624,N_13673);
and U13960 (N_13960,N_13521,N_13697);
or U13961 (N_13961,N_13561,N_13756);
xnor U13962 (N_13962,N_13765,N_13749);
and U13963 (N_13963,N_13566,N_13759);
xnor U13964 (N_13964,N_13650,N_13646);
or U13965 (N_13965,N_13533,N_13629);
nor U13966 (N_13966,N_13620,N_13735);
or U13967 (N_13967,N_13595,N_13638);
and U13968 (N_13968,N_13515,N_13661);
nor U13969 (N_13969,N_13775,N_13718);
and U13970 (N_13970,N_13758,N_13608);
and U13971 (N_13971,N_13633,N_13677);
or U13972 (N_13972,N_13514,N_13533);
and U13973 (N_13973,N_13601,N_13714);
and U13974 (N_13974,N_13702,N_13626);
and U13975 (N_13975,N_13641,N_13510);
nor U13976 (N_13976,N_13527,N_13704);
xor U13977 (N_13977,N_13738,N_13660);
nand U13978 (N_13978,N_13604,N_13675);
and U13979 (N_13979,N_13624,N_13724);
nand U13980 (N_13980,N_13757,N_13668);
or U13981 (N_13981,N_13535,N_13613);
and U13982 (N_13982,N_13516,N_13501);
nor U13983 (N_13983,N_13678,N_13786);
nor U13984 (N_13984,N_13663,N_13625);
nor U13985 (N_13985,N_13701,N_13604);
or U13986 (N_13986,N_13506,N_13673);
nand U13987 (N_13987,N_13706,N_13595);
and U13988 (N_13988,N_13541,N_13743);
and U13989 (N_13989,N_13641,N_13770);
xor U13990 (N_13990,N_13577,N_13750);
and U13991 (N_13991,N_13763,N_13743);
and U13992 (N_13992,N_13794,N_13552);
nor U13993 (N_13993,N_13700,N_13611);
nor U13994 (N_13994,N_13758,N_13593);
and U13995 (N_13995,N_13629,N_13513);
xnor U13996 (N_13996,N_13663,N_13594);
xor U13997 (N_13997,N_13735,N_13544);
or U13998 (N_13998,N_13535,N_13758);
and U13999 (N_13999,N_13698,N_13521);
nor U14000 (N_14000,N_13542,N_13584);
and U14001 (N_14001,N_13760,N_13574);
and U14002 (N_14002,N_13752,N_13608);
and U14003 (N_14003,N_13687,N_13571);
and U14004 (N_14004,N_13530,N_13787);
nor U14005 (N_14005,N_13626,N_13707);
nand U14006 (N_14006,N_13719,N_13773);
xor U14007 (N_14007,N_13554,N_13686);
nand U14008 (N_14008,N_13599,N_13660);
or U14009 (N_14009,N_13536,N_13701);
nand U14010 (N_14010,N_13751,N_13771);
and U14011 (N_14011,N_13744,N_13542);
or U14012 (N_14012,N_13698,N_13792);
xor U14013 (N_14013,N_13735,N_13673);
or U14014 (N_14014,N_13629,N_13546);
nand U14015 (N_14015,N_13657,N_13748);
xnor U14016 (N_14016,N_13531,N_13713);
or U14017 (N_14017,N_13592,N_13620);
and U14018 (N_14018,N_13584,N_13713);
and U14019 (N_14019,N_13658,N_13541);
nor U14020 (N_14020,N_13790,N_13603);
xnor U14021 (N_14021,N_13700,N_13629);
xnor U14022 (N_14022,N_13548,N_13728);
nor U14023 (N_14023,N_13771,N_13519);
or U14024 (N_14024,N_13639,N_13702);
nand U14025 (N_14025,N_13596,N_13795);
nor U14026 (N_14026,N_13518,N_13575);
or U14027 (N_14027,N_13745,N_13583);
and U14028 (N_14028,N_13723,N_13779);
nand U14029 (N_14029,N_13682,N_13507);
nand U14030 (N_14030,N_13799,N_13656);
or U14031 (N_14031,N_13744,N_13692);
nand U14032 (N_14032,N_13663,N_13763);
xnor U14033 (N_14033,N_13746,N_13729);
nor U14034 (N_14034,N_13709,N_13725);
xnor U14035 (N_14035,N_13505,N_13506);
and U14036 (N_14036,N_13757,N_13649);
xor U14037 (N_14037,N_13774,N_13671);
nor U14038 (N_14038,N_13719,N_13677);
nor U14039 (N_14039,N_13610,N_13561);
nor U14040 (N_14040,N_13601,N_13610);
xnor U14041 (N_14041,N_13762,N_13794);
or U14042 (N_14042,N_13616,N_13566);
and U14043 (N_14043,N_13549,N_13562);
or U14044 (N_14044,N_13665,N_13722);
and U14045 (N_14045,N_13647,N_13611);
xor U14046 (N_14046,N_13786,N_13620);
and U14047 (N_14047,N_13640,N_13603);
or U14048 (N_14048,N_13579,N_13588);
nand U14049 (N_14049,N_13617,N_13702);
or U14050 (N_14050,N_13740,N_13661);
and U14051 (N_14051,N_13537,N_13767);
nor U14052 (N_14052,N_13651,N_13642);
or U14053 (N_14053,N_13617,N_13594);
xnor U14054 (N_14054,N_13758,N_13767);
and U14055 (N_14055,N_13749,N_13763);
nor U14056 (N_14056,N_13599,N_13565);
nand U14057 (N_14057,N_13589,N_13657);
xor U14058 (N_14058,N_13580,N_13678);
nor U14059 (N_14059,N_13686,N_13714);
xor U14060 (N_14060,N_13744,N_13507);
or U14061 (N_14061,N_13731,N_13697);
and U14062 (N_14062,N_13731,N_13621);
or U14063 (N_14063,N_13507,N_13741);
and U14064 (N_14064,N_13573,N_13705);
nand U14065 (N_14065,N_13761,N_13625);
nand U14066 (N_14066,N_13701,N_13627);
nor U14067 (N_14067,N_13545,N_13617);
xor U14068 (N_14068,N_13515,N_13758);
xor U14069 (N_14069,N_13606,N_13696);
xor U14070 (N_14070,N_13739,N_13648);
nor U14071 (N_14071,N_13528,N_13693);
xnor U14072 (N_14072,N_13797,N_13727);
or U14073 (N_14073,N_13593,N_13640);
nor U14074 (N_14074,N_13574,N_13636);
xnor U14075 (N_14075,N_13638,N_13566);
and U14076 (N_14076,N_13762,N_13639);
xnor U14077 (N_14077,N_13738,N_13669);
and U14078 (N_14078,N_13781,N_13527);
and U14079 (N_14079,N_13647,N_13579);
and U14080 (N_14080,N_13793,N_13761);
xor U14081 (N_14081,N_13706,N_13773);
or U14082 (N_14082,N_13772,N_13637);
nand U14083 (N_14083,N_13728,N_13730);
or U14084 (N_14084,N_13710,N_13751);
xnor U14085 (N_14085,N_13776,N_13629);
xor U14086 (N_14086,N_13597,N_13668);
or U14087 (N_14087,N_13711,N_13668);
nand U14088 (N_14088,N_13788,N_13530);
and U14089 (N_14089,N_13541,N_13575);
or U14090 (N_14090,N_13659,N_13742);
and U14091 (N_14091,N_13567,N_13724);
or U14092 (N_14092,N_13620,N_13777);
or U14093 (N_14093,N_13707,N_13619);
nor U14094 (N_14094,N_13557,N_13751);
nand U14095 (N_14095,N_13730,N_13707);
xor U14096 (N_14096,N_13660,N_13764);
nand U14097 (N_14097,N_13749,N_13584);
and U14098 (N_14098,N_13661,N_13643);
and U14099 (N_14099,N_13648,N_13539);
xor U14100 (N_14100,N_13829,N_13899);
nor U14101 (N_14101,N_13981,N_14022);
nand U14102 (N_14102,N_13892,N_13898);
nor U14103 (N_14103,N_13983,N_14069);
and U14104 (N_14104,N_14016,N_13968);
and U14105 (N_14105,N_14094,N_13942);
or U14106 (N_14106,N_14006,N_14003);
nand U14107 (N_14107,N_13906,N_14049);
or U14108 (N_14108,N_14051,N_14055);
xor U14109 (N_14109,N_13919,N_13973);
nand U14110 (N_14110,N_13812,N_13807);
nand U14111 (N_14111,N_13834,N_14089);
and U14112 (N_14112,N_13816,N_13963);
nand U14113 (N_14113,N_13847,N_13970);
nand U14114 (N_14114,N_13914,N_14031);
or U14115 (N_14115,N_13949,N_13991);
nor U14116 (N_14116,N_14024,N_13947);
nand U14117 (N_14117,N_14054,N_13854);
or U14118 (N_14118,N_13868,N_13818);
or U14119 (N_14119,N_14078,N_13999);
nor U14120 (N_14120,N_13875,N_14068);
and U14121 (N_14121,N_14010,N_13945);
and U14122 (N_14122,N_13996,N_13946);
nor U14123 (N_14123,N_13993,N_13822);
xnor U14124 (N_14124,N_13851,N_13846);
nor U14125 (N_14125,N_13910,N_14039);
or U14126 (N_14126,N_13828,N_14047);
nand U14127 (N_14127,N_14075,N_14057);
and U14128 (N_14128,N_14040,N_13915);
nor U14129 (N_14129,N_13870,N_13921);
and U14130 (N_14130,N_13986,N_14044);
nor U14131 (N_14131,N_14045,N_14065);
nor U14132 (N_14132,N_13920,N_13841);
and U14133 (N_14133,N_13853,N_13957);
nor U14134 (N_14134,N_14020,N_13948);
or U14135 (N_14135,N_13858,N_14005);
nand U14136 (N_14136,N_14082,N_13863);
and U14137 (N_14137,N_14001,N_13872);
and U14138 (N_14138,N_14028,N_13844);
or U14139 (N_14139,N_14025,N_13940);
nand U14140 (N_14140,N_14015,N_13825);
nand U14141 (N_14141,N_13902,N_13843);
nand U14142 (N_14142,N_14096,N_13802);
nor U14143 (N_14143,N_13953,N_13839);
and U14144 (N_14144,N_13939,N_13956);
nand U14145 (N_14145,N_13985,N_13903);
and U14146 (N_14146,N_14070,N_13893);
nor U14147 (N_14147,N_14009,N_14095);
and U14148 (N_14148,N_13900,N_14077);
and U14149 (N_14149,N_13979,N_13980);
xor U14150 (N_14150,N_13880,N_14093);
nand U14151 (N_14151,N_14038,N_13992);
or U14152 (N_14152,N_14026,N_14059);
and U14153 (N_14153,N_13808,N_13855);
and U14154 (N_14154,N_13813,N_14076);
and U14155 (N_14155,N_13929,N_13852);
and U14156 (N_14156,N_14036,N_13937);
nor U14157 (N_14157,N_13938,N_14084);
nor U14158 (N_14158,N_13804,N_13826);
nor U14159 (N_14159,N_14032,N_14046);
xnor U14160 (N_14160,N_14098,N_14058);
xnor U14161 (N_14161,N_13801,N_13998);
and U14162 (N_14162,N_14037,N_13982);
nor U14163 (N_14163,N_13856,N_13909);
or U14164 (N_14164,N_13995,N_13864);
nand U14165 (N_14165,N_13809,N_14023);
or U14166 (N_14166,N_13972,N_13806);
or U14167 (N_14167,N_13971,N_13926);
nor U14168 (N_14168,N_13944,N_13974);
or U14169 (N_14169,N_13859,N_13827);
and U14170 (N_14170,N_14099,N_13886);
nand U14171 (N_14171,N_14083,N_13924);
xor U14172 (N_14172,N_13833,N_13918);
or U14173 (N_14173,N_14066,N_13836);
nor U14174 (N_14174,N_13842,N_13913);
nor U14175 (N_14175,N_14086,N_13876);
and U14176 (N_14176,N_14063,N_14017);
xnor U14177 (N_14177,N_13862,N_13881);
and U14178 (N_14178,N_14061,N_13907);
nand U14179 (N_14179,N_13933,N_14090);
xor U14180 (N_14180,N_13901,N_13960);
nand U14181 (N_14181,N_14073,N_14011);
nand U14182 (N_14182,N_13962,N_13819);
xor U14183 (N_14183,N_14050,N_13873);
nor U14184 (N_14184,N_13984,N_13821);
xnor U14185 (N_14185,N_13925,N_13800);
or U14186 (N_14186,N_13930,N_14072);
nor U14187 (N_14187,N_13958,N_13976);
nor U14188 (N_14188,N_14019,N_14034);
nand U14189 (N_14189,N_13917,N_13871);
xnor U14190 (N_14190,N_13865,N_13928);
xnor U14191 (N_14191,N_14064,N_14053);
nand U14192 (N_14192,N_14043,N_13883);
xor U14193 (N_14193,N_13987,N_13954);
nand U14194 (N_14194,N_13815,N_13850);
nor U14195 (N_14195,N_14021,N_13869);
xor U14196 (N_14196,N_13994,N_13931);
and U14197 (N_14197,N_13959,N_13837);
nor U14198 (N_14198,N_13814,N_13882);
nor U14199 (N_14199,N_14079,N_13967);
nand U14200 (N_14200,N_14048,N_13922);
or U14201 (N_14201,N_13817,N_14097);
and U14202 (N_14202,N_13890,N_14004);
or U14203 (N_14203,N_13989,N_14085);
nand U14204 (N_14204,N_13912,N_13884);
xnor U14205 (N_14205,N_13990,N_14014);
or U14206 (N_14206,N_13988,N_13810);
nand U14207 (N_14207,N_14018,N_13952);
nor U14208 (N_14208,N_13877,N_14041);
nand U14209 (N_14209,N_13831,N_14062);
nor U14210 (N_14210,N_14007,N_13923);
nor U14211 (N_14211,N_13845,N_13905);
xnor U14212 (N_14212,N_13965,N_13889);
nor U14213 (N_14213,N_13832,N_13977);
xor U14214 (N_14214,N_13803,N_13895);
xnor U14215 (N_14215,N_13874,N_13997);
xnor U14216 (N_14216,N_14088,N_14071);
xor U14217 (N_14217,N_14091,N_13835);
nand U14218 (N_14218,N_13861,N_14081);
or U14219 (N_14219,N_13934,N_13955);
xnor U14220 (N_14220,N_13830,N_13823);
nor U14221 (N_14221,N_14029,N_14087);
nand U14222 (N_14222,N_13911,N_13978);
nor U14223 (N_14223,N_14027,N_13961);
nand U14224 (N_14224,N_13811,N_13943);
or U14225 (N_14225,N_13927,N_13840);
or U14226 (N_14226,N_13896,N_13820);
and U14227 (N_14227,N_13824,N_13969);
xnor U14228 (N_14228,N_13950,N_13888);
nor U14229 (N_14229,N_13916,N_14092);
and U14230 (N_14230,N_13857,N_13867);
and U14231 (N_14231,N_14042,N_13932);
and U14232 (N_14232,N_13805,N_13966);
or U14233 (N_14233,N_13866,N_14052);
nand U14234 (N_14234,N_14035,N_14033);
nand U14235 (N_14235,N_13885,N_14030);
and U14236 (N_14236,N_13860,N_13879);
and U14237 (N_14237,N_14056,N_13941);
or U14238 (N_14238,N_13935,N_13951);
nor U14239 (N_14239,N_13936,N_14067);
nand U14240 (N_14240,N_13849,N_13848);
nand U14241 (N_14241,N_13908,N_13964);
nand U14242 (N_14242,N_13891,N_14080);
and U14243 (N_14243,N_14074,N_14008);
xor U14244 (N_14244,N_13878,N_14060);
nor U14245 (N_14245,N_14000,N_13894);
xor U14246 (N_14246,N_13838,N_13904);
nor U14247 (N_14247,N_14013,N_14002);
xor U14248 (N_14248,N_13897,N_14012);
xor U14249 (N_14249,N_13887,N_13975);
and U14250 (N_14250,N_14015,N_13800);
xor U14251 (N_14251,N_13869,N_13879);
nor U14252 (N_14252,N_13968,N_13937);
or U14253 (N_14253,N_13843,N_13946);
xnor U14254 (N_14254,N_14071,N_13924);
xor U14255 (N_14255,N_13825,N_13840);
nand U14256 (N_14256,N_13906,N_13974);
nor U14257 (N_14257,N_13863,N_13887);
nor U14258 (N_14258,N_13923,N_13992);
or U14259 (N_14259,N_14089,N_13993);
and U14260 (N_14260,N_13937,N_13919);
nor U14261 (N_14261,N_13970,N_13913);
nand U14262 (N_14262,N_13907,N_14070);
nor U14263 (N_14263,N_13952,N_13935);
nor U14264 (N_14264,N_13934,N_13939);
xor U14265 (N_14265,N_14026,N_14024);
nor U14266 (N_14266,N_13989,N_14069);
or U14267 (N_14267,N_13810,N_13848);
xor U14268 (N_14268,N_14099,N_13840);
nand U14269 (N_14269,N_14041,N_14034);
nand U14270 (N_14270,N_13883,N_13812);
xnor U14271 (N_14271,N_13825,N_13932);
nor U14272 (N_14272,N_14038,N_13868);
and U14273 (N_14273,N_14030,N_13865);
xnor U14274 (N_14274,N_13908,N_13832);
or U14275 (N_14275,N_13917,N_13913);
and U14276 (N_14276,N_13829,N_14020);
nand U14277 (N_14277,N_13987,N_13900);
and U14278 (N_14278,N_14063,N_14068);
and U14279 (N_14279,N_13853,N_14025);
and U14280 (N_14280,N_14026,N_14093);
nor U14281 (N_14281,N_14098,N_13866);
xnor U14282 (N_14282,N_13962,N_13918);
and U14283 (N_14283,N_13811,N_13822);
nor U14284 (N_14284,N_13807,N_13941);
xor U14285 (N_14285,N_13928,N_13812);
nand U14286 (N_14286,N_14018,N_13852);
and U14287 (N_14287,N_14021,N_14067);
nor U14288 (N_14288,N_13921,N_13987);
or U14289 (N_14289,N_13994,N_13899);
or U14290 (N_14290,N_14009,N_13887);
xnor U14291 (N_14291,N_13891,N_14072);
xor U14292 (N_14292,N_14000,N_14087);
nor U14293 (N_14293,N_13848,N_13865);
nor U14294 (N_14294,N_13975,N_13971);
nor U14295 (N_14295,N_13839,N_13957);
nor U14296 (N_14296,N_13995,N_13918);
xnor U14297 (N_14297,N_14042,N_14076);
xor U14298 (N_14298,N_13975,N_14062);
xor U14299 (N_14299,N_13803,N_13987);
nand U14300 (N_14300,N_13887,N_14075);
nor U14301 (N_14301,N_13858,N_13895);
or U14302 (N_14302,N_14024,N_13878);
xor U14303 (N_14303,N_13813,N_14089);
nor U14304 (N_14304,N_13843,N_14045);
xnor U14305 (N_14305,N_13995,N_14050);
nor U14306 (N_14306,N_13859,N_13868);
xor U14307 (N_14307,N_14039,N_14049);
xor U14308 (N_14308,N_13921,N_13810);
nor U14309 (N_14309,N_14009,N_13892);
or U14310 (N_14310,N_13806,N_13890);
and U14311 (N_14311,N_13840,N_13983);
nor U14312 (N_14312,N_14087,N_13824);
and U14313 (N_14313,N_14022,N_13819);
xnor U14314 (N_14314,N_13838,N_14004);
nand U14315 (N_14315,N_13820,N_13934);
or U14316 (N_14316,N_13982,N_13842);
nand U14317 (N_14317,N_14039,N_14051);
nand U14318 (N_14318,N_13992,N_14020);
or U14319 (N_14319,N_13991,N_14018);
and U14320 (N_14320,N_14024,N_13898);
or U14321 (N_14321,N_13906,N_13893);
or U14322 (N_14322,N_14040,N_13991);
nor U14323 (N_14323,N_14062,N_14039);
or U14324 (N_14324,N_13915,N_14046);
and U14325 (N_14325,N_13955,N_13800);
and U14326 (N_14326,N_14098,N_13855);
nor U14327 (N_14327,N_14023,N_14086);
nor U14328 (N_14328,N_14097,N_13967);
nor U14329 (N_14329,N_14029,N_14064);
nand U14330 (N_14330,N_13905,N_14017);
and U14331 (N_14331,N_13965,N_13860);
xor U14332 (N_14332,N_14046,N_14097);
nor U14333 (N_14333,N_14047,N_13841);
xor U14334 (N_14334,N_13869,N_13841);
and U14335 (N_14335,N_13838,N_13863);
nand U14336 (N_14336,N_14034,N_13905);
nor U14337 (N_14337,N_13888,N_13921);
and U14338 (N_14338,N_14053,N_13992);
or U14339 (N_14339,N_14073,N_14038);
and U14340 (N_14340,N_13891,N_13905);
nor U14341 (N_14341,N_13910,N_13880);
nand U14342 (N_14342,N_14077,N_14091);
or U14343 (N_14343,N_14065,N_13817);
or U14344 (N_14344,N_13847,N_13967);
nand U14345 (N_14345,N_13818,N_13824);
nor U14346 (N_14346,N_14041,N_13839);
and U14347 (N_14347,N_14010,N_13898);
or U14348 (N_14348,N_13852,N_14026);
nor U14349 (N_14349,N_13865,N_14007);
xor U14350 (N_14350,N_14000,N_13978);
or U14351 (N_14351,N_14053,N_13809);
or U14352 (N_14352,N_13937,N_14015);
and U14353 (N_14353,N_14068,N_13894);
xnor U14354 (N_14354,N_14070,N_13832);
or U14355 (N_14355,N_13864,N_13863);
and U14356 (N_14356,N_14035,N_13846);
or U14357 (N_14357,N_13904,N_13808);
xor U14358 (N_14358,N_14080,N_13897);
xnor U14359 (N_14359,N_13849,N_14016);
nor U14360 (N_14360,N_14066,N_13859);
or U14361 (N_14361,N_14051,N_13906);
xnor U14362 (N_14362,N_13906,N_14095);
xnor U14363 (N_14363,N_13845,N_13858);
and U14364 (N_14364,N_13941,N_13999);
nand U14365 (N_14365,N_14095,N_13815);
or U14366 (N_14366,N_13825,N_13991);
nand U14367 (N_14367,N_13938,N_13959);
or U14368 (N_14368,N_13963,N_13840);
xor U14369 (N_14369,N_14047,N_13922);
and U14370 (N_14370,N_14082,N_13800);
or U14371 (N_14371,N_14019,N_13954);
and U14372 (N_14372,N_14044,N_13810);
xnor U14373 (N_14373,N_13926,N_13859);
and U14374 (N_14374,N_13867,N_13858);
nand U14375 (N_14375,N_14028,N_13813);
nor U14376 (N_14376,N_14033,N_14059);
nor U14377 (N_14377,N_13829,N_13930);
nor U14378 (N_14378,N_14095,N_13827);
xnor U14379 (N_14379,N_14027,N_13921);
xnor U14380 (N_14380,N_13993,N_14057);
nor U14381 (N_14381,N_14050,N_14066);
nor U14382 (N_14382,N_13823,N_13974);
or U14383 (N_14383,N_13828,N_13814);
nor U14384 (N_14384,N_13862,N_13982);
nand U14385 (N_14385,N_13976,N_13968);
or U14386 (N_14386,N_13924,N_13953);
nor U14387 (N_14387,N_13802,N_13947);
nand U14388 (N_14388,N_13871,N_13920);
xnor U14389 (N_14389,N_14098,N_13944);
nand U14390 (N_14390,N_13879,N_14043);
xnor U14391 (N_14391,N_13808,N_13974);
nor U14392 (N_14392,N_13824,N_14011);
nand U14393 (N_14393,N_13895,N_13919);
xnor U14394 (N_14394,N_13984,N_13995);
or U14395 (N_14395,N_13885,N_14074);
xnor U14396 (N_14396,N_13924,N_14035);
nor U14397 (N_14397,N_13865,N_14080);
nand U14398 (N_14398,N_13863,N_13951);
nor U14399 (N_14399,N_13887,N_14010);
xor U14400 (N_14400,N_14263,N_14342);
or U14401 (N_14401,N_14312,N_14199);
nor U14402 (N_14402,N_14144,N_14382);
and U14403 (N_14403,N_14393,N_14316);
xor U14404 (N_14404,N_14142,N_14127);
or U14405 (N_14405,N_14201,N_14138);
or U14406 (N_14406,N_14205,N_14307);
nand U14407 (N_14407,N_14198,N_14213);
nor U14408 (N_14408,N_14306,N_14166);
nand U14409 (N_14409,N_14167,N_14285);
xnor U14410 (N_14410,N_14126,N_14243);
nand U14411 (N_14411,N_14208,N_14270);
or U14412 (N_14412,N_14294,N_14105);
or U14413 (N_14413,N_14154,N_14183);
and U14414 (N_14414,N_14257,N_14239);
and U14415 (N_14415,N_14268,N_14356);
nor U14416 (N_14416,N_14140,N_14241);
nor U14417 (N_14417,N_14273,N_14321);
xnor U14418 (N_14418,N_14373,N_14326);
xor U14419 (N_14419,N_14182,N_14170);
nor U14420 (N_14420,N_14113,N_14139);
nand U14421 (N_14421,N_14180,N_14130);
xor U14422 (N_14422,N_14339,N_14129);
xor U14423 (N_14423,N_14278,N_14293);
xnor U14424 (N_14424,N_14381,N_14394);
nand U14425 (N_14425,N_14203,N_14301);
and U14426 (N_14426,N_14189,N_14334);
and U14427 (N_14427,N_14264,N_14360);
or U14428 (N_14428,N_14128,N_14319);
or U14429 (N_14429,N_14341,N_14192);
and U14430 (N_14430,N_14379,N_14132);
nor U14431 (N_14431,N_14358,N_14350);
nand U14432 (N_14432,N_14186,N_14240);
and U14433 (N_14433,N_14322,N_14300);
or U14434 (N_14434,N_14115,N_14367);
nor U14435 (N_14435,N_14390,N_14204);
and U14436 (N_14436,N_14124,N_14317);
nand U14437 (N_14437,N_14308,N_14274);
and U14438 (N_14438,N_14384,N_14175);
xnor U14439 (N_14439,N_14254,N_14385);
or U14440 (N_14440,N_14149,N_14296);
and U14441 (N_14441,N_14258,N_14229);
or U14442 (N_14442,N_14399,N_14188);
and U14443 (N_14443,N_14344,N_14354);
or U14444 (N_14444,N_14256,N_14153);
nor U14445 (N_14445,N_14295,N_14315);
and U14446 (N_14446,N_14232,N_14152);
nand U14447 (N_14447,N_14174,N_14260);
xnor U14448 (N_14448,N_14106,N_14185);
xnor U14449 (N_14449,N_14378,N_14158);
and U14450 (N_14450,N_14346,N_14365);
nor U14451 (N_14451,N_14348,N_14216);
xnor U14452 (N_14452,N_14242,N_14218);
nor U14453 (N_14453,N_14195,N_14271);
nand U14454 (N_14454,N_14112,N_14235);
and U14455 (N_14455,N_14212,N_14250);
xnor U14456 (N_14456,N_14340,N_14297);
or U14457 (N_14457,N_14333,N_14147);
nor U14458 (N_14458,N_14221,N_14200);
nand U14459 (N_14459,N_14347,N_14374);
nor U14460 (N_14460,N_14364,N_14332);
xnor U14461 (N_14461,N_14287,N_14209);
or U14462 (N_14462,N_14249,N_14190);
nand U14463 (N_14463,N_14236,N_14161);
xor U14464 (N_14464,N_14159,N_14122);
nor U14465 (N_14465,N_14336,N_14318);
xnor U14466 (N_14466,N_14119,N_14118);
nor U14467 (N_14467,N_14359,N_14101);
or U14468 (N_14468,N_14357,N_14369);
and U14469 (N_14469,N_14234,N_14143);
nor U14470 (N_14470,N_14237,N_14179);
nand U14471 (N_14471,N_14109,N_14255);
nor U14472 (N_14472,N_14377,N_14193);
or U14473 (N_14473,N_14137,N_14135);
xor U14474 (N_14474,N_14397,N_14310);
nand U14475 (N_14475,N_14362,N_14288);
nor U14476 (N_14476,N_14168,N_14338);
nand U14477 (N_14477,N_14325,N_14206);
and U14478 (N_14478,N_14392,N_14372);
nand U14479 (N_14479,N_14395,N_14353);
xor U14480 (N_14480,N_14245,N_14145);
xnor U14481 (N_14481,N_14352,N_14313);
nand U14482 (N_14482,N_14156,N_14177);
and U14483 (N_14483,N_14355,N_14160);
nand U14484 (N_14484,N_14184,N_14290);
nor U14485 (N_14485,N_14314,N_14202);
nand U14486 (N_14486,N_14171,N_14335);
or U14487 (N_14487,N_14169,N_14226);
or U14488 (N_14488,N_14280,N_14197);
nand U14489 (N_14489,N_14329,N_14247);
and U14490 (N_14490,N_14351,N_14162);
nand U14491 (N_14491,N_14214,N_14269);
nand U14492 (N_14492,N_14225,N_14230);
or U14493 (N_14493,N_14211,N_14272);
and U14494 (N_14494,N_14330,N_14151);
or U14495 (N_14495,N_14121,N_14187);
and U14496 (N_14496,N_14117,N_14387);
nand U14497 (N_14497,N_14146,N_14102);
nor U14498 (N_14498,N_14246,N_14328);
or U14499 (N_14499,N_14238,N_14303);
nand U14500 (N_14500,N_14155,N_14210);
xnor U14501 (N_14501,N_14116,N_14194);
xor U14502 (N_14502,N_14133,N_14207);
and U14503 (N_14503,N_14244,N_14262);
and U14504 (N_14504,N_14252,N_14291);
or U14505 (N_14505,N_14259,N_14125);
nand U14506 (N_14506,N_14289,N_14227);
nor U14507 (N_14507,N_14370,N_14222);
xnor U14508 (N_14508,N_14228,N_14327);
or U14509 (N_14509,N_14324,N_14337);
xor U14510 (N_14510,N_14380,N_14100);
nor U14511 (N_14511,N_14275,N_14286);
nor U14512 (N_14512,N_14396,N_14172);
nand U14513 (N_14513,N_14323,N_14388);
or U14514 (N_14514,N_14104,N_14345);
or U14515 (N_14515,N_14368,N_14181);
nand U14516 (N_14516,N_14361,N_14331);
or U14517 (N_14517,N_14111,N_14215);
nor U14518 (N_14518,N_14157,N_14248);
nand U14519 (N_14519,N_14389,N_14108);
nand U14520 (N_14520,N_14178,N_14253);
nand U14521 (N_14521,N_14299,N_14309);
nand U14522 (N_14522,N_14120,N_14220);
and U14523 (N_14523,N_14283,N_14191);
or U14524 (N_14524,N_14302,N_14265);
or U14525 (N_14525,N_14376,N_14103);
or U14526 (N_14526,N_14224,N_14261);
nor U14527 (N_14527,N_14298,N_14131);
nor U14528 (N_14528,N_14284,N_14217);
nand U14529 (N_14529,N_14349,N_14231);
xor U14530 (N_14530,N_14148,N_14383);
nand U14531 (N_14531,N_14398,N_14107);
or U14532 (N_14532,N_14266,N_14123);
nand U14533 (N_14533,N_14173,N_14136);
and U14534 (N_14534,N_14304,N_14251);
nand U14535 (N_14535,N_14196,N_14292);
and U14536 (N_14536,N_14219,N_14163);
nor U14537 (N_14537,N_14282,N_14165);
or U14538 (N_14538,N_14110,N_14343);
nand U14539 (N_14539,N_14267,N_14363);
or U14540 (N_14540,N_14164,N_14276);
xnor U14541 (N_14541,N_14366,N_14281);
nand U14542 (N_14542,N_14141,N_14375);
and U14543 (N_14543,N_14176,N_14311);
nand U14544 (N_14544,N_14233,N_14305);
xnor U14545 (N_14545,N_14150,N_14371);
or U14546 (N_14546,N_14277,N_14223);
or U14547 (N_14547,N_14386,N_14320);
xnor U14548 (N_14548,N_14114,N_14391);
and U14549 (N_14549,N_14279,N_14134);
nor U14550 (N_14550,N_14153,N_14358);
nand U14551 (N_14551,N_14297,N_14242);
nor U14552 (N_14552,N_14310,N_14323);
xor U14553 (N_14553,N_14334,N_14127);
nor U14554 (N_14554,N_14357,N_14146);
or U14555 (N_14555,N_14230,N_14292);
nand U14556 (N_14556,N_14308,N_14110);
nor U14557 (N_14557,N_14129,N_14222);
and U14558 (N_14558,N_14243,N_14180);
xnor U14559 (N_14559,N_14394,N_14319);
nor U14560 (N_14560,N_14397,N_14236);
xor U14561 (N_14561,N_14108,N_14146);
or U14562 (N_14562,N_14358,N_14367);
or U14563 (N_14563,N_14278,N_14101);
nor U14564 (N_14564,N_14337,N_14198);
nor U14565 (N_14565,N_14183,N_14297);
nand U14566 (N_14566,N_14230,N_14151);
or U14567 (N_14567,N_14355,N_14279);
nor U14568 (N_14568,N_14129,N_14234);
and U14569 (N_14569,N_14209,N_14294);
or U14570 (N_14570,N_14354,N_14291);
nand U14571 (N_14571,N_14273,N_14282);
or U14572 (N_14572,N_14218,N_14119);
and U14573 (N_14573,N_14291,N_14310);
or U14574 (N_14574,N_14304,N_14140);
or U14575 (N_14575,N_14116,N_14373);
and U14576 (N_14576,N_14337,N_14246);
nand U14577 (N_14577,N_14332,N_14109);
nand U14578 (N_14578,N_14128,N_14363);
nor U14579 (N_14579,N_14234,N_14140);
nor U14580 (N_14580,N_14207,N_14217);
and U14581 (N_14581,N_14351,N_14130);
or U14582 (N_14582,N_14263,N_14181);
or U14583 (N_14583,N_14270,N_14301);
and U14584 (N_14584,N_14171,N_14305);
xor U14585 (N_14585,N_14280,N_14148);
nand U14586 (N_14586,N_14219,N_14304);
xor U14587 (N_14587,N_14386,N_14142);
nand U14588 (N_14588,N_14189,N_14205);
or U14589 (N_14589,N_14250,N_14159);
xnor U14590 (N_14590,N_14215,N_14345);
xnor U14591 (N_14591,N_14328,N_14396);
and U14592 (N_14592,N_14316,N_14314);
or U14593 (N_14593,N_14300,N_14328);
nor U14594 (N_14594,N_14355,N_14275);
or U14595 (N_14595,N_14397,N_14122);
or U14596 (N_14596,N_14342,N_14362);
nand U14597 (N_14597,N_14386,N_14374);
xnor U14598 (N_14598,N_14272,N_14114);
or U14599 (N_14599,N_14164,N_14269);
nand U14600 (N_14600,N_14312,N_14284);
or U14601 (N_14601,N_14218,N_14343);
nand U14602 (N_14602,N_14275,N_14222);
or U14603 (N_14603,N_14191,N_14137);
or U14604 (N_14604,N_14121,N_14362);
or U14605 (N_14605,N_14239,N_14375);
xor U14606 (N_14606,N_14287,N_14276);
and U14607 (N_14607,N_14320,N_14399);
nand U14608 (N_14608,N_14204,N_14241);
and U14609 (N_14609,N_14148,N_14351);
or U14610 (N_14610,N_14323,N_14121);
nand U14611 (N_14611,N_14165,N_14194);
and U14612 (N_14612,N_14322,N_14204);
and U14613 (N_14613,N_14271,N_14264);
nand U14614 (N_14614,N_14210,N_14100);
nand U14615 (N_14615,N_14161,N_14184);
and U14616 (N_14616,N_14353,N_14192);
xnor U14617 (N_14617,N_14206,N_14237);
xor U14618 (N_14618,N_14108,N_14217);
nand U14619 (N_14619,N_14141,N_14102);
and U14620 (N_14620,N_14134,N_14147);
nand U14621 (N_14621,N_14268,N_14325);
or U14622 (N_14622,N_14265,N_14240);
and U14623 (N_14623,N_14305,N_14122);
nor U14624 (N_14624,N_14168,N_14318);
nor U14625 (N_14625,N_14167,N_14293);
nand U14626 (N_14626,N_14329,N_14236);
xnor U14627 (N_14627,N_14201,N_14159);
nand U14628 (N_14628,N_14111,N_14307);
nor U14629 (N_14629,N_14253,N_14147);
xnor U14630 (N_14630,N_14299,N_14274);
nor U14631 (N_14631,N_14161,N_14238);
and U14632 (N_14632,N_14270,N_14227);
nor U14633 (N_14633,N_14229,N_14245);
nand U14634 (N_14634,N_14275,N_14310);
and U14635 (N_14635,N_14139,N_14379);
and U14636 (N_14636,N_14365,N_14239);
xnor U14637 (N_14637,N_14207,N_14377);
or U14638 (N_14638,N_14172,N_14350);
or U14639 (N_14639,N_14290,N_14159);
or U14640 (N_14640,N_14242,N_14323);
and U14641 (N_14641,N_14223,N_14270);
and U14642 (N_14642,N_14153,N_14241);
xor U14643 (N_14643,N_14319,N_14396);
and U14644 (N_14644,N_14315,N_14210);
xor U14645 (N_14645,N_14188,N_14378);
and U14646 (N_14646,N_14281,N_14154);
nand U14647 (N_14647,N_14191,N_14206);
or U14648 (N_14648,N_14344,N_14298);
or U14649 (N_14649,N_14340,N_14204);
or U14650 (N_14650,N_14196,N_14125);
xnor U14651 (N_14651,N_14305,N_14389);
nor U14652 (N_14652,N_14231,N_14113);
and U14653 (N_14653,N_14233,N_14246);
or U14654 (N_14654,N_14199,N_14156);
and U14655 (N_14655,N_14215,N_14360);
or U14656 (N_14656,N_14279,N_14109);
and U14657 (N_14657,N_14147,N_14243);
and U14658 (N_14658,N_14221,N_14184);
or U14659 (N_14659,N_14232,N_14315);
and U14660 (N_14660,N_14357,N_14259);
nor U14661 (N_14661,N_14142,N_14162);
and U14662 (N_14662,N_14300,N_14246);
nor U14663 (N_14663,N_14362,N_14211);
nor U14664 (N_14664,N_14218,N_14371);
and U14665 (N_14665,N_14173,N_14155);
or U14666 (N_14666,N_14265,N_14368);
or U14667 (N_14667,N_14218,N_14126);
xor U14668 (N_14668,N_14100,N_14127);
xor U14669 (N_14669,N_14171,N_14249);
nand U14670 (N_14670,N_14202,N_14336);
and U14671 (N_14671,N_14330,N_14197);
or U14672 (N_14672,N_14118,N_14117);
and U14673 (N_14673,N_14222,N_14268);
xor U14674 (N_14674,N_14314,N_14182);
nor U14675 (N_14675,N_14279,N_14242);
nand U14676 (N_14676,N_14112,N_14344);
nor U14677 (N_14677,N_14350,N_14386);
or U14678 (N_14678,N_14243,N_14267);
nor U14679 (N_14679,N_14268,N_14382);
nand U14680 (N_14680,N_14125,N_14328);
or U14681 (N_14681,N_14108,N_14162);
xor U14682 (N_14682,N_14123,N_14235);
nand U14683 (N_14683,N_14250,N_14246);
xor U14684 (N_14684,N_14347,N_14143);
or U14685 (N_14685,N_14111,N_14293);
xnor U14686 (N_14686,N_14391,N_14121);
xor U14687 (N_14687,N_14322,N_14159);
or U14688 (N_14688,N_14387,N_14306);
and U14689 (N_14689,N_14317,N_14248);
nor U14690 (N_14690,N_14119,N_14196);
or U14691 (N_14691,N_14353,N_14232);
xnor U14692 (N_14692,N_14310,N_14294);
nor U14693 (N_14693,N_14346,N_14336);
or U14694 (N_14694,N_14192,N_14392);
nor U14695 (N_14695,N_14242,N_14102);
xor U14696 (N_14696,N_14178,N_14293);
and U14697 (N_14697,N_14204,N_14179);
xnor U14698 (N_14698,N_14159,N_14279);
nand U14699 (N_14699,N_14145,N_14307);
xnor U14700 (N_14700,N_14698,N_14403);
and U14701 (N_14701,N_14672,N_14490);
nor U14702 (N_14702,N_14625,N_14520);
and U14703 (N_14703,N_14539,N_14687);
and U14704 (N_14704,N_14410,N_14559);
xnor U14705 (N_14705,N_14467,N_14401);
xor U14706 (N_14706,N_14680,N_14523);
or U14707 (N_14707,N_14453,N_14430);
nor U14708 (N_14708,N_14650,N_14437);
nand U14709 (N_14709,N_14540,N_14555);
or U14710 (N_14710,N_14411,N_14530);
nor U14711 (N_14711,N_14588,N_14564);
xnor U14712 (N_14712,N_14451,N_14684);
or U14713 (N_14713,N_14491,N_14648);
and U14714 (N_14714,N_14528,N_14614);
or U14715 (N_14715,N_14507,N_14518);
or U14716 (N_14716,N_14612,N_14638);
or U14717 (N_14717,N_14547,N_14488);
and U14718 (N_14718,N_14603,N_14461);
nor U14719 (N_14719,N_14502,N_14423);
or U14720 (N_14720,N_14541,N_14569);
nor U14721 (N_14721,N_14594,N_14419);
nor U14722 (N_14722,N_14532,N_14450);
xnor U14723 (N_14723,N_14416,N_14605);
and U14724 (N_14724,N_14439,N_14481);
and U14725 (N_14725,N_14571,N_14484);
xor U14726 (N_14726,N_14560,N_14557);
or U14727 (N_14727,N_14601,N_14441);
xor U14728 (N_14728,N_14658,N_14435);
nand U14729 (N_14729,N_14427,N_14476);
and U14730 (N_14730,N_14630,N_14534);
nor U14731 (N_14731,N_14667,N_14677);
or U14732 (N_14732,N_14619,N_14431);
nand U14733 (N_14733,N_14600,N_14568);
or U14734 (N_14734,N_14485,N_14682);
nand U14735 (N_14735,N_14636,N_14606);
xnor U14736 (N_14736,N_14514,N_14543);
or U14737 (N_14737,N_14621,N_14611);
or U14738 (N_14738,N_14574,N_14400);
nand U14739 (N_14739,N_14660,N_14622);
nor U14740 (N_14740,N_14604,N_14512);
nand U14741 (N_14741,N_14581,N_14692);
xor U14742 (N_14742,N_14644,N_14402);
nand U14743 (N_14743,N_14546,N_14527);
or U14744 (N_14744,N_14506,N_14688);
xnor U14745 (N_14745,N_14616,N_14444);
and U14746 (N_14746,N_14428,N_14538);
and U14747 (N_14747,N_14550,N_14639);
xor U14748 (N_14748,N_14478,N_14694);
xnor U14749 (N_14749,N_14627,N_14406);
nand U14750 (N_14750,N_14666,N_14641);
nand U14751 (N_14751,N_14548,N_14623);
nor U14752 (N_14752,N_14609,N_14697);
xnor U14753 (N_14753,N_14699,N_14524);
or U14754 (N_14754,N_14468,N_14679);
nor U14755 (N_14755,N_14533,N_14575);
and U14756 (N_14756,N_14448,N_14469);
and U14757 (N_14757,N_14498,N_14492);
nor U14758 (N_14758,N_14563,N_14509);
nand U14759 (N_14759,N_14495,N_14521);
nor U14760 (N_14760,N_14649,N_14407);
xnor U14761 (N_14761,N_14493,N_14519);
nor U14762 (N_14762,N_14598,N_14417);
nor U14763 (N_14763,N_14654,N_14565);
nand U14764 (N_14764,N_14561,N_14477);
and U14765 (N_14765,N_14434,N_14631);
or U14766 (N_14766,N_14551,N_14695);
or U14767 (N_14767,N_14586,N_14497);
or U14768 (N_14768,N_14577,N_14470);
or U14769 (N_14769,N_14443,N_14635);
xnor U14770 (N_14770,N_14589,N_14657);
nand U14771 (N_14771,N_14661,N_14473);
or U14772 (N_14772,N_14691,N_14633);
or U14773 (N_14773,N_14554,N_14531);
nor U14774 (N_14774,N_14647,N_14580);
or U14775 (N_14775,N_14583,N_14620);
or U14776 (N_14776,N_14637,N_14504);
and U14777 (N_14777,N_14420,N_14617);
xnor U14778 (N_14778,N_14446,N_14452);
nand U14779 (N_14779,N_14670,N_14696);
and U14780 (N_14780,N_14607,N_14662);
nand U14781 (N_14781,N_14513,N_14664);
nor U14782 (N_14782,N_14408,N_14414);
nor U14783 (N_14783,N_14425,N_14421);
or U14784 (N_14784,N_14429,N_14653);
and U14785 (N_14785,N_14458,N_14579);
or U14786 (N_14786,N_14632,N_14545);
nand U14787 (N_14787,N_14505,N_14447);
nand U14788 (N_14788,N_14693,N_14608);
or U14789 (N_14789,N_14573,N_14659);
nor U14790 (N_14790,N_14438,N_14613);
nand U14791 (N_14791,N_14466,N_14681);
xor U14792 (N_14792,N_14676,N_14412);
xnor U14793 (N_14793,N_14440,N_14462);
and U14794 (N_14794,N_14494,N_14454);
or U14795 (N_14795,N_14642,N_14405);
nor U14796 (N_14796,N_14433,N_14460);
nor U14797 (N_14797,N_14516,N_14675);
nand U14798 (N_14798,N_14590,N_14629);
xnor U14799 (N_14799,N_14517,N_14669);
nor U14800 (N_14800,N_14671,N_14496);
or U14801 (N_14801,N_14562,N_14500);
or U14802 (N_14802,N_14415,N_14455);
nor U14803 (N_14803,N_14424,N_14449);
xor U14804 (N_14804,N_14529,N_14436);
or U14805 (N_14805,N_14503,N_14413);
nand U14806 (N_14806,N_14422,N_14549);
nand U14807 (N_14807,N_14651,N_14510);
nand U14808 (N_14808,N_14572,N_14542);
and U14809 (N_14809,N_14634,N_14442);
nand U14810 (N_14810,N_14686,N_14483);
nand U14811 (N_14811,N_14553,N_14656);
and U14812 (N_14812,N_14432,N_14566);
xnor U14813 (N_14813,N_14499,N_14570);
xnor U14814 (N_14814,N_14585,N_14487);
nand U14815 (N_14815,N_14618,N_14597);
or U14816 (N_14816,N_14567,N_14457);
xor U14817 (N_14817,N_14652,N_14584);
nand U14818 (N_14818,N_14456,N_14599);
xor U14819 (N_14819,N_14418,N_14515);
and U14820 (N_14820,N_14591,N_14445);
xnor U14821 (N_14821,N_14643,N_14610);
and U14822 (N_14822,N_14587,N_14426);
and U14823 (N_14823,N_14482,N_14474);
nor U14824 (N_14824,N_14471,N_14537);
xnor U14825 (N_14825,N_14595,N_14683);
and U14826 (N_14826,N_14536,N_14674);
nand U14827 (N_14827,N_14525,N_14596);
nor U14828 (N_14828,N_14646,N_14535);
nand U14829 (N_14829,N_14592,N_14463);
xnor U14830 (N_14830,N_14526,N_14628);
nor U14831 (N_14831,N_14615,N_14673);
nand U14832 (N_14832,N_14602,N_14552);
or U14833 (N_14833,N_14668,N_14578);
xor U14834 (N_14834,N_14645,N_14404);
or U14835 (N_14835,N_14489,N_14508);
nor U14836 (N_14836,N_14459,N_14640);
nor U14837 (N_14837,N_14558,N_14655);
and U14838 (N_14838,N_14665,N_14544);
or U14839 (N_14839,N_14479,N_14480);
or U14840 (N_14840,N_14472,N_14624);
nand U14841 (N_14841,N_14689,N_14593);
xor U14842 (N_14842,N_14576,N_14685);
nand U14843 (N_14843,N_14409,N_14690);
or U14844 (N_14844,N_14464,N_14582);
nand U14845 (N_14845,N_14663,N_14556);
and U14846 (N_14846,N_14626,N_14678);
nand U14847 (N_14847,N_14475,N_14465);
or U14848 (N_14848,N_14511,N_14522);
and U14849 (N_14849,N_14501,N_14486);
and U14850 (N_14850,N_14508,N_14613);
nor U14851 (N_14851,N_14613,N_14480);
and U14852 (N_14852,N_14648,N_14452);
nor U14853 (N_14853,N_14606,N_14614);
nor U14854 (N_14854,N_14663,N_14549);
nand U14855 (N_14855,N_14659,N_14625);
nand U14856 (N_14856,N_14431,N_14436);
or U14857 (N_14857,N_14400,N_14448);
or U14858 (N_14858,N_14581,N_14688);
nand U14859 (N_14859,N_14624,N_14674);
nand U14860 (N_14860,N_14513,N_14540);
nor U14861 (N_14861,N_14603,N_14417);
xnor U14862 (N_14862,N_14431,N_14449);
and U14863 (N_14863,N_14573,N_14417);
nand U14864 (N_14864,N_14544,N_14698);
or U14865 (N_14865,N_14538,N_14481);
nand U14866 (N_14866,N_14556,N_14460);
and U14867 (N_14867,N_14501,N_14617);
xor U14868 (N_14868,N_14432,N_14630);
and U14869 (N_14869,N_14653,N_14408);
xor U14870 (N_14870,N_14429,N_14451);
nand U14871 (N_14871,N_14689,N_14433);
and U14872 (N_14872,N_14554,N_14609);
and U14873 (N_14873,N_14617,N_14620);
and U14874 (N_14874,N_14404,N_14566);
nand U14875 (N_14875,N_14461,N_14632);
xnor U14876 (N_14876,N_14492,N_14553);
xor U14877 (N_14877,N_14489,N_14473);
nor U14878 (N_14878,N_14449,N_14480);
or U14879 (N_14879,N_14572,N_14677);
xor U14880 (N_14880,N_14504,N_14555);
nand U14881 (N_14881,N_14486,N_14511);
or U14882 (N_14882,N_14626,N_14618);
and U14883 (N_14883,N_14555,N_14424);
xor U14884 (N_14884,N_14491,N_14447);
or U14885 (N_14885,N_14401,N_14473);
and U14886 (N_14886,N_14686,N_14601);
or U14887 (N_14887,N_14628,N_14465);
or U14888 (N_14888,N_14661,N_14458);
nor U14889 (N_14889,N_14492,N_14679);
and U14890 (N_14890,N_14680,N_14480);
or U14891 (N_14891,N_14660,N_14567);
nand U14892 (N_14892,N_14614,N_14625);
or U14893 (N_14893,N_14512,N_14639);
and U14894 (N_14894,N_14697,N_14485);
xnor U14895 (N_14895,N_14523,N_14691);
nand U14896 (N_14896,N_14414,N_14405);
or U14897 (N_14897,N_14415,N_14593);
and U14898 (N_14898,N_14633,N_14631);
nor U14899 (N_14899,N_14434,N_14463);
and U14900 (N_14900,N_14687,N_14682);
xnor U14901 (N_14901,N_14562,N_14485);
or U14902 (N_14902,N_14515,N_14621);
and U14903 (N_14903,N_14611,N_14647);
nand U14904 (N_14904,N_14495,N_14475);
xor U14905 (N_14905,N_14678,N_14479);
xor U14906 (N_14906,N_14669,N_14690);
nand U14907 (N_14907,N_14444,N_14673);
nor U14908 (N_14908,N_14526,N_14522);
xor U14909 (N_14909,N_14445,N_14688);
nand U14910 (N_14910,N_14550,N_14617);
xor U14911 (N_14911,N_14656,N_14571);
xor U14912 (N_14912,N_14459,N_14568);
nand U14913 (N_14913,N_14574,N_14469);
nand U14914 (N_14914,N_14497,N_14431);
nor U14915 (N_14915,N_14451,N_14602);
nand U14916 (N_14916,N_14459,N_14602);
and U14917 (N_14917,N_14547,N_14461);
nor U14918 (N_14918,N_14485,N_14447);
and U14919 (N_14919,N_14636,N_14588);
or U14920 (N_14920,N_14698,N_14683);
and U14921 (N_14921,N_14553,N_14400);
nand U14922 (N_14922,N_14648,N_14493);
and U14923 (N_14923,N_14495,N_14516);
or U14924 (N_14924,N_14627,N_14650);
or U14925 (N_14925,N_14496,N_14492);
and U14926 (N_14926,N_14665,N_14641);
or U14927 (N_14927,N_14515,N_14411);
xor U14928 (N_14928,N_14443,N_14681);
and U14929 (N_14929,N_14513,N_14410);
and U14930 (N_14930,N_14575,N_14615);
and U14931 (N_14931,N_14433,N_14550);
and U14932 (N_14932,N_14462,N_14406);
or U14933 (N_14933,N_14683,N_14569);
nor U14934 (N_14934,N_14671,N_14505);
and U14935 (N_14935,N_14561,N_14499);
nor U14936 (N_14936,N_14555,N_14573);
nor U14937 (N_14937,N_14539,N_14592);
and U14938 (N_14938,N_14602,N_14684);
nor U14939 (N_14939,N_14520,N_14611);
and U14940 (N_14940,N_14674,N_14590);
nand U14941 (N_14941,N_14509,N_14559);
or U14942 (N_14942,N_14686,N_14430);
nor U14943 (N_14943,N_14585,N_14544);
nand U14944 (N_14944,N_14515,N_14567);
nand U14945 (N_14945,N_14699,N_14667);
and U14946 (N_14946,N_14427,N_14428);
or U14947 (N_14947,N_14594,N_14606);
nor U14948 (N_14948,N_14530,N_14562);
xor U14949 (N_14949,N_14514,N_14453);
xnor U14950 (N_14950,N_14559,N_14478);
and U14951 (N_14951,N_14402,N_14531);
xor U14952 (N_14952,N_14563,N_14613);
or U14953 (N_14953,N_14594,N_14566);
or U14954 (N_14954,N_14682,N_14582);
nand U14955 (N_14955,N_14409,N_14513);
or U14956 (N_14956,N_14616,N_14515);
xnor U14957 (N_14957,N_14510,N_14586);
or U14958 (N_14958,N_14696,N_14555);
and U14959 (N_14959,N_14632,N_14602);
nand U14960 (N_14960,N_14511,N_14599);
nor U14961 (N_14961,N_14610,N_14457);
nor U14962 (N_14962,N_14462,N_14451);
nand U14963 (N_14963,N_14514,N_14446);
and U14964 (N_14964,N_14476,N_14516);
and U14965 (N_14965,N_14621,N_14610);
nand U14966 (N_14966,N_14464,N_14454);
or U14967 (N_14967,N_14671,N_14423);
and U14968 (N_14968,N_14522,N_14617);
or U14969 (N_14969,N_14555,N_14519);
nor U14970 (N_14970,N_14610,N_14546);
nor U14971 (N_14971,N_14496,N_14469);
xnor U14972 (N_14972,N_14503,N_14466);
nand U14973 (N_14973,N_14608,N_14480);
or U14974 (N_14974,N_14537,N_14641);
nor U14975 (N_14975,N_14591,N_14550);
nand U14976 (N_14976,N_14688,N_14602);
or U14977 (N_14977,N_14435,N_14483);
or U14978 (N_14978,N_14461,N_14567);
and U14979 (N_14979,N_14606,N_14666);
and U14980 (N_14980,N_14447,N_14525);
nand U14981 (N_14981,N_14695,N_14429);
nor U14982 (N_14982,N_14669,N_14494);
xnor U14983 (N_14983,N_14461,N_14404);
or U14984 (N_14984,N_14503,N_14552);
xor U14985 (N_14985,N_14508,N_14531);
xor U14986 (N_14986,N_14629,N_14606);
nor U14987 (N_14987,N_14401,N_14689);
nand U14988 (N_14988,N_14582,N_14425);
nand U14989 (N_14989,N_14666,N_14433);
or U14990 (N_14990,N_14426,N_14576);
nor U14991 (N_14991,N_14620,N_14678);
and U14992 (N_14992,N_14596,N_14407);
xor U14993 (N_14993,N_14589,N_14525);
nand U14994 (N_14994,N_14495,N_14606);
xnor U14995 (N_14995,N_14603,N_14693);
nor U14996 (N_14996,N_14553,N_14446);
or U14997 (N_14997,N_14678,N_14490);
and U14998 (N_14998,N_14567,N_14673);
xnor U14999 (N_14999,N_14575,N_14500);
nand UO_0 (O_0,N_14903,N_14705);
nor UO_1 (O_1,N_14778,N_14863);
nor UO_2 (O_2,N_14885,N_14779);
xnor UO_3 (O_3,N_14988,N_14898);
nor UO_4 (O_4,N_14743,N_14809);
and UO_5 (O_5,N_14973,N_14919);
and UO_6 (O_6,N_14733,N_14747);
or UO_7 (O_7,N_14785,N_14766);
xor UO_8 (O_8,N_14897,N_14707);
and UO_9 (O_9,N_14940,N_14794);
or UO_10 (O_10,N_14920,N_14822);
or UO_11 (O_11,N_14726,N_14955);
and UO_12 (O_12,N_14929,N_14839);
nand UO_13 (O_13,N_14811,N_14717);
nor UO_14 (O_14,N_14770,N_14964);
or UO_15 (O_15,N_14953,N_14710);
and UO_16 (O_16,N_14819,N_14891);
xnor UO_17 (O_17,N_14798,N_14928);
nor UO_18 (O_18,N_14909,N_14817);
nor UO_19 (O_19,N_14951,N_14886);
xor UO_20 (O_20,N_14744,N_14915);
nand UO_21 (O_21,N_14758,N_14737);
or UO_22 (O_22,N_14847,N_14944);
or UO_23 (O_23,N_14876,N_14760);
or UO_24 (O_24,N_14967,N_14948);
nand UO_25 (O_25,N_14816,N_14712);
nand UO_26 (O_26,N_14983,N_14856);
nor UO_27 (O_27,N_14959,N_14804);
and UO_28 (O_28,N_14729,N_14939);
xnor UO_29 (O_29,N_14889,N_14751);
and UO_30 (O_30,N_14767,N_14974);
or UO_31 (O_31,N_14802,N_14880);
or UO_32 (O_32,N_14957,N_14949);
or UO_33 (O_33,N_14821,N_14986);
nand UO_34 (O_34,N_14810,N_14771);
and UO_35 (O_35,N_14888,N_14952);
nand UO_36 (O_36,N_14947,N_14950);
nand UO_37 (O_37,N_14818,N_14987);
or UO_38 (O_38,N_14812,N_14994);
xnor UO_39 (O_39,N_14901,N_14725);
xnor UO_40 (O_40,N_14752,N_14993);
and UO_41 (O_41,N_14713,N_14941);
or UO_42 (O_42,N_14746,N_14872);
nor UO_43 (O_43,N_14899,N_14700);
nor UO_44 (O_44,N_14765,N_14956);
nand UO_45 (O_45,N_14851,N_14735);
or UO_46 (O_46,N_14775,N_14991);
xnor UO_47 (O_47,N_14908,N_14721);
xnor UO_48 (O_48,N_14756,N_14992);
and UO_49 (O_49,N_14861,N_14722);
nand UO_50 (O_50,N_14706,N_14926);
nand UO_51 (O_51,N_14893,N_14784);
and UO_52 (O_52,N_14961,N_14946);
and UO_53 (O_53,N_14868,N_14931);
and UO_54 (O_54,N_14971,N_14764);
or UO_55 (O_55,N_14724,N_14792);
nor UO_56 (O_56,N_14836,N_14815);
nor UO_57 (O_57,N_14843,N_14846);
nor UO_58 (O_58,N_14989,N_14823);
and UO_59 (O_59,N_14854,N_14966);
and UO_60 (O_60,N_14984,N_14832);
and UO_61 (O_61,N_14896,N_14921);
and UO_62 (O_62,N_14781,N_14871);
or UO_63 (O_63,N_14910,N_14795);
nor UO_64 (O_64,N_14783,N_14938);
nand UO_65 (O_65,N_14867,N_14805);
nor UO_66 (O_66,N_14808,N_14803);
or UO_67 (O_67,N_14999,N_14776);
xor UO_68 (O_68,N_14845,N_14906);
xnor UO_69 (O_69,N_14933,N_14954);
or UO_70 (O_70,N_14749,N_14895);
xor UO_71 (O_71,N_14780,N_14934);
or UO_72 (O_72,N_14719,N_14978);
nand UO_73 (O_73,N_14820,N_14790);
or UO_74 (O_74,N_14761,N_14740);
nand UO_75 (O_75,N_14985,N_14890);
xor UO_76 (O_76,N_14828,N_14741);
and UO_77 (O_77,N_14731,N_14704);
nand UO_78 (O_78,N_14745,N_14757);
or UO_79 (O_79,N_14976,N_14945);
and UO_80 (O_80,N_14918,N_14972);
nor UO_81 (O_81,N_14701,N_14981);
and UO_82 (O_82,N_14883,N_14807);
nand UO_83 (O_83,N_14936,N_14734);
nor UO_84 (O_84,N_14777,N_14924);
or UO_85 (O_85,N_14869,N_14727);
and UO_86 (O_86,N_14716,N_14732);
nand UO_87 (O_87,N_14904,N_14759);
nand UO_88 (O_88,N_14848,N_14857);
xnor UO_89 (O_89,N_14997,N_14742);
nor UO_90 (O_90,N_14878,N_14830);
or UO_91 (O_91,N_14937,N_14858);
xnor UO_92 (O_92,N_14942,N_14838);
or UO_93 (O_93,N_14873,N_14962);
xnor UO_94 (O_94,N_14927,N_14907);
and UO_95 (O_95,N_14827,N_14958);
and UO_96 (O_96,N_14829,N_14826);
or UO_97 (O_97,N_14702,N_14894);
nand UO_98 (O_98,N_14849,N_14865);
nand UO_99 (O_99,N_14835,N_14975);
nand UO_100 (O_100,N_14853,N_14916);
xnor UO_101 (O_101,N_14968,N_14750);
nor UO_102 (O_102,N_14960,N_14982);
nor UO_103 (O_103,N_14925,N_14738);
or UO_104 (O_104,N_14754,N_14862);
xnor UO_105 (O_105,N_14844,N_14806);
xnor UO_106 (O_106,N_14730,N_14748);
nand UO_107 (O_107,N_14753,N_14833);
nand UO_108 (O_108,N_14932,N_14789);
xnor UO_109 (O_109,N_14902,N_14814);
xnor UO_110 (O_110,N_14892,N_14917);
xor UO_111 (O_111,N_14728,N_14980);
or UO_112 (O_112,N_14723,N_14739);
or UO_113 (O_113,N_14793,N_14990);
nand UO_114 (O_114,N_14841,N_14720);
nor UO_115 (O_115,N_14996,N_14905);
nor UO_116 (O_116,N_14773,N_14995);
xnor UO_117 (O_117,N_14879,N_14866);
nor UO_118 (O_118,N_14840,N_14922);
or UO_119 (O_119,N_14970,N_14969);
nand UO_120 (O_120,N_14837,N_14800);
xnor UO_121 (O_121,N_14887,N_14703);
or UO_122 (O_122,N_14979,N_14855);
or UO_123 (O_123,N_14755,N_14786);
or UO_124 (O_124,N_14965,N_14852);
and UO_125 (O_125,N_14762,N_14782);
and UO_126 (O_126,N_14963,N_14831);
nor UO_127 (O_127,N_14774,N_14875);
or UO_128 (O_128,N_14714,N_14881);
and UO_129 (O_129,N_14711,N_14912);
nand UO_130 (O_130,N_14882,N_14797);
nor UO_131 (O_131,N_14736,N_14718);
or UO_132 (O_132,N_14860,N_14801);
or UO_133 (O_133,N_14850,N_14791);
nand UO_134 (O_134,N_14842,N_14799);
and UO_135 (O_135,N_14877,N_14813);
xnor UO_136 (O_136,N_14769,N_14900);
or UO_137 (O_137,N_14923,N_14768);
nand UO_138 (O_138,N_14998,N_14709);
and UO_139 (O_139,N_14874,N_14796);
nand UO_140 (O_140,N_14935,N_14763);
nand UO_141 (O_141,N_14825,N_14787);
xor UO_142 (O_142,N_14943,N_14715);
xor UO_143 (O_143,N_14864,N_14870);
nor UO_144 (O_144,N_14772,N_14930);
nand UO_145 (O_145,N_14859,N_14824);
nor UO_146 (O_146,N_14788,N_14884);
or UO_147 (O_147,N_14913,N_14914);
nor UO_148 (O_148,N_14977,N_14834);
nor UO_149 (O_149,N_14911,N_14708);
xor UO_150 (O_150,N_14753,N_14771);
and UO_151 (O_151,N_14993,N_14861);
nand UO_152 (O_152,N_14967,N_14987);
or UO_153 (O_153,N_14752,N_14875);
or UO_154 (O_154,N_14789,N_14968);
or UO_155 (O_155,N_14994,N_14948);
or UO_156 (O_156,N_14754,N_14890);
xor UO_157 (O_157,N_14712,N_14838);
xnor UO_158 (O_158,N_14816,N_14740);
and UO_159 (O_159,N_14739,N_14957);
nor UO_160 (O_160,N_14836,N_14741);
or UO_161 (O_161,N_14700,N_14770);
xnor UO_162 (O_162,N_14883,N_14967);
xnor UO_163 (O_163,N_14838,N_14722);
nand UO_164 (O_164,N_14927,N_14774);
nor UO_165 (O_165,N_14871,N_14979);
nand UO_166 (O_166,N_14958,N_14742);
xor UO_167 (O_167,N_14849,N_14789);
xnor UO_168 (O_168,N_14740,N_14951);
nor UO_169 (O_169,N_14763,N_14890);
and UO_170 (O_170,N_14992,N_14887);
and UO_171 (O_171,N_14930,N_14831);
and UO_172 (O_172,N_14723,N_14996);
xor UO_173 (O_173,N_14974,N_14764);
xnor UO_174 (O_174,N_14950,N_14823);
nand UO_175 (O_175,N_14981,N_14819);
xnor UO_176 (O_176,N_14911,N_14875);
nand UO_177 (O_177,N_14720,N_14739);
xnor UO_178 (O_178,N_14865,N_14916);
nand UO_179 (O_179,N_14858,N_14792);
or UO_180 (O_180,N_14989,N_14873);
and UO_181 (O_181,N_14766,N_14984);
and UO_182 (O_182,N_14994,N_14959);
nand UO_183 (O_183,N_14733,N_14867);
and UO_184 (O_184,N_14972,N_14818);
and UO_185 (O_185,N_14943,N_14817);
and UO_186 (O_186,N_14985,N_14940);
and UO_187 (O_187,N_14959,N_14992);
or UO_188 (O_188,N_14903,N_14841);
or UO_189 (O_189,N_14725,N_14880);
nand UO_190 (O_190,N_14884,N_14782);
or UO_191 (O_191,N_14949,N_14829);
or UO_192 (O_192,N_14834,N_14835);
nand UO_193 (O_193,N_14850,N_14977);
xor UO_194 (O_194,N_14864,N_14929);
nand UO_195 (O_195,N_14992,N_14856);
xnor UO_196 (O_196,N_14931,N_14901);
xor UO_197 (O_197,N_14787,N_14903);
and UO_198 (O_198,N_14839,N_14819);
xor UO_199 (O_199,N_14734,N_14744);
nand UO_200 (O_200,N_14787,N_14745);
xor UO_201 (O_201,N_14855,N_14707);
nand UO_202 (O_202,N_14845,N_14766);
nor UO_203 (O_203,N_14840,N_14848);
xnor UO_204 (O_204,N_14989,N_14905);
nor UO_205 (O_205,N_14765,N_14992);
and UO_206 (O_206,N_14931,N_14774);
nand UO_207 (O_207,N_14980,N_14811);
or UO_208 (O_208,N_14837,N_14790);
and UO_209 (O_209,N_14880,N_14967);
or UO_210 (O_210,N_14799,N_14986);
nand UO_211 (O_211,N_14733,N_14761);
nor UO_212 (O_212,N_14851,N_14865);
nor UO_213 (O_213,N_14828,N_14726);
nor UO_214 (O_214,N_14790,N_14850);
or UO_215 (O_215,N_14846,N_14927);
nor UO_216 (O_216,N_14845,N_14774);
and UO_217 (O_217,N_14846,N_14866);
or UO_218 (O_218,N_14887,N_14755);
nand UO_219 (O_219,N_14701,N_14891);
xnor UO_220 (O_220,N_14812,N_14848);
xor UO_221 (O_221,N_14919,N_14989);
and UO_222 (O_222,N_14824,N_14971);
nor UO_223 (O_223,N_14823,N_14786);
nand UO_224 (O_224,N_14920,N_14841);
xor UO_225 (O_225,N_14849,N_14980);
xnor UO_226 (O_226,N_14858,N_14892);
nor UO_227 (O_227,N_14709,N_14959);
nor UO_228 (O_228,N_14901,N_14719);
xnor UO_229 (O_229,N_14819,N_14820);
and UO_230 (O_230,N_14787,N_14885);
or UO_231 (O_231,N_14722,N_14783);
or UO_232 (O_232,N_14812,N_14767);
or UO_233 (O_233,N_14725,N_14732);
or UO_234 (O_234,N_14906,N_14798);
nor UO_235 (O_235,N_14929,N_14977);
nand UO_236 (O_236,N_14735,N_14954);
nand UO_237 (O_237,N_14894,N_14995);
xor UO_238 (O_238,N_14926,N_14959);
and UO_239 (O_239,N_14829,N_14966);
xor UO_240 (O_240,N_14856,N_14728);
or UO_241 (O_241,N_14874,N_14839);
xor UO_242 (O_242,N_14969,N_14914);
or UO_243 (O_243,N_14782,N_14806);
nand UO_244 (O_244,N_14753,N_14985);
xnor UO_245 (O_245,N_14714,N_14931);
or UO_246 (O_246,N_14993,N_14826);
or UO_247 (O_247,N_14706,N_14747);
or UO_248 (O_248,N_14855,N_14829);
or UO_249 (O_249,N_14843,N_14738);
or UO_250 (O_250,N_14924,N_14864);
or UO_251 (O_251,N_14738,N_14742);
nor UO_252 (O_252,N_14859,N_14729);
or UO_253 (O_253,N_14921,N_14803);
or UO_254 (O_254,N_14763,N_14932);
and UO_255 (O_255,N_14960,N_14838);
nand UO_256 (O_256,N_14867,N_14760);
xnor UO_257 (O_257,N_14720,N_14952);
nor UO_258 (O_258,N_14915,N_14812);
nor UO_259 (O_259,N_14967,N_14989);
xor UO_260 (O_260,N_14914,N_14800);
and UO_261 (O_261,N_14823,N_14814);
nand UO_262 (O_262,N_14782,N_14879);
xor UO_263 (O_263,N_14881,N_14922);
nor UO_264 (O_264,N_14794,N_14978);
nand UO_265 (O_265,N_14890,N_14785);
nand UO_266 (O_266,N_14709,N_14873);
or UO_267 (O_267,N_14702,N_14876);
nand UO_268 (O_268,N_14890,N_14819);
nand UO_269 (O_269,N_14765,N_14983);
nor UO_270 (O_270,N_14962,N_14989);
nor UO_271 (O_271,N_14941,N_14873);
nand UO_272 (O_272,N_14855,N_14830);
xor UO_273 (O_273,N_14994,N_14727);
nor UO_274 (O_274,N_14967,N_14930);
nor UO_275 (O_275,N_14944,N_14935);
and UO_276 (O_276,N_14817,N_14803);
xnor UO_277 (O_277,N_14924,N_14819);
nand UO_278 (O_278,N_14850,N_14933);
or UO_279 (O_279,N_14761,N_14714);
xnor UO_280 (O_280,N_14713,N_14760);
and UO_281 (O_281,N_14851,N_14997);
xnor UO_282 (O_282,N_14865,N_14909);
nor UO_283 (O_283,N_14701,N_14877);
or UO_284 (O_284,N_14930,N_14724);
and UO_285 (O_285,N_14987,N_14883);
nor UO_286 (O_286,N_14774,N_14778);
nor UO_287 (O_287,N_14798,N_14749);
nand UO_288 (O_288,N_14789,N_14921);
nor UO_289 (O_289,N_14804,N_14737);
nand UO_290 (O_290,N_14799,N_14843);
or UO_291 (O_291,N_14835,N_14727);
or UO_292 (O_292,N_14724,N_14987);
and UO_293 (O_293,N_14889,N_14855);
or UO_294 (O_294,N_14900,N_14747);
and UO_295 (O_295,N_14807,N_14948);
and UO_296 (O_296,N_14742,N_14701);
nand UO_297 (O_297,N_14750,N_14839);
and UO_298 (O_298,N_14981,N_14835);
xnor UO_299 (O_299,N_14827,N_14862);
nand UO_300 (O_300,N_14824,N_14735);
nand UO_301 (O_301,N_14839,N_14907);
nand UO_302 (O_302,N_14855,N_14905);
nand UO_303 (O_303,N_14800,N_14769);
nand UO_304 (O_304,N_14957,N_14869);
xnor UO_305 (O_305,N_14999,N_14952);
nor UO_306 (O_306,N_14864,N_14787);
and UO_307 (O_307,N_14795,N_14728);
or UO_308 (O_308,N_14901,N_14912);
or UO_309 (O_309,N_14898,N_14998);
or UO_310 (O_310,N_14889,N_14794);
or UO_311 (O_311,N_14899,N_14957);
nand UO_312 (O_312,N_14773,N_14775);
nor UO_313 (O_313,N_14994,N_14831);
and UO_314 (O_314,N_14998,N_14920);
nand UO_315 (O_315,N_14827,N_14822);
or UO_316 (O_316,N_14940,N_14814);
xnor UO_317 (O_317,N_14714,N_14743);
and UO_318 (O_318,N_14941,N_14903);
nor UO_319 (O_319,N_14773,N_14785);
and UO_320 (O_320,N_14720,N_14842);
and UO_321 (O_321,N_14980,N_14751);
nor UO_322 (O_322,N_14768,N_14919);
xor UO_323 (O_323,N_14996,N_14975);
nand UO_324 (O_324,N_14894,N_14751);
nor UO_325 (O_325,N_14713,N_14969);
nand UO_326 (O_326,N_14756,N_14790);
and UO_327 (O_327,N_14836,N_14841);
or UO_328 (O_328,N_14900,N_14784);
xnor UO_329 (O_329,N_14897,N_14755);
nor UO_330 (O_330,N_14895,N_14727);
nand UO_331 (O_331,N_14924,N_14862);
nor UO_332 (O_332,N_14793,N_14839);
and UO_333 (O_333,N_14838,N_14743);
xor UO_334 (O_334,N_14993,N_14809);
nand UO_335 (O_335,N_14789,N_14797);
nor UO_336 (O_336,N_14825,N_14829);
and UO_337 (O_337,N_14813,N_14796);
or UO_338 (O_338,N_14719,N_14836);
nor UO_339 (O_339,N_14879,N_14703);
nand UO_340 (O_340,N_14954,N_14729);
nor UO_341 (O_341,N_14710,N_14820);
or UO_342 (O_342,N_14894,N_14780);
xnor UO_343 (O_343,N_14808,N_14825);
nand UO_344 (O_344,N_14903,N_14966);
nand UO_345 (O_345,N_14825,N_14939);
nor UO_346 (O_346,N_14942,N_14857);
and UO_347 (O_347,N_14714,N_14735);
or UO_348 (O_348,N_14801,N_14755);
nand UO_349 (O_349,N_14823,N_14959);
xnor UO_350 (O_350,N_14862,N_14912);
or UO_351 (O_351,N_14974,N_14914);
nand UO_352 (O_352,N_14955,N_14821);
xnor UO_353 (O_353,N_14712,N_14878);
nand UO_354 (O_354,N_14927,N_14819);
nor UO_355 (O_355,N_14929,N_14701);
nor UO_356 (O_356,N_14736,N_14721);
nand UO_357 (O_357,N_14956,N_14952);
xor UO_358 (O_358,N_14956,N_14999);
nor UO_359 (O_359,N_14726,N_14717);
xnor UO_360 (O_360,N_14919,N_14740);
nand UO_361 (O_361,N_14746,N_14844);
nand UO_362 (O_362,N_14958,N_14780);
xor UO_363 (O_363,N_14999,N_14841);
nor UO_364 (O_364,N_14758,N_14700);
nand UO_365 (O_365,N_14797,N_14844);
or UO_366 (O_366,N_14786,N_14803);
or UO_367 (O_367,N_14801,N_14913);
xor UO_368 (O_368,N_14863,N_14937);
and UO_369 (O_369,N_14915,N_14955);
nor UO_370 (O_370,N_14777,N_14887);
xor UO_371 (O_371,N_14747,N_14838);
or UO_372 (O_372,N_14702,N_14994);
nor UO_373 (O_373,N_14792,N_14980);
xor UO_374 (O_374,N_14720,N_14722);
nand UO_375 (O_375,N_14809,N_14979);
xnor UO_376 (O_376,N_14853,N_14714);
nor UO_377 (O_377,N_14976,N_14831);
xnor UO_378 (O_378,N_14907,N_14883);
xor UO_379 (O_379,N_14766,N_14875);
or UO_380 (O_380,N_14875,N_14888);
nor UO_381 (O_381,N_14893,N_14923);
xor UO_382 (O_382,N_14895,N_14918);
nand UO_383 (O_383,N_14902,N_14904);
and UO_384 (O_384,N_14871,N_14829);
nor UO_385 (O_385,N_14894,N_14820);
and UO_386 (O_386,N_14742,N_14894);
xnor UO_387 (O_387,N_14895,N_14863);
xor UO_388 (O_388,N_14858,N_14822);
nand UO_389 (O_389,N_14733,N_14712);
and UO_390 (O_390,N_14977,N_14739);
xnor UO_391 (O_391,N_14937,N_14998);
or UO_392 (O_392,N_14931,N_14884);
or UO_393 (O_393,N_14805,N_14745);
and UO_394 (O_394,N_14826,N_14972);
xnor UO_395 (O_395,N_14871,N_14948);
xnor UO_396 (O_396,N_14882,N_14731);
xnor UO_397 (O_397,N_14802,N_14894);
and UO_398 (O_398,N_14940,N_14990);
nor UO_399 (O_399,N_14942,N_14727);
nand UO_400 (O_400,N_14979,N_14733);
xor UO_401 (O_401,N_14756,N_14906);
and UO_402 (O_402,N_14830,N_14764);
xor UO_403 (O_403,N_14831,N_14700);
xor UO_404 (O_404,N_14880,N_14731);
xor UO_405 (O_405,N_14843,N_14965);
nor UO_406 (O_406,N_14744,N_14837);
and UO_407 (O_407,N_14829,N_14742);
xnor UO_408 (O_408,N_14993,N_14784);
nand UO_409 (O_409,N_14899,N_14988);
nor UO_410 (O_410,N_14750,N_14944);
and UO_411 (O_411,N_14965,N_14912);
nor UO_412 (O_412,N_14963,N_14900);
or UO_413 (O_413,N_14836,N_14863);
nor UO_414 (O_414,N_14932,N_14873);
xnor UO_415 (O_415,N_14853,N_14829);
nor UO_416 (O_416,N_14890,N_14817);
nand UO_417 (O_417,N_14852,N_14879);
or UO_418 (O_418,N_14908,N_14865);
xnor UO_419 (O_419,N_14930,N_14883);
and UO_420 (O_420,N_14866,N_14783);
nand UO_421 (O_421,N_14795,N_14862);
nor UO_422 (O_422,N_14733,N_14784);
nand UO_423 (O_423,N_14922,N_14720);
nand UO_424 (O_424,N_14995,N_14861);
or UO_425 (O_425,N_14749,N_14887);
nand UO_426 (O_426,N_14711,N_14816);
or UO_427 (O_427,N_14793,N_14988);
nand UO_428 (O_428,N_14842,N_14731);
nand UO_429 (O_429,N_14973,N_14980);
xnor UO_430 (O_430,N_14972,N_14910);
nand UO_431 (O_431,N_14902,N_14711);
xor UO_432 (O_432,N_14779,N_14724);
and UO_433 (O_433,N_14889,N_14947);
or UO_434 (O_434,N_14983,N_14708);
and UO_435 (O_435,N_14757,N_14989);
xor UO_436 (O_436,N_14845,N_14773);
nand UO_437 (O_437,N_14885,N_14826);
xor UO_438 (O_438,N_14963,N_14955);
and UO_439 (O_439,N_14884,N_14774);
and UO_440 (O_440,N_14727,N_14930);
xnor UO_441 (O_441,N_14862,N_14958);
and UO_442 (O_442,N_14811,N_14777);
nor UO_443 (O_443,N_14827,N_14879);
nand UO_444 (O_444,N_14932,N_14927);
nand UO_445 (O_445,N_14990,N_14782);
nand UO_446 (O_446,N_14957,N_14711);
and UO_447 (O_447,N_14739,N_14747);
nor UO_448 (O_448,N_14789,N_14722);
nor UO_449 (O_449,N_14791,N_14992);
and UO_450 (O_450,N_14934,N_14969);
or UO_451 (O_451,N_14757,N_14996);
nor UO_452 (O_452,N_14818,N_14721);
and UO_453 (O_453,N_14771,N_14750);
xnor UO_454 (O_454,N_14871,N_14958);
and UO_455 (O_455,N_14954,N_14977);
xor UO_456 (O_456,N_14926,N_14794);
and UO_457 (O_457,N_14917,N_14713);
and UO_458 (O_458,N_14781,N_14987);
xnor UO_459 (O_459,N_14823,N_14996);
and UO_460 (O_460,N_14833,N_14923);
nor UO_461 (O_461,N_14717,N_14902);
xor UO_462 (O_462,N_14778,N_14855);
or UO_463 (O_463,N_14725,N_14857);
nand UO_464 (O_464,N_14901,N_14996);
nor UO_465 (O_465,N_14927,N_14999);
nand UO_466 (O_466,N_14953,N_14764);
nand UO_467 (O_467,N_14870,N_14894);
and UO_468 (O_468,N_14971,N_14834);
xnor UO_469 (O_469,N_14712,N_14722);
and UO_470 (O_470,N_14712,N_14736);
or UO_471 (O_471,N_14757,N_14952);
or UO_472 (O_472,N_14857,N_14893);
nor UO_473 (O_473,N_14983,N_14864);
xor UO_474 (O_474,N_14726,N_14744);
and UO_475 (O_475,N_14796,N_14754);
and UO_476 (O_476,N_14873,N_14864);
nor UO_477 (O_477,N_14828,N_14952);
xor UO_478 (O_478,N_14940,N_14901);
or UO_479 (O_479,N_14703,N_14797);
or UO_480 (O_480,N_14995,N_14842);
xor UO_481 (O_481,N_14703,N_14956);
nand UO_482 (O_482,N_14979,N_14836);
and UO_483 (O_483,N_14866,N_14882);
or UO_484 (O_484,N_14943,N_14706);
nand UO_485 (O_485,N_14754,N_14865);
or UO_486 (O_486,N_14876,N_14966);
or UO_487 (O_487,N_14715,N_14724);
xor UO_488 (O_488,N_14924,N_14725);
and UO_489 (O_489,N_14829,N_14752);
nand UO_490 (O_490,N_14836,N_14881);
nor UO_491 (O_491,N_14852,N_14863);
nor UO_492 (O_492,N_14954,N_14866);
xor UO_493 (O_493,N_14832,N_14913);
and UO_494 (O_494,N_14785,N_14779);
nor UO_495 (O_495,N_14917,N_14968);
and UO_496 (O_496,N_14854,N_14897);
xnor UO_497 (O_497,N_14944,N_14842);
nand UO_498 (O_498,N_14880,N_14799);
xor UO_499 (O_499,N_14920,N_14849);
xor UO_500 (O_500,N_14810,N_14991);
and UO_501 (O_501,N_14728,N_14764);
nand UO_502 (O_502,N_14731,N_14945);
or UO_503 (O_503,N_14728,N_14868);
and UO_504 (O_504,N_14833,N_14721);
and UO_505 (O_505,N_14831,N_14884);
nor UO_506 (O_506,N_14778,N_14875);
or UO_507 (O_507,N_14943,N_14927);
nand UO_508 (O_508,N_14961,N_14970);
xor UO_509 (O_509,N_14918,N_14866);
xor UO_510 (O_510,N_14758,N_14878);
and UO_511 (O_511,N_14972,N_14932);
xnor UO_512 (O_512,N_14819,N_14857);
xnor UO_513 (O_513,N_14859,N_14920);
or UO_514 (O_514,N_14941,N_14926);
nor UO_515 (O_515,N_14840,N_14830);
nand UO_516 (O_516,N_14872,N_14948);
nor UO_517 (O_517,N_14852,N_14833);
xor UO_518 (O_518,N_14898,N_14985);
nand UO_519 (O_519,N_14916,N_14840);
nand UO_520 (O_520,N_14751,N_14748);
nand UO_521 (O_521,N_14798,N_14756);
xnor UO_522 (O_522,N_14771,N_14756);
and UO_523 (O_523,N_14950,N_14839);
or UO_524 (O_524,N_14919,N_14991);
or UO_525 (O_525,N_14984,N_14925);
nand UO_526 (O_526,N_14990,N_14767);
nand UO_527 (O_527,N_14834,N_14945);
xor UO_528 (O_528,N_14863,N_14886);
nand UO_529 (O_529,N_14815,N_14911);
or UO_530 (O_530,N_14862,N_14896);
nor UO_531 (O_531,N_14796,N_14824);
and UO_532 (O_532,N_14757,N_14868);
nand UO_533 (O_533,N_14749,N_14826);
and UO_534 (O_534,N_14767,N_14880);
nand UO_535 (O_535,N_14905,N_14732);
xor UO_536 (O_536,N_14735,N_14718);
xnor UO_537 (O_537,N_14770,N_14858);
nor UO_538 (O_538,N_14822,N_14767);
or UO_539 (O_539,N_14704,N_14887);
nor UO_540 (O_540,N_14846,N_14971);
nor UO_541 (O_541,N_14747,N_14817);
nand UO_542 (O_542,N_14839,N_14806);
xnor UO_543 (O_543,N_14758,N_14847);
and UO_544 (O_544,N_14751,N_14865);
and UO_545 (O_545,N_14780,N_14870);
or UO_546 (O_546,N_14902,N_14915);
or UO_547 (O_547,N_14994,N_14910);
and UO_548 (O_548,N_14982,N_14967);
or UO_549 (O_549,N_14734,N_14849);
or UO_550 (O_550,N_14790,N_14766);
xor UO_551 (O_551,N_14894,N_14781);
nor UO_552 (O_552,N_14810,N_14760);
xor UO_553 (O_553,N_14902,N_14724);
nor UO_554 (O_554,N_14846,N_14946);
nor UO_555 (O_555,N_14961,N_14706);
or UO_556 (O_556,N_14875,N_14898);
or UO_557 (O_557,N_14919,N_14722);
or UO_558 (O_558,N_14820,N_14837);
xor UO_559 (O_559,N_14972,N_14864);
nand UO_560 (O_560,N_14766,N_14737);
xnor UO_561 (O_561,N_14949,N_14734);
or UO_562 (O_562,N_14900,N_14998);
xor UO_563 (O_563,N_14926,N_14854);
or UO_564 (O_564,N_14938,N_14725);
xnor UO_565 (O_565,N_14705,N_14763);
xor UO_566 (O_566,N_14721,N_14916);
and UO_567 (O_567,N_14992,N_14710);
and UO_568 (O_568,N_14992,N_14748);
nor UO_569 (O_569,N_14838,N_14898);
nand UO_570 (O_570,N_14948,N_14766);
nor UO_571 (O_571,N_14911,N_14987);
and UO_572 (O_572,N_14977,N_14941);
nand UO_573 (O_573,N_14803,N_14802);
or UO_574 (O_574,N_14966,N_14938);
nand UO_575 (O_575,N_14738,N_14934);
nor UO_576 (O_576,N_14903,N_14973);
xor UO_577 (O_577,N_14775,N_14929);
nor UO_578 (O_578,N_14936,N_14872);
or UO_579 (O_579,N_14722,N_14868);
nor UO_580 (O_580,N_14956,N_14725);
or UO_581 (O_581,N_14993,N_14713);
and UO_582 (O_582,N_14991,N_14970);
nor UO_583 (O_583,N_14983,N_14975);
nor UO_584 (O_584,N_14960,N_14834);
nand UO_585 (O_585,N_14862,N_14718);
nand UO_586 (O_586,N_14908,N_14938);
xnor UO_587 (O_587,N_14979,N_14837);
or UO_588 (O_588,N_14744,N_14787);
nand UO_589 (O_589,N_14931,N_14850);
xnor UO_590 (O_590,N_14734,N_14755);
or UO_591 (O_591,N_14734,N_14906);
nor UO_592 (O_592,N_14707,N_14941);
and UO_593 (O_593,N_14813,N_14936);
and UO_594 (O_594,N_14824,N_14871);
xor UO_595 (O_595,N_14703,N_14993);
nor UO_596 (O_596,N_14929,N_14805);
nor UO_597 (O_597,N_14971,N_14719);
or UO_598 (O_598,N_14930,N_14885);
nor UO_599 (O_599,N_14963,N_14787);
xor UO_600 (O_600,N_14868,N_14782);
or UO_601 (O_601,N_14737,N_14935);
and UO_602 (O_602,N_14857,N_14856);
and UO_603 (O_603,N_14881,N_14733);
or UO_604 (O_604,N_14831,N_14868);
or UO_605 (O_605,N_14922,N_14899);
or UO_606 (O_606,N_14812,N_14755);
nor UO_607 (O_607,N_14850,N_14741);
nand UO_608 (O_608,N_14860,N_14847);
nor UO_609 (O_609,N_14838,N_14794);
xor UO_610 (O_610,N_14773,N_14977);
and UO_611 (O_611,N_14913,N_14964);
or UO_612 (O_612,N_14791,N_14835);
xnor UO_613 (O_613,N_14780,N_14885);
xnor UO_614 (O_614,N_14901,N_14836);
or UO_615 (O_615,N_14753,N_14823);
nand UO_616 (O_616,N_14756,N_14736);
xor UO_617 (O_617,N_14865,N_14788);
or UO_618 (O_618,N_14743,N_14833);
or UO_619 (O_619,N_14977,N_14764);
xnor UO_620 (O_620,N_14894,N_14757);
or UO_621 (O_621,N_14794,N_14752);
xor UO_622 (O_622,N_14958,N_14767);
and UO_623 (O_623,N_14872,N_14781);
or UO_624 (O_624,N_14973,N_14965);
nand UO_625 (O_625,N_14924,N_14921);
or UO_626 (O_626,N_14732,N_14901);
nor UO_627 (O_627,N_14987,N_14896);
or UO_628 (O_628,N_14853,N_14721);
and UO_629 (O_629,N_14850,N_14920);
xnor UO_630 (O_630,N_14977,N_14986);
nor UO_631 (O_631,N_14892,N_14870);
and UO_632 (O_632,N_14981,N_14769);
xor UO_633 (O_633,N_14885,N_14742);
xnor UO_634 (O_634,N_14931,N_14904);
or UO_635 (O_635,N_14713,N_14926);
or UO_636 (O_636,N_14720,N_14957);
or UO_637 (O_637,N_14940,N_14821);
nor UO_638 (O_638,N_14922,N_14975);
nand UO_639 (O_639,N_14982,N_14763);
nand UO_640 (O_640,N_14891,N_14965);
nor UO_641 (O_641,N_14970,N_14997);
nand UO_642 (O_642,N_14883,N_14823);
nand UO_643 (O_643,N_14813,N_14994);
xor UO_644 (O_644,N_14915,N_14876);
xor UO_645 (O_645,N_14763,N_14807);
and UO_646 (O_646,N_14814,N_14818);
or UO_647 (O_647,N_14879,N_14744);
xor UO_648 (O_648,N_14742,N_14938);
nor UO_649 (O_649,N_14859,N_14895);
nand UO_650 (O_650,N_14785,N_14953);
nand UO_651 (O_651,N_14919,N_14931);
nor UO_652 (O_652,N_14828,N_14918);
or UO_653 (O_653,N_14891,N_14795);
nor UO_654 (O_654,N_14898,N_14797);
nand UO_655 (O_655,N_14911,N_14822);
xor UO_656 (O_656,N_14970,N_14852);
nand UO_657 (O_657,N_14901,N_14840);
and UO_658 (O_658,N_14798,N_14752);
xor UO_659 (O_659,N_14736,N_14935);
xor UO_660 (O_660,N_14794,N_14793);
xnor UO_661 (O_661,N_14996,N_14733);
xor UO_662 (O_662,N_14984,N_14887);
nand UO_663 (O_663,N_14763,N_14746);
nor UO_664 (O_664,N_14980,N_14755);
or UO_665 (O_665,N_14878,N_14902);
xnor UO_666 (O_666,N_14837,N_14729);
nand UO_667 (O_667,N_14721,N_14941);
nor UO_668 (O_668,N_14735,N_14867);
or UO_669 (O_669,N_14720,N_14761);
xnor UO_670 (O_670,N_14799,N_14887);
xnor UO_671 (O_671,N_14987,N_14878);
xor UO_672 (O_672,N_14746,N_14938);
nand UO_673 (O_673,N_14954,N_14875);
or UO_674 (O_674,N_14967,N_14915);
xor UO_675 (O_675,N_14779,N_14742);
and UO_676 (O_676,N_14880,N_14712);
or UO_677 (O_677,N_14889,N_14806);
and UO_678 (O_678,N_14996,N_14726);
nor UO_679 (O_679,N_14810,N_14946);
nor UO_680 (O_680,N_14849,N_14805);
and UO_681 (O_681,N_14902,N_14992);
xor UO_682 (O_682,N_14793,N_14728);
nand UO_683 (O_683,N_14828,N_14824);
nand UO_684 (O_684,N_14729,N_14927);
or UO_685 (O_685,N_14743,N_14754);
nor UO_686 (O_686,N_14711,N_14960);
or UO_687 (O_687,N_14751,N_14858);
nand UO_688 (O_688,N_14805,N_14865);
and UO_689 (O_689,N_14749,N_14900);
nand UO_690 (O_690,N_14709,N_14738);
nor UO_691 (O_691,N_14788,N_14719);
and UO_692 (O_692,N_14742,N_14936);
xnor UO_693 (O_693,N_14989,N_14752);
or UO_694 (O_694,N_14991,N_14824);
nor UO_695 (O_695,N_14826,N_14776);
or UO_696 (O_696,N_14725,N_14937);
and UO_697 (O_697,N_14912,N_14991);
xnor UO_698 (O_698,N_14778,N_14776);
or UO_699 (O_699,N_14724,N_14865);
or UO_700 (O_700,N_14825,N_14975);
nand UO_701 (O_701,N_14886,N_14745);
xor UO_702 (O_702,N_14837,N_14861);
xnor UO_703 (O_703,N_14912,N_14700);
or UO_704 (O_704,N_14976,N_14949);
nand UO_705 (O_705,N_14954,N_14726);
or UO_706 (O_706,N_14952,N_14759);
nand UO_707 (O_707,N_14833,N_14723);
nand UO_708 (O_708,N_14849,N_14905);
and UO_709 (O_709,N_14749,N_14868);
or UO_710 (O_710,N_14807,N_14851);
nand UO_711 (O_711,N_14803,N_14964);
and UO_712 (O_712,N_14734,N_14964);
nor UO_713 (O_713,N_14877,N_14796);
xnor UO_714 (O_714,N_14757,N_14715);
nor UO_715 (O_715,N_14836,N_14764);
and UO_716 (O_716,N_14914,N_14779);
nand UO_717 (O_717,N_14731,N_14733);
and UO_718 (O_718,N_14937,N_14952);
nand UO_719 (O_719,N_14897,N_14902);
and UO_720 (O_720,N_14709,N_14978);
xnor UO_721 (O_721,N_14806,N_14878);
xnor UO_722 (O_722,N_14924,N_14784);
and UO_723 (O_723,N_14911,N_14725);
and UO_724 (O_724,N_14711,N_14745);
or UO_725 (O_725,N_14973,N_14768);
or UO_726 (O_726,N_14959,N_14874);
xnor UO_727 (O_727,N_14887,N_14896);
or UO_728 (O_728,N_14903,N_14770);
and UO_729 (O_729,N_14839,N_14739);
nor UO_730 (O_730,N_14765,N_14931);
xor UO_731 (O_731,N_14967,N_14885);
and UO_732 (O_732,N_14704,N_14929);
nand UO_733 (O_733,N_14790,N_14987);
and UO_734 (O_734,N_14868,N_14899);
nor UO_735 (O_735,N_14744,N_14916);
nor UO_736 (O_736,N_14700,N_14774);
or UO_737 (O_737,N_14967,N_14886);
xor UO_738 (O_738,N_14828,N_14739);
xor UO_739 (O_739,N_14835,N_14813);
nor UO_740 (O_740,N_14846,N_14886);
and UO_741 (O_741,N_14898,N_14976);
or UO_742 (O_742,N_14970,N_14700);
and UO_743 (O_743,N_14877,N_14972);
nor UO_744 (O_744,N_14989,N_14956);
or UO_745 (O_745,N_14993,N_14983);
nor UO_746 (O_746,N_14713,N_14882);
and UO_747 (O_747,N_14731,N_14863);
nand UO_748 (O_748,N_14906,N_14825);
nor UO_749 (O_749,N_14774,N_14767);
nand UO_750 (O_750,N_14805,N_14871);
nor UO_751 (O_751,N_14782,N_14987);
nand UO_752 (O_752,N_14978,N_14703);
xor UO_753 (O_753,N_14841,N_14843);
xor UO_754 (O_754,N_14712,N_14989);
nor UO_755 (O_755,N_14877,N_14815);
and UO_756 (O_756,N_14719,N_14959);
nor UO_757 (O_757,N_14929,N_14951);
and UO_758 (O_758,N_14800,N_14725);
and UO_759 (O_759,N_14936,N_14833);
nand UO_760 (O_760,N_14936,N_14968);
xor UO_761 (O_761,N_14790,N_14928);
nor UO_762 (O_762,N_14913,N_14825);
nand UO_763 (O_763,N_14890,N_14792);
nand UO_764 (O_764,N_14739,N_14999);
and UO_765 (O_765,N_14847,N_14811);
or UO_766 (O_766,N_14706,N_14972);
nor UO_767 (O_767,N_14870,N_14767);
or UO_768 (O_768,N_14980,N_14754);
nor UO_769 (O_769,N_14812,N_14870);
nor UO_770 (O_770,N_14828,N_14719);
nand UO_771 (O_771,N_14868,N_14720);
nand UO_772 (O_772,N_14832,N_14742);
nand UO_773 (O_773,N_14762,N_14765);
nor UO_774 (O_774,N_14826,N_14998);
or UO_775 (O_775,N_14881,N_14801);
nor UO_776 (O_776,N_14959,N_14763);
nor UO_777 (O_777,N_14840,N_14942);
xor UO_778 (O_778,N_14968,N_14876);
nor UO_779 (O_779,N_14878,N_14952);
nand UO_780 (O_780,N_14896,N_14746);
nand UO_781 (O_781,N_14886,N_14895);
nand UO_782 (O_782,N_14830,N_14792);
nand UO_783 (O_783,N_14913,N_14837);
nor UO_784 (O_784,N_14774,N_14819);
or UO_785 (O_785,N_14952,N_14816);
and UO_786 (O_786,N_14937,N_14886);
or UO_787 (O_787,N_14816,N_14905);
nand UO_788 (O_788,N_14970,N_14776);
nand UO_789 (O_789,N_14823,N_14829);
xor UO_790 (O_790,N_14801,N_14756);
nand UO_791 (O_791,N_14904,N_14923);
nor UO_792 (O_792,N_14702,N_14863);
nand UO_793 (O_793,N_14968,N_14872);
and UO_794 (O_794,N_14920,N_14743);
nor UO_795 (O_795,N_14774,N_14925);
nor UO_796 (O_796,N_14930,N_14969);
or UO_797 (O_797,N_14851,N_14940);
or UO_798 (O_798,N_14907,N_14753);
and UO_799 (O_799,N_14975,N_14981);
xor UO_800 (O_800,N_14779,N_14746);
xor UO_801 (O_801,N_14948,N_14865);
and UO_802 (O_802,N_14895,N_14728);
xnor UO_803 (O_803,N_14892,N_14850);
and UO_804 (O_804,N_14786,N_14898);
and UO_805 (O_805,N_14828,N_14882);
xnor UO_806 (O_806,N_14874,N_14816);
xor UO_807 (O_807,N_14962,N_14909);
nor UO_808 (O_808,N_14895,N_14783);
nor UO_809 (O_809,N_14925,N_14955);
or UO_810 (O_810,N_14854,N_14759);
and UO_811 (O_811,N_14935,N_14914);
nor UO_812 (O_812,N_14927,N_14921);
xnor UO_813 (O_813,N_14922,N_14847);
or UO_814 (O_814,N_14928,N_14890);
nor UO_815 (O_815,N_14889,N_14904);
nor UO_816 (O_816,N_14974,N_14996);
and UO_817 (O_817,N_14792,N_14718);
nor UO_818 (O_818,N_14749,N_14944);
nand UO_819 (O_819,N_14731,N_14745);
nand UO_820 (O_820,N_14857,N_14997);
or UO_821 (O_821,N_14884,N_14906);
xnor UO_822 (O_822,N_14837,N_14814);
xnor UO_823 (O_823,N_14825,N_14817);
and UO_824 (O_824,N_14909,N_14876);
nor UO_825 (O_825,N_14975,N_14978);
nand UO_826 (O_826,N_14935,N_14963);
or UO_827 (O_827,N_14783,N_14758);
nor UO_828 (O_828,N_14997,N_14941);
nand UO_829 (O_829,N_14980,N_14753);
nand UO_830 (O_830,N_14889,N_14742);
or UO_831 (O_831,N_14876,N_14814);
and UO_832 (O_832,N_14975,N_14745);
or UO_833 (O_833,N_14848,N_14720);
nor UO_834 (O_834,N_14995,N_14766);
or UO_835 (O_835,N_14792,N_14992);
nand UO_836 (O_836,N_14900,N_14737);
and UO_837 (O_837,N_14785,N_14956);
or UO_838 (O_838,N_14905,N_14883);
nor UO_839 (O_839,N_14929,N_14974);
xnor UO_840 (O_840,N_14796,N_14782);
nand UO_841 (O_841,N_14806,N_14728);
or UO_842 (O_842,N_14733,N_14995);
nor UO_843 (O_843,N_14816,N_14914);
nor UO_844 (O_844,N_14975,N_14989);
xor UO_845 (O_845,N_14918,N_14996);
or UO_846 (O_846,N_14910,N_14773);
nand UO_847 (O_847,N_14914,N_14889);
or UO_848 (O_848,N_14980,N_14978);
and UO_849 (O_849,N_14947,N_14957);
xor UO_850 (O_850,N_14982,N_14959);
nor UO_851 (O_851,N_14780,N_14809);
or UO_852 (O_852,N_14755,N_14791);
xnor UO_853 (O_853,N_14810,N_14886);
nor UO_854 (O_854,N_14855,N_14921);
nor UO_855 (O_855,N_14812,N_14824);
nor UO_856 (O_856,N_14738,N_14827);
or UO_857 (O_857,N_14873,N_14749);
xor UO_858 (O_858,N_14809,N_14760);
xor UO_859 (O_859,N_14912,N_14774);
nand UO_860 (O_860,N_14962,N_14893);
and UO_861 (O_861,N_14997,N_14823);
nand UO_862 (O_862,N_14809,N_14961);
and UO_863 (O_863,N_14791,N_14944);
xor UO_864 (O_864,N_14756,N_14864);
or UO_865 (O_865,N_14835,N_14967);
xnor UO_866 (O_866,N_14730,N_14969);
xor UO_867 (O_867,N_14778,N_14986);
nand UO_868 (O_868,N_14723,N_14913);
and UO_869 (O_869,N_14761,N_14804);
xor UO_870 (O_870,N_14909,N_14866);
or UO_871 (O_871,N_14768,N_14959);
and UO_872 (O_872,N_14704,N_14848);
nor UO_873 (O_873,N_14882,N_14864);
xor UO_874 (O_874,N_14769,N_14754);
and UO_875 (O_875,N_14792,N_14804);
or UO_876 (O_876,N_14873,N_14743);
xnor UO_877 (O_877,N_14961,N_14965);
or UO_878 (O_878,N_14835,N_14755);
xor UO_879 (O_879,N_14783,N_14813);
nor UO_880 (O_880,N_14874,N_14947);
and UO_881 (O_881,N_14988,N_14788);
nor UO_882 (O_882,N_14918,N_14980);
and UO_883 (O_883,N_14803,N_14856);
xor UO_884 (O_884,N_14763,N_14724);
nand UO_885 (O_885,N_14834,N_14883);
xor UO_886 (O_886,N_14857,N_14798);
nor UO_887 (O_887,N_14848,N_14877);
and UO_888 (O_888,N_14910,N_14987);
and UO_889 (O_889,N_14893,N_14944);
or UO_890 (O_890,N_14757,N_14991);
and UO_891 (O_891,N_14714,N_14871);
nand UO_892 (O_892,N_14708,N_14969);
nand UO_893 (O_893,N_14890,N_14712);
or UO_894 (O_894,N_14839,N_14873);
nand UO_895 (O_895,N_14774,N_14803);
nand UO_896 (O_896,N_14739,N_14886);
or UO_897 (O_897,N_14725,N_14735);
nand UO_898 (O_898,N_14805,N_14939);
nand UO_899 (O_899,N_14894,N_14854);
or UO_900 (O_900,N_14850,N_14970);
and UO_901 (O_901,N_14731,N_14868);
nor UO_902 (O_902,N_14854,N_14992);
nand UO_903 (O_903,N_14736,N_14765);
or UO_904 (O_904,N_14943,N_14819);
nand UO_905 (O_905,N_14943,N_14839);
or UO_906 (O_906,N_14720,N_14798);
xnor UO_907 (O_907,N_14958,N_14765);
nand UO_908 (O_908,N_14973,N_14811);
and UO_909 (O_909,N_14738,N_14848);
or UO_910 (O_910,N_14807,N_14866);
nor UO_911 (O_911,N_14882,N_14799);
nand UO_912 (O_912,N_14701,N_14855);
nand UO_913 (O_913,N_14947,N_14721);
nand UO_914 (O_914,N_14916,N_14875);
nor UO_915 (O_915,N_14943,N_14962);
or UO_916 (O_916,N_14724,N_14929);
xor UO_917 (O_917,N_14861,N_14833);
nand UO_918 (O_918,N_14857,N_14832);
xor UO_919 (O_919,N_14981,N_14962);
or UO_920 (O_920,N_14868,N_14976);
xnor UO_921 (O_921,N_14908,N_14889);
and UO_922 (O_922,N_14960,N_14740);
and UO_923 (O_923,N_14797,N_14801);
or UO_924 (O_924,N_14804,N_14822);
nand UO_925 (O_925,N_14714,N_14934);
nor UO_926 (O_926,N_14721,N_14821);
and UO_927 (O_927,N_14761,N_14998);
and UO_928 (O_928,N_14715,N_14718);
xor UO_929 (O_929,N_14937,N_14846);
nor UO_930 (O_930,N_14797,N_14913);
nor UO_931 (O_931,N_14763,N_14922);
nor UO_932 (O_932,N_14730,N_14832);
nand UO_933 (O_933,N_14767,N_14925);
nor UO_934 (O_934,N_14968,N_14700);
nor UO_935 (O_935,N_14988,N_14886);
nor UO_936 (O_936,N_14748,N_14844);
or UO_937 (O_937,N_14746,N_14800);
xnor UO_938 (O_938,N_14955,N_14780);
nor UO_939 (O_939,N_14784,N_14873);
or UO_940 (O_940,N_14901,N_14957);
xnor UO_941 (O_941,N_14838,N_14732);
nor UO_942 (O_942,N_14999,N_14855);
and UO_943 (O_943,N_14787,N_14803);
or UO_944 (O_944,N_14837,N_14717);
and UO_945 (O_945,N_14881,N_14742);
nor UO_946 (O_946,N_14743,N_14986);
nand UO_947 (O_947,N_14738,N_14785);
or UO_948 (O_948,N_14814,N_14862);
nor UO_949 (O_949,N_14981,N_14893);
and UO_950 (O_950,N_14751,N_14760);
nor UO_951 (O_951,N_14830,N_14717);
xnor UO_952 (O_952,N_14859,N_14843);
and UO_953 (O_953,N_14814,N_14774);
and UO_954 (O_954,N_14937,N_14842);
xnor UO_955 (O_955,N_14867,N_14739);
nor UO_956 (O_956,N_14799,N_14725);
or UO_957 (O_957,N_14758,N_14793);
nor UO_958 (O_958,N_14991,N_14702);
xnor UO_959 (O_959,N_14821,N_14854);
nor UO_960 (O_960,N_14776,N_14809);
nand UO_961 (O_961,N_14778,N_14741);
and UO_962 (O_962,N_14877,N_14724);
nand UO_963 (O_963,N_14885,N_14729);
nand UO_964 (O_964,N_14987,N_14789);
xor UO_965 (O_965,N_14704,N_14706);
or UO_966 (O_966,N_14978,N_14758);
nor UO_967 (O_967,N_14899,N_14790);
nand UO_968 (O_968,N_14809,N_14764);
nand UO_969 (O_969,N_14758,N_14770);
nand UO_970 (O_970,N_14877,N_14816);
nand UO_971 (O_971,N_14738,N_14981);
nand UO_972 (O_972,N_14846,N_14885);
nor UO_973 (O_973,N_14720,N_14875);
nor UO_974 (O_974,N_14934,N_14815);
nand UO_975 (O_975,N_14711,N_14713);
and UO_976 (O_976,N_14765,N_14861);
and UO_977 (O_977,N_14826,N_14997);
xor UO_978 (O_978,N_14897,N_14709);
xnor UO_979 (O_979,N_14912,N_14726);
xor UO_980 (O_980,N_14711,N_14720);
nor UO_981 (O_981,N_14935,N_14843);
and UO_982 (O_982,N_14777,N_14813);
nor UO_983 (O_983,N_14875,N_14759);
xor UO_984 (O_984,N_14704,N_14930);
and UO_985 (O_985,N_14731,N_14836);
xor UO_986 (O_986,N_14922,N_14751);
or UO_987 (O_987,N_14871,N_14816);
xor UO_988 (O_988,N_14706,N_14745);
nor UO_989 (O_989,N_14966,N_14897);
or UO_990 (O_990,N_14924,N_14832);
and UO_991 (O_991,N_14724,N_14909);
nand UO_992 (O_992,N_14705,N_14930);
or UO_993 (O_993,N_14761,N_14896);
or UO_994 (O_994,N_14992,N_14908);
xor UO_995 (O_995,N_14826,N_14788);
or UO_996 (O_996,N_14753,N_14725);
and UO_997 (O_997,N_14927,N_14802);
nand UO_998 (O_998,N_14743,N_14939);
xor UO_999 (O_999,N_14732,N_14987);
or UO_1000 (O_1000,N_14820,N_14857);
and UO_1001 (O_1001,N_14983,N_14731);
or UO_1002 (O_1002,N_14935,N_14762);
or UO_1003 (O_1003,N_14715,N_14953);
and UO_1004 (O_1004,N_14915,N_14842);
or UO_1005 (O_1005,N_14878,N_14897);
and UO_1006 (O_1006,N_14770,N_14809);
xnor UO_1007 (O_1007,N_14915,N_14917);
nand UO_1008 (O_1008,N_14719,N_14887);
or UO_1009 (O_1009,N_14867,N_14839);
and UO_1010 (O_1010,N_14957,N_14961);
nand UO_1011 (O_1011,N_14824,N_14949);
or UO_1012 (O_1012,N_14715,N_14809);
nand UO_1013 (O_1013,N_14756,N_14953);
or UO_1014 (O_1014,N_14970,N_14737);
and UO_1015 (O_1015,N_14860,N_14832);
nand UO_1016 (O_1016,N_14711,N_14783);
or UO_1017 (O_1017,N_14972,N_14763);
and UO_1018 (O_1018,N_14941,N_14989);
nand UO_1019 (O_1019,N_14933,N_14893);
xor UO_1020 (O_1020,N_14868,N_14737);
and UO_1021 (O_1021,N_14757,N_14857);
nor UO_1022 (O_1022,N_14970,N_14929);
nand UO_1023 (O_1023,N_14946,N_14800);
nor UO_1024 (O_1024,N_14779,N_14859);
and UO_1025 (O_1025,N_14795,N_14794);
and UO_1026 (O_1026,N_14893,N_14880);
or UO_1027 (O_1027,N_14844,N_14737);
xnor UO_1028 (O_1028,N_14728,N_14959);
xnor UO_1029 (O_1029,N_14907,N_14961);
and UO_1030 (O_1030,N_14834,N_14953);
xnor UO_1031 (O_1031,N_14710,N_14702);
or UO_1032 (O_1032,N_14746,N_14889);
xnor UO_1033 (O_1033,N_14880,N_14709);
and UO_1034 (O_1034,N_14824,N_14958);
nor UO_1035 (O_1035,N_14825,N_14999);
or UO_1036 (O_1036,N_14863,N_14959);
or UO_1037 (O_1037,N_14735,N_14732);
nand UO_1038 (O_1038,N_14994,N_14996);
and UO_1039 (O_1039,N_14859,N_14900);
xor UO_1040 (O_1040,N_14866,N_14892);
xor UO_1041 (O_1041,N_14729,N_14763);
nand UO_1042 (O_1042,N_14840,N_14872);
nand UO_1043 (O_1043,N_14915,N_14962);
xnor UO_1044 (O_1044,N_14859,N_14850);
and UO_1045 (O_1045,N_14785,N_14939);
and UO_1046 (O_1046,N_14830,N_14782);
or UO_1047 (O_1047,N_14792,N_14864);
and UO_1048 (O_1048,N_14951,N_14963);
or UO_1049 (O_1049,N_14908,N_14944);
or UO_1050 (O_1050,N_14964,N_14831);
nor UO_1051 (O_1051,N_14908,N_14793);
nand UO_1052 (O_1052,N_14755,N_14761);
or UO_1053 (O_1053,N_14868,N_14996);
or UO_1054 (O_1054,N_14747,N_14773);
nand UO_1055 (O_1055,N_14934,N_14794);
and UO_1056 (O_1056,N_14781,N_14891);
xnor UO_1057 (O_1057,N_14894,N_14886);
xor UO_1058 (O_1058,N_14898,N_14757);
nor UO_1059 (O_1059,N_14793,N_14832);
xor UO_1060 (O_1060,N_14750,N_14964);
nor UO_1061 (O_1061,N_14896,N_14819);
or UO_1062 (O_1062,N_14867,N_14806);
or UO_1063 (O_1063,N_14923,N_14924);
xnor UO_1064 (O_1064,N_14872,N_14748);
or UO_1065 (O_1065,N_14731,N_14991);
nand UO_1066 (O_1066,N_14793,N_14883);
xor UO_1067 (O_1067,N_14765,N_14869);
nand UO_1068 (O_1068,N_14868,N_14732);
xor UO_1069 (O_1069,N_14801,N_14796);
nand UO_1070 (O_1070,N_14739,N_14711);
or UO_1071 (O_1071,N_14986,N_14796);
or UO_1072 (O_1072,N_14896,N_14886);
and UO_1073 (O_1073,N_14868,N_14723);
xnor UO_1074 (O_1074,N_14772,N_14975);
or UO_1075 (O_1075,N_14819,N_14919);
and UO_1076 (O_1076,N_14784,N_14958);
nand UO_1077 (O_1077,N_14719,N_14911);
nand UO_1078 (O_1078,N_14742,N_14708);
and UO_1079 (O_1079,N_14860,N_14726);
or UO_1080 (O_1080,N_14924,N_14778);
or UO_1081 (O_1081,N_14877,N_14719);
and UO_1082 (O_1082,N_14855,N_14723);
xnor UO_1083 (O_1083,N_14778,N_14810);
and UO_1084 (O_1084,N_14886,N_14878);
xor UO_1085 (O_1085,N_14955,N_14858);
nand UO_1086 (O_1086,N_14950,N_14752);
xnor UO_1087 (O_1087,N_14818,N_14936);
nor UO_1088 (O_1088,N_14806,N_14904);
xor UO_1089 (O_1089,N_14711,N_14999);
xnor UO_1090 (O_1090,N_14904,N_14728);
nand UO_1091 (O_1091,N_14747,N_14946);
xor UO_1092 (O_1092,N_14870,N_14772);
nand UO_1093 (O_1093,N_14905,N_14784);
or UO_1094 (O_1094,N_14917,N_14780);
and UO_1095 (O_1095,N_14944,N_14757);
nand UO_1096 (O_1096,N_14746,N_14886);
nand UO_1097 (O_1097,N_14900,N_14731);
and UO_1098 (O_1098,N_14830,N_14774);
xnor UO_1099 (O_1099,N_14979,N_14842);
or UO_1100 (O_1100,N_14789,N_14795);
nand UO_1101 (O_1101,N_14919,N_14796);
or UO_1102 (O_1102,N_14838,N_14905);
or UO_1103 (O_1103,N_14743,N_14878);
nand UO_1104 (O_1104,N_14909,N_14732);
nor UO_1105 (O_1105,N_14823,N_14977);
nor UO_1106 (O_1106,N_14716,N_14846);
xnor UO_1107 (O_1107,N_14836,N_14700);
nand UO_1108 (O_1108,N_14796,N_14881);
xor UO_1109 (O_1109,N_14740,N_14724);
or UO_1110 (O_1110,N_14748,N_14913);
nand UO_1111 (O_1111,N_14873,N_14872);
or UO_1112 (O_1112,N_14819,N_14720);
and UO_1113 (O_1113,N_14714,N_14814);
nand UO_1114 (O_1114,N_14925,N_14788);
or UO_1115 (O_1115,N_14758,N_14979);
nor UO_1116 (O_1116,N_14743,N_14981);
or UO_1117 (O_1117,N_14869,N_14903);
nor UO_1118 (O_1118,N_14835,N_14719);
nand UO_1119 (O_1119,N_14982,N_14729);
and UO_1120 (O_1120,N_14773,N_14800);
or UO_1121 (O_1121,N_14900,N_14729);
or UO_1122 (O_1122,N_14727,N_14757);
nor UO_1123 (O_1123,N_14907,N_14795);
xor UO_1124 (O_1124,N_14842,N_14901);
and UO_1125 (O_1125,N_14877,N_14707);
nor UO_1126 (O_1126,N_14872,N_14858);
nor UO_1127 (O_1127,N_14980,N_14784);
nand UO_1128 (O_1128,N_14776,N_14768);
nor UO_1129 (O_1129,N_14934,N_14881);
and UO_1130 (O_1130,N_14761,N_14729);
nor UO_1131 (O_1131,N_14971,N_14826);
xnor UO_1132 (O_1132,N_14713,N_14990);
nand UO_1133 (O_1133,N_14975,N_14783);
xnor UO_1134 (O_1134,N_14984,N_14810);
and UO_1135 (O_1135,N_14759,N_14785);
xor UO_1136 (O_1136,N_14974,N_14810);
xor UO_1137 (O_1137,N_14811,N_14835);
xnor UO_1138 (O_1138,N_14702,N_14904);
xnor UO_1139 (O_1139,N_14811,N_14771);
and UO_1140 (O_1140,N_14736,N_14944);
nor UO_1141 (O_1141,N_14884,N_14950);
nand UO_1142 (O_1142,N_14763,N_14751);
and UO_1143 (O_1143,N_14927,N_14708);
or UO_1144 (O_1144,N_14952,N_14736);
nand UO_1145 (O_1145,N_14717,N_14734);
xor UO_1146 (O_1146,N_14816,N_14862);
or UO_1147 (O_1147,N_14740,N_14702);
xnor UO_1148 (O_1148,N_14790,N_14847);
nand UO_1149 (O_1149,N_14718,N_14967);
and UO_1150 (O_1150,N_14858,N_14945);
nor UO_1151 (O_1151,N_14970,N_14751);
xor UO_1152 (O_1152,N_14935,N_14796);
xor UO_1153 (O_1153,N_14853,N_14946);
or UO_1154 (O_1154,N_14858,N_14995);
xor UO_1155 (O_1155,N_14872,N_14827);
nand UO_1156 (O_1156,N_14765,N_14945);
and UO_1157 (O_1157,N_14703,N_14866);
or UO_1158 (O_1158,N_14763,N_14991);
nor UO_1159 (O_1159,N_14978,N_14929);
nor UO_1160 (O_1160,N_14990,N_14797);
xnor UO_1161 (O_1161,N_14984,N_14874);
and UO_1162 (O_1162,N_14759,N_14702);
and UO_1163 (O_1163,N_14915,N_14903);
nand UO_1164 (O_1164,N_14835,N_14880);
xnor UO_1165 (O_1165,N_14947,N_14966);
nor UO_1166 (O_1166,N_14884,N_14740);
or UO_1167 (O_1167,N_14784,N_14725);
nor UO_1168 (O_1168,N_14988,N_14843);
or UO_1169 (O_1169,N_14703,N_14782);
or UO_1170 (O_1170,N_14747,N_14934);
nor UO_1171 (O_1171,N_14819,N_14925);
or UO_1172 (O_1172,N_14806,N_14871);
nor UO_1173 (O_1173,N_14787,N_14713);
xor UO_1174 (O_1174,N_14844,N_14907);
nand UO_1175 (O_1175,N_14947,N_14863);
nor UO_1176 (O_1176,N_14716,N_14715);
or UO_1177 (O_1177,N_14884,N_14747);
nand UO_1178 (O_1178,N_14940,N_14734);
nor UO_1179 (O_1179,N_14850,N_14855);
or UO_1180 (O_1180,N_14955,N_14848);
or UO_1181 (O_1181,N_14916,N_14864);
or UO_1182 (O_1182,N_14931,N_14814);
or UO_1183 (O_1183,N_14995,N_14918);
nand UO_1184 (O_1184,N_14952,N_14895);
xnor UO_1185 (O_1185,N_14777,N_14760);
nand UO_1186 (O_1186,N_14983,N_14736);
xor UO_1187 (O_1187,N_14785,N_14706);
nand UO_1188 (O_1188,N_14780,N_14763);
and UO_1189 (O_1189,N_14757,N_14812);
nor UO_1190 (O_1190,N_14968,N_14841);
or UO_1191 (O_1191,N_14737,N_14946);
nand UO_1192 (O_1192,N_14961,N_14782);
nor UO_1193 (O_1193,N_14965,N_14904);
and UO_1194 (O_1194,N_14983,N_14838);
xor UO_1195 (O_1195,N_14889,N_14935);
or UO_1196 (O_1196,N_14911,N_14761);
nor UO_1197 (O_1197,N_14782,N_14805);
or UO_1198 (O_1198,N_14708,N_14772);
nand UO_1199 (O_1199,N_14780,N_14807);
and UO_1200 (O_1200,N_14862,N_14797);
nand UO_1201 (O_1201,N_14917,N_14881);
or UO_1202 (O_1202,N_14872,N_14972);
xor UO_1203 (O_1203,N_14723,N_14842);
or UO_1204 (O_1204,N_14995,N_14978);
nand UO_1205 (O_1205,N_14960,N_14787);
nor UO_1206 (O_1206,N_14723,N_14705);
and UO_1207 (O_1207,N_14812,N_14785);
xor UO_1208 (O_1208,N_14946,N_14745);
nor UO_1209 (O_1209,N_14881,N_14765);
xnor UO_1210 (O_1210,N_14756,N_14796);
nand UO_1211 (O_1211,N_14832,N_14870);
or UO_1212 (O_1212,N_14810,N_14852);
xor UO_1213 (O_1213,N_14714,N_14728);
xnor UO_1214 (O_1214,N_14855,N_14859);
xor UO_1215 (O_1215,N_14921,N_14737);
nor UO_1216 (O_1216,N_14814,N_14941);
or UO_1217 (O_1217,N_14904,N_14807);
nor UO_1218 (O_1218,N_14878,N_14990);
or UO_1219 (O_1219,N_14918,N_14795);
xnor UO_1220 (O_1220,N_14757,N_14842);
or UO_1221 (O_1221,N_14925,N_14892);
xor UO_1222 (O_1222,N_14952,N_14876);
nand UO_1223 (O_1223,N_14774,N_14738);
nand UO_1224 (O_1224,N_14705,N_14811);
nand UO_1225 (O_1225,N_14861,N_14936);
and UO_1226 (O_1226,N_14709,N_14741);
nand UO_1227 (O_1227,N_14767,N_14860);
and UO_1228 (O_1228,N_14964,N_14979);
and UO_1229 (O_1229,N_14989,N_14940);
and UO_1230 (O_1230,N_14742,N_14818);
or UO_1231 (O_1231,N_14985,N_14941);
or UO_1232 (O_1232,N_14803,N_14846);
xor UO_1233 (O_1233,N_14938,N_14710);
nor UO_1234 (O_1234,N_14875,N_14870);
nor UO_1235 (O_1235,N_14970,N_14769);
or UO_1236 (O_1236,N_14966,N_14962);
or UO_1237 (O_1237,N_14940,N_14748);
and UO_1238 (O_1238,N_14771,N_14852);
nand UO_1239 (O_1239,N_14841,N_14784);
and UO_1240 (O_1240,N_14987,N_14868);
or UO_1241 (O_1241,N_14733,N_14925);
nand UO_1242 (O_1242,N_14828,N_14974);
or UO_1243 (O_1243,N_14845,N_14813);
nand UO_1244 (O_1244,N_14760,N_14705);
and UO_1245 (O_1245,N_14846,N_14769);
xnor UO_1246 (O_1246,N_14813,N_14787);
xor UO_1247 (O_1247,N_14796,N_14711);
nand UO_1248 (O_1248,N_14816,N_14954);
xor UO_1249 (O_1249,N_14795,N_14915);
nor UO_1250 (O_1250,N_14795,N_14822);
xnor UO_1251 (O_1251,N_14929,N_14998);
xor UO_1252 (O_1252,N_14974,N_14954);
or UO_1253 (O_1253,N_14960,N_14733);
nand UO_1254 (O_1254,N_14990,N_14824);
nand UO_1255 (O_1255,N_14711,N_14992);
or UO_1256 (O_1256,N_14840,N_14959);
nor UO_1257 (O_1257,N_14986,N_14957);
xnor UO_1258 (O_1258,N_14779,N_14784);
nand UO_1259 (O_1259,N_14896,N_14967);
nor UO_1260 (O_1260,N_14894,N_14733);
and UO_1261 (O_1261,N_14938,N_14994);
or UO_1262 (O_1262,N_14881,N_14806);
or UO_1263 (O_1263,N_14795,N_14819);
nor UO_1264 (O_1264,N_14903,N_14859);
xnor UO_1265 (O_1265,N_14760,N_14784);
nor UO_1266 (O_1266,N_14850,N_14811);
and UO_1267 (O_1267,N_14790,N_14781);
nand UO_1268 (O_1268,N_14734,N_14750);
nand UO_1269 (O_1269,N_14757,N_14878);
or UO_1270 (O_1270,N_14775,N_14888);
nor UO_1271 (O_1271,N_14977,N_14771);
xor UO_1272 (O_1272,N_14985,N_14919);
or UO_1273 (O_1273,N_14879,N_14712);
xor UO_1274 (O_1274,N_14913,N_14842);
nor UO_1275 (O_1275,N_14966,N_14777);
xor UO_1276 (O_1276,N_14725,N_14789);
nand UO_1277 (O_1277,N_14730,N_14779);
nor UO_1278 (O_1278,N_14872,N_14947);
and UO_1279 (O_1279,N_14995,N_14823);
nor UO_1280 (O_1280,N_14725,N_14704);
or UO_1281 (O_1281,N_14862,N_14856);
nor UO_1282 (O_1282,N_14787,N_14725);
xnor UO_1283 (O_1283,N_14777,N_14790);
and UO_1284 (O_1284,N_14857,N_14985);
nand UO_1285 (O_1285,N_14787,N_14953);
and UO_1286 (O_1286,N_14719,N_14793);
and UO_1287 (O_1287,N_14876,N_14963);
and UO_1288 (O_1288,N_14758,N_14984);
xor UO_1289 (O_1289,N_14905,N_14828);
or UO_1290 (O_1290,N_14720,N_14889);
nand UO_1291 (O_1291,N_14752,N_14708);
or UO_1292 (O_1292,N_14945,N_14711);
xor UO_1293 (O_1293,N_14817,N_14809);
or UO_1294 (O_1294,N_14874,N_14732);
and UO_1295 (O_1295,N_14895,N_14949);
or UO_1296 (O_1296,N_14887,N_14762);
and UO_1297 (O_1297,N_14778,N_14708);
nor UO_1298 (O_1298,N_14797,N_14832);
or UO_1299 (O_1299,N_14727,N_14839);
or UO_1300 (O_1300,N_14875,N_14950);
xnor UO_1301 (O_1301,N_14900,N_14708);
and UO_1302 (O_1302,N_14713,N_14927);
and UO_1303 (O_1303,N_14795,N_14817);
xor UO_1304 (O_1304,N_14965,N_14953);
nand UO_1305 (O_1305,N_14925,N_14714);
nor UO_1306 (O_1306,N_14906,N_14702);
xor UO_1307 (O_1307,N_14893,N_14748);
and UO_1308 (O_1308,N_14815,N_14914);
xnor UO_1309 (O_1309,N_14716,N_14810);
and UO_1310 (O_1310,N_14975,N_14728);
and UO_1311 (O_1311,N_14936,N_14810);
and UO_1312 (O_1312,N_14928,N_14745);
and UO_1313 (O_1313,N_14932,N_14997);
nand UO_1314 (O_1314,N_14826,N_14878);
or UO_1315 (O_1315,N_14859,N_14722);
or UO_1316 (O_1316,N_14845,N_14835);
nor UO_1317 (O_1317,N_14719,N_14962);
nand UO_1318 (O_1318,N_14725,N_14968);
or UO_1319 (O_1319,N_14845,N_14779);
nand UO_1320 (O_1320,N_14977,N_14865);
and UO_1321 (O_1321,N_14906,N_14847);
nor UO_1322 (O_1322,N_14914,N_14875);
and UO_1323 (O_1323,N_14990,N_14810);
nand UO_1324 (O_1324,N_14918,N_14714);
nand UO_1325 (O_1325,N_14707,N_14809);
or UO_1326 (O_1326,N_14783,N_14735);
or UO_1327 (O_1327,N_14794,N_14858);
or UO_1328 (O_1328,N_14834,N_14708);
and UO_1329 (O_1329,N_14993,N_14835);
and UO_1330 (O_1330,N_14847,N_14981);
nor UO_1331 (O_1331,N_14759,N_14886);
or UO_1332 (O_1332,N_14945,N_14714);
nor UO_1333 (O_1333,N_14706,N_14967);
nor UO_1334 (O_1334,N_14807,N_14942);
or UO_1335 (O_1335,N_14771,N_14850);
and UO_1336 (O_1336,N_14920,N_14915);
and UO_1337 (O_1337,N_14786,N_14862);
nand UO_1338 (O_1338,N_14885,N_14817);
nand UO_1339 (O_1339,N_14761,N_14847);
and UO_1340 (O_1340,N_14723,N_14909);
and UO_1341 (O_1341,N_14964,N_14860);
nand UO_1342 (O_1342,N_14772,N_14738);
nor UO_1343 (O_1343,N_14926,N_14755);
xor UO_1344 (O_1344,N_14769,N_14772);
nor UO_1345 (O_1345,N_14806,N_14834);
or UO_1346 (O_1346,N_14894,N_14900);
nand UO_1347 (O_1347,N_14967,N_14969);
nor UO_1348 (O_1348,N_14720,N_14881);
and UO_1349 (O_1349,N_14857,N_14920);
or UO_1350 (O_1350,N_14838,N_14950);
or UO_1351 (O_1351,N_14887,N_14750);
or UO_1352 (O_1352,N_14906,N_14801);
xnor UO_1353 (O_1353,N_14724,N_14893);
nor UO_1354 (O_1354,N_14806,N_14747);
nor UO_1355 (O_1355,N_14995,N_14961);
nor UO_1356 (O_1356,N_14838,N_14790);
nand UO_1357 (O_1357,N_14971,N_14783);
xor UO_1358 (O_1358,N_14736,N_14803);
nor UO_1359 (O_1359,N_14997,N_14812);
nand UO_1360 (O_1360,N_14937,N_14922);
xnor UO_1361 (O_1361,N_14856,N_14936);
and UO_1362 (O_1362,N_14777,N_14820);
and UO_1363 (O_1363,N_14708,N_14754);
nand UO_1364 (O_1364,N_14882,N_14792);
and UO_1365 (O_1365,N_14805,N_14972);
nor UO_1366 (O_1366,N_14858,N_14969);
and UO_1367 (O_1367,N_14726,N_14856);
xor UO_1368 (O_1368,N_14770,N_14830);
or UO_1369 (O_1369,N_14979,N_14900);
nand UO_1370 (O_1370,N_14886,N_14938);
and UO_1371 (O_1371,N_14807,N_14951);
nand UO_1372 (O_1372,N_14810,N_14831);
or UO_1373 (O_1373,N_14955,N_14830);
and UO_1374 (O_1374,N_14813,N_14988);
xnor UO_1375 (O_1375,N_14803,N_14784);
or UO_1376 (O_1376,N_14728,N_14939);
xor UO_1377 (O_1377,N_14923,N_14702);
or UO_1378 (O_1378,N_14801,N_14892);
xor UO_1379 (O_1379,N_14753,N_14755);
nor UO_1380 (O_1380,N_14819,N_14763);
xnor UO_1381 (O_1381,N_14739,N_14718);
nand UO_1382 (O_1382,N_14838,N_14845);
or UO_1383 (O_1383,N_14876,N_14851);
or UO_1384 (O_1384,N_14754,N_14751);
nand UO_1385 (O_1385,N_14739,N_14750);
and UO_1386 (O_1386,N_14726,N_14733);
or UO_1387 (O_1387,N_14913,N_14943);
and UO_1388 (O_1388,N_14922,N_14759);
nand UO_1389 (O_1389,N_14917,N_14845);
nand UO_1390 (O_1390,N_14939,N_14765);
nand UO_1391 (O_1391,N_14902,N_14812);
nor UO_1392 (O_1392,N_14894,N_14917);
and UO_1393 (O_1393,N_14830,N_14914);
nand UO_1394 (O_1394,N_14705,N_14707);
nand UO_1395 (O_1395,N_14773,N_14856);
xor UO_1396 (O_1396,N_14839,N_14729);
or UO_1397 (O_1397,N_14883,N_14794);
and UO_1398 (O_1398,N_14923,N_14758);
or UO_1399 (O_1399,N_14795,N_14791);
and UO_1400 (O_1400,N_14786,N_14767);
or UO_1401 (O_1401,N_14823,N_14731);
or UO_1402 (O_1402,N_14886,N_14740);
or UO_1403 (O_1403,N_14931,N_14831);
or UO_1404 (O_1404,N_14843,N_14984);
nor UO_1405 (O_1405,N_14884,N_14840);
nor UO_1406 (O_1406,N_14741,N_14906);
xor UO_1407 (O_1407,N_14973,N_14742);
nand UO_1408 (O_1408,N_14753,N_14844);
xor UO_1409 (O_1409,N_14829,N_14735);
xor UO_1410 (O_1410,N_14779,N_14823);
and UO_1411 (O_1411,N_14731,N_14760);
xor UO_1412 (O_1412,N_14708,N_14753);
nor UO_1413 (O_1413,N_14979,N_14711);
or UO_1414 (O_1414,N_14884,N_14830);
nor UO_1415 (O_1415,N_14995,N_14752);
or UO_1416 (O_1416,N_14777,N_14801);
nand UO_1417 (O_1417,N_14926,N_14730);
and UO_1418 (O_1418,N_14962,N_14747);
nor UO_1419 (O_1419,N_14870,N_14921);
nand UO_1420 (O_1420,N_14721,N_14793);
and UO_1421 (O_1421,N_14715,N_14891);
xnor UO_1422 (O_1422,N_14913,N_14897);
and UO_1423 (O_1423,N_14978,N_14917);
nor UO_1424 (O_1424,N_14767,N_14868);
xnor UO_1425 (O_1425,N_14828,N_14857);
xnor UO_1426 (O_1426,N_14877,N_14957);
xnor UO_1427 (O_1427,N_14974,N_14970);
nand UO_1428 (O_1428,N_14919,N_14913);
xor UO_1429 (O_1429,N_14843,N_14766);
and UO_1430 (O_1430,N_14706,N_14878);
nand UO_1431 (O_1431,N_14721,N_14799);
xnor UO_1432 (O_1432,N_14874,N_14908);
or UO_1433 (O_1433,N_14738,N_14870);
nand UO_1434 (O_1434,N_14736,N_14706);
or UO_1435 (O_1435,N_14769,N_14850);
nand UO_1436 (O_1436,N_14741,N_14835);
xor UO_1437 (O_1437,N_14985,N_14957);
and UO_1438 (O_1438,N_14756,N_14926);
nand UO_1439 (O_1439,N_14952,N_14927);
nand UO_1440 (O_1440,N_14853,N_14809);
nand UO_1441 (O_1441,N_14840,N_14709);
and UO_1442 (O_1442,N_14772,N_14729);
or UO_1443 (O_1443,N_14980,N_14819);
or UO_1444 (O_1444,N_14990,N_14988);
nand UO_1445 (O_1445,N_14794,N_14984);
xnor UO_1446 (O_1446,N_14900,N_14877);
xor UO_1447 (O_1447,N_14782,N_14750);
or UO_1448 (O_1448,N_14773,N_14957);
and UO_1449 (O_1449,N_14711,N_14927);
nor UO_1450 (O_1450,N_14751,N_14702);
or UO_1451 (O_1451,N_14970,N_14785);
nand UO_1452 (O_1452,N_14764,N_14762);
or UO_1453 (O_1453,N_14923,N_14795);
or UO_1454 (O_1454,N_14969,N_14786);
or UO_1455 (O_1455,N_14846,N_14983);
or UO_1456 (O_1456,N_14975,N_14763);
xnor UO_1457 (O_1457,N_14878,N_14983);
nor UO_1458 (O_1458,N_14826,N_14901);
nand UO_1459 (O_1459,N_14810,N_14732);
or UO_1460 (O_1460,N_14763,N_14985);
nand UO_1461 (O_1461,N_14784,N_14878);
or UO_1462 (O_1462,N_14976,N_14909);
and UO_1463 (O_1463,N_14715,N_14820);
nor UO_1464 (O_1464,N_14979,N_14902);
and UO_1465 (O_1465,N_14765,N_14897);
and UO_1466 (O_1466,N_14743,N_14883);
or UO_1467 (O_1467,N_14968,N_14810);
xor UO_1468 (O_1468,N_14778,N_14887);
nor UO_1469 (O_1469,N_14807,N_14857);
xor UO_1470 (O_1470,N_14866,N_14946);
or UO_1471 (O_1471,N_14827,N_14988);
nand UO_1472 (O_1472,N_14970,N_14915);
xor UO_1473 (O_1473,N_14816,N_14719);
and UO_1474 (O_1474,N_14983,N_14923);
xor UO_1475 (O_1475,N_14825,N_14848);
xor UO_1476 (O_1476,N_14985,N_14800);
and UO_1477 (O_1477,N_14706,N_14817);
and UO_1478 (O_1478,N_14771,N_14754);
or UO_1479 (O_1479,N_14841,N_14824);
nor UO_1480 (O_1480,N_14724,N_14964);
or UO_1481 (O_1481,N_14758,N_14958);
or UO_1482 (O_1482,N_14757,N_14769);
xor UO_1483 (O_1483,N_14949,N_14984);
xor UO_1484 (O_1484,N_14953,N_14860);
xnor UO_1485 (O_1485,N_14897,N_14716);
xor UO_1486 (O_1486,N_14946,N_14740);
xor UO_1487 (O_1487,N_14954,N_14984);
nand UO_1488 (O_1488,N_14884,N_14837);
and UO_1489 (O_1489,N_14787,N_14736);
and UO_1490 (O_1490,N_14763,N_14715);
and UO_1491 (O_1491,N_14769,N_14832);
xnor UO_1492 (O_1492,N_14737,N_14922);
nor UO_1493 (O_1493,N_14804,N_14985);
or UO_1494 (O_1494,N_14970,N_14950);
or UO_1495 (O_1495,N_14977,N_14980);
xnor UO_1496 (O_1496,N_14722,N_14744);
and UO_1497 (O_1497,N_14896,N_14754);
xor UO_1498 (O_1498,N_14968,N_14821);
or UO_1499 (O_1499,N_14745,N_14950);
xor UO_1500 (O_1500,N_14983,N_14991);
or UO_1501 (O_1501,N_14906,N_14999);
xnor UO_1502 (O_1502,N_14953,N_14851);
nand UO_1503 (O_1503,N_14738,N_14782);
xor UO_1504 (O_1504,N_14720,N_14781);
nor UO_1505 (O_1505,N_14840,N_14766);
and UO_1506 (O_1506,N_14944,N_14987);
or UO_1507 (O_1507,N_14932,N_14738);
nor UO_1508 (O_1508,N_14957,N_14933);
xnor UO_1509 (O_1509,N_14850,N_14782);
nor UO_1510 (O_1510,N_14860,N_14902);
and UO_1511 (O_1511,N_14776,N_14845);
and UO_1512 (O_1512,N_14888,N_14891);
and UO_1513 (O_1513,N_14936,N_14839);
or UO_1514 (O_1514,N_14762,N_14744);
xnor UO_1515 (O_1515,N_14736,N_14754);
nand UO_1516 (O_1516,N_14965,N_14772);
nor UO_1517 (O_1517,N_14866,N_14753);
nor UO_1518 (O_1518,N_14826,N_14973);
nor UO_1519 (O_1519,N_14770,N_14941);
nor UO_1520 (O_1520,N_14823,N_14887);
xor UO_1521 (O_1521,N_14916,N_14860);
nand UO_1522 (O_1522,N_14716,N_14972);
or UO_1523 (O_1523,N_14924,N_14750);
xor UO_1524 (O_1524,N_14851,N_14961);
and UO_1525 (O_1525,N_14968,N_14728);
nand UO_1526 (O_1526,N_14949,N_14858);
and UO_1527 (O_1527,N_14907,N_14972);
nand UO_1528 (O_1528,N_14732,N_14828);
or UO_1529 (O_1529,N_14719,N_14815);
nand UO_1530 (O_1530,N_14700,N_14733);
nand UO_1531 (O_1531,N_14896,N_14712);
xor UO_1532 (O_1532,N_14860,N_14719);
or UO_1533 (O_1533,N_14874,N_14716);
nor UO_1534 (O_1534,N_14784,N_14976);
or UO_1535 (O_1535,N_14834,N_14877);
or UO_1536 (O_1536,N_14720,N_14747);
and UO_1537 (O_1537,N_14923,N_14844);
and UO_1538 (O_1538,N_14830,N_14897);
or UO_1539 (O_1539,N_14802,N_14774);
and UO_1540 (O_1540,N_14935,N_14916);
xor UO_1541 (O_1541,N_14794,N_14941);
nor UO_1542 (O_1542,N_14761,N_14775);
and UO_1543 (O_1543,N_14776,N_14989);
nor UO_1544 (O_1544,N_14980,N_14939);
and UO_1545 (O_1545,N_14929,N_14706);
nor UO_1546 (O_1546,N_14898,N_14897);
and UO_1547 (O_1547,N_14709,N_14734);
nor UO_1548 (O_1548,N_14803,N_14888);
nor UO_1549 (O_1549,N_14822,N_14727);
nor UO_1550 (O_1550,N_14829,N_14895);
nor UO_1551 (O_1551,N_14966,N_14856);
nor UO_1552 (O_1552,N_14930,N_14710);
and UO_1553 (O_1553,N_14784,N_14986);
or UO_1554 (O_1554,N_14717,N_14864);
and UO_1555 (O_1555,N_14704,N_14760);
nand UO_1556 (O_1556,N_14944,N_14913);
or UO_1557 (O_1557,N_14734,N_14702);
nor UO_1558 (O_1558,N_14920,N_14766);
nor UO_1559 (O_1559,N_14973,N_14948);
and UO_1560 (O_1560,N_14733,N_14956);
or UO_1561 (O_1561,N_14917,N_14949);
xnor UO_1562 (O_1562,N_14932,N_14823);
xor UO_1563 (O_1563,N_14875,N_14907);
xor UO_1564 (O_1564,N_14762,N_14941);
and UO_1565 (O_1565,N_14814,N_14806);
nand UO_1566 (O_1566,N_14748,N_14939);
or UO_1567 (O_1567,N_14965,N_14767);
xor UO_1568 (O_1568,N_14947,N_14883);
or UO_1569 (O_1569,N_14794,N_14801);
and UO_1570 (O_1570,N_14835,N_14745);
nand UO_1571 (O_1571,N_14907,N_14988);
and UO_1572 (O_1572,N_14774,N_14964);
nor UO_1573 (O_1573,N_14855,N_14759);
and UO_1574 (O_1574,N_14859,N_14791);
xor UO_1575 (O_1575,N_14780,N_14820);
xnor UO_1576 (O_1576,N_14918,N_14747);
nand UO_1577 (O_1577,N_14705,N_14970);
nor UO_1578 (O_1578,N_14955,N_14784);
or UO_1579 (O_1579,N_14866,N_14942);
and UO_1580 (O_1580,N_14908,N_14749);
xor UO_1581 (O_1581,N_14890,N_14823);
nor UO_1582 (O_1582,N_14749,N_14706);
or UO_1583 (O_1583,N_14934,N_14799);
xor UO_1584 (O_1584,N_14885,N_14857);
nand UO_1585 (O_1585,N_14709,N_14838);
and UO_1586 (O_1586,N_14781,N_14978);
or UO_1587 (O_1587,N_14847,N_14782);
and UO_1588 (O_1588,N_14852,N_14937);
nand UO_1589 (O_1589,N_14721,N_14954);
nand UO_1590 (O_1590,N_14729,N_14812);
and UO_1591 (O_1591,N_14849,N_14728);
nor UO_1592 (O_1592,N_14902,N_14702);
nor UO_1593 (O_1593,N_14974,N_14893);
nand UO_1594 (O_1594,N_14757,N_14984);
or UO_1595 (O_1595,N_14910,N_14793);
nand UO_1596 (O_1596,N_14892,N_14913);
nor UO_1597 (O_1597,N_14748,N_14816);
or UO_1598 (O_1598,N_14775,N_14747);
or UO_1599 (O_1599,N_14708,N_14729);
xor UO_1600 (O_1600,N_14914,N_14955);
nand UO_1601 (O_1601,N_14836,N_14770);
nor UO_1602 (O_1602,N_14888,N_14898);
or UO_1603 (O_1603,N_14733,N_14853);
or UO_1604 (O_1604,N_14836,N_14944);
or UO_1605 (O_1605,N_14705,N_14908);
or UO_1606 (O_1606,N_14832,N_14750);
or UO_1607 (O_1607,N_14813,N_14747);
xnor UO_1608 (O_1608,N_14762,N_14823);
and UO_1609 (O_1609,N_14886,N_14811);
xnor UO_1610 (O_1610,N_14987,N_14992);
nor UO_1611 (O_1611,N_14973,N_14966);
xor UO_1612 (O_1612,N_14701,N_14811);
or UO_1613 (O_1613,N_14944,N_14731);
nand UO_1614 (O_1614,N_14820,N_14722);
nand UO_1615 (O_1615,N_14767,N_14927);
nor UO_1616 (O_1616,N_14965,N_14992);
nor UO_1617 (O_1617,N_14729,N_14801);
xnor UO_1618 (O_1618,N_14944,N_14964);
and UO_1619 (O_1619,N_14935,N_14918);
or UO_1620 (O_1620,N_14740,N_14994);
nor UO_1621 (O_1621,N_14905,N_14949);
xor UO_1622 (O_1622,N_14938,N_14778);
nand UO_1623 (O_1623,N_14794,N_14896);
or UO_1624 (O_1624,N_14791,N_14731);
xor UO_1625 (O_1625,N_14845,N_14952);
nand UO_1626 (O_1626,N_14756,N_14715);
xnor UO_1627 (O_1627,N_14986,N_14773);
nor UO_1628 (O_1628,N_14721,N_14819);
or UO_1629 (O_1629,N_14753,N_14871);
nand UO_1630 (O_1630,N_14774,N_14894);
nor UO_1631 (O_1631,N_14990,N_14846);
or UO_1632 (O_1632,N_14789,N_14957);
nand UO_1633 (O_1633,N_14772,N_14723);
nor UO_1634 (O_1634,N_14806,N_14905);
xor UO_1635 (O_1635,N_14841,N_14953);
xor UO_1636 (O_1636,N_14732,N_14881);
or UO_1637 (O_1637,N_14774,N_14863);
and UO_1638 (O_1638,N_14849,N_14778);
and UO_1639 (O_1639,N_14731,N_14730);
nand UO_1640 (O_1640,N_14826,N_14910);
xnor UO_1641 (O_1641,N_14902,N_14730);
nor UO_1642 (O_1642,N_14949,N_14915);
nand UO_1643 (O_1643,N_14878,N_14728);
xnor UO_1644 (O_1644,N_14888,N_14832);
and UO_1645 (O_1645,N_14771,N_14859);
nor UO_1646 (O_1646,N_14817,N_14854);
or UO_1647 (O_1647,N_14976,N_14712);
nand UO_1648 (O_1648,N_14718,N_14871);
nor UO_1649 (O_1649,N_14797,N_14925);
xor UO_1650 (O_1650,N_14974,N_14930);
and UO_1651 (O_1651,N_14746,N_14790);
nand UO_1652 (O_1652,N_14701,N_14820);
and UO_1653 (O_1653,N_14998,N_14813);
nand UO_1654 (O_1654,N_14859,N_14935);
and UO_1655 (O_1655,N_14898,N_14893);
and UO_1656 (O_1656,N_14925,N_14790);
xnor UO_1657 (O_1657,N_14903,N_14884);
or UO_1658 (O_1658,N_14908,N_14751);
and UO_1659 (O_1659,N_14772,N_14818);
nor UO_1660 (O_1660,N_14996,N_14826);
and UO_1661 (O_1661,N_14988,N_14736);
nand UO_1662 (O_1662,N_14779,N_14855);
and UO_1663 (O_1663,N_14767,N_14785);
or UO_1664 (O_1664,N_14919,N_14779);
and UO_1665 (O_1665,N_14702,N_14724);
xor UO_1666 (O_1666,N_14858,N_14722);
xor UO_1667 (O_1667,N_14757,N_14772);
nor UO_1668 (O_1668,N_14895,N_14971);
nand UO_1669 (O_1669,N_14864,N_14798);
nand UO_1670 (O_1670,N_14942,N_14725);
xor UO_1671 (O_1671,N_14708,N_14771);
xnor UO_1672 (O_1672,N_14834,N_14797);
nor UO_1673 (O_1673,N_14815,N_14752);
xnor UO_1674 (O_1674,N_14910,N_14947);
nor UO_1675 (O_1675,N_14873,N_14844);
or UO_1676 (O_1676,N_14750,N_14933);
and UO_1677 (O_1677,N_14985,N_14708);
and UO_1678 (O_1678,N_14968,N_14973);
xor UO_1679 (O_1679,N_14809,N_14741);
xnor UO_1680 (O_1680,N_14882,N_14923);
nor UO_1681 (O_1681,N_14923,N_14888);
and UO_1682 (O_1682,N_14770,N_14993);
xor UO_1683 (O_1683,N_14877,N_14861);
and UO_1684 (O_1684,N_14775,N_14746);
and UO_1685 (O_1685,N_14799,N_14988);
nor UO_1686 (O_1686,N_14742,N_14737);
or UO_1687 (O_1687,N_14782,N_14723);
nor UO_1688 (O_1688,N_14901,N_14730);
xnor UO_1689 (O_1689,N_14862,N_14768);
nand UO_1690 (O_1690,N_14981,N_14747);
or UO_1691 (O_1691,N_14944,N_14815);
or UO_1692 (O_1692,N_14788,N_14879);
xor UO_1693 (O_1693,N_14926,N_14740);
nor UO_1694 (O_1694,N_14729,N_14762);
nand UO_1695 (O_1695,N_14835,N_14710);
nor UO_1696 (O_1696,N_14880,N_14852);
nand UO_1697 (O_1697,N_14961,N_14700);
or UO_1698 (O_1698,N_14966,N_14964);
nor UO_1699 (O_1699,N_14932,N_14852);
nand UO_1700 (O_1700,N_14810,N_14953);
nor UO_1701 (O_1701,N_14745,N_14724);
nand UO_1702 (O_1702,N_14814,N_14921);
nor UO_1703 (O_1703,N_14809,N_14862);
nor UO_1704 (O_1704,N_14877,N_14993);
and UO_1705 (O_1705,N_14744,N_14969);
nor UO_1706 (O_1706,N_14716,N_14830);
nand UO_1707 (O_1707,N_14991,N_14921);
xor UO_1708 (O_1708,N_14975,N_14954);
or UO_1709 (O_1709,N_14837,N_14953);
nand UO_1710 (O_1710,N_14877,N_14954);
nand UO_1711 (O_1711,N_14931,N_14739);
and UO_1712 (O_1712,N_14980,N_14707);
xnor UO_1713 (O_1713,N_14776,N_14986);
xor UO_1714 (O_1714,N_14816,N_14812);
nor UO_1715 (O_1715,N_14829,N_14928);
xnor UO_1716 (O_1716,N_14796,N_14748);
and UO_1717 (O_1717,N_14899,N_14987);
nand UO_1718 (O_1718,N_14728,N_14708);
nand UO_1719 (O_1719,N_14959,N_14975);
xnor UO_1720 (O_1720,N_14725,N_14930);
nand UO_1721 (O_1721,N_14904,N_14723);
nor UO_1722 (O_1722,N_14802,N_14892);
or UO_1723 (O_1723,N_14938,N_14839);
xor UO_1724 (O_1724,N_14951,N_14781);
nor UO_1725 (O_1725,N_14827,N_14897);
nor UO_1726 (O_1726,N_14860,N_14742);
and UO_1727 (O_1727,N_14702,N_14789);
and UO_1728 (O_1728,N_14988,N_14994);
nand UO_1729 (O_1729,N_14979,N_14742);
or UO_1730 (O_1730,N_14788,N_14827);
nor UO_1731 (O_1731,N_14816,N_14786);
nor UO_1732 (O_1732,N_14945,N_14837);
and UO_1733 (O_1733,N_14803,N_14885);
and UO_1734 (O_1734,N_14722,N_14728);
nor UO_1735 (O_1735,N_14752,N_14746);
or UO_1736 (O_1736,N_14708,N_14746);
xnor UO_1737 (O_1737,N_14906,N_14844);
nand UO_1738 (O_1738,N_14820,N_14946);
nor UO_1739 (O_1739,N_14802,N_14872);
nor UO_1740 (O_1740,N_14930,N_14736);
and UO_1741 (O_1741,N_14948,N_14844);
nor UO_1742 (O_1742,N_14859,N_14795);
xnor UO_1743 (O_1743,N_14989,N_14888);
nor UO_1744 (O_1744,N_14764,N_14841);
xnor UO_1745 (O_1745,N_14896,N_14959);
nand UO_1746 (O_1746,N_14865,N_14966);
and UO_1747 (O_1747,N_14783,N_14855);
or UO_1748 (O_1748,N_14795,N_14754);
and UO_1749 (O_1749,N_14943,N_14720);
and UO_1750 (O_1750,N_14946,N_14700);
nand UO_1751 (O_1751,N_14863,N_14919);
nand UO_1752 (O_1752,N_14812,N_14865);
or UO_1753 (O_1753,N_14829,N_14858);
or UO_1754 (O_1754,N_14717,N_14753);
and UO_1755 (O_1755,N_14892,N_14710);
nor UO_1756 (O_1756,N_14776,N_14761);
nor UO_1757 (O_1757,N_14995,N_14747);
or UO_1758 (O_1758,N_14745,N_14737);
nand UO_1759 (O_1759,N_14884,N_14995);
or UO_1760 (O_1760,N_14711,N_14929);
or UO_1761 (O_1761,N_14782,N_14943);
nor UO_1762 (O_1762,N_14877,N_14836);
and UO_1763 (O_1763,N_14738,N_14990);
and UO_1764 (O_1764,N_14948,N_14822);
or UO_1765 (O_1765,N_14958,N_14965);
nand UO_1766 (O_1766,N_14887,N_14938);
or UO_1767 (O_1767,N_14845,N_14929);
or UO_1768 (O_1768,N_14846,N_14777);
nand UO_1769 (O_1769,N_14808,N_14793);
nor UO_1770 (O_1770,N_14860,N_14704);
and UO_1771 (O_1771,N_14897,N_14769);
xor UO_1772 (O_1772,N_14736,N_14927);
nand UO_1773 (O_1773,N_14816,N_14847);
and UO_1774 (O_1774,N_14908,N_14732);
nor UO_1775 (O_1775,N_14727,N_14854);
xor UO_1776 (O_1776,N_14742,N_14800);
or UO_1777 (O_1777,N_14868,N_14816);
nor UO_1778 (O_1778,N_14980,N_14968);
or UO_1779 (O_1779,N_14755,N_14928);
nor UO_1780 (O_1780,N_14973,N_14728);
nor UO_1781 (O_1781,N_14857,N_14734);
and UO_1782 (O_1782,N_14870,N_14781);
or UO_1783 (O_1783,N_14929,N_14872);
xor UO_1784 (O_1784,N_14910,N_14899);
nand UO_1785 (O_1785,N_14795,N_14727);
and UO_1786 (O_1786,N_14713,N_14857);
and UO_1787 (O_1787,N_14830,N_14978);
nor UO_1788 (O_1788,N_14975,N_14948);
and UO_1789 (O_1789,N_14783,N_14931);
or UO_1790 (O_1790,N_14826,N_14870);
or UO_1791 (O_1791,N_14964,N_14815);
nand UO_1792 (O_1792,N_14972,N_14779);
xor UO_1793 (O_1793,N_14844,N_14778);
nand UO_1794 (O_1794,N_14701,N_14935);
xor UO_1795 (O_1795,N_14844,N_14837);
and UO_1796 (O_1796,N_14805,N_14863);
nor UO_1797 (O_1797,N_14853,N_14734);
nor UO_1798 (O_1798,N_14700,N_14914);
nor UO_1799 (O_1799,N_14836,N_14735);
or UO_1800 (O_1800,N_14701,N_14934);
nand UO_1801 (O_1801,N_14880,N_14770);
nand UO_1802 (O_1802,N_14828,N_14811);
nand UO_1803 (O_1803,N_14876,N_14783);
nand UO_1804 (O_1804,N_14850,N_14911);
nor UO_1805 (O_1805,N_14975,N_14947);
xor UO_1806 (O_1806,N_14963,N_14885);
nand UO_1807 (O_1807,N_14825,N_14789);
nor UO_1808 (O_1808,N_14878,N_14979);
nand UO_1809 (O_1809,N_14904,N_14873);
xor UO_1810 (O_1810,N_14914,N_14839);
and UO_1811 (O_1811,N_14945,N_14701);
nand UO_1812 (O_1812,N_14728,N_14949);
xnor UO_1813 (O_1813,N_14746,N_14979);
and UO_1814 (O_1814,N_14964,N_14703);
and UO_1815 (O_1815,N_14710,N_14913);
nand UO_1816 (O_1816,N_14954,N_14762);
nand UO_1817 (O_1817,N_14922,N_14723);
xor UO_1818 (O_1818,N_14903,N_14897);
and UO_1819 (O_1819,N_14908,N_14782);
nand UO_1820 (O_1820,N_14964,N_14891);
and UO_1821 (O_1821,N_14929,N_14703);
nand UO_1822 (O_1822,N_14747,N_14988);
nor UO_1823 (O_1823,N_14755,N_14979);
or UO_1824 (O_1824,N_14850,N_14827);
and UO_1825 (O_1825,N_14962,N_14814);
xnor UO_1826 (O_1826,N_14848,N_14722);
nor UO_1827 (O_1827,N_14850,N_14882);
nand UO_1828 (O_1828,N_14869,N_14843);
xor UO_1829 (O_1829,N_14928,N_14797);
xor UO_1830 (O_1830,N_14908,N_14722);
or UO_1831 (O_1831,N_14915,N_14869);
nor UO_1832 (O_1832,N_14882,N_14751);
or UO_1833 (O_1833,N_14730,N_14712);
and UO_1834 (O_1834,N_14897,N_14976);
xor UO_1835 (O_1835,N_14952,N_14976);
nand UO_1836 (O_1836,N_14726,N_14932);
nand UO_1837 (O_1837,N_14731,N_14747);
nand UO_1838 (O_1838,N_14993,N_14711);
and UO_1839 (O_1839,N_14967,N_14976);
and UO_1840 (O_1840,N_14912,N_14717);
nor UO_1841 (O_1841,N_14916,N_14717);
and UO_1842 (O_1842,N_14869,N_14929);
xor UO_1843 (O_1843,N_14727,N_14871);
and UO_1844 (O_1844,N_14962,N_14850);
or UO_1845 (O_1845,N_14845,N_14974);
and UO_1846 (O_1846,N_14926,N_14979);
nor UO_1847 (O_1847,N_14892,N_14799);
or UO_1848 (O_1848,N_14858,N_14916);
nor UO_1849 (O_1849,N_14835,N_14859);
and UO_1850 (O_1850,N_14843,N_14711);
nand UO_1851 (O_1851,N_14817,N_14753);
nor UO_1852 (O_1852,N_14793,N_14712);
and UO_1853 (O_1853,N_14973,N_14712);
nand UO_1854 (O_1854,N_14957,N_14992);
and UO_1855 (O_1855,N_14825,N_14891);
nor UO_1856 (O_1856,N_14936,N_14785);
nor UO_1857 (O_1857,N_14747,N_14889);
xnor UO_1858 (O_1858,N_14969,N_14977);
nand UO_1859 (O_1859,N_14917,N_14814);
nand UO_1860 (O_1860,N_14701,N_14933);
and UO_1861 (O_1861,N_14930,N_14921);
nand UO_1862 (O_1862,N_14735,N_14962);
and UO_1863 (O_1863,N_14868,N_14805);
and UO_1864 (O_1864,N_14779,N_14865);
xor UO_1865 (O_1865,N_14917,N_14994);
nor UO_1866 (O_1866,N_14805,N_14836);
xor UO_1867 (O_1867,N_14998,N_14838);
nand UO_1868 (O_1868,N_14924,N_14799);
xnor UO_1869 (O_1869,N_14709,N_14792);
or UO_1870 (O_1870,N_14817,N_14938);
xnor UO_1871 (O_1871,N_14767,N_14764);
or UO_1872 (O_1872,N_14941,N_14760);
nand UO_1873 (O_1873,N_14904,N_14906);
and UO_1874 (O_1874,N_14967,N_14773);
xnor UO_1875 (O_1875,N_14857,N_14766);
or UO_1876 (O_1876,N_14770,N_14908);
or UO_1877 (O_1877,N_14976,N_14844);
and UO_1878 (O_1878,N_14878,N_14783);
nor UO_1879 (O_1879,N_14977,N_14962);
or UO_1880 (O_1880,N_14831,N_14947);
or UO_1881 (O_1881,N_14802,N_14911);
nand UO_1882 (O_1882,N_14740,N_14721);
nand UO_1883 (O_1883,N_14933,N_14854);
nor UO_1884 (O_1884,N_14757,N_14874);
or UO_1885 (O_1885,N_14906,N_14948);
nand UO_1886 (O_1886,N_14834,N_14874);
and UO_1887 (O_1887,N_14785,N_14920);
and UO_1888 (O_1888,N_14978,N_14792);
and UO_1889 (O_1889,N_14885,N_14739);
or UO_1890 (O_1890,N_14795,N_14780);
or UO_1891 (O_1891,N_14902,N_14818);
nand UO_1892 (O_1892,N_14934,N_14912);
or UO_1893 (O_1893,N_14883,N_14780);
and UO_1894 (O_1894,N_14764,N_14807);
nor UO_1895 (O_1895,N_14775,N_14878);
or UO_1896 (O_1896,N_14782,N_14954);
nand UO_1897 (O_1897,N_14954,N_14897);
xor UO_1898 (O_1898,N_14941,N_14849);
nor UO_1899 (O_1899,N_14701,N_14918);
nand UO_1900 (O_1900,N_14830,N_14888);
or UO_1901 (O_1901,N_14755,N_14813);
xnor UO_1902 (O_1902,N_14754,N_14884);
or UO_1903 (O_1903,N_14983,N_14915);
nand UO_1904 (O_1904,N_14725,N_14823);
nand UO_1905 (O_1905,N_14857,N_14811);
nand UO_1906 (O_1906,N_14957,N_14749);
nor UO_1907 (O_1907,N_14715,N_14788);
nand UO_1908 (O_1908,N_14825,N_14921);
nand UO_1909 (O_1909,N_14723,N_14916);
or UO_1910 (O_1910,N_14749,N_14790);
nor UO_1911 (O_1911,N_14902,N_14755);
nand UO_1912 (O_1912,N_14709,N_14991);
nand UO_1913 (O_1913,N_14875,N_14960);
nand UO_1914 (O_1914,N_14775,N_14703);
nor UO_1915 (O_1915,N_14737,N_14862);
and UO_1916 (O_1916,N_14869,N_14973);
xor UO_1917 (O_1917,N_14788,N_14753);
nor UO_1918 (O_1918,N_14787,N_14836);
or UO_1919 (O_1919,N_14747,N_14727);
xnor UO_1920 (O_1920,N_14810,N_14779);
nand UO_1921 (O_1921,N_14815,N_14726);
nand UO_1922 (O_1922,N_14739,N_14941);
nor UO_1923 (O_1923,N_14730,N_14828);
xor UO_1924 (O_1924,N_14783,N_14888);
nand UO_1925 (O_1925,N_14878,N_14872);
or UO_1926 (O_1926,N_14864,N_14794);
nor UO_1927 (O_1927,N_14800,N_14768);
or UO_1928 (O_1928,N_14833,N_14882);
xnor UO_1929 (O_1929,N_14737,N_14886);
xnor UO_1930 (O_1930,N_14915,N_14968);
nor UO_1931 (O_1931,N_14969,N_14869);
xor UO_1932 (O_1932,N_14939,N_14900);
nand UO_1933 (O_1933,N_14731,N_14708);
or UO_1934 (O_1934,N_14761,N_14712);
and UO_1935 (O_1935,N_14893,N_14881);
and UO_1936 (O_1936,N_14941,N_14884);
and UO_1937 (O_1937,N_14712,N_14786);
or UO_1938 (O_1938,N_14800,N_14969);
nor UO_1939 (O_1939,N_14903,N_14907);
xor UO_1940 (O_1940,N_14784,N_14817);
nor UO_1941 (O_1941,N_14728,N_14753);
and UO_1942 (O_1942,N_14727,N_14940);
nand UO_1943 (O_1943,N_14711,N_14876);
nand UO_1944 (O_1944,N_14756,N_14910);
xor UO_1945 (O_1945,N_14913,N_14729);
or UO_1946 (O_1946,N_14779,N_14729);
nand UO_1947 (O_1947,N_14717,N_14763);
or UO_1948 (O_1948,N_14752,N_14842);
nand UO_1949 (O_1949,N_14749,N_14888);
and UO_1950 (O_1950,N_14757,N_14816);
and UO_1951 (O_1951,N_14713,N_14984);
xor UO_1952 (O_1952,N_14969,N_14897);
and UO_1953 (O_1953,N_14922,N_14870);
xnor UO_1954 (O_1954,N_14773,N_14713);
xor UO_1955 (O_1955,N_14762,N_14981);
and UO_1956 (O_1956,N_14728,N_14923);
nor UO_1957 (O_1957,N_14785,N_14733);
or UO_1958 (O_1958,N_14895,N_14714);
and UO_1959 (O_1959,N_14785,N_14805);
nand UO_1960 (O_1960,N_14861,N_14916);
and UO_1961 (O_1961,N_14787,N_14887);
xor UO_1962 (O_1962,N_14975,N_14860);
nand UO_1963 (O_1963,N_14797,N_14857);
nor UO_1964 (O_1964,N_14994,N_14909);
xnor UO_1965 (O_1965,N_14797,N_14717);
or UO_1966 (O_1966,N_14882,N_14715);
and UO_1967 (O_1967,N_14929,N_14990);
and UO_1968 (O_1968,N_14890,N_14978);
xor UO_1969 (O_1969,N_14948,N_14773);
nor UO_1970 (O_1970,N_14923,N_14743);
and UO_1971 (O_1971,N_14821,N_14773);
or UO_1972 (O_1972,N_14731,N_14856);
xor UO_1973 (O_1973,N_14752,N_14934);
nor UO_1974 (O_1974,N_14965,N_14774);
and UO_1975 (O_1975,N_14899,N_14827);
or UO_1976 (O_1976,N_14997,N_14964);
and UO_1977 (O_1977,N_14996,N_14998);
xnor UO_1978 (O_1978,N_14754,N_14948);
and UO_1979 (O_1979,N_14993,N_14781);
and UO_1980 (O_1980,N_14844,N_14805);
and UO_1981 (O_1981,N_14896,N_14844);
nor UO_1982 (O_1982,N_14727,N_14730);
and UO_1983 (O_1983,N_14886,N_14801);
nor UO_1984 (O_1984,N_14976,N_14783);
nand UO_1985 (O_1985,N_14869,N_14762);
nor UO_1986 (O_1986,N_14994,N_14722);
or UO_1987 (O_1987,N_14707,N_14868);
and UO_1988 (O_1988,N_14868,N_14748);
and UO_1989 (O_1989,N_14897,N_14823);
and UO_1990 (O_1990,N_14832,N_14755);
and UO_1991 (O_1991,N_14848,N_14887);
and UO_1992 (O_1992,N_14829,N_14713);
xor UO_1993 (O_1993,N_14954,N_14967);
and UO_1994 (O_1994,N_14793,N_14730);
xor UO_1995 (O_1995,N_14915,N_14809);
and UO_1996 (O_1996,N_14720,N_14713);
or UO_1997 (O_1997,N_14777,N_14944);
nand UO_1998 (O_1998,N_14939,N_14824);
and UO_1999 (O_1999,N_14961,N_14905);
endmodule